
module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, NorthIn, SouthIn, 
    EastIn, WestIn, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] SouthIn;
input  [7:0] ScanIn;
output [7:0] Out;
output [7:0] ScanOut;
input  [7:0] NorthIn;
input  [7:0] WestIn;
input  [7:0] EastIn;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[7] , \ScanOut[5]1 , \ScanOut[4]1 , n185, n182, \ScanOut[1]1 , 
        n184, \ScanOut[0]1 , n183, \ScanOut[6]1 , \ScanOut[3]1 , n176, 
        \ScanOut[2]1 , n181, n186, n178, n179, n177, n180;
    assign ScanOut[7] = \ScanOut[7] ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[7] = \ScanOut[7] ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO22 U28 ( .A(ScanIn[1]), .B(n176), .C(\ScanOut[1]1 ), .D(n177), .Z(
        n185) );
    VMW_AO22 U33 ( .A(ScanIn[6]), .B(n176), .C(\ScanOut[6]1 ), .D(n177), .Z(
        n180) );
    VMW_AO22 U34 ( .A(ScanIn[7]), .B(n176), .C(\ScanOut[7] ), .D(n177), .Z(
        n179) );
    VMW_NOR2 U35 ( .A(ScanEnable), .B(Reset), .Z(n177) );
    VMW_AO22 U27 ( .A(ScanIn[0]), .B(n176), .C(\ScanOut[0]1 ), .D(n177), .Z(
        n186) );
    VMW_FD \Out_reg[5]  ( .D(n181), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO22 U29 ( .A(ScanIn[2]), .B(n176), .C(\ScanOut[2]1 ), .D(n177), .Z(
        n184) );
    VMW_FD \Out_reg[7]  ( .D(n179), .CP(Clk), .Q(\ScanOut[7] ) );
    VMW_FD \Out_reg[3]  ( .D(n183), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n185), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_AO22 U32 ( .A(ScanIn[5]), .B(n176), .C(\ScanOut[5]1 ), .D(n177), .Z(
        n181) );
    VMW_AO22 U30 ( .A(ScanIn[3]), .B(n176), .C(\ScanOut[3]1 ), .D(n177), .Z(
        n183) );
    VMW_FD \Out_reg[6]  ( .D(n180), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U31 ( .A(ScanIn[4]), .B(n176), .C(\ScanOut[4]1 ), .D(n177), .Z(
        n182) );
    VMW_NOR2 U36 ( .A(n178), .B(Reset), .Z(n176) );
    VMW_INV U37 ( .A(ScanEnable), .Z(n178) );
    VMW_FD \Out_reg[2]  ( .D(n184), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_FD \Out_reg[4]  ( .D(n182), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n186), .CP(Clk), .Q(\ScanOut[0]1 ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_2 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n1, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_1 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_AND2 U1 ( .A(A[0]), .B(B[0]), .Z(\carry[1] ) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .CO(\carry[2] ) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .CO(\carry[7] ), .S(
        SUM[6]) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .CO(\carry[3] ), .S(
        SUM[2]) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .CO(\carry[4] ), .S(
        SUM[3]) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .CO(\carry[5] ), .S(
        SUM[4]) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .CO(\carry[6] ), .S(
        SUM[5]) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_0 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n3, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n3) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n3), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, NorthIn, SouthIn, 
    EastIn, WestIn, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] SouthIn;
input  [7:0] ScanIn;
output [7:0] Out;
output [7:0] ScanOut;
input  [7:0] NorthIn;
input  [7:0] WestIn;
input  [7:0] EastIn;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[7] , \ScanOut[5]1 , \ScanOut[4]1 , n222, n217, n225, n219, 
        n210, \ScanOut[6]1 , n224, \a184[4] , \n161[4] , \ScanOut[1]1 , n218, 
        \n158[4] , \ScanOut[0]1 , n211, n216, \n158[2] , n223, \n161[2] , 
        \n158[6] , \a184[6] , \n161[6] , \ScanOut[3]1 , \n158[7] , n214, 
        \n161[7] , \a184[7] , n206, n221, \n158[3] , \ScanOut[2]1 , \a184[3] , 
        \n161[3] , \n161[1] , \n158[8] , n226, \a184[8] , \n161[8] , \n158[1] , 
        n213, \a184[5] , n208, \n161[5] , \n158[5] , n209, n212, n215, n207, 
        n220;
    wire UNCONNECTED_1 , UNCONNECTED_2 ;
    assign ScanOut[7] = \ScanOut[7] ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[7] = \ScanOut[7] ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO21 U33 ( .A(\ScanOut[0]1 ), .B(n206), .C(n207), .Z(n223) );
    VMW_AO21 U34 ( .A(\ScanOut[1]1 ), .B(n206), .C(n208), .Z(n222) );
    VMW_NOR2 U41 ( .A(n214), .B(Reset), .Z(n213) );
    VMW_AO22 U46 ( .A(ScanIn[3]), .B(n213), .C(\a184[6] ), .D(n215), .Z(n210)
         );
    VMW_AO21 U35 ( .A(\ScanOut[2]1 ), .B(n206), .C(n209), .Z(n221) );
    VMW_AO22 U48 ( .A(ScanIn[1]), .B(n213), .C(\a184[4] ), .D(n215), .Z(n208)
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_1 add_98 ( .A({
        \n158[1] , \n158[2] , \n158[3] , \n158[4] , \n158[5] , \n158[6] , 
        \n158[7] , \n158[8] }), .B(WestIn), .CI(n225), .SUM({\a184[8] , 
        \a184[7] , \a184[6] , \a184[5] , \a184[4] , \a184[3] , UNCONNECTED_1, 
        UNCONNECTED_2}) );
    VMW_PULLDOWN U32 ( .Z(n224) );
    VMW_AO22 U40 ( .A(\ScanOut[7] ), .B(n206), .C(ScanIn[7]), .D(n213), .Z(
        n216) );
    VMW_FD \Out_reg[5]  ( .D(n218), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO22 U47 ( .A(ScanIn[2]), .B(n213), .C(\a184[5] ), .D(n215), .Z(n209)
         );
    VMW_AO22 U49 ( .A(ScanIn[0]), .B(n213), .C(\a184[3] ), .D(n215), .Z(n207)
         );
    VMW_FD \Out_reg[1]  ( .D(n222), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_FD \Out_reg[7]  ( .D(n216), .CP(Clk), .Q(\ScanOut[7] ) );
    VMW_FD \Out_reg[3]  ( .D(n220), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_PULLDOWN U30 ( .Z(n225) );
    VMW_AO22 U39 ( .A(\ScanOut[6]1 ), .B(n206), .C(ScanIn[6]), .D(n213), .Z(
        n217) );
    VMW_FD \Out_reg[6]  ( .D(n217), .CP(Clk), .Q(\ScanOut[6]1 ) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_0 add_98_2 ( .A(
        NorthIn), .B(SouthIn), .CI(n224), .SUM({\n161[1] , \n161[2] , 
        \n161[3] , \n161[4] , \n161[5] , \n161[6] , \n161[7] , \n161[8] }) );
    VMW_PULLDOWN U31 ( .Z(n226) );
    VMW_AO21 U36 ( .A(\ScanOut[3]1 ), .B(n206), .C(n210), .Z(n220) );
    VMW_AO21 U37 ( .A(\ScanOut[4]1 ), .B(n206), .C(n211), .Z(n219) );
    VMW_NOR3 U42 ( .A(ScanEnable), .B(Reset), .C(Enable), .Z(n206) );
    VMW_AO22 U45 ( .A(ScanIn[4]), .B(n213), .C(\a184[7] ), .D(n215), .Z(n211)
         );
    VMW_FD \Out_reg[2]  ( .D(n221), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_INV U50 ( .A(ScanEnable), .Z(n214) );
    VMW_FD \Out_reg[4]  ( .D(n219), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n223), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_AO21 U38 ( .A(\ScanOut[5]1 ), .B(n206), .C(n212), .Z(n218) );
    VMW_NOR3 U43 ( .A(Reset), .B(ScanEnable), .C(n206), .Z(n215) );
    VMW_AO22 U44 ( .A(ScanIn[5]), .B(n213), .C(\a184[8] ), .D(n215), .Z(n212)
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_2 add_98_1 ( .A({
        \n161[1] , \n161[2] , \n161[3] , \n161[4] , \n161[5] , \n161[6] , 
        \n161[7] , \n161[8] }), .B(EastIn), .CI(n226), .SUM({\n158[1] , 
        \n158[2] , \n158[3] , \n158[4] , \n158[5] , \n158[6] , \n158[7] , 
        \n158[8] }) );
endmodule


module Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 ( A, SUM );
input  [6:0] A;
output [6:0] SUM;
    wire n5, n9, n7, n12, n6, n13, n8, n10, n11;
    VMW_AO21 U3 ( .A(n5), .B(A[2]), .C(n6), .Z(SUM[2]) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(n9), .Z(SUM[1]) );
    VMW_INV U6 ( .A(A[0]), .Z(SUM[0]) );
    VMW_AO22 U14 ( .A(A[5]), .B(n13), .C(n12), .D(n10), .Z(SUM[5]) );
    VMW_AO21 U7 ( .A(n8), .B(A[4]), .C(n10), .Z(SUM[4]) );
    VMW_AND2 U8 ( .A(n10), .B(n12), .Z(n11) );
    VMW_XOR2 U13 ( .A(A[6]), .B(n11), .Z(SUM[6]) );
    VMW_OR2 U9 ( .A(A[0]), .B(A[1]), .Z(n5) );
    VMW_NOR2 U12 ( .A(n8), .B(A[4]), .Z(n10) );
    VMW_INV U15 ( .A(A[5]), .Z(n12) );
    VMW_INV U17 ( .A(A[3]), .Z(n7) );
    VMW_NOR2 U10 ( .A(n5), .B(A[2]), .Z(n6) );
    VMW_NAND2 U11 ( .A(n6), .B(n7), .Z(n8) );
    VMW_OAI21 U4 ( .A(n6), .B(n7), .C(n8), .Z(SUM[3]) );
    VMW_INV U18 ( .A(n5), .Z(n9) );
    VMW_INV U16 ( .A(n10), .Z(n13) );
endmodule


module Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, ScanId, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] ScanIn;
output [7:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire n379, \count[2] , n387, n362, n406, n395, \count[6] , n370, n389, 
        n408, n377, n392, \count[4] , n380, n401, n365, \count[0] , n393, n376, 
        \ScanReg[2] , n409, \count260[3] , n388, n364, n400, n381, 
        \ScanReg[6] , n386, n407, \ScanReg[4] , n363, \count260[5] , n378, 
        \count260[1] , \ScanReg[0] , n371, n394, \count260[0] , \ScanReg[1] , 
        \ScanReg[7] , n405, n384, \ScanReg[5] , \count260[4] , n396, n373, 
        n368, n374, \count260[6] , n383, n391, n410, n402, n366, n390, n398, 
        \count260[2] , \ScanReg[3] , n411, n375, \count[1] , n399, n367, n382, 
        n403, n385, \count[5] , n404, n369, \count[3] , n372, n397;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_PULLDOWN U54 ( .Z(n372) );
    VMW_PULLDOWN U73 ( .Z(n399) );
    VMW_INV U113 ( .A(n370), .Z(ScanEnable) );
    VMW_BUFIZ U134 ( .A(n393), .E(n377), .Z(\arr[3] ) );
    VMW_PULLDOWN U68 ( .Z(n391) );
    VMW_AND2 U96 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_AO22 U108 ( .A(\count[0] ), .B(n366), .C(\ScanReg[0] ), .D(n365), .Z(
        n373) );
    VMW_BUFIZ U141 ( .A(n400), .E(n377), .Z(\arr[18] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \count_reg[6]  ( .D(n405), .CP(Clk), .Q(\count[6] ) );
    VMW_PULLDOWN U61 ( .Z(n382) );
    VMW_AO22 U84 ( .A(ScanOut[4]), .B(n363), .C(\count260[4] ), .D(n364), .Z(
        n407) );
    VMW_FD \count_reg[2]  ( .D(n409), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_PULLDOWN U66 ( .Z(n389) );
    VMW_XNOR2 U101 ( .A(Addr[0]), .B(ScanId), .Z(n371) );
    VMW_AO22 U106 ( .A(\count[2] ), .B(n366), .C(\ScanReg[2] ), .D(n365), .Z(
        n388) );
    VMW_BUFIZ U121 ( .A(n380), .E(n377), .Z(\arr[14] ) );
    VMW_BUFIZ U126 ( .A(n385), .E(n377), .Z(\arr[31] ) );
    VMW_PULLDOWN U74 ( .Z(n400) );
    VMW_AO22 U83 ( .A(ScanOut[3]), .B(n363), .C(\count260[3] ), .D(n364), .Z(
        n408) );
    VMW_FD \count_reg[0]  ( .D(n411), .CP(Clk), .Q(\count[0] ) );
    VMW_NOR2 U91 ( .A(n367), .B(n368), .Z(n364) );
    VMW_AND2 U98 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_BUFIZ U128 ( .A(n387), .E(n377), .Z(\arr[28] ) );
    VMW_FD \count_reg[4]  ( .D(n407), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U114 ( .A(n372), .E(n377), .Z(\arr[19] ) );
    VMW_BUFIZ U133 ( .A(n392), .E(n377), .Z(\arr[20] ) );
    VMW_AND2 U99 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_PULLDOWN U55 ( .Z(n374) );
    VMW_PULLDOWN U67 ( .Z(n390) );
    VMW_AO22 U82 ( .A(ScanOut[2]), .B(n363), .C(\count260[2] ), .D(n364), .Z(
        n409) );
    VMW_AO22 U107 ( .A(\count[1] ), .B(n366), .C(\ScanReg[1] ), .D(n365), .Z(
        n403) );
    VMW_BUFIZ U120 ( .A(n379), .E(n377), .Z(\arr[27] ) );
    VMW_PULLDOWN U69 ( .Z(n392) );
    VMW_PULLDOWN U75 ( .Z(n401) );
    VMW_BUFIZ U115 ( .A(n373), .E(n377), .Z(\arr[0] ) );
    VMW_BUFIZ U132 ( .A(n391), .E(n377), .Z(\arr[29] ) );
    VMW_OAI21 U90 ( .A(n368), .B(Enable), .C(n369), .Z(n367) );
    VMW_OR4 U109 ( .A(\count[3] ), .B(\count[4] ), .C(\count[5] ), .D(
        \count[6] ), .Z(n362) );
    VMW_BUFIZ U129 ( .A(n388), .E(n377), .Z(\arr[2] ) );
    VMW_PULLDOWN U72 ( .Z(n398) );
    VMW_AND2 U97 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_BUFIZ U140 ( .A(n399), .E(n377), .Z(\arr[15] ) );
    VMW_INV U112 ( .A(Reset), .Z(n369) );
    VMW_BUFIZ U135 ( .A(n394), .E(n377), .Z(\arr[24] ) );
    VMW_PULLDOWN U60 ( .Z(n381) );
    VMW_AO22 U85 ( .A(ScanOut[5]), .B(n363), .C(\count260[5] ), .D(n364), .Z(
        n406) );
    VMW_OAI21 U100 ( .A(WR), .B(RD), .C(n371), .Z(n370) );
    VMW_BUFIZ U127 ( .A(n386), .E(n377), .Z(\arr[21] ) );
    VMW_PULLDOWN U56 ( .Z(n375) );
    VMW_PULLDOWN U57 ( .Z(n376) );
    VMW_BUFIZ U137 ( .A(n396), .E(n377), .Z(\arr[7] ) );
    VMW_PULLDOWN U58 ( .Z(n379) );
    VMW_PULLDOWN U59 ( .Z(n380) );
    VMW_PULLDOWN U62 ( .Z(n383) );
    VMW_PULLDOWN U70 ( .Z(n394) );
    VMW_AND2 U79 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_AND2 U95 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AND2 U110 ( .A(n366), .B(WR), .Z(n368) );
    VMW_BUFIZ U119 ( .A(n378), .E(n377), .Z(\arr[4] ) );
    VMW_BUFIZ U142 ( .A(n401), .E(n377), .Z(\arr[22] ) );
    VMW_AND2 U87 ( .A(\ScanReg[7] ), .B(n365), .Z(n396) );
    VMW_BUFIZ U125 ( .A(n384), .E(n377), .Z(\arr[6] ) );
    VMW_PULLDOWN U65 ( .Z(n387) );
    VMW_AO22 U102 ( .A(\count[6] ), .B(n366), .C(\ScanReg[6] ), .D(n365), .Z(
        n384) );
    VMW_AO22 U105 ( .A(\count[3] ), .B(n366), .C(\ScanReg[3] ), .D(n365), .Z(
        n393) );
    VMW_AO22 U80 ( .A(ScanOut[0]), .B(n363), .C(\count260[0] ), .D(n364), .Z(
        n411) );
    VMW_BUFIZ U122 ( .A(n381), .E(n377), .Z(\arr[25] ) );
    Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 sub_189 ( .A({
        \count[6] , \count[5] , \count[4] , \count[3] , \count[2] , \count[1] , 
        \count[0] }), .SUM({\count260[6] , \count260[5] , \count260[4] , 
        \count260[3] , \count260[2] , \count260[1] , \count260[0] }) );
    VMW_BUFIZ U139 ( .A(n398), .E(n377), .Z(\arr[26] ) );
    VMW_PULLDOWN U77 ( .Z(n404) );
    VMW_XOR2 U89 ( .A(Addr[0]), .B(Id), .Z(n365) );
    VMW_NOR2 U92 ( .A(n367), .B(n365), .Z(n363) );
    VMW_BUFIZ U145 ( .A(n404), .E(n377), .Z(\arr[8] ) );
    VMW_BUFIZ U117 ( .A(n375), .E(n377), .Z(\arr[10] ) );
    VMW_BUFIZ U130 ( .A(n389), .E(n377), .Z(\arr[13] ) );
    VMW_BUFIZ U138 ( .A(n397), .E(n377), .Z(\arr[5] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n406), .CP(Clk), .Q(\count[5] ) );
    VMW_PULLDOWN U64 ( .Z(n386) );
    VMW_AO22 U81 ( .A(ScanOut[1]), .B(n363), .C(\count260[1] ), .D(n364), .Z(
        n410) );
    VMW_AO22 U104 ( .A(\count[4] ), .B(n366), .C(\ScanReg[4] ), .D(n365), .Z(
        n378) );
    VMW_PULLDOWN U76 ( .Z(n402) );
    VMW_BUFIZ U116 ( .A(n374), .E(n377), .Z(\arr[23] ) );
    VMW_BUFIZ U123 ( .A(n382), .E(n377), .Z(\arr[16] ) );
    VMW_AO21 U88 ( .A(RD), .B(ScanEnable), .C(n366), .Z(n377) );
    VMW_AND2 U93 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_BUFIZ U131 ( .A(n390), .E(n377), .Z(\arr[30] ) );
    VMW_FD \count_reg[1]  ( .D(n410), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_BUFIZ U143 ( .A(n402), .E(n377), .Z(\arr[11] ) );
    VMW_BUFIZ U144 ( .A(n403), .E(n377), .Z(\arr[1] ) );
    VMW_FD \count_reg[3]  ( .D(n408), .CP(Clk), .Q(\count[3] ) );
    VMW_BUFIZ U136 ( .A(n395), .E(n377), .Z(\arr[17] ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_PULLDOWN U63 ( .Z(n385) );
    VMW_PULLDOWN U71 ( .Z(n395) );
    VMW_INV U111 ( .A(n365), .Z(n366) );
    VMW_BUFIZ U124 ( .A(n383), .E(n377), .Z(\arr[12] ) );
    VMW_OR4 U78 ( .A(\count[1] ), .B(\count[2] ), .C(\count[0] ), .D(n362), 
        .Z(Enable) );
    VMW_AO22 U86 ( .A(ScanOut[6]), .B(n363), .C(\count260[6] ), .D(n364), .Z(
        n405) );
    VMW_AO22 U103 ( .A(\count[5] ), .B(n366), .C(\ScanReg[5] ), .D(n365), .Z(
        n397) );
    VMW_BUFIZ U118 ( .A(n376), .E(n377), .Z(\arr[9] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \nOut1_20[5] , \nOut8_10[4] , \nOut9_31[2] , \nOut2_15[3] , 
        \nOut1_23[6] , \nOut8_13[7] , \nScanOut268[5] , \nOut10_29[0] , 
        \nOut15_15[7] , \nOut26_21[6] , \nOut30_19[1] , \nOut31_1[0] , 
        \nOut15_16[4] , \nOut19_19[1] , \nScanOut869[0] , \nOut26_22[5] , 
        \nScanOut1019[6] , \nScanOut108[0] , \nScanOut708[4] , 
        \nScanOut468[1] , \nOut31_2[3] , \nScanOut689[6] , \nOut0_1[1] , 
        \nOut0_2[2] , \nScanOut4[1] , \nScanOut7[2] , \nScanOut11[1] , 
        \nOut2_16[0] , \nOut7_29[4] , \nScanOut338[2] , \nOut16_20[1] , 
        \nOut25_14[0] , \nScanOut658[3] , \nOut16_23[2] , \nScanOut538[6] , 
        \nOut20_28[7] , \nOut25_17[3] , \nOut29_18[6] , \nScanOut939[7] , 
        \nScanOut396[2] , \nScanOut871[2] , \nOut31_23[6] , \nScanOut12[2] , 
        \nOut0_19[1] , \nScanOut110[2] , \nOut5_25[6] , \nScanOut270[7] , 
        \nOut11_10[4] , \nOut18_20[5] , \nOut22_24[5] , \nScanOut945[1] , 
        \nOut10_31[2] , \nScanOut596[6] , \nScanOut1001[4] , \nScanOut344[4] , 
        \nScanOut624[5] , \nScanOut710[6] , \nScanOut997[7] , \nScanOut470[3] , 
        \nScanOut544[0] , \nScanOut627[6] , \nScanOut113[1] , \nOut5_26[5] , 
        \nScanOut273[4] , \nScanOut713[5] , \nScanOut994[4] , \nOut9_29[0] , 
        \nScanOut347[7] , \nScanOut473[0] , \nScanOut547[3] , \nOut18_8[6] , 
        \nScanOut872[1] , \nScanOut946[2] , \nOut1_9[6] , \nOut12_9[3] , 
        \nOut31_20[5] , \nScanOut52[0] , \nScanOut75[5] , \nOut6_10[0] , 
        \nScanOut174[6] , \nOut7_9[2] , \nOut11_13[7] , \nScanOut395[1] , 
        \nOut27_18[2] , \nScanOut214[3] , \nOut14_9[7] , \nScanOut595[5] , 
        \nScanOut1002[7] , \nOut18_23[6] , \nScanOut640[1] , \nOut22_27[6] , 
        \nScanOut774[2] , \nScanOut320[0] , \nOut12_25[2] , \nScanOut414[7] , 
        \nScanOut520[4] , \nOut20_30[5] , \nOut21_11[3] , \nOut28_21[2] , 
        \nScanOut692[7] , \nScanOut815[6] , \nOut7_31[6] , \nScanOut921[5] , 
        \nScanOut76[6] , \nScanOut691[4] , \nScanOut816[5] , \nOut29_9[3] , 
        \nOut6_13[3] , \nScanOut177[5] , \nScanOut217[0] , \nOut23_8[6] , 
        \nScanOut922[6] , \nScanOut323[3] , \nScanOut643[2] , \nScanOut777[1] , 
        \nOut28_22[1] , \nScanOut181[5] , \nOut12_26[1] , \nScanOut417[4] , 
        \nScanOut523[7] , \nOut17_19[5] , \nOut21_12[0] , \nOut25_8[2] , 
        \nOut7_16[3] , \nScanOut832[3] , \nScanOut781[1] , \nScanOut906[0] , 
        \nOut2_29[7] , \nScanOut153[3] , \nOut13_23[1] , \nScanOut433[2] , 
        \nScanOut507[1] , \nOut20_17[0] , \nOut25_28[4] , \nOut29_27[1] , 
        \nScanOut80[6] , \nScanOut667[4] , \nScanOut753[7] , \nScanOut150[0] , 
        \nScanOut233[6] , \nScanOut307[5] , \nScanOut35[7] , \nScanOut36[4] , 
        \nScanOut51[3] , \nScanOut83[5] , \nScanOut230[5] , \nOut13_20[2] , 
        \nOut29_24[2] , \nScanOut430[1] , \nScanOut504[2] , \nOut20_14[3] , 
        \nScanOut304[6] , \nScanOut664[7] , \nScanOut750[4] , \nScanOut182[6] , 
        \nScanOut782[2] , \nScanOut831[0] , \nOut4_23[5] , \nScanOut137[7] , 
        \nOut7_15[0] , \nScanOut905[3] , \nScanOut257[2] , \nScanOut457[6] , 
        \nScanOut563[5] , \nOut30_9[7] , \nScanOut363[1] , \nScanOut285[4] , 
        \nOut10_16[7] , \nOut15_29[3] , \nScanOut603[0] , \nScanOut884[1] , 
        \nScanOut737[3] , \nOut19_26[6] , \nOut23_22[6] , \nScanOut485[0] , 
        \nScanOut856[7] , \nOut30_25[5] , \nOut10_15[4] , \nScanOut962[4] , 
        \nScanOut486[3] , \nOut19_25[5] , \nOut23_21[5] , \nScanOut855[4] , 
        \nScanOut961[7] , \nScanOut49[1] , \nOut3_6[3] , \nOut4_20[6] , 
        \nScanOut134[4] , \nScanOut286[7] , \nScanOut454[5] , \nScanOut560[6] , 
        \nOut30_26[6] , \nScanOut254[1] , \nScanOut600[3] , \nScanOut734[0] , 
        \nScanOut887[2] , \nScanOut360[2] , \nScanOut148[2] , \nOut12_19[6] , 
        \nOut24_12[3] , \nScanOut228[7] , \nOut9_7[6] , \nOut24_3[6] , 
        \nScanOut428[3] , \nOut17_26[2] , \nOut22_3[2] , \nScanOut748[6] , 
        \nOut3_13[0] , \nOut10_6[6] , \nOut5_6[7] , \nOut16_6[2] , 
        \nScanOut829[2] , \nOut3_5[0] , \nScanOut199[7] , \nOut10_5[5] , 
        \nOut28_2[7] , \nOut3_10[3] , \nOut2_31[5] , \nOut5_5[4] , 
        \nScanOut799[3] , \nOut28_1[4] , \nScanOut98[4] , \nOut9_4[5] , 
        \nOut16_5[1] , \nOut24_0[5] , \nOut17_25[1] , \nOut24_11[0] , 
        \nOut25_30[6] , \nOut6_2[6] , \nOut22_0[1] , \nOut27_27[5] , 
        \nOut13_2[7] , \nOut14_13[4] , \nOut22_18[1] , \nOut15_2[3] , 
        \nScanOut979[5] , \nOut0_25[5] , \nOut0_26[6] , \nScanOut578[4] , 
        \nOut21_7[3] , \nOut5_19[2] , \nOut9_16[7] , \nOut19_3[2] , 
        \nScanOut618[1] , \nOut27_7[7] , \nOut9_15[4] , \nScanOut378[0] , 
        \nOut19_0[1] , \nOut21_4[0] , \nOut27_4[4] , \nOut6_1[5] , 
        \nOut14_10[7] , \nOut15_1[0] , \nOut15_31[1] , \nOut27_24[6] , 
        \nScanOut9[4] , \nOut0_30[2] , \nScanOut38[2] , \nOut10_18[1] , 
        \nOut13_1[4] , \nOut15_27[5] , \nOut19_28[0] , \nOut26_13[4] , 
        \nScanOut858[1] , \nOut1_12[7] , \nScanOut139[1] , \nOut30_7[1] , 
        \nOut8_22[6] , \nScanOut259[4] , \nScanOut459[0] , \nScanOut739[5] , 
        \nOut30_4[2] , \nOut1_11[4] , \nScanOut889[4] , \nOut8_21[5] , 
        \nScanOut288[1] , \nOut15_24[6] , \nScanOut488[5] , \nOut26_10[7] , 
        \nOut27_31[1] , \nOut16_12[3] , \nScanOut509[7] , \nOut30_28[0] , 
        \nOut20_19[6] , \nOut29_29[7] , \nOut0_14[4] , \nScanOut20[0] , 
        \nScanOut23[3] , \nOut0_28[0] , \nOut2_24[2] , \nOut2_27[1] , 
        \nOut7_18[5] , \nScanOut309[3] , \nScanOut669[2] , \nOut25_26[2] , 
        \nScanOut908[6] , \nScanOut122[0] , \nScanOut442[1] , \nOut16_11[0] , 
        \nOut17_30[6] , \nOut25_25[1] , \nScanOut576[2] , \nScanOut616[7] , 
        \nOut21_9[5] , \nOut5_17[4] , \nScanOut242[5] , \nScanOut722[4] , 
        \nOut27_9[1] , \nScanOut891[6] , \nOut9_18[1] , \nScanOut376[6] , 
        \nOut11_22[6] , \nScanOut490[7] , \nOut27_29[3] , \nOut18_12[7] , 
        \nOut22_16[7] , \nScanOut843[0] , \nScanOut977[3] , \nScanOut290[3] , 
        \nScanOut293[0] , \nOut11_21[5] , \nOut18_11[4] , \nOut22_15[4] , 
        \nOut30_30[2] , \nOut31_11[4] , \nOut19_30[2] , \nScanOut493[4] , 
        \nScanOut840[3] , \nOut31_12[7] , \nOut2_3[1] , \nScanOut44[4] , 
        \nScanOut47[7] , \nOut3_8[5] , \nScanOut121[3] , \nScanOut974[0] , 
        \nOut5_14[7] , \nScanOut241[6] , \nScanOut441[2] , \nScanOut575[1] , 
        \nScanOut194[2] , \nScanOut375[5] , \nScanOut615[4] , \nScanOut892[5] , 
        \nScanOut721[7] , \nOut5_8[1] , \nOut10_8[0] , \nOut16_8[4] , 
        \nScanOut794[6] , \nScanOut827[4] , \nScanOut95[1] , \nScanOut146[4] , 
        \nOut6_22[2] , \nScanOut913[7] , \nScanOut226[1] , \nOut9_9[0] , 
        \nOut12_17[0] , \nOut28_13[0] , \nScanOut512[6] , \nScanOut426[5] , 
        \nOut17_28[4] , \nOut21_23[1] , \nScanOut312[2] , \nScanOut672[3] , 
        \nScanOut746[0] , \nScanOut96[2] , \nScanOut145[7] , \nOut12_14[3] , 
        \nScanOut425[6] , \nScanOut511[5] , \nOut21_20[2] , \nScanOut671[0] , 
        \nOut28_10[3] , \nOut29_31[5] , \nScanOut745[3] , \nOut6_21[1] , 
        \nScanOut197[1] , \nScanOut225[2] , \nScanOut311[1] , \nScanOut824[7] , 
        \nScanOut797[5] , \nScanOut910[4] , \nOut2_18[6] , \nScanOut60[2] , 
        \nScanOut161[1] , \nScanOut201[4] , \nScanOut335[7] , \nScanOut655[6] , 
        \nScanOut761[5] , \nOut12_30[5] , \nOut13_11[3] , \nOut29_15[3] , 
        \nScanOut401[0] , \nScanOut535[3] , \nOut20_25[2] , \nScanOut687[0] , 
        \nScanOut800[1] , \nScanOut63[1] , \nOut7_24[1] , \nScanOut934[2] , 
        \nOut7_27[2] , \nScanOut684[3] , \nScanOut803[2] , \nScanOut937[1] , 
        \nOut2_0[2] , \nOut3_21[2] , \nScanOut105[5] , \nOut4_11[7] , 
        \nScanOut162[2] , \nScanOut202[7] , \nScanOut656[5] , \nScanOut762[6] , 
        \nScanOut336[4] , \nOut13_12[0] , \nScanOut402[3] , \nScanOut536[0] , 
        \nOut20_26[1] , \nOut25_19[5] , \nScanOut265[0] , \nOut10_24[5] , 
        \nScanOut383[5] , \nScanOut864[5] , \nOut29_16[0] , \nOut30_17[7] , 
        \nScanOut950[6] , \nScanOut583[1] , \nOut19_14[4] , \nScanOut1014[3] , 
        \nScanOut631[2] , \nOut23_10[4] , \nOut22_31[2] , \nScanOut705[1] , 
        \nScanOut982[0] , \nOut5_30[1] , \nScanOut351[3] , \nScanOut465[4] , 
        \nScanOut551[7] , \nScanOut106[6] , \nOut4_12[4] , \nScanOut266[3] , 
        \nScanOut352[0] , \nScanOut632[1] , \nScanOut706[2] , \nScanOut981[3] , 
        \nOut4_0[6] , \nOut10_27[6] , \nScanOut380[6] , \nScanOut466[7] , 
        \nScanOut552[4] , \nOut15_18[2] , \nOut23_13[7] , \nScanOut867[6] , 
        \nOut30_14[4] , \nScanOut953[5] , \nOut19_17[7] , \nScanOut580[2] , 
        \nScanOut1017[0] , \nOut29_4[6] , \nOut11_0[7] , \nOut17_0[3] , 
        \nScanOut78[0] , \nOut3_22[1] , \nScanOut179[3] , \nScanOut219[6] , 
        \nOut8_1[7] , \nOut17_14[0] , \nOut23_5[3] , \nOut25_5[7] , 
        \nOut24_20[1] , \nOut12_28[7] , \nOut23_6[0] , \nOut24_23[2] , 
        \nScanOut779[7] , \nOut8_2[4] , \nOut25_6[4] , \nScanOut419[2] , 
        \nOut17_17[3] , \nOut17_3[0] , \nOut4_3[5] , \nScanOut818[3] , 
        \nOut29_7[5] , \nOut9_24[5] , \nOut11_3[4] , \nOut18_5[3] , 
        \nOut1_4[3] , \nOut20_1[2] , \nOut26_1[6] , \nScanOut999[1] , 
        \nScanOut398[4] , \nOut0_9[0] , \nOut0_17[7] , \nOut1_7[0] , 
        \nOut7_4[7] , \nOut12_4[6] , \nOut14_4[2] , \nOut14_21[6] , 
        \nOut12_7[5] , \nScanOut598[0] , \nOut27_15[7] , \nScanOut948[4] , 
        \nOut7_7[4] , \nOut27_16[4] , \nOut14_7[1] , \nOut14_22[5] , 
        \nOut22_29[0] , \nScanOut25[4] , \nScanOut41[0] , \nOut1_14[0] , 
        \nOut2_21[6] , \nScanOut88[7] , \nOut5_28[3] , \nOut9_27[6] , 
        \nScanOut629[0] , \nOut26_2[5] , \nOut18_6[0] , \nScanOut349[1] , 
        \nScanOut549[5] , \nOut20_2[1] , \nOut16_14[4] , \nOut25_20[5] , 
        \nOut2_22[5] , \nScanOut59[2] , \nScanOut189[4] , \nScanOut789[0] , 
        \nScanOut839[1] , \nScanOut158[1] , \nScanOut238[4] , \nScanOut758[5] , 
        \nOut13_28[3] , \nScanOut438[0] , \nOut16_17[7] , \nOut25_23[6] , 
        \nOut15_21[2] , \nOut26_15[3] , \nOut1_17[3] , \nOut4_28[7] , 
        \nOut8_24[1] , \nOut8_27[2] , \nOut30_1[6] , \nScanOut368[3] , 
        \nOut15_22[1] , \nScanOut568[7] , \nScanOut608[2] , \nOut30_2[5] , 
        \nOut23_29[4] , \nScanOut969[6] , \nScanOut792[1] , \nOut26_16[0] , 
        \nScanOut821[3] , \nScanOut42[3] , \nOut3_18[2] , \nScanOut90[5] , 
        \nScanOut93[6] , \nOut6_24[5] , \nScanOut192[5] , \nScanOut915[0] , 
        \nScanOut674[4] , \nScanOut740[7] , \nScanOut140[3] , \nScanOut220[6] , 
        \nScanOut314[5] , \nScanOut420[2] , \nScanOut514[1] , \nOut21_25[6] , 
        \nScanOut223[5] , \nOut12_11[7] , \nOut28_15[7] , \nOut13_30[1] , 
        \nScanOut317[6] , \nScanOut677[7] , \nOut22_8[0] , \nScanOut743[4] , 
        \nScanOut143[0] , \nOut12_12[4] , \nOut24_19[1] , \nScanOut423[1] , 
        \nScanOut517[2] , \nOut24_8[4] , \nOut28_16[4] , \nOut21_26[5] , 
        \nOut6_27[6] , \nScanOut822[0] , \nScanOut791[2] , \nScanOut916[3] , 
        \nOut28_9[5] , \nScanOut124[7] , \nOut4_30[5] , \nOut5_11[3] , 
        \nScanOut191[6] , \nScanOut244[2] , \nScanOut370[1] , \nScanOut610[0] , 
        \nScanOut724[3] , \nScanOut897[1] , \nScanOut296[4] , \nScanOut444[6] , 
        \nScanOut570[5] , \nScanOut845[7] , \nOut31_17[3] , \nScanOut971[4] , 
        \nScanOut26[7] , \nOut11_24[1] , \nOut18_14[0] , \nOut22_10[0] , 
        \nOut23_31[6] , \nOut13_9[5] , \nScanOut496[0] , \nScanOut846[4] , 
        \nScanOut972[7] , \nOut0_11[0] , \nOut0_12[3] , \nOut1_28[4] , 
        \nScanOut103[2] , \nScanOut127[4] , \nOut5_12[0] , \nOut6_9[4] , 
        \nScanOut295[7] , \nOut11_27[2] , \nOut31_14[0] , \nScanOut247[1] , 
        \nOut14_18[6] , \nScanOut495[3] , \nOut15_9[1] , \nOut18_17[3] , 
        \nOut22_13[3] , \nOut19_8[0] , \nScanOut613[3] , \nScanOut894[2] , 
        \nScanOut727[0] , \nScanOut373[2] , \nScanOut447[5] , \nScanOut573[6] , 
        \nOut10_22[2] , \nScanOut585[6] , \nOut19_12[3] , \nOut23_16[3] , 
        \nOut26_29[7] , \nScanOut385[2] , \nOut30_11[0] , \nScanOut1012[4] , 
        \nOut31_30[6] , \nScanOut862[2] , \nScanOut956[1] , \nOut4_17[0] , 
        \nScanOut263[7] , \nScanOut463[3] , \nScanOut557[0] , \nOut31_9[1] , 
        \nOut8_18[5] , \nScanOut357[4] , \nScanOut637[5] , \nScanOut65[6] , 
        \nScanOut66[5] , \nScanOut100[1] , \nScanOut460[0] , \nScanOut554[3] , 
        \nScanOut703[6] , \nScanOut984[7] , \nOut4_14[3] , \nScanOut260[4] , 
        \nScanOut634[6] , \nScanOut700[5] , \nScanOut987[4] , \nScanOut167[6] , 
        \nOut10_21[1] , \nScanOut354[7] , \nScanOut386[1] , \nOut18_30[6] , 
        \nScanOut586[5] , \nOut19_11[0] , \nOut23_15[0] , \nScanOut1011[7] , 
        \nScanOut861[1] , \nScanOut955[2] , \nScanOut407[7] , \nOut16_28[0] , 
        \nScanOut533[4] , \nOut30_12[3] , \nOut20_23[5] , \nScanOut207[3] , 
        \nOut13_17[4] , \nOut29_13[4] , \nScanOut653[1] , \nScanOut767[2] , 
        \nScanOut333[0] , \nScanOut681[7] , \nScanOut806[6] , \nOut7_21[5] , 
        \nOut7_22[6] , \nScanOut932[5] , \nScanOut682[4] , \nScanOut805[5] , 
        \nScanOut931[6] , \nScanOut118[3] , \nScanOut164[5] , \nOut13_14[7] , 
        \nOut28_31[1] , \nScanOut204[0] , \nScanOut404[4] , \nScanOut530[7] , 
        \nOut29_10[7] , \nOut20_20[6] , \nScanOut330[3] , \nScanOut478[2] , 
        \nScanOut650[2] , \nScanOut764[1] , \nOut20_7[5] , \nScanOut19[0] , 
        \nOut7_2[0] , \nScanOut278[6] , \nScanOut718[7] , \nOut26_7[1] , 
        \nOut9_22[2] , \nOut11_18[5] , \nOut18_3[4] , \nOut12_2[1] , 
        \nOut14_2[5] , \nOut27_13[0] , \nScanOut1009[5] , \nOut14_27[1] , 
        \nOut18_28[4] , \nScanOut879[3] , \nOut1_1[7] , \nOut1_2[4] , 
        \nOut7_1[3] , \nOut14_1[6] , \nOut14_24[2] , \nOut27_10[3] , 
        \nOut26_31[5] , \nOut1_30[6] , \nOut9_21[1] , \nOut12_1[2] , 
        \nOut31_28[4] , \nOut20_4[6] , \nOut18_0[7] , \nScanOut14[5] , 
        \nScanOut17[6] , \nOut2_5[6] , \nOut2_6[5] , \nOut26_4[2] , 
        \nOut3_27[5] , \nOut11_6[0] , \nOut4_6[1] , \nOut17_6[4] , 
        \nOut6_18[1] , \nOut29_2[1] , \nOut8_4[3] , \nOut8_7[0] , 
        \nOut17_12[7] , \nScanOut528[5] , \nOut24_26[6] , \nOut28_29[3] , 
        \nScanOut929[4] , \nOut21_19[2] , \nOut25_3[0] , \nScanOut328[1] , 
        \nOut23_3[4] , \nScanOut648[0] , \nOut25_0[3] , \nOut11_5[3] , 
        \nOut16_30[2] , \nOut17_11[4] , \nOut23_0[7] , \nOut24_25[5] , 
        \nOut2_8[3] , \nOut2_10[7] , \nOut2_13[4] , \nScanOut68[3] , 
        \nOut3_24[6] , \nOut4_5[2] , \nScanOut699[5] , \nOut17_5[7] , 
        \nOut29_1[2] , \nScanOut808[0] , \nOut3_31[1] , \nScanOut169[0] , 
        \nOut13_19[2] , \nScanOut409[1] , \nOut16_26[6] , \nOut25_12[7] , 
        \nScanOut209[5] , \nScanOut769[4] , \nOut16_25[5] , \nOut24_30[2] , 
        \nOut25_11[4] , \nOut1_25[1] , \nOut1_26[2] , \nOut4_19[6] , 
        \nOut8_16[3] , \nScanOut559[6] , \nOut31_7[7] , \nScanOut359[2] , 
        \nScanOut388[7] , \nOut15_10[3] , \nOut15_13[0] , \nScanOut639[3] , 
        \nOut14_31[5] , \nScanOut588[3] , \nOut23_18[5] , \nOut26_24[2] , 
        \nOut26_27[1] , \nScanOut958[7] , \nOut31_4[4] , \nScanOut172[1] , 
        \nOut8_15[0] , \nScanOut989[2] , \nOut12_23[5] , \nOut24_28[0] , 
        \nOut28_27[5] , \nScanOut212[4] , \nOut8_9[6] , \nScanOut526[3] , 
        \nScanOut412[0] , \nOut21_17[4] , \nScanOut326[7] , \nScanOut646[6] , 
        \nScanOut772[5] , \nScanOut70[1] , \nScanOut73[2] , \nOut3_29[3] , 
        \nOut11_8[6] , \nOut4_8[7] , \nOut17_8[2] , \nScanOut694[0] , 
        \nScanOut813[1] , \nOut6_16[7] , \nScanOut927[2] , \nScanOut697[3] , 
        \nScanOut810[2] , \nScanOut171[2] , \nOut6_15[4] , \nScanOut411[3] , 
        \nScanOut525[0] , \nScanOut924[1] , \nOut21_14[7] , \nOut28_24[6] , 
        \nScanOut211[7] , \nOut12_20[6] , \nScanOut645[5] , \nScanOut771[6] , 
        \nScanOut325[4] , \nOut11_16[3] , \nOut14_29[7] , \nScanOut590[1] , 
        \nOut22_22[2] , \nScanOut1007[3] , \nOut18_26[2] , \nScanOut877[5] , 
        \nScanOut115[6] , \nScanOut116[5] , \nScanOut390[5] , \nScanOut943[6] , 
        \nScanOut476[4] , \nScanOut542[7] , \nOut31_25[1] , \nOut5_23[1] , 
        \nScanOut276[0] , \nOut20_9[3] , \nScanOut622[2] , \nScanOut716[1] , 
        \nOut26_9[7] , \nScanOut991[0] , \nScanOut342[3] , \nOut5_20[2] , 
        \nScanOut275[3] , \nScanOut475[7] , \nScanOut541[4] , \nOut11_15[0] , 
        \nScanOut341[0] , \nOut18_25[1] , \nScanOut621[1] , \nScanOut715[2] , 
        \nScanOut992[3] , \nOut22_21[1] , \nScanOut393[6] , \nScanOut593[2] , 
        \nOut31_26[2] , \nScanOut1004[0] , \nScanOut874[6] , \nScanOut940[5] , 
        \nScanOut30[3] , \nOut4_25[2] , \nScanOut251[5] , \nScanOut605[7] , 
        \nScanOut882[6] , \nScanOut731[4] , \nScanOut365[6] , \nScanOut131[0] , 
        \nScanOut451[1] , \nScanOut565[2] , \nScanOut850[0] , \nScanOut33[0] , 
        \nScanOut280[0] , \nScanOut283[3] , \nScanOut964[3] , \nOut10_10[0] , 
        \nOut30_23[2] , \nOut11_31[6] , \nScanOut483[7] , \nScanOut1020[6] , 
        \nOut19_20[1] , \nOut23_24[1] , \nScanOut853[3] , \nOut30_20[1] , 
        \nScanOut967[0] , \nOut1_19[5] , \nOut4_26[1] , \nScanOut252[6] , 
        \nOut10_13[3] , \nOut19_23[2] , \nOut23_27[2] , \nScanOut480[4] , 
        \nOut26_18[6] , \nScanOut1023[5] , \nScanOut366[5] , \nOut8_29[4] , 
        \nScanOut606[4] , \nScanOut881[5] , \nScanOut54[7] , \nScanOut132[3] , 
        \nScanOut732[7] , \nOut7_10[4] , \nScanOut452[2] , \nScanOut566[1] , 
        \nScanOut834[4] , \nOut6_31[2] , \nScanOut787[6] , \nScanOut900[7] , 
        \nScanOut187[2] , \nScanOut235[1] , \nScanOut301[2] , \nScanOut1[5] , 
        \nScanOut86[1] , \nScanOut661[3] , \nScanOut755[0] , \nScanOut155[4] , 
        \nOut13_25[6] , \nOut29_21[6] , \nScanOut2[6] , \nScanOut85[2] , 
        \nScanOut435[5] , \nScanOut501[6] , \nOut20_11[7] , \nOut21_30[1] , 
        \nScanOut662[0] , \nScanOut756[3] , \nScanOut156[7] , \nScanOut236[2] , 
        \nScanOut302[1] , \nScanOut436[6] , \nScanOut502[5] , \nOut16_19[1] , 
        \nOut20_12[4] , \nOut0_4[5] , \nScanOut57[4] , \nOut13_26[5] , 
        \nOut29_22[5] , \nScanOut784[5] , \nScanOut837[7] , \nScanOut184[1] , 
        \nOut7_13[7] , \nScanOut903[4] , \nOut0_7[6] , \nOut0_20[1] , 
        \nOut6_4[1] , \nScanOut298[2] , \nOut13_4[0] , \nOut31_19[5] , 
        \nOut14_15[3] , \nOut15_4[4] , \nOut27_21[2] , \nOut9_10[0] , 
        \nOut8_31[6] , \nScanOut498[6] , \nOut19_5[5] , \nOut0_23[2] , 
        \nOut21_1[4] , \nOut27_1[0] , \nScanOut899[7] , \nOut27_2[3] , 
        \nScanOut28[1] , \nScanOut129[2] , \nScanOut249[7] , \nScanOut729[6] , 
        \nOut9_13[3] , \nOut19_6[6] , \nScanOut449[3] , \nOut13_7[3] , 
        \nOut21_2[7] , \nScanOut848[2] , \nOut0_17[3] , \nOut2_3[5] , 
        \nOut3_3[7] , \nOut3_15[7] , \nOut5_0[0] , \nOut6_7[2] , 
        \nOut11_29[4] , \nOut27_22[1] , \nOut9_1[1] , \nOut14_16[0] , 
        \nOut15_7[7] , \nOut18_19[5] , \nOut22_5[5] , \nOut24_5[1] , 
        \nOut17_20[5] , \nOut24_14[4] , \nOut28_4[0] , \nOut3_16[4] , 
        \nOut3_0[4] , \nOut10_0[1] , \nOut16_0[5] , \nOut5_3[3] , 
        \nOut16_3[6] , \nOut6_29[0] , \nOut28_7[3] , \nScanOut918[5] , 
        \nOut9_2[2] , \nOut10_3[2] , \nScanOut319[0] , \nOut22_6[6] , 
        \nScanOut519[4] , \nScanOut679[1] , \nOut24_17[7] , \nOut28_18[2] , 
        \nOut24_6[2] , \nOut11_3[0] , \nOut17_23[6] , \nOut21_28[3] , 
        \nOut2_0[6] , \nScanOut78[4] , \nOut4_3[1] , \nScanOut818[7] , 
        \nOut29_7[1] , \nOut3_22[5] , \nScanOut179[7] , \nOut8_2[0] , 
        \nOut17_3[4] , \nOut25_6[0] , \nOut12_28[3] , \nScanOut419[6] , 
        \nOut17_17[7] , \nOut24_23[6] , \nScanOut219[2] , \nScanOut779[3] , 
        \nOut8_1[3] , \nOut17_14[4] , \nOut23_6[4] , \nOut24_20[5] , 
        \nOut25_5[3] , \nOut23_5[7] , \nOut3_21[6] , \nOut11_0[3] , 
        \nOut17_0[7] , \nOut4_0[2] , \nOut5_28[7] , \nOut9_27[2] , 
        \nScanOut549[1] , \nOut20_2[5] , \nOut29_4[2] , \nOut18_6[4] , 
        \nScanOut349[5] , \nOut1_7[4] , \nOut7_7[0] , \nOut14_7[5] , 
        \nScanOut629[4] , \nOut26_2[1] , \nOut14_22[1] , \nOut22_29[4] , 
        \nOut27_16[0] , \nOut7_4[3] , \nOut12_7[1] , \nOut27_15[3] , 
        \nScanOut948[0] , \nOut14_4[6] , \nScanOut598[4] , \nOut14_21[2] , 
        \nOut0_14[0] , \nOut1_4[7] , \nOut12_4[2] , \nScanOut398[0] , 
        \nOut20_1[6] , \nOut9_24[1] , \nOut26_1[2] , \nScanOut999[5] , 
        \nOut13_12[4] , \nOut18_5[7] , \nOut25_19[1] , \nOut0_1[5] , 
        \nScanOut9[0] , \nScanOut20[4] , \nOut2_18[2] , \nScanOut162[6] , 
        \nScanOut202[3] , \nScanOut402[7] , \nScanOut536[4] , \nOut29_16[4] , 
        \nOut20_26[5] , \nScanOut336[0] , \nScanOut656[1] , \nScanOut762[2] , 
        \nScanOut60[6] , \nScanOut63[5] , \nOut7_27[6] , \nScanOut684[7] , 
        \nScanOut803[6] , \nScanOut937[5] , \nScanOut687[4] , \nScanOut800[5] , 
        \nScanOut105[1] , \nScanOut106[2] , \nScanOut161[5] , \nOut7_24[5] , 
        \nScanOut934[6] , \nScanOut401[4] , \nScanOut535[7] , \nOut20_25[6] , 
        \nScanOut201[0] , \nOut12_30[1] , \nOut13_11[7] , \nOut29_15[7] , 
        \nScanOut655[2] , \nScanOut761[1] , \nOut10_27[2] , \nScanOut335[3] , 
        \nScanOut580[6] , \nScanOut380[2] , \nOut15_18[6] , \nScanOut1017[4] , 
        \nOut19_17[3] , \nOut23_13[3] , \nScanOut867[2] , \nScanOut953[1] , 
        \nScanOut466[3] , \nScanOut552[0] , \nOut30_14[0] , \nOut4_12[0] , 
        \nScanOut266[7] , \nScanOut632[5] , \nScanOut706[6] , \nScanOut981[7] , 
        \nScanOut352[4] , \nOut4_11[3] , \nScanOut265[4] , \nScanOut465[0] , 
        \nScanOut551[3] , \nScanOut121[7] , \nOut5_14[3] , \nOut5_30[5] , 
        \nScanOut241[2] , \nOut10_24[1] , \nScanOut351[7] , \nOut19_14[0] , 
        \nScanOut631[6] , \nScanOut705[5] , \nScanOut982[4] , \nOut23_10[0] , 
        \nOut22_31[6] , \nScanOut383[1] , \nScanOut583[5] , \nOut30_17[3] , 
        \nScanOut1014[7] , \nScanOut615[0] , \nScanOut864[1] , 
        \nScanOut892[1] , \nScanOut950[2] , \nScanOut721[3] , \nScanOut375[1] , 
        \nScanOut441[6] , \nScanOut575[5] , \nScanOut840[7] , \nScanOut23[7] , 
        \nScanOut290[7] , \nScanOut293[4] , \nScanOut974[4] , \nOut11_21[1] , 
        \nOut31_12[3] , \nScanOut493[0] , \nOut18_11[0] , \nOut22_15[0] , 
        \nOut19_30[6] , \nScanOut843[4] , \nOut30_30[6] , \nOut31_11[0] , 
        \nScanOut977[7] , \nOut0_28[4] , \nOut5_17[0] , \nScanOut242[1] , 
        \nOut11_22[2] , \nOut18_12[3] , \nOut22_16[3] , \nOut27_29[7] , 
        \nScanOut490[3] , \nOut9_18[5] , \nScanOut376[2] , \nScanOut616[3] , 
        \nOut27_9[5] , \nOut0_30[6] , \nScanOut44[0] , \nScanOut122[4] , 
        \nScanOut722[0] , \nScanOut891[2] , \nOut6_21[5] , \nScanOut442[5] , 
        \nScanOut576[6] , \nOut21_9[1] , \nScanOut824[3] , \nScanOut797[1] , 
        \nScanOut910[0] , \nScanOut47[3] , \nScanOut95[5] , \nScanOut96[6] , 
        \nScanOut197[5] , \nScanOut225[6] , \nScanOut311[5] , \nScanOut671[4] , 
        \nScanOut745[7] , \nScanOut145[3] , \nOut12_14[7] , \nScanOut425[2] , 
        \nScanOut511[1] , \nOut28_10[7] , \nOut29_31[1] , \nOut21_20[6] , 
        \nScanOut672[7] , \nScanOut746[4] , \nOut5_8[5] , \nScanOut146[0] , 
        \nScanOut226[5] , \nOut9_9[4] , \nScanOut312[6] , \nScanOut512[2] , 
        \nScanOut426[1] , \nOut17_28[0] , \nOut21_23[5] , \nOut12_17[4] , 
        \nOut28_13[4] , \nScanOut794[2] , \nScanOut827[0] , \nOut3_8[1] , 
        \nOut6_22[6] , \nScanOut194[6] , \nOut10_8[4] , \nOut16_8[0] , 
        \nScanOut913[3] , \nOut8_21[1] , \nScanOut288[5] , \nOut15_24[2] , 
        \nOut30_28[4] , \nScanOut488[1] , \nOut26_10[3] , \nOut27_31[5] , 
        \nScanOut38[6] , \nOut1_11[0] , \nScanOut889[0] , \nOut1_12[3] , 
        \nOut30_4[6] , \nScanOut139[5] , \nOut8_22[2] , \nScanOut259[0] , 
        \nScanOut739[1] , \nScanOut459[4] , \nOut30_7[5] , \nScanOut858[5] , 
        \nOut2_24[6] , \nOut10_18[5] , \nOut15_27[1] , \nOut19_28[4] , 
        \nOut26_13[0] , \nOut16_11[4] , \nOut17_30[2] , \nOut25_25[5] , 
        \nOut2_27[5] , \nOut7_18[1] , \nScanOut309[7] , \nScanOut908[2] , 
        \nScanOut669[6] , \nScanOut49[5] , \nOut3_5[4] , \nOut3_10[7] , 
        \nOut2_31[1] , \nScanOut98[0] , \nOut16_12[7] , \nScanOut509[3] , 
        \nOut25_26[6] , \nOut29_29[3] , \nOut20_19[2] , \nOut22_0[5] , 
        \nOut9_4[1] , \nOut24_11[4] , \nOut24_0[1] , \nOut25_30[2] , 
        \nOut17_25[5] , \nOut5_5[0] , \nOut16_5[5] , \nScanOut799[7] , 
        \nScanOut199[3] , \nOut28_1[0] , \nOut5_6[3] , \nOut10_5[1] , 
        \nScanOut829[6] , \nOut28_2[3] , \nOut3_6[7] , \nOut3_13[4] , 
        \nOut10_6[2] , \nOut16_6[6] , \nScanOut148[6] , \nScanOut228[3] , 
        \nScanOut748[2] , \nOut9_7[2] , \nOut22_3[6] , \nOut24_3[2] , 
        \nOut12_19[2] , \nScanOut428[7] , \nOut17_26[6] , \nOut24_12[7] , 
        \nOut13_1[0] , \nOut0_2[6] , \nOut0_25[1] , \nOut6_1[1] , 
        \nOut27_24[2] , \nOut14_10[3] , \nOut15_1[4] , \nOut15_31[5] , 
        \nOut0_26[2] , \nOut5_19[6] , \nOut9_15[0] , \nOut19_0[5] , 
        \nOut27_4[0] , \nOut9_16[3] , \nOut19_3[6] , \nOut21_4[4] , 
        \nScanOut378[4] , \nOut27_7[3] , \nScanOut578[0] , \nScanOut618[5] , 
        \nOut21_7[7] , \nScanOut4[5] , \nScanOut51[7] , \nOut6_2[2] , 
        \nOut13_2[3] , \nOut14_13[0] , \nScanOut979[1] , \nOut15_2[7] , 
        \nOut22_18[5] , \nOut27_27[1] , \nScanOut782[6] , \nScanOut831[4] , 
        \nScanOut83[1] , \nScanOut182[2] , \nOut7_15[4] , \nScanOut905[7] , 
        \nScanOut664[3] , \nScanOut750[0] , \nScanOut150[4] , \nScanOut230[1] , 
        \nScanOut304[2] , \nScanOut430[5] , \nScanOut504[6] , \nOut20_14[7] , 
        \nOut29_24[6] , \nScanOut7[6] , \nScanOut80[2] , \nScanOut233[2] , 
        \nOut13_20[6] , \nScanOut307[1] , \nScanOut667[0] , \nScanOut753[3] , 
        \nScanOut153[7] , \nOut13_23[5] , \nOut25_28[0] , \nScanOut11[5] , 
        \nScanOut12[6] , \nScanOut35[3] , \nScanOut52[4] , \nOut2_29[3] , 
        \nScanOut433[6] , \nScanOut507[5] , \nOut29_27[5] , \nOut20_17[4] , 
        \nOut7_16[7] , \nScanOut832[7] , \nScanOut781[5] , \nScanOut906[4] , 
        \nOut4_20[2] , \nScanOut181[1] , \nScanOut254[5] , \nScanOut360[6] , 
        \nScanOut134[0] , \nScanOut600[7] , \nScanOut734[4] , \nScanOut887[6] , 
        \nScanOut286[3] , \nScanOut454[1] , \nScanOut560[2] , \nScanOut855[0] , 
        \nOut30_26[2] , \nScanOut961[3] , \nScanOut36[0] , \nOut10_15[0] , 
        \nOut19_25[1] , \nOut23_21[1] , \nScanOut486[7] , \nScanOut856[3] , 
        \nOut1_9[2] , \nOut4_23[1] , \nScanOut257[6] , \nScanOut285[0] , 
        \nScanOut962[0] , \nOut10_16[3] , \nOut30_25[1] , \nOut15_29[7] , 
        \nScanOut485[4] , \nOut23_22[2] , \nOut19_26[2] , \nScanOut603[4] , 
        \nScanOut884[5] , \nScanOut737[7] , \nScanOut363[5] , \nScanOut137[3] , 
        \nScanOut457[2] , \nScanOut563[1] , \nOut7_9[6] , \nOut11_13[3] , 
        \nOut14_9[3] , \nOut30_9[3] , \nOut18_23[2] , \nOut22_27[2] , 
        \nScanOut595[1] , \nOut27_18[6] , \nOut31_20[1] , \nScanOut1002[3] , 
        \nOut12_9[7] , \nScanOut395[5] , \nScanOut872[5] , \nScanOut946[6] , 
        \nOut0_19[5] , \nScanOut113[5] , \nOut5_26[1] , \nScanOut273[0] , 
        \nScanOut473[4] , \nScanOut547[7] , \nOut9_29[4] , \nScanOut347[3] , 
        \nOut18_8[2] , \nScanOut627[2] , \nScanOut110[6] , \nScanOut470[7] , 
        \nScanOut544[4] , \nScanOut713[1] , \nScanOut994[0] , \nOut5_25[2] , 
        \nScanOut270[3] , \nScanOut624[1] , \nScanOut710[2] , \nScanOut997[3] , 
        \nOut11_10[0] , \nScanOut344[0] , \nOut10_31[6] , \nScanOut596[2] , 
        \nOut18_20[1] , \nOut22_24[1] , \nScanOut1001[0] , \nScanOut871[6] , 
        \nOut1_23[2] , \nScanOut75[1] , \nScanOut76[2] , \nScanOut177[1] , 
        \nScanOut396[6] , \nScanOut945[5] , \nScanOut417[0] , \nScanOut523[3] , 
        \nOut31_23[2] , \nOut17_19[1] , \nOut21_12[4] , \nOut25_8[6] , 
        \nOut28_22[5] , \nScanOut217[4] , \nOut12_26[5] , \nScanOut643[6] , 
        \nOut23_8[2] , \nScanOut777[5] , \nScanOut323[7] , \nScanOut691[0] , 
        \nScanOut816[1] , \nOut29_9[7] , \nOut6_10[4] , \nOut6_13[7] , 
        \nScanOut692[3] , \nScanOut815[2] , \nScanOut922[2] , \nOut7_31[2] , 
        \nScanOut921[1] , \nScanOut108[4] , \nScanOut174[2] , \nOut12_25[6] , 
        \nOut28_21[6] , \nScanOut214[7] , \nScanOut414[3] , \nScanOut520[0] , 
        \nOut20_30[1] , \nOut21_11[7] , \nScanOut320[4] , \nScanOut468[5] , 
        \nScanOut640[5] , \nScanOut774[6] , \nOut31_2[7] , \nOut8_13[3] , 
        \nScanOut268[1] , \nScanOut708[0] , \nOut10_29[4] , \nOut26_22[1] , 
        \nOut15_15[3] , \nOut15_16[0] , \nOut19_19[5] , \nScanOut1019[2] , 
        \nScanOut869[4] , \nOut26_21[2] , \nOut30_19[5] , \nOut2_16[4] , 
        \nOut1_20[1] , \nOut8_10[0] , \nOut9_31[6] , \nOut31_1[4] , 
        \nOut7_29[0] , \nScanOut939[3] , \nScanOut338[6] , \nOut16_23[6] , 
        \nScanOut538[2] , \nOut25_17[7] , \nOut29_18[2] , \nOut20_28[3] , 
        \nOut16_20[5] , \nScanOut658[7] , \nOut25_14[4] , \nScanOut1[1] , 
        \nScanOut2[2] , \nOut0_4[1] , \nOut0_7[2] , \nOut2_15[7] , 
        \nScanOut689[2] , \nOut6_7[6] , \nOut11_29[0] , \nOut14_16[4] , 
        \nOut15_7[3] , \nOut18_19[1] , \nOut27_22[5] , \nOut0_20[5] , 
        \nOut0_23[6] , \nScanOut28[5] , \nOut13_7[7] , \nScanOut848[6] , 
        \nScanOut129[6] , \nScanOut249[3] , \nScanOut449[7] , \nOut21_2[3] , 
        \nOut9_13[7] , \nOut19_6[2] , \nOut21_1[0] , \nScanOut729[2] , 
        \nOut27_2[7] , \nOut27_1[4] , \nOut6_4[5] , \nOut9_10[4] , 
        \nOut8_31[2] , \nOut19_5[1] , \nScanOut899[3] , \nOut27_21[6] , 
        \nOut13_4[4] , \nOut14_15[7] , \nScanOut498[2] , \nOut15_4[0] , 
        \nScanOut30[7] , \nScanOut33[4] , \nOut1_19[1] , \nOut3_3[3] , 
        \nOut9_2[6] , \nScanOut298[6] , \nScanOut519[0] , \nOut31_19[1] , 
        \nOut24_6[6] , \nOut10_3[6] , \nScanOut319[4] , \nOut17_23[2] , 
        \nOut21_28[7] , \nOut22_6[2] , \nScanOut679[5] , \nOut24_17[3] , 
        \nOut28_18[6] , \nOut3_15[3] , \nOut3_16[0] , \nOut5_3[7] , 
        \nOut6_29[4] , \nOut28_7[7] , \nScanOut918[1] , \nOut3_0[0] , 
        \nOut16_3[2] , \nOut10_0[5] , \nScanOut132[7] , \nOut5_0[4] , 
        \nOut16_0[1] , \nOut9_1[5] , \nOut24_5[5] , \nOut24_14[0] , 
        \nOut28_4[4] , \nScanOut452[6] , \nOut17_20[1] , \nScanOut566[5] , 
        \nOut22_5[1] , \nScanOut606[0] , \nScanOut881[1] , \nOut4_26[5] , 
        \nScanOut252[2] , \nScanOut732[3] , \nScanOut366[1] , \nOut8_29[0] , 
        \nOut10_13[7] , \nOut26_18[2] , \nScanOut480[0] , \nOut19_23[6] , 
        \nScanOut1023[1] , \nOut23_27[6] , \nScanOut853[7] , \nScanOut967[4] , 
        \nScanOut280[4] , \nScanOut283[7] , \nOut10_10[4] , \nOut19_20[5] , 
        \nOut23_24[5] , \nOut30_20[5] , \nOut11_31[2] , \nScanOut483[3] , 
        \nScanOut1020[2] , \nScanOut850[4] , \nOut30_23[6] , \nScanOut57[0] , 
        \nOut4_25[6] , \nScanOut131[4] , \nScanOut964[7] , \nScanOut251[1] , 
        \nScanOut451[5] , \nScanOut565[6] , \nScanOut365[2] , \nScanOut184[5] , 
        \nScanOut605[3] , \nScanOut882[2] , \nScanOut731[0] , \nScanOut784[1] , 
        \nScanOut837[3] , \nScanOut156[3] , \nOut7_13[3] , \nScanOut903[0] , 
        \nOut29_22[1] , \nScanOut85[6] , \nScanOut236[6] , \nOut13_26[1] , 
        \nScanOut436[2] , \nScanOut502[1] , \nOut16_19[5] , \nOut20_12[0] , 
        \nScanOut302[5] , \nScanOut662[4] , \nScanOut756[7] , \nScanOut155[0] , 
        \nOut13_25[2] , \nScanOut435[1] , \nScanOut501[2] , \nOut20_11[3] , 
        \nOut21_30[5] , \nScanOut54[3] , \nScanOut86[5] , \nScanOut661[7] , 
        \nOut29_21[2] , \nScanOut755[4] , \nScanOut187[6] , \nScanOut235[5] , 
        \nScanOut301[6] , \nOut7_10[0] , \nScanOut834[0] , \nOut6_31[6] , 
        \nScanOut787[2] , \nScanOut900[3] , \nScanOut70[5] , \nScanOut171[6] , 
        \nScanOut211[3] , \nScanOut325[0] , \nScanOut645[1] , \nScanOut771[2] , 
        \nOut28_24[2] , \nOut12_20[2] , \nScanOut411[7] , \nScanOut525[4] , 
        \nOut21_14[3] , \nScanOut697[7] , \nScanOut810[6] , \nScanOut73[6] , 
        \nOut4_8[3] , \nOut6_15[0] , \nScanOut694[4] , \nScanOut813[5] , 
        \nScanOut924[5] , \nOut6_16[3] , \nScanOut927[6] , \nOut0_11[4] , 
        \nScanOut14[1] , \nOut2_8[7] , \nOut3_29[7] , \nOut17_8[6] , 
        \nOut11_8[2] , \nScanOut172[5] , \nScanOut212[0] , \nScanOut646[2] , 
        \nScanOut772[1] , \nOut8_9[2] , \nScanOut326[3] , \nScanOut526[7] , 
        \nOut12_23[1] , \nScanOut412[4] , \nOut21_17[0] , \nOut24_28[4] , 
        \nOut28_27[1] , \nScanOut874[2] , \nScanOut940[1] , \nScanOut17[2] , 
        \nScanOut115[2] , \nOut5_20[6] , \nScanOut275[7] , \nOut11_15[4] , 
        \nScanOut393[2] , \nOut31_26[6] , \nOut18_25[5] , \nScanOut593[6] , 
        \nScanOut1004[4] , \nScanOut621[5] , \nOut22_21[5] , \nScanOut715[6] , 
        \nScanOut992[7] , \nScanOut341[4] , \nScanOut475[3] , \nScanOut541[0] , 
        \nScanOut116[1] , \nOut5_23[5] , \nScanOut276[4] , \nScanOut342[7] , 
        \nScanOut622[6] , \nScanOut716[5] , \nOut26_9[3] , \nScanOut991[4] , 
        \nScanOut390[1] , \nScanOut476[0] , \nScanOut542[3] , \nOut20_9[7] , 
        \nScanOut877[1] , \nOut31_25[5] , \nOut2_10[3] , \nOut3_31[5] , 
        \nOut11_16[7] , \nOut14_29[3] , \nScanOut943[2] , \nOut18_26[6] , 
        \nOut22_22[6] , \nScanOut590[5] , \nScanOut1007[7] , \nOut2_13[0] , 
        \nScanOut169[4] , \nScanOut209[1] , \nOut16_25[1] , \nOut24_30[6] , 
        \nOut25_11[0] , \nOut13_19[6] , \nScanOut769[0] , \nOut25_12[3] , 
        \nScanOut409[5] , \nOut16_26[2] , \nOut1_25[5] , \nScanOut68[7] , 
        \nScanOut808[4] , \nOut8_15[4] , \nOut1_26[6] , \nScanOut388[3] , 
        \nOut31_4[0] , \nScanOut989[6] , \nOut15_10[7] , \nOut14_31[1] , 
        \nOut15_13[4] , \nScanOut588[7] , \nOut26_24[6] , \nOut23_18[1] , 
        \nOut26_27[5] , \nScanOut958[3] , \nOut1_30[2] , \nOut4_19[2] , 
        \nOut8_16[7] , \nScanOut639[7] , \nScanOut359[6] , \nScanOut559[2] , 
        \nOut31_7[3] , \nOut0_12[7] , \nScanOut19[4] , \nOut1_1[3] , 
        \nOut9_21[5] , \nOut26_4[6] , \nOut12_1[6] , \nOut18_0[3] , 
        \nOut20_4[2] , \nOut1_2[0] , \nOut7_1[7] , \nOut31_28[0] , 
        \nOut14_1[2] , \nOut27_10[7] , \nOut26_31[1] , \nOut14_24[6] , 
        \nScanOut879[7] , \nOut7_2[4] , \nOut11_18[1] , \nOut12_2[5] , 
        \nOut14_2[1] , \nOut14_27[5] , \nOut18_28[0] , \nOut27_13[4] , 
        \nScanOut278[2] , \nScanOut1009[1] , \nOut9_22[6] , \nOut18_3[0] , 
        \nOut2_5[2] , \nOut3_24[2] , \nScanOut118[7] , \nOut20_7[1] , 
        \nScanOut718[3] , \nOut26_7[5] , \nScanOut478[6] , \nOut4_5[6] , 
        \nOut17_5[3] , \nScanOut699[1] , \nOut29_1[6] , \nOut2_6[1] , 
        \nOut3_27[1] , \nOut4_6[5] , \nOut8_4[7] , \nOut11_5[7] , 
        \nOut23_0[3] , \nOut24_25[1] , \nOut25_0[7] , \nOut8_7[4] , 
        \nScanOut328[5] , \nOut16_30[6] , \nOut17_11[0] , \nScanOut648[4] , 
        \nOut23_3[0] , \nOut17_12[3] , \nScanOut528[1] , \nOut21_19[6] , 
        \nOut25_3[4] , \nOut24_26[2] , \nOut28_29[7] , \nOut6_18[5] , 
        \nOut29_2[5] , \nOut17_6[0] , \nScanOut929[0] , \nOut11_6[4] , 
        \nScanOut100[5] , \nOut4_14[7] , \nScanOut260[0] , \nOut10_21[5] , 
        \nScanOut386[5] , \nOut18_30[2] , \nOut19_11[4] , \nOut23_15[4] , 
        \nScanOut861[5] , \nOut30_12[7] , \nScanOut955[6] , \nScanOut586[1] , 
        \nScanOut1011[3] , \nScanOut354[3] , \nScanOut634[2] , 
        \nScanOut700[1] , \nScanOut987[0] , \nScanOut460[4] , \nScanOut554[7] , 
        \nScanOut1[3] , \nOut0_4[3] , \nOut0_9[6] , \nOut0_9[4] , 
        \nScanOut41[4] , \nScanOut42[7] , \nOut1_28[0] , \nScanOut637[1] , 
        \nScanOut65[2] , \nScanOut103[6] , \nOut4_17[4] , \nScanOut263[3] , 
        \nScanOut703[2] , \nScanOut984[3] , \nOut8_18[1] , \nScanOut357[0] , 
        \nScanOut463[7] , \nScanOut557[4] , \nScanOut164[1] , \nScanOut204[4] , 
        \nOut10_22[6] , \nScanOut385[6] , \nScanOut862[6] , \nOut31_9[5] , 
        \nOut30_11[4] , \nScanOut956[5] , \nOut31_30[2] , \nScanOut585[2] , 
        \nOut26_29[3] , \nOut19_12[7] , \nScanOut1012[0] , \nScanOut650[6] , 
        \nOut23_16[7] , \nScanOut764[5] , \nScanOut330[7] , \nOut13_14[3] , 
        \nScanOut404[0] , \nScanOut530[3] , \nOut20_20[2] , \nOut28_31[5] , 
        \nOut7_21[1] , \nScanOut682[0] , \nScanOut805[1] , \nOut29_10[3] , 
        \nScanOut931[2] , \nScanOut66[1] , \nScanOut681[3] , \nScanOut806[2] , 
        \nScanOut167[2] , \nScanOut207[7] , \nOut7_22[2] , \nScanOut932[1] , 
        \nScanOut333[4] , \nScanOut653[5] , \nScanOut767[6] , \nOut6_27[2] , 
        \nScanOut191[2] , \nOut13_17[0] , \nOut29_13[0] , \nScanOut407[3] , 
        \nOut16_28[4] , \nScanOut533[0] , \nOut20_23[1] , \nScanOut822[4] , 
        \nScanOut791[6] , \nScanOut916[7] , \nOut3_18[6] , \nOut28_9[1] , 
        \nScanOut90[1] , \nScanOut143[4] , \nOut12_12[0] , \nScanOut423[5] , 
        \nScanOut517[6] , \nOut24_8[0] , \nOut21_26[1] , \nOut24_19[5] , 
        \nScanOut677[3] , \nOut28_16[0] , \nScanOut743[0] , \nScanOut93[2] , 
        \nScanOut140[7] , \nScanOut223[1] , \nScanOut317[2] , \nOut22_8[4] , 
        \nScanOut220[2] , \nOut12_11[3] , \nOut28_15[3] , \nOut13_30[5] , 
        \nScanOut420[6] , \nScanOut514[5] , \nOut21_25[2] , \nScanOut314[1] , 
        \nScanOut674[0] , \nScanOut740[3] , \nScanOut192[1] , \nScanOut792[5] , 
        \nScanOut821[7] , \nScanOut127[0] , \nOut6_24[1] , \nScanOut915[4] , 
        \nOut5_12[4] , \nScanOut247[5] , \nScanOut447[1] , \nScanOut573[2] , 
        \nOut19_8[4] , \nOut6_9[0] , \nOut11_27[6] , \nScanOut373[6] , 
        \nOut14_18[2] , \nScanOut613[7] , \nScanOut894[6] , \nOut22_13[7] , 
        \nScanOut727[4] , \nOut15_9[5] , \nOut18_17[7] , \nScanOut495[7] , 
        \nOut0_11[6] , \nOut0_12[5] , \nScanOut25[0] , \nScanOut26[3] , 
        \nScanOut295[3] , \nOut13_9[1] , \nOut31_14[4] , \nScanOut846[0] , 
        \nOut11_24[5] , \nScanOut972[3] , \nScanOut496[4] , \nOut18_14[4] , 
        \nOut22_10[4] , \nOut23_31[2] , \nScanOut845[3] , \nScanOut971[0] , 
        \nOut1_14[4] , \nOut1_17[7] , \nOut2_21[2] , \nOut2_22[1] , 
        \nScanOut124[3] , \nScanOut296[0] , \nScanOut444[2] , \nScanOut570[1] , 
        \nOut31_17[7] , \nOut4_30[1] , \nOut5_11[7] , \nScanOut244[6] , 
        \nScanOut610[4] , \nScanOut724[7] , \nScanOut897[5] , \nScanOut370[5] , 
        \nScanOut158[5] , \nOut13_28[7] , \nOut25_23[2] , \nScanOut238[0] , 
        \nScanOut438[4] , \nOut16_17[3] , \nScanOut758[1] , \nScanOut59[6] , 
        \nScanOut839[5] , \nScanOut189[0] , \nScanOut789[4] , \nScanOut88[3] , 
        \nOut16_14[0] , \nOut25_20[1] , \nOut15_22[5] , \nOut26_16[4] , 
        \nScanOut568[3] , \nOut23_29[0] , \nScanOut969[2] , \nOut30_2[1] , 
        \nOut4_28[3] , \nOut8_27[6] , \nScanOut608[6] , \nScanOut368[7] , 
        \nOut8_24[5] , \nOut30_1[2] , \nScanOut118[5] , \nOut15_21[6] , 
        \nOut20_7[3] , \nOut26_15[7] , \nScanOut278[0] , \nOut9_22[4] , 
        \nScanOut478[4] , \nOut18_3[2] , \nScanOut718[1] , \nOut26_7[7] , 
        \nScanOut19[6] , \nOut1_2[2] , \nOut7_2[6] , \nOut14_2[3] , 
        \nOut14_27[7] , \nOut18_28[2] , \nScanOut1009[3] , \nOut11_18[3] , 
        \nOut27_13[6] , \nOut12_2[7] , \nOut1_1[1] , \nOut7_1[5] , 
        \nOut27_10[5] , \nOut26_31[3] , \nScanOut879[5] , \nOut12_1[4] , 
        \nOut14_1[0] , \nOut14_24[4] , \nOut20_4[0] , \nOut31_28[2] , 
        \nOut26_4[4] , \nScanOut25[2] , \nOut2_5[0] , \nOut2_6[3] , 
        \nOut1_30[0] , \nOut9_21[7] , \nOut18_0[1] , \nOut11_6[6] , 
        \nOut3_27[3] , \nOut4_6[7] , \nOut6_18[7] , \nScanOut929[2] , 
        \nOut29_2[7] , \nOut8_4[5] , \nOut8_7[6] , \nOut17_6[2] , 
        \nOut17_12[1] , \nOut21_19[4] , \nScanOut328[7] , \nScanOut528[3] , 
        \nOut25_3[6] , \nScanOut648[6] , \nOut24_26[0] , \nOut28_29[5] , 
        \nOut23_3[2] , \nOut24_25[3] , \nOut16_30[4] , \nOut17_11[2] , 
        \nOut25_0[5] , \nOut23_0[1] , \nScanOut41[6] , \nOut1_28[2] , 
        \nOut3_24[0] , \nOut11_5[5] , \nOut17_5[1] , \nOut4_5[4] , 
        \nOut29_1[4] , \nScanOut103[4] , \nOut10_22[4] , \nScanOut585[0] , 
        \nScanOut699[3] , \nScanOut1012[2] , \nOut26_29[1] , \nScanOut385[4] , 
        \nOut19_12[5] , \nOut23_16[5] , \nScanOut862[4] , \nScanOut956[7] , 
        \nOut30_11[6] , \nOut31_30[0] , \nScanOut463[5] , \nScanOut557[6] , 
        \nOut31_9[7] , \nScanOut637[3] , \nScanOut703[0] , \nScanOut984[1] , 
        \nScanOut65[0] , \nScanOut66[3] , \nScanOut100[7] , \nOut4_17[6] , 
        \nScanOut357[2] , \nOut8_18[3] , \nScanOut263[1] , \nOut4_14[5] , 
        \nScanOut354[1] , \nScanOut460[6] , \nScanOut554[5] , \nScanOut167[0] , 
        \nScanOut260[2] , \nOut10_21[7] , \nOut18_30[0] , \nScanOut634[0] , 
        \nScanOut700[3] , \nScanOut987[2] , \nOut23_15[6] , \nOut19_11[6] , 
        \nScanOut1011[1] , \nScanOut386[7] , \nScanOut586[3] , 
        \nScanOut861[7] , \nOut30_12[5] , \nScanOut955[4] , \nOut29_13[2] , 
        \nScanOut207[5] , \nScanOut333[6] , \nOut13_17[2] , \nScanOut407[1] , 
        \nOut16_28[6] , \nScanOut533[2] , \nOut20_23[3] , \nScanOut653[7] , 
        \nScanOut767[4] , \nOut7_21[3] , \nOut7_22[0] , \nScanOut681[1] , 
        \nScanOut932[3] , \nScanOut806[0] , \nScanOut931[0] , \nScanOut164[3] , 
        \nOut13_14[1] , \nScanOut404[2] , \nScanOut682[2] , \nScanOut805[3] , 
        \nScanOut530[1] , \nOut20_20[0] , \nOut29_10[1] , \nScanOut204[6] , 
        \nScanOut330[5] , \nScanOut650[4] , \nScanOut764[7] , \nOut28_31[7] , 
        \nScanOut42[5] , \nScanOut90[3] , \nScanOut93[0] , \nOut6_24[3] , 
        \nScanOut792[7] , \nScanOut915[6] , \nScanOut192[3] , \nScanOut821[5] , 
        \nScanOut220[0] , \nScanOut314[3] , \nScanOut140[5] , \nScanOut674[2] , 
        \nScanOut740[1] , \nOut28_15[1] , \nOut12_11[1] , \nOut13_30[7] , 
        \nScanOut420[4] , \nOut21_25[0] , \nScanOut514[7] , \nScanOut143[6] , 
        \nScanOut223[3] , \nScanOut317[0] , \nScanOut677[1] , \nScanOut743[2] , 
        \nOut22_8[6] , \nOut12_12[2] , \nScanOut423[7] , \nOut21_26[3] , 
        \nScanOut517[4] , \nOut24_8[2] , \nOut24_19[7] , \nOut28_16[2] , 
        \nOut6_27[0] , \nScanOut916[5] , \nOut28_9[3] , \nOut3_18[4] , 
        \nScanOut791[4] , \nScanOut822[6] , \nScanOut124[1] , \nOut4_30[3] , 
        \nScanOut191[0] , \nScanOut610[6] , \nScanOut724[5] , \nScanOut897[7] , 
        \nOut5_11[5] , \nScanOut370[7] , \nScanOut244[4] , \nScanOut444[0] , 
        \nScanOut570[3] , \nScanOut971[2] , \nScanOut295[1] , \nScanOut296[2] , 
        \nScanOut845[1] , \nOut31_17[5] , \nOut11_24[7] , \nScanOut496[6] , 
        \nOut18_14[6] , \nOut22_10[6] , \nOut23_31[0] , \nOut31_14[6] , 
        \nScanOut26[1] , \nOut1_14[6] , \nOut2_21[0] , \nScanOut88[1] , 
        \nScanOut127[2] , \nOut5_12[6] , \nOut6_9[2] , \nOut13_9[3] , 
        \nScanOut972[1] , \nOut14_18[0] , \nScanOut846[2] , \nOut15_9[7] , 
        \nOut22_13[5] , \nScanOut495[5] , \nOut18_17[5] , \nOut11_27[4] , 
        \nScanOut373[4] , \nScanOut247[7] , \nOut19_8[6] , \nScanOut613[5] , 
        \nScanOut727[6] , \nScanOut894[4] , \nScanOut447[3] , \nScanOut573[0] , 
        \nOut16_14[2] , \nOut25_20[3] , \nScanOut789[6] , \nOut2_22[3] , 
        \nScanOut189[2] , \nScanOut59[4] , \nScanOut158[7] , \nScanOut238[2] , 
        \nScanOut839[7] , \nOut13_28[5] , \nScanOut758[3] , \nOut25_23[0] , 
        \nOut8_24[7] , \nScanOut438[6] , \nOut16_17[1] , \nOut15_21[4] , 
        \nOut26_15[5] , \nOut1_17[5] , \nOut30_1[0] , \nOut4_28[1] , 
        \nOut8_27[4] , \nScanOut608[4] , \nScanOut298[4] , \nScanOut368[5] , 
        \nOut13_4[6] , \nOut15_22[7] , \nScanOut568[1] , \nOut23_29[2] , 
        \nOut26_16[6] , \nOut30_2[3] , \nScanOut969[0] , \nOut31_19[3] , 
        \nOut0_7[0] , \nOut0_20[7] , \nOut6_4[7] , \nScanOut498[0] , 
        \nOut14_15[5] , \nOut27_21[4] , \nOut15_4[2] , \nScanOut899[1] , 
        \nOut0_23[4] , \nScanOut249[1] , \nOut9_10[6] , \nOut27_1[6] , 
        \nOut9_13[5] , \nOut8_31[0] , \nOut19_5[3] , \nOut21_1[2] , 
        \nOut19_6[0] , \nScanOut729[0] , \nOut27_2[5] , \nScanOut129[4] , 
        \nOut21_2[1] , \nScanOut449[5] , \nScanOut28[7] , \nScanOut30[5] , 
        \nOut3_3[1] , \nOut3_15[1] , \nOut6_7[4] , \nOut13_7[5] , 
        \nScanOut848[4] , \nOut14_16[6] , \nOut15_7[1] , \nOut18_19[3] , 
        \nOut9_1[7] , \nOut11_29[2] , \nOut27_22[7] , \nOut17_20[3] , 
        \nOut22_5[3] , \nOut24_14[2] , \nOut16_0[3] , \nOut24_5[7] , 
        \nOut3_16[2] , \nOut3_0[2] , \nOut5_0[6] , \nOut28_4[6] , \nOut5_3[5] , 
        \nOut10_0[7] , \nOut28_7[5] , \nOut6_29[6] , \nScanOut918[3] , 
        \nOut16_3[0] , \nOut10_3[4] , \nOut4_25[4] , \nOut9_2[4] , 
        \nScanOut319[6] , \nOut22_6[0] , \nScanOut679[7] , \nScanOut519[2] , 
        \nOut17_23[0] , \nOut21_28[5] , \nOut24_6[4] , \nOut24_17[1] , 
        \nOut28_18[4] , \nScanOut131[6] , \nScanOut251[3] , \nScanOut365[0] , 
        \nScanOut605[1] , \nScanOut731[2] , \nScanOut882[0] , \nScanOut283[5] , 
        \nScanOut451[7] , \nScanOut565[4] , \nOut30_23[4] , \nScanOut33[6] , 
        \nOut10_10[6] , \nOut11_31[0] , \nScanOut483[1] , \nOut19_20[7] , 
        \nOut23_24[7] , \nScanOut850[6] , \nScanOut964[5] , \nScanOut1020[0] , 
        \nScanOut967[6] , \nOut1_19[3] , \nScanOut280[6] , \nScanOut853[5] , 
        \nOut30_20[7] , \nOut10_13[5] , \nScanOut480[2] , \nScanOut1023[3] , 
        \nOut19_23[4] , \nOut26_18[0] , \nScanOut606[2] , \nOut23_27[4] , 
        \nScanOut732[1] , \nScanOut54[1] , \nOut4_26[7] , \nScanOut881[3] , 
        \nScanOut132[5] , \nScanOut252[0] , \nOut8_29[2] , \nScanOut366[3] , 
        \nScanOut452[4] , \nScanOut566[7] , \nOut7_10[2] , \nOut6_31[4] , 
        \nScanOut900[1] , \nScanOut86[7] , \nScanOut187[4] , \nScanOut787[0] , 
        \nScanOut834[2] , \nScanOut235[7] , \nScanOut301[4] , \nScanOut661[5] , 
        \nScanOut755[6] , \nOut13_25[0] , \nScanOut435[3] , \nOut20_11[1] , 
        \nOut21_30[7] , \nScanOut501[0] , \nOut29_21[0] , \nScanOut2[0] , 
        \nScanOut85[4] , \nScanOut155[2] , \nScanOut236[4] , \nScanOut302[7] , 
        \nScanOut662[6] , \nScanOut756[5] , \nOut2_8[5] , \nScanOut57[2] , 
        \nScanOut156[1] , \nOut29_22[3] , \nOut13_26[3] , \nScanOut436[0] , 
        \nOut16_19[7] , \nOut20_12[2] , \nScanOut502[3] , \nScanOut172[7] , 
        \nScanOut184[7] , \nOut7_13[1] , \nScanOut784[3] , \nScanOut903[2] , 
        \nScanOut837[1] , \nOut8_9[0] , \nOut12_23[3] , \nScanOut412[6] , 
        \nOut21_17[2] , \nScanOut526[5] , \nOut24_28[6] , \nScanOut212[2] , 
        \nScanOut326[1] , \nScanOut646[0] , \nScanOut772[3] , \nOut28_27[3] , 
        \nOut11_8[0] , \nScanOut70[7] , \nScanOut73[4] , \nOut6_16[1] , 
        \nScanOut927[4] , \nOut3_29[5] , \nOut4_8[1] , \nScanOut813[7] , 
        \nScanOut694[6] , \nOut17_8[4] , \nScanOut171[4] , \nOut6_15[2] , 
        \nScanOut924[7] , \nScanOut697[5] , \nScanOut810[4] , \nScanOut211[1] , 
        \nScanOut325[2] , \nOut12_20[0] , \nOut28_24[0] , \nScanOut411[5] , 
        \nOut21_14[1] , \nScanOut525[6] , \nOut14_29[1] , \nScanOut645[3] , 
        \nScanOut771[0] , \nOut22_22[4] , \nOut18_26[4] , \nOut11_16[5] , 
        \nScanOut590[7] , \nScanOut1007[5] , \nScanEnable[0] , \nScanOut14[3] , 
        \nScanOut17[0] , \nScanOut390[3] , \nOut31_25[7] , \nScanOut115[0] , 
        \nScanOut116[3] , \nScanOut877[3] , \nScanOut943[0] , \nOut5_23[7] , 
        \nScanOut342[5] , \nScanOut476[2] , \nOut20_9[5] , \nScanOut542[1] , 
        \nScanOut276[6] , \nScanOut475[1] , \nScanOut622[4] , \nScanOut716[7] , 
        \nOut26_9[1] , \nScanOut991[6] , \nScanOut541[2] , \nOut5_20[4] , 
        \nScanOut341[6] , \nScanOut621[7] , \nScanOut715[4] , \nScanOut992[5] , 
        \nScanOut275[5] , \nOut11_15[6] , \nScanOut593[4] , \nScanOut1004[6] , 
        \nOut18_25[7] , \nOut22_21[7] , \nScanOut940[3] , \nOut2_10[1] , 
        \nOut2_13[2] , \nScanOut393[0] , \nScanOut874[0] , \nOut31_26[4] , 
        \nScanOut68[5] , \nScanOut169[6] , \nOut13_19[4] , \nOut25_12[1] , 
        \nScanOut808[6] , \nScanOut209[3] , \nScanOut409[7] , \nOut16_26[0] , 
        \nOut16_25[3] , \nScanOut769[2] , \nOut24_30[4] , \nOut25_11[2] , 
        \nScanOut49[7] , \nOut1_25[7] , \nOut1_26[4] , \nOut3_31[7] , 
        \nScanOut559[0] , \nOut31_7[1] , \nOut4_19[0] , \nOut8_16[5] , 
        \nScanOut639[5] , \nScanOut359[4] , \nOut8_15[6] , \nScanOut388[1] , 
        \nOut15_10[5] , \nOut15_13[6] , \nOut26_27[7] , \nOut23_18[3] , 
        \nScanOut958[1] , \nOut14_31[3] , \nScanOut588[5] , \nOut26_24[4] , 
        \nOut31_4[2] , \nScanOut989[4] , \nOut3_6[5] , \nScanOut148[4] , 
        \nOut9_7[0] , \nScanOut428[5] , \nOut17_26[4] , \nOut12_19[0] , 
        \nOut24_3[0] , \nOut24_12[5] , \nScanOut228[1] , \nOut22_3[4] , 
        \nScanOut748[0] , \nOut10_6[0] , \nOut3_5[6] , \nOut3_13[6] , 
        \nOut5_6[1] , \nOut28_2[1] , \nOut16_6[4] , \nScanOut829[4] , 
        \nOut3_10[5] , \nScanOut199[1] , \nOut10_5[3] , \nOut16_5[7] , 
        \nOut2_31[3] , \nOut0_1[7] , \nOut0_2[4] , \nScanOut98[2] , 
        \nOut5_5[2] , \nOut28_1[2] , \nOut9_4[3] , \nOut17_25[7] , 
        \nOut24_11[6] , \nOut25_30[0] , \nScanOut799[5] , \nOut22_0[7] , 
        \nOut24_0[3] , \nOut6_2[0] , \nOut14_13[2] , \nOut22_18[7] , 
        \nOut15_2[5] , \nOut27_27[3] , \nOut0_25[3] , \nOut0_26[0] , 
        \nOut5_19[4] , \nOut9_16[1] , \nOut13_2[1] , \nScanOut979[3] , 
        \nScanOut578[2] , \nOut21_7[5] , \nScanOut378[6] , \nOut19_3[4] , 
        \nScanOut618[7] , \nOut27_7[1] , \nOut21_4[6] , \nOut27_4[2] , 
        \nOut6_1[3] , \nOut9_15[2] , \nOut19_0[7] , \nOut13_1[2] , 
        \nOut14_10[1] , \nOut15_1[6] , \nOut27_24[0] , \nOut15_31[7] , 
        \nScanOut4[7] , \nScanOut7[4] , \nScanOut52[6] , \nOut2_29[1] , 
        \nScanOut181[3] , \nOut7_16[5] , \nScanOut906[6] , \nOut13_23[7] , 
        \nScanOut781[7] , \nOut25_28[2] , \nScanOut832[5] , \nOut29_27[7] , 
        \nScanOut80[0] , \nScanOut153[5] , \nScanOut233[0] , \nScanOut307[3] , 
        \nScanOut433[4] , \nOut20_17[6] , \nScanOut507[7] , \nScanOut430[7] , 
        \nOut20_14[5] , \nScanOut667[2] , \nScanOut753[1] , \nScanOut504[4] , 
        \nScanOut11[7] , \nScanOut35[1] , \nScanOut36[2] , \nScanOut51[5] , 
        \nScanOut83[3] , \nScanOut150[6] , \nOut29_24[4] , \nOut13_20[4] , 
        \nScanOut182[0] , \nScanOut230[3] , \nScanOut304[0] , \nScanOut664[1] , 
        \nScanOut750[2] , \nOut4_23[3] , \nScanOut137[1] , \nOut7_15[6] , 
        \nScanOut782[4] , \nScanOut905[5] , \nScanOut457[0] , \nScanOut831[6] , 
        \nScanOut563[3] , \nScanOut603[6] , \nScanOut737[5] , \nOut30_9[1] , 
        \nScanOut884[7] , \nScanOut257[4] , \nScanOut363[7] , \nOut10_16[1] , 
        \nScanOut485[6] , \nOut15_29[5] , \nOut19_26[0] , \nOut23_22[0] , 
        \nScanOut285[2] , \nScanOut856[1] , \nScanOut962[2] , \nOut30_25[3] , 
        \nScanOut286[1] , \nOut10_15[2] , \nScanOut486[5] , \nOut19_25[3] , 
        \nOut23_21[3] , \nOut30_26[0] , \nScanOut961[1] , \nOut4_20[0] , 
        \nScanOut134[2] , \nScanOut855[2] , \nScanOut454[3] , \nScanOut560[0] , 
        \nScanOut254[7] , \nScanOut360[4] , \nScanOut600[5] , \nScanOut734[6] , 
        \nScanOut887[4] , \nScanOut12[4] , \nOut0_19[7] , \nScanOut110[4] , 
        \nOut5_25[0] , \nOut11_10[2] , \nOut10_31[4] , \nScanOut396[4] , 
        \nScanOut871[4] , \nScanOut945[7] , \nOut31_23[0] , \nScanOut1001[2] , 
        \nScanOut596[0] , \nScanOut344[2] , \nOut18_20[3] , \nOut22_24[3] , 
        \nScanOut624[3] , \nScanOut710[0] , \nScanOut997[1] , \nScanOut270[1] , 
        \nScanOut470[5] , \nScanOut544[6] , \nOut5_26[3] , \nScanOut347[1] , 
        \nScanOut273[2] , \nOut9_29[6] , \nOut18_8[0] , \nScanOut627[0] , 
        \nScanOut713[3] , \nScanOut994[2] , \nOut1_9[0] , \nScanOut113[7] , 
        \nScanOut395[7] , \nScanOut473[6] , \nScanOut547[5] , \nOut31_20[3] , 
        \nScanOut946[4] , \nOut1_20[3] , \nScanOut75[3] , \nOut6_10[6] , 
        \nScanOut174[0] , \nOut7_9[4] , \nOut12_9[5] , \nOut14_9[1] , 
        \nOut18_23[0] , \nScanOut872[7] , \nOut22_27[0] , \nScanOut595[3] , 
        \nScanOut1002[1] , \nOut27_18[4] , \nScanOut214[5] , \nScanOut320[6] , 
        \nOut11_13[1] , \nOut12_25[4] , \nScanOut640[7] , \nScanOut774[4] , 
        \nOut7_31[0] , \nScanOut414[1] , \nOut21_11[5] , \nOut28_21[4] , 
        \nScanOut520[2] , \nOut20_30[3] , \nScanOut921[3] , \nScanOut76[0] , 
        \nScanOut692[1] , \nScanOut815[0] , \nOut6_13[5] , \nScanOut922[0] , 
        \nScanOut177[3] , \nScanOut217[6] , \nScanOut323[5] , \nScanOut643[4] , 
        \nScanOut691[2] , \nOut29_9[5] , \nScanOut777[7] , \nScanOut816[3] , 
        \nOut23_8[0] , \nScanOut417[2] , \nOut17_19[3] , \nOut21_12[6] , 
        \nScanOut523[1] , \nOut25_8[4] , \nOut8_10[2] , \nOut12_26[7] , 
        \nOut28_22[7] , \nOut9_31[4] , \nOut31_1[6] , \nOut2_15[5] , 
        \nOut1_23[0] , \nOut10_29[6] , \nOut15_15[1] , \nOut30_19[7] , 
        \nOut26_21[0] , \nScanOut869[6] , \nScanOut1019[0] , \nOut15_16[2] , 
        \nOut19_19[7] , \nOut26_22[3] , \nScanOut708[2] , \nScanOut108[6] , 
        \nOut8_13[1] , \nScanOut268[3] , \nScanOut468[7] , \nOut31_2[5] , 
        \nScanOut689[0] , \nOut0_14[2] , \nOut2_3[7] , \nOut2_16[6] , 
        \nScanOut338[4] , \nOut16_20[7] , \nOut25_14[6] , \nOut16_23[4] , 
        \nOut20_28[1] , \nScanOut658[5] , \nOut25_17[5] , \nOut29_18[0] , 
        \nScanOut538[0] , \nOut2_0[4] , \nOut3_21[4] , \nOut7_29[2] , 
        \nScanOut939[1] , \nOut4_0[0] , \nOut17_0[5] , \nOut29_4[0] , 
        \nScanOut78[6] , \nScanOut179[5] , \nScanOut219[0] , \nOut8_1[1] , 
        \nOut11_0[1] , \nOut17_14[6] , \nOut23_5[5] , \nOut24_20[7] , 
        \nOut25_5[1] , \nScanOut779[1] , \nOut8_2[2] , \nOut23_6[6] , 
        \nOut12_28[1] , \nScanOut419[4] , \nOut17_17[5] , \nOut25_6[2] , 
        \nOut24_23[4] , \nOut3_22[7] , \nOut4_3[3] , \nScanOut818[5] , 
        \nOut29_7[3] , \nOut17_3[6] , \nOut11_3[2] , \nOut26_1[0] , 
        \nScanOut999[7] , \nOut9_24[3] , \nOut18_5[5] , \nOut12_4[0] , 
        \nOut20_1[4] , \nScanOut1[7] , \nScanOut2[4] , \nScanOut9[2] , 
        \nOut0_17[1] , \nOut1_4[5] , \nScanOut398[2] , \nOut1_7[6] , 
        \nOut7_4[1] , \nScanOut598[6] , \nOut14_4[4] , \nOut14_21[0] , 
        \nOut27_15[1] , \nOut5_28[5] , \nOut7_7[2] , \nOut12_7[3] , 
        \nOut14_7[7] , \nOut14_22[3] , \nScanOut948[2] , \nOut22_29[6] , 
        \nOut27_16[2] , \nOut9_27[0] , \nOut18_6[6] , \nScanOut349[7] , 
        \nOut26_2[3] , \nScanOut20[6] , \nScanOut23[5] , \nOut0_28[6] , 
        \nOut2_18[0] , \nScanOut60[4] , \nScanOut161[7] , \nScanOut201[2] , 
        \nScanOut335[1] , \nScanOut549[3] , \nOut20_2[7] , \nScanOut629[6] , 
        \nScanOut655[0] , \nScanOut761[3] , \nScanOut401[6] , \nScanOut535[5] , 
        \nOut20_25[4] , \nOut29_15[5] , \nOut12_30[3] , \nOut13_11[5] , 
        \nOut7_24[7] , \nScanOut687[6] , \nScanOut934[4] , \nScanOut800[7] , 
        \nScanOut63[7] , \nOut7_27[4] , \nScanOut937[7] , \nScanOut105[3] , 
        \nOut4_11[1] , \nOut5_30[7] , \nScanOut162[4] , \nScanOut202[1] , 
        \nScanOut336[2] , \nScanOut684[5] , \nScanOut803[4] , \nOut13_12[6] , 
        \nScanOut656[3] , \nScanOut762[0] , \nOut25_19[3] , \nOut29_16[6] , 
        \nOut10_24[3] , \nScanOut383[3] , \nScanOut402[5] , \nScanOut536[6] , 
        \nOut20_26[7] , \nOut30_17[1] , \nScanOut583[7] , \nOut19_14[2] , 
        \nScanOut864[3] , \nScanOut950[0] , \nOut23_10[2] , \nOut22_31[4] , 
        \nScanOut1014[5] , \nScanOut351[5] , \nScanOut265[6] , 
        \nScanOut631[4] , \nScanOut705[7] , \nScanOut982[6] , \nScanOut106[0] , 
        \nOut4_12[2] , \nScanOut352[6] , \nScanOut465[2] , \nScanOut551[1] , 
        \nScanOut632[7] , \nScanOut706[4] , \nScanOut981[5] , \nScanOut266[5] , 
        \nScanOut466[1] , \nScanOut552[2] , \nScanOut122[6] , \nOut10_27[0] , 
        \nScanOut380[0] , \nScanOut867[0] , \nScanOut953[3] , \nOut30_14[2] , 
        \nScanOut1017[6] , \nOut15_18[4] , \nScanOut580[4] , \nOut23_13[1] , 
        \nOut19_17[1] , \nOut21_9[3] , \nOut5_17[2] , \nScanOut376[0] , 
        \nScanOut442[7] , \nScanOut576[4] , \nScanOut242[3] , \nOut9_18[7] , 
        \nScanOut616[1] , \nScanOut722[2] , \nScanOut891[0] , \nScanOut290[5] , 
        \nOut11_22[0] , \nScanOut490[1] , \nOut18_12[1] , \nOut27_9[7] , 
        \nOut22_16[1] , \nOut27_29[5] , \nOut30_30[4] , \nOut31_11[2] , 
        \nScanOut977[5] , \nOut11_21[3] , \nScanOut493[2] , \nScanOut843[6] , 
        \nOut18_11[2] , \nOut19_30[4] , \nOut22_15[2] , \nOut0_30[4] , 
        \nScanOut38[4] , \nScanOut44[2] , \nScanOut47[1] , \nOut3_8[3] , 
        \nScanOut121[5] , \nScanOut293[6] , \nScanOut840[5] , \nScanOut974[6] , 
        \nOut31_12[1] , \nScanOut441[4] , \nScanOut575[7] , \nOut5_14[1] , 
        \nScanOut375[3] , \nScanOut615[2] , \nScanOut721[1] , \nScanOut892[3] , 
        \nScanOut241[0] , \nOut10_8[6] , \nScanOut194[4] , \nScanOut95[7] , 
        \nOut5_8[7] , \nScanOut146[2] , \nOut6_22[4] , \nScanOut794[0] , 
        \nScanOut913[1] , \nOut9_9[6] , \nScanOut426[3] , \nOut16_8[2] , 
        \nScanOut827[2] , \nOut21_23[7] , \nScanOut512[0] , \nOut17_28[2] , 
        \nOut28_13[6] , \nOut12_17[6] , \nScanOut96[4] , \nScanOut145[1] , 
        \nScanOut226[7] , \nScanOut312[4] , \nScanOut672[5] , \nScanOut746[6] , 
        \nOut12_14[5] , \nOut28_10[5] , \nOut29_31[3] , \nScanOut225[4] , 
        \nScanOut311[7] , \nScanOut425[0] , \nOut21_20[4] , \nScanOut511[3] , 
        \nOut6_21[7] , \nScanOut197[7] , \nScanOut671[6] , \nScanOut745[5] , 
        \nScanOut910[2] , \nOut10_18[7] , \nScanOut797[3] , \nOut26_13[2] , 
        \nScanOut824[1] , \nOut15_27[3] , \nOut19_28[6] , \nOut1_11[2] , 
        \nOut1_12[1] , \nScanOut139[7] , \nScanOut459[6] , \nScanOut858[7] , 
        \nOut30_7[7] , \nScanOut739[3] , \nOut8_21[3] , \nOut8_22[0] , 
        \nScanOut259[2] , \nOut30_4[4] , \nScanOut889[2] , \nScanOut288[7] , 
        \nOut15_24[0] , \nScanOut488[3] , \nOut26_10[1] , \nOut27_31[7] , 
        \nOut30_28[6] , \nOut29_29[1] , \nScanOut14[7] , \nOut2_8[1] , 
        \nOut2_10[5] , \nOut2_24[4] , \nOut2_27[7] , \nScanOut309[5] , 
        \nOut16_12[5] , \nOut25_26[4] , \nScanOut509[1] , \nOut20_19[0] , 
        \nScanOut669[4] , \nOut7_18[3] , \nScanOut908[0] , \nOut16_11[6] , 
        \nOut17_30[0] , \nOut25_25[7] , \nOut2_13[6] , \nScanOut68[1] , 
        \nOut3_31[3] , \nScanOut169[2] , \nScanOut209[7] , \nOut16_25[7] , 
        \nOut24_30[0] , \nOut25_11[6] , \nScanOut769[6] , \nOut13_19[0] , 
        \nScanOut409[3] , \nOut16_26[4] , \nOut25_12[5] , \nScanOut808[2] , 
        \nOut1_25[3] , \nScanOut989[0] , \nOut1_26[0] , \nOut4_19[4] , 
        \nOut8_15[2] , \nOut8_16[1] , \nScanOut388[5] , \nOut31_4[6] , 
        \nOut15_10[1] , \nScanOut588[1] , \nOut26_24[0] , \nOut15_13[2] , 
        \nOut14_31[7] , \nOut23_18[7] , \nScanOut958[5] , \nOut26_27[3] , 
        \nScanOut359[0] , \nScanOut70[3] , \nScanOut171[0] , \nScanOut211[5] , 
        \nScanOut325[6] , \nScanOut559[4] , \nScanOut639[1] , \nOut31_7[5] , 
        \nScanOut645[7] , \nScanOut771[4] , \nScanOut411[1] , \nOut21_14[5] , 
        \nScanOut525[2] , \nOut12_20[4] , \nOut28_24[4] , \nScanOut73[0] , 
        \nOut3_29[1] , \nOut6_15[6] , \nScanOut924[3] , \nOut17_8[0] , 
        \nScanOut697[1] , \nScanOut810[0] , \nOut6_16[5] , \nScanOut927[0] , 
        \nOut4_8[5] , \nScanOut813[3] , \nScanOut694[2] , \nScanOut172[3] , 
        \nScanOut212[6] , \nScanOut326[5] , \nOut11_8[4] , \nOut12_23[7] , 
        \nScanOut646[4] , \nScanOut772[7] , \nOut24_28[2] , \nOut8_9[4] , 
        \nOut28_27[7] , \nScanOut393[4] , \nScanOut412[2] , \nOut21_17[6] , 
        \nScanOut526[1] , \nOut31_26[0] , \nScanOut940[7] , \nScanOut17[4] , 
        \nScanOut115[4] , \nOut5_20[0] , \nOut11_15[2] , \nOut18_25[3] , 
        \nScanOut874[4] , \nScanOut593[0] , \nOut22_21[3] , \nScanOut1004[2] , 
        \nScanOut341[2] , \nScanOut275[1] , \nScanOut621[3] , \nScanOut715[0] , 
        \nScanOut992[1] , \nScanOut116[7] , \nOut5_23[3] , \nScanOut342[1] , 
        \nScanOut475[5] , \nScanOut541[6] , \nScanOut622[0] , \nScanOut716[3] , 
        \nOut26_9[5] , \nScanOut991[2] , \nScanOut276[2] , \nScanOut476[6] , 
        \nScanOut542[5] , \nOut20_9[1] , \nScanOut30[1] , \nScanOut33[2] , 
        \nOut1_19[7] , \nOut4_26[3] , \nScanOut132[1] , \nOut11_16[1] , 
        \nScanOut390[7] , \nScanOut877[7] , \nScanOut943[4] , \nScanOut590[3] , 
        \nOut31_25[3] , \nScanOut1007[1] , \nOut14_29[5] , \nOut18_26[0] , 
        \nOut22_22[0] , \nScanOut452[0] , \nScanOut566[3] , \nScanOut252[4] , 
        \nOut8_29[6] , \nScanOut366[7] , \nScanOut606[6] , \nScanOut732[5] , 
        \nScanOut280[2] , \nOut10_13[1] , \nScanOut480[6] , \nOut19_23[0] , 
        \nScanOut881[7] , \nOut23_27[0] , \nOut26_18[4] , \nScanOut1023[7] , 
        \nOut30_20[3] , \nScanOut967[2] , \nOut10_10[2] , \nOut11_31[4] , 
        \nScanOut483[5] , \nScanOut853[1] , \nScanOut1020[4] , \nOut19_20[3] , 
        \nOut23_24[3] , \nScanOut57[6] , \nOut4_25[0] , \nScanOut131[2] , 
        \nScanOut283[1] , \nScanOut850[2] , \nScanOut964[1] , \nOut30_23[0] , 
        \nScanOut451[3] , \nScanOut565[0] , \nScanOut605[5] , \nScanOut731[6] , 
        \nScanOut882[4] , \nScanOut184[3] , \nScanOut251[7] , \nScanOut365[4] , 
        \nOut7_13[5] , \nScanOut784[7] , \nScanOut903[6] , \nScanOut436[4] , 
        \nOut16_19[3] , \nScanOut837[5] , \nOut20_12[6] , \nScanOut502[7] , 
        \nOut29_22[7] , \nScanOut85[0] , \nScanOut156[5] , \nOut13_26[7] , 
        \nScanOut236[0] , \nScanOut302[3] , \nScanOut662[2] , \nScanOut756[1] , 
        \nOut13_25[4] , \nScanOut155[6] , \nOut29_21[4] , \nScanOut301[0] , 
        \nScanOut435[7] , \nOut20_11[5] , \nOut21_30[3] , \nScanOut501[4] , 
        \nOut0_4[7] , \nOut0_7[4] , \nScanOut28[3] , \nScanOut54[5] , 
        \nScanOut86[3] , \nScanOut235[3] , \nScanOut187[0] , \nScanOut661[1] , 
        \nScanOut755[2] , \nOut7_10[6] , \nOut6_31[0] , \nScanOut900[5] , 
        \nOut6_7[0] , \nScanOut787[4] , \nScanOut834[6] , \nOut11_29[6] , 
        \nOut14_16[2] , \nOut15_7[5] , \nOut27_22[3] , \nOut18_19[7] , 
        \nOut13_7[1] , \nScanOut848[0] , \nOut0_20[3] , \nOut0_23[0] , 
        \nScanOut129[0] , \nScanOut449[1] , \nOut21_2[5] , \nScanOut729[4] , 
        \nScanOut249[5] , \nOut9_13[1] , \nOut27_2[1] , \nOut9_10[2] , 
        \nOut19_6[4] , \nOut21_1[6] , \nOut8_31[4] , \nOut19_5[7] , 
        \nOut27_1[2] , \nScanOut899[5] , \nOut6_4[3] , \nOut14_15[1] , 
        \nOut15_4[6] , \nScanOut498[4] , \nScanOut298[0] , \nOut27_21[0] , 
        \nOut31_19[7] , \nScanOut9[6] , \nOut0_9[2] , \nScanOut26[5] , 
        \nScanOut41[2] , \nScanOut42[1] , \nOut1_14[2] , \nOut1_17[1] , 
        \nOut2_21[4] , \nOut2_22[7] , \nScanOut59[0] , \nOut3_3[5] , 
        \nOut9_2[0] , \nOut13_4[2] , \nScanOut519[6] , \nOut17_23[4] , 
        \nOut21_28[1] , \nOut24_17[5] , \nOut28_18[0] , \nScanOut319[2] , 
        \nOut22_6[4] , \nOut24_6[0] , \nScanOut679[3] , \nOut3_15[5] , 
        \nOut3_16[6] , \nOut10_3[0] , \nOut16_3[4] , \nOut3_0[6] , 
        \nOut5_3[1] , \nOut28_7[1] , \nOut6_29[2] , \nScanOut918[7] , 
        \nOut10_0[3] , \nOut5_0[2] , \nOut28_4[2] , \nOut16_0[7] , 
        \nScanOut158[3] , \nOut9_1[3] , \nOut17_20[7] , \nOut13_28[1] , 
        \nScanOut438[2] , \nOut16_17[5] , \nOut22_5[7] , \nOut24_5[3] , 
        \nOut24_14[6] , \nOut25_23[4] , \nScanOut238[6] , \nScanOut758[7] , 
        \nScanOut839[3] , \nScanOut189[6] , \nScanOut88[5] , \nOut16_14[6] , 
        \nOut25_20[7] , \nScanOut789[2] , \nOut4_28[5] , \nOut8_27[0] , 
        \nOut15_22[3] , \nScanOut568[5] , \nOut23_29[6] , \nOut26_16[2] , 
        \nOut30_2[7] , \nScanOut969[4] , \nScanOut368[1] , \nScanOut608[0] , 
        \nOut30_1[4] , \nOut3_18[0] , \nScanOut191[4] , \nOut8_24[3] , 
        \nOut15_21[0] , \nOut26_15[1] , \nOut6_27[4] , \nScanOut916[1] , 
        \nScanOut90[7] , \nScanOut143[2] , \nOut12_12[6] , \nScanOut791[0] , 
        \nOut28_9[7] , \nScanOut822[2] , \nOut24_19[3] , \nOut28_16[6] , 
        \nScanOut223[7] , \nScanOut317[4] , \nScanOut423[3] , \nOut21_26[7] , 
        \nScanOut517[0] , \nOut24_8[6] , \nOut22_8[2] , \nScanOut93[4] , 
        \nScanOut140[1] , \nScanOut420[0] , \nOut21_25[4] , \nScanOut677[5] , 
        \nScanOut743[6] , \nScanOut514[3] , \nOut28_15[5] , \nOut12_11[5] , 
        \nOut13_30[3] , \nScanOut192[7] , \nScanOut220[4] , \nScanOut314[7] , 
        \nScanOut674[6] , \nScanOut740[5] , \nScanOut127[6] , \nOut6_24[7] , 
        \nScanOut792[3] , \nScanOut915[2] , \nScanOut447[7] , \nScanOut821[1] , 
        \nScanOut573[4] , \nOut5_12[2] , \nScanOut373[0] , \nScanOut613[1] , 
        \nScanOut727[2] , \nScanOut894[0] , \nOut6_9[6] , \nScanOut247[3] , 
        \nOut19_8[2] , \nScanOut495[1] , \nOut11_27[0] , \nOut14_18[4] , 
        \nOut22_13[1] , \nOut15_9[3] , \nOut18_17[1] , \nScanOut295[5] , 
        \nOut13_9[7] , \nScanOut972[5] , \nScanOut846[6] , \nOut31_14[2] , 
        \nOut0_11[2] , \nScanOut25[6] , \nScanOut296[6] , \nOut11_24[3] , 
        \nScanOut496[2] , \nOut18_14[2] , \nOut22_10[2] , \nOut23_31[4] , 
        \nOut31_17[1] , \nScanOut971[6] , \nOut1_28[6] , \nScanOut100[3] , 
        \nOut4_14[1] , \nScanOut124[5] , \nScanOut845[5] , \nOut4_30[7] , 
        \nScanOut444[4] , \nScanOut570[7] , \nOut5_11[1] , \nScanOut370[3] , 
        \nScanOut244[0] , \nOut10_21[3] , \nScanOut386[3] , \nScanOut610[2] , 
        \nScanOut724[1] , \nScanOut861[3] , \nScanOut897[3] , \nScanOut955[0] , 
        \nScanOut586[7] , \nOut30_12[1] , \nScanOut1011[5] , \nScanOut354[5] , 
        \nOut18_30[4] , \nOut23_15[2] , \nOut19_11[2] , \nScanOut634[4] , 
        \nScanOut700[7] , \nScanOut987[6] , \nScanOut260[6] , \nScanOut460[2] , 
        \nScanOut554[1] , \nOut4_17[2] , \nScanOut357[6] , \nOut8_18[7] , 
        \nScanOut263[5] , \nScanOut637[7] , \nScanOut703[4] , \nScanOut984[5] , 
        \nScanOut65[4] , \nScanOut103[0] , \nOut31_9[3] , \nScanOut164[7] , 
        \nScanOut204[2] , \nOut10_22[0] , \nScanOut385[0] , \nScanOut463[1] , 
        \nScanOut557[2] , \nOut30_11[2] , \nOut31_30[4] , \nOut19_12[1] , 
        \nScanOut862[0] , \nScanOut956[3] , \nOut23_16[1] , \nScanOut1012[6] , 
        \nScanOut330[1] , \nScanOut585[4] , \nOut26_29[5] , \nOut13_14[5] , 
        \nScanOut650[0] , \nScanOut764[3] , \nOut29_10[5] , \nOut7_21[7] , 
        \nScanOut404[6] , \nOut28_31[3] , \nScanOut530[5] , \nOut20_20[4] , 
        \nScanOut931[4] , \nScanOut66[7] , \nScanOut682[6] , \nScanOut805[7] , 
        \nScanOut167[4] , \nScanOut207[1] , \nOut7_22[4] , \nScanOut333[2] , 
        \nScanOut653[3] , \nScanOut681[5] , \nScanOut932[7] , \nScanOut767[0] , 
        \nScanOut806[4] , \nScanOut407[5] , \nOut16_28[2] , \nOut20_23[7] , 
        \nScanOut533[6] , \nOut29_13[6] , \nOut9_21[3] , \nOut13_17[6] , 
        \nOut18_0[5] , \nOut26_4[0] , \nOut0_12[1] , \nScanOut19[2] , 
        \nOut1_1[5] , \nOut1_30[4] , \nOut20_4[4] , \nOut7_1[1] , 
        \nOut12_1[0] , \nOut31_28[6] , \nOut14_1[4] , \nOut14_24[0] , 
        \nOut26_31[7] , \nOut27_10[1] , \nOut1_2[6] , \nOut12_2[3] , 
        \nScanOut879[1] , \nOut7_2[2] , \nOut27_13[2] , \nScanOut1009[7] , 
        \nOut11_18[7] , \nOut14_2[7] , \nOut14_27[3] , \nOut18_28[6] , 
        \nScanOut718[5] , \nOut26_7[3] , \nOut0_30[0] , \nOut2_5[4] , 
        \nOut3_24[4] , \nOut4_5[0] , \nScanOut118[1] , \nScanOut278[4] , 
        \nOut9_22[0] , \nOut18_3[6] , \nScanOut478[0] , \nOut20_7[7] , 
        \nOut29_1[0] , \nScanOut699[7] , \nOut11_5[1] , \nOut17_5[5] , 
        \nOut2_6[7] , \nOut3_27[7] , \nOut8_4[1] , \nOut23_0[5] , \nOut8_7[2] , 
        \nScanOut328[3] , \nOut16_30[0] , \nOut17_11[6] , \nOut25_0[1] , 
        \nOut24_25[7] , \nOut17_12[5] , \nScanOut648[2] , \nOut23_3[6] , 
        \nOut24_26[4] , \nOut28_29[1] , \nOut21_19[0] , \nOut17_6[6] , 
        \nScanOut528[7] , \nOut25_3[2] , \nOut4_6[3] , \nOut6_18[3] , 
        \nScanOut929[6] , \nOut29_2[3] , \nOut1_11[6] , \nScanOut288[3] , 
        \nOut11_6[2] , \nOut30_28[2] , \nOut15_24[4] , \nScanOut488[7] , 
        \nOut26_10[5] , \nOut27_31[3] , \nScanOut889[6] , \nScanOut38[0] , 
        \nOut1_12[5] , \nOut8_21[7] , \nOut8_22[4] , \nOut30_4[0] , 
        \nScanOut259[6] , \nScanOut739[7] , \nScanOut139[3] , \nOut30_7[3] , 
        \nScanOut459[2] , \nOut2_24[0] , \nOut10_18[3] , \nOut15_27[7] , 
        \nOut19_28[2] , \nScanOut858[3] , \nOut16_11[2] , \nOut25_25[3] , 
        \nOut26_13[6] , \nOut17_30[4] , \nOut2_27[3] , \nOut7_18[7] , 
        \nScanOut908[4] , \nScanOut309[1] , \nScanOut669[0] , \nOut16_12[1] , 
        \nOut20_19[4] , \nScanOut509[5] , \nOut0_17[5] , \nScanOut20[2] , 
        \nScanOut121[1] , \nOut5_14[5] , \nScanOut375[7] , \nOut25_26[0] , 
        \nOut29_29[5] , \nScanOut241[4] , \nScanOut615[6] , \nScanOut721[5] , 
        \nScanOut892[7] , \nScanOut293[2] , \nScanOut441[0] , \nScanOut575[3] , 
        \nOut31_12[5] , \nScanOut23[1] , \nOut11_21[7] , \nScanOut493[6] , 
        \nOut18_11[6] , \nOut19_30[0] , \nOut22_15[6] , \nScanOut840[1] , 
        \nScanOut974[2] , \nScanOut977[1] , \nOut0_28[2] , \nScanOut290[1] , 
        \nScanOut843[2] , \nOut30_30[0] , \nOut31_11[6] , \nOut11_22[4] , 
        \nScanOut490[5] , \nOut27_29[1] , \nOut18_12[5] , \nScanOut616[5] , 
        \nOut22_16[5] , \nScanOut722[6] , \nOut27_9[3] , \nScanOut891[4] , 
        \nOut2_3[3] , \nScanOut44[6] , \nScanOut122[2] , \nOut5_17[6] , 
        \nScanOut376[4] , \nScanOut242[7] , \nOut9_18[3] , \nScanOut442[3] , 
        \nScanOut576[0] , \nOut21_9[7] , \nOut6_21[3] , \nScanOut910[6] , 
        \nScanOut47[5] , \nScanOut95[3] , \nScanOut96[0] , \nScanOut197[3] , 
        \nScanOut797[7] , \nScanOut824[5] , \nScanOut145[5] , \nScanOut225[0] , 
        \nScanOut311[3] , \nScanOut671[2] , \nScanOut745[1] , \nOut12_14[1] , 
        \nScanOut425[4] , \nOut21_20[0] , \nScanOut511[7] , \nOut28_10[1] , 
        \nOut29_31[7] , \nScanOut226[3] , \nScanOut312[0] , \nScanOut146[6] , 
        \nScanOut672[1] , \nScanOut746[2] , \nOut28_13[2] , \nOut9_9[2] , 
        \nOut12_17[2] , \nScanOut426[7] , \nOut17_28[6] , \nOut21_23[3] , 
        \nScanOut512[4] , \nOut16_8[6] , \nOut2_18[4] , \nScanOut63[3] , 
        \nOut3_8[7] , \nOut5_8[3] , \nOut6_22[0] , \nScanOut794[4] , 
        \nScanOut913[5] , \nScanOut827[6] , \nScanOut162[0] , \nScanOut194[0] , 
        \nOut10_8[2] , \nOut13_12[2] , \nScanOut402[1] , \nScanOut536[2] , 
        \nOut20_26[3] , \nOut25_19[7] , \nOut29_16[2] , \nScanOut202[5] , 
        \nScanOut336[6] , \nScanOut656[7] , \nScanOut762[4] , \nOut7_27[0] , 
        \nScanOut937[3] , \nScanOut684[1] , \nScanOut803[0] , \nScanOut60[0] , 
        \nScanOut105[7] , \nScanOut106[4] , \nScanOut161[3] , \nOut7_24[3] , 
        \nScanOut687[2] , \nScanOut934[0] , \nScanOut800[3] , \nOut29_15[1] , 
        \nScanOut201[6] , \nScanOut335[5] , \nOut12_30[7] , \nOut13_11[1] , 
        \nScanOut401[2] , \nScanOut535[1] , \nOut20_25[0] , \nOut10_27[4] , 
        \nOut15_18[0] , \nScanOut655[4] , \nScanOut761[7] , \nScanOut580[0] , 
        \nOut19_17[5] , \nOut23_13[5] , \nScanOut1017[2] , \nScanOut380[4] , 
        \nScanOut867[4] , \nOut30_14[6] , \nScanOut953[7] , \nOut4_12[6] , 
        \nScanOut352[2] , \nScanOut466[5] , \nScanOut552[6] , \nScanOut266[1] , 
        \nScanOut465[6] , \nScanOut632[3] , \nScanOut706[0] , \nScanOut981[1] , 
        \nScanOut551[5] , \nOut4_11[5] , \nOut5_30[3] , \nScanOut351[1] , 
        \nScanOut631[0] , \nScanOut705[3] , \nScanOut982[2] , \nScanOut265[2] , 
        \nOut10_24[7] , \nScanOut1014[1] , \nScanOut383[7] , \nScanOut583[3] , 
        \nOut19_14[6] , \nOut23_10[6] , \nOut22_31[0] , \nScanOut864[7] , 
        \nScanOut950[4] , \nOut30_17[5] , \nOut2_0[0] , \nScanOut78[2] , 
        \nOut3_22[3] , \nOut11_3[6] , \nOut17_3[2] , \nOut4_3[7] , 
        \nScanOut818[1] , \nOut29_7[7] , \nScanOut179[1] , \nOut12_28[5] , 
        \nOut24_23[0] , \nScanOut219[4] , \nOut8_2[6] , \nScanOut419[0] , 
        \nOut25_6[6] , \nOut17_17[1] , \nOut8_1[5] , \nOut17_14[2] , 
        \nOut23_6[2] , \nScanOut779[5] , \nOut11_0[5] , \nOut23_5[1] , 
        \nOut24_20[3] , \nOut25_5[5] , \nOut3_21[0] , \nOut4_0[4] , 
        \nOut29_4[4] , \nOut17_0[1] , \nScanOut549[7] , \nOut20_2[3] , 
        \nOut26_2[7] , \nOut1_4[1] , \nOut1_7[2] , \nOut5_28[1] , 
        \nOut9_27[4] , \nOut18_6[2] , \nScanOut629[2] , \nScanOut349[3] , 
        \nOut7_7[6] , \nOut12_7[7] , \nOut14_7[3] , \nOut14_22[7] , 
        \nOut22_29[2] , \nOut27_16[6] , \nScanOut948[6] , \nOut7_4[5] , 
        \nOut14_4[0] , \nOut14_21[4] , \nScanOut598[2] , \nOut27_15[5] , 
        \nScanOut398[6] , \nOut12_4[4] , \nOut0_14[6] , \nOut9_24[7] , 
        \nOut18_5[1] , \nOut20_1[0] , \nOut26_1[4] , \nScanOut999[3] , 
        \nOut1_23[4] , \nScanOut108[2] , \nOut31_2[1] , \nOut8_13[5] , 
        \nScanOut468[3] , \nScanOut268[7] , \nScanOut708[6] , \nOut10_29[2] , 
        \nOut15_16[6] , \nOut19_19[3] , \nOut26_22[7] , \nScanOut1019[4] , 
        \nOut15_15[5] , \nOut26_21[4] , \nScanOut869[2] , \nOut30_19[3] , 
        \nOut31_1[2] , \nOut2_16[2] , \nOut1_20[7] , \nOut7_29[6] , 
        \nOut8_10[6] , \nOut9_31[0] , \nScanOut939[5] , \nScanOut338[0] , 
        \nOut16_23[0] , \nScanOut538[4] , \nOut20_28[5] , \nScanOut658[1] , 
        \nOut25_17[1] , \nOut29_18[4] , \nOut16_20[3] , \nOut25_14[2] , 
        \nScanOut0[3] , \nOut0_1[3] , \nScanOut4[3] , \nScanOut11[3] , 
        \nScanOut12[0] , \nOut2_15[1] , \nOut7_9[0] , \nScanOut595[7] , 
        \nScanOut689[4] , \nScanOut1002[5] , \nOut11_13[5] , \nOut12_9[1] , 
        \nOut14_9[5] , \nOut18_23[4] , \nOut27_18[0] , \nOut22_27[4] , 
        \nScanOut946[0] , \nOut0_19[3] , \nOut1_9[4] , \nScanOut395[3] , 
        \nScanOut872[3] , \nOut31_20[7] , \nScanOut113[3] , \nScanOut473[2] , 
        \nScanOut547[1] , \nScanOut627[4] , \nScanOut713[7] , \nScanOut994[6] , 
        \nScanOut110[0] , \nOut5_26[7] , \nScanOut347[5] , \nScanOut273[6] , 
        \nOut9_29[2] , \nOut18_8[4] , \nOut5_25[4] , \nScanOut344[6] , 
        \nScanOut470[1] , \nScanOut544[2] , \nScanOut270[5] , \nOut11_10[6] , 
        \nOut10_31[0] , \nOut18_20[7] , \nScanOut624[7] , \nScanOut710[4] , 
        \nScanOut997[5] , \nOut22_24[7] , \nScanOut596[4] , \nScanOut1001[6] , 
        \nScanOut396[0] , \nOut31_23[4] , \nScanOut51[1] , \nScanOut75[7] , 
        \nScanOut76[4] , \nScanOut177[7] , \nScanOut871[0] , \nScanOut945[3] , 
        \nScanOut217[2] , \nScanOut323[1] , \nOut12_26[3] , \nOut28_22[3] , 
        \nScanOut417[6] , \nOut21_12[2] , \nScanOut523[5] , \nOut17_19[7] , 
        \nOut25_8[0] , \nOut23_8[4] , \nScanOut643[0] , \nScanOut777[3] , 
        \nOut6_10[2] , \nOut6_13[1] , \nScanOut922[4] , \nOut7_31[4] , 
        \nScanOut691[6] , \nOut29_9[1] , \nScanOut816[7] , \nScanOut921[7] , 
        \nScanOut174[4] , \nOut12_25[0] , \nScanOut414[5] , \nOut21_11[1] , 
        \nScanOut692[5] , \nScanOut815[4] , \nScanOut520[6] , \nOut20_30[7] , 
        \nScanOut214[1] , \nScanOut320[2] , \nScanOut640[3] , \nScanOut774[0] , 
        \nOut28_21[0] , \nScanOut83[7] , \nScanOut182[4] , \nOut7_15[2] , 
        \nScanOut782[0] , \nScanOut905[1] , \nScanOut831[2] , \nScanOut230[7] , 
        \nScanOut304[4] , \nScanOut664[5] , \nScanOut750[6] , \nOut29_24[0] , 
        \nScanOut7[0] , \nScanOut80[4] , \nScanOut150[2] , \nOut13_20[0] , 
        \nScanOut430[3] , \nOut20_14[1] , \nScanOut504[0] , \nScanOut233[4] , 
        \nScanOut307[7] , \nScanOut667[6] , \nScanOut753[5] , \nOut13_23[3] , 
        \nScanOut433[0] , \nOut20_17[2] , \nScanOut507[3] , \nOut25_28[6] , 
        \nScanOut35[5] , \nScanOut52[2] , \nScanOut153[1] , \nOut29_27[3] , 
        \nOut7_16[1] , \nScanOut906[2] , \nOut2_29[5] , \nScanOut781[3] , 
        \nScanOut832[1] , \nOut4_20[4] , \nScanOut181[7] , \nScanOut600[1] , 
        \nScanOut734[2] , \nScanOut887[0] , \nScanOut134[6] , \nScanOut254[3] , 
        \nScanOut360[0] , \nScanOut454[7] , \nScanOut560[4] , \nScanOut961[5] , 
        \nScanOut36[6] , \nScanOut285[6] , \nScanOut286[5] , \nScanOut855[6] , 
        \nOut30_26[4] , \nOut10_15[6] , \nScanOut486[1] , \nOut19_25[7] , 
        \nOut23_21[7] , \nOut30_25[7] , \nScanOut49[3] , \nOut3_5[2] , 
        \nOut3_10[1] , \nScanOut98[6] , \nOut4_23[7] , \nOut10_16[5] , 
        \nOut15_29[1] , \nOut23_22[4] , \nScanOut856[5] , \nScanOut962[6] , 
        \nScanOut485[2] , \nOut19_26[4] , \nScanOut137[5] , \nScanOut257[0] , 
        \nScanOut363[3] , \nScanOut603[2] , \nScanOut737[1] , \nScanOut884[3] , 
        \nScanOut457[4] , \nOut30_9[5] , \nScanOut563[7] , \nOut5_5[6] , 
        \nOut9_4[7] , \nOut17_25[3] , \nOut22_0[3] , \nOut24_11[2] , 
        \nOut24_0[7] , \nOut25_30[4] , \nOut28_1[6] , \nOut16_5[3] , 
        \nScanOut799[1] , \nOut2_31[7] , \nOut10_5[7] , \nOut3_13[2] , 
        \nScanOut199[5] , \nOut16_6[0] , \nOut28_2[5] , \nOut3_6[1] , 
        \nOut5_6[5] , \nScanOut829[0] , \nScanOut148[0] , \nScanOut228[5] , 
        \nOut10_6[4] , \nOut22_3[0] , \nOut12_19[4] , \nScanOut748[4] , 
        \nOut24_12[1] , \nOut9_7[4] , \nScanOut428[1] , \nOut17_26[0] , 
        \nOut24_3[4] , \nOut0_2[0] , \nOut0_25[7] , \nOut6_1[7] , 
        \nOut13_1[6] , \nOut14_10[5] , \nOut15_1[2] , \nOut15_31[3] , 
        \nOut9_15[6] , \nOut27_24[4] , \nOut19_0[3] , \nOut0_26[4] , 
        \nOut21_4[2] , \nOut27_4[6] , \nOut27_7[5] , \nOut5_19[0] , 
        \nOut9_16[5] , \nScanOut618[3] , \nScanOut378[2] , \nOut13_2[5] , 
        \nScanOut578[6] , \nOut19_3[0] , \nOut21_7[1] , \nScanOut979[7] , 
        \nScanOut3[0] , \nOut0_5[3] , \nOut0_6[0] , \nOut0_22[4] , 
        \nOut3_1[2] , \nOut3_2[1] , \nOut3_17[2] , \nOut5_2[5] , \nOut6_2[4] , 
        \nOut6_28[6] , \nOut14_13[6] , \nOut27_27[7] , \nOut15_2[1] , 
        \nOut22_18[3] , \nScanOut919[3] , \nOut16_2[0] , \nOut28_6[5] , 
        \nOut10_2[4] , \nOut3_14[1] , \nOut9_3[4] , \nScanOut318[6] , 
        \nScanOut678[7] , \nOut17_22[0] , \nOut22_7[0] , \nOut21_29[5] , 
        \nOut24_7[4] , \nOut9_0[7] , \nScanOut518[2] , \nOut17_21[3] , 
        \nOut22_4[3] , \nOut24_16[1] , \nOut28_19[4] , \nOut24_15[2] , 
        \nOut24_4[7] , \nOut16_1[3] , \nOut5_1[6] , \nOut28_5[6] , 
        \nScanOut248[1] , \nOut9_12[5] , \nOut10_1[7] , \nOut19_7[0] , 
        \nScanOut728[0] , \nOut27_3[5] , \nScanOut128[4] , \nOut21_3[1] , 
        \nScanOut448[5] , \nScanOut29[7] , \nOut6_6[4] , \nOut13_6[5] , 
        \nOut14_17[6] , \nScanOut849[4] , \nOut15_6[1] , \nOut18_18[3] , 
        \nScanOut299[4] , \nOut11_28[2] , \nOut27_23[7] , \nOut13_5[6] , 
        \nOut31_18[3] , \nOut0_21[7] , \nOut6_5[7] , \nScanOut499[0] , 
        \nOut14_14[5] , \nOut15_5[2] , \nOut27_20[4] , \nScanOut898[1] , 
        \nScanOut84[4] , \nScanOut237[4] , \nOut8_30[0] , \nOut9_11[6] , 
        \nOut27_0[6] , \nScanOut303[7] , \nOut19_4[3] , \nOut21_0[2] , 
        \nScanOut157[1] , \nOut13_27[3] , \nScanOut663[6] , \nScanOut757[5] , 
        \nScanOut55[1] , \nScanOut56[2] , \nOut7_12[1] , \nScanOut437[0] , 
        \nOut16_18[7] , \nOut20_13[2] , \nOut29_23[3] , \nScanOut503[3] , 
        \nScanOut902[2] , \nScanOut185[7] , \nScanOut785[3] , \nScanOut836[1] , 
        \nScanOut87[7] , \nScanOut186[4] , \nOut6_30[4] , \nScanOut786[0] , 
        \nOut7_11[2] , \nScanOut901[1] , \nScanOut835[2] , \nScanOut154[2] , 
        \nScanOut234[7] , \nScanOut300[4] , \nScanOut660[5] , \nScanOut754[6] , 
        \nScanOut434[3] , \nOut20_10[1] , \nScanOut500[0] , \nOut21_31[7] , 
        \nOut29_20[0] , \nScanOut15[3] , \nScanOut31[5] , \nScanOut32[6] , 
        \nOut13_24[0] , \nOut1_18[3] , \nScanOut281[6] , \nScanOut852[5] , 
        \nScanOut966[6] , \nOut30_21[7] , \nOut10_12[5] , \nScanOut481[2] , 
        \nScanOut1022[3] , \nOut19_22[4] , \nOut23_26[4] , \nOut26_19[0] , 
        \nScanOut733[1] , \nScanOut880[3] , \nOut4_24[4] , \nOut4_27[7] , 
        \nOut8_28[2] , \nScanOut607[2] , \nScanOut133[5] , \nScanOut253[0] , 
        \nScanOut367[3] , \nScanOut453[4] , \nScanOut567[7] , \nScanOut130[6] , 
        \nScanOut250[3] , \nScanOut364[0] , \nScanOut604[1] , \nScanOut730[2] , 
        \nScanOut883[0] , \nScanOut282[5] , \nScanOut450[7] , \nScanOut564[4] , 
        \nOut30_22[4] , \nScanOut965[5] , \nScanOut114[0] , \nOut10_11[6] , 
        \nOut11_30[0] , \nScanOut482[1] , \nOut19_21[7] , \nScanOut851[6] , 
        \nOut23_25[7] , \nScanOut1021[0] , \nScanOut474[1] , \nScanOut540[2] , 
        \nOut5_21[4] , \nScanOut620[7] , \nScanOut714[4] , \nScanOut993[5] , 
        \nScanOut274[5] , \nScanOut340[6] , \nOut11_14[6] , \nScanOut592[4] , 
        \nScanOut1005[6] , \nOut18_24[7] , \nOut22_20[7] , \nScanOut16[0] , 
        \nOut11_17[5] , \nScanOut392[0] , \nScanOut875[0] , \nScanOut941[3] , 
        \nOut14_28[1] , \nOut18_27[4] , \nOut31_27[4] , \nOut22_23[4] , 
        \nScanOut591[7] , \nScanOut1006[5] , \nScanOut391[3] , \nOut31_24[7] , 
        \nScanOut942[0] , \nOut2_9[5] , \nScanOut71[7] , \nScanOut117[3] , 
        \nOut20_8[5] , \nScanOut876[3] , \nOut5_22[7] , \nScanOut477[2] , 
        \nScanOut543[1] , \nOut6_14[2] , \nScanOut277[6] , \nScanOut343[5] , 
        \nScanOut623[4] , \nScanOut717[7] , \nOut26_8[1] , \nScanOut990[6] , 
        \nScanOut925[7] , \nScanOut170[4] , \nOut12_21[0] , \nScanOut696[5] , 
        \nScanOut811[4] , \nScanOut173[7] , \nScanOut210[1] , \nScanOut324[2] , 
        \nScanOut410[5] , \nOut28_25[0] , \nScanOut524[6] , \nOut21_15[1] , 
        \nOut8_8[0] , \nScanOut413[6] , \nScanOut644[3] , \nScanOut770[0] , 
        \nOut21_16[2] , \nScanOut527[5] , \nScanOut213[2] , \nScanOut327[1] , 
        \nOut12_22[3] , \nOut28_26[3] , \nScanOut647[0] , \nOut24_29[6] , 
        \nScanOut773[3] , \nOut11_9[0] , \nOut1_24[7] , \nScanOut72[4] , 
        \nOut3_28[5] , \nOut4_9[1] , \nOut6_17[1] , \nScanOut926[4] , 
        \nScanOut695[6] , \nScanOut812[7] , \nOut8_14[6] , \nScanOut389[1] , 
        \nOut14_30[3] , \nOut15_11[5] , \nOut17_9[4] , \nScanOut589[5] , 
        \nOut26_25[4] , \nOut31_5[2] , \nScanOut988[4] , \nOut1_27[4] , 
        \nScanOut558[0] , \nScanOut638[5] , \nOut31_6[1] , \nOut4_18[0] , 
        \nScanOut358[4] , \nOut8_17[5] , \nOut15_12[6] , \nOut26_26[7] , 
        \nOut16_24[3] , \nOut23_19[3] , \nScanOut959[1] , \nOut25_10[2] , 
        \nOut24_31[4] , \nOut0_10[6] , \nOut1_0[1] , \nOut2_4[0] , 
        \nOut2_11[1] , \nOut2_12[2] , \nOut3_30[7] , \nScanOut69[5] , 
        \nScanOut168[6] , \nScanOut809[6] , \nScanOut208[3] , \nOut13_18[4] , 
        \nOut25_13[1] , \nScanOut408[7] , \nOut16_27[0] , \nOut8_5[5] , 
        \nOut17_10[2] , \nOut24_24[3] , \nScanOut768[2] , \nOut16_31[4] , 
        \nOut25_1[5] , \nOut23_1[1] , \nOut2_7[3] , \nOut3_25[0] , 
        \nOut11_4[5] , \nOut17_4[1] , \nOut4_4[4] , \nOut11_7[6] , 
        \nScanOut698[3] , \nOut29_0[4] , \nOut3_26[3] , \nOut4_7[7] , 
        \nOut6_19[7] , \nScanOut928[2] , \nOut29_3[7] , \nOut7_0[5] , 
        \nOut8_6[6] , \nOut17_7[2] , \nOut25_2[6] , \nScanOut329[7] , 
        \nOut17_13[1] , \nOut21_18[4] , \nScanOut529[3] , \nScanOut649[6] , 
        \nOut24_27[0] , \nOut28_28[5] , \nOut23_2[2] , \nOut26_30[3] , 
        \nOut27_11[5] , \nOut12_0[4] , \nOut14_25[4] , \nOut14_0[0] , 
        \nOut31_29[2] , \nOut20_5[0] , \nOut26_5[4] , \nOut0_13[5] , 
        \nOut1_31[0] , \nScanOut119[5] , \nOut9_20[7] , \nOut18_1[1] , 
        \nScanOut279[0] , \nOut9_23[4] , \nScanOut479[4] , \nOut20_6[3] , 
        \nOut18_2[2] , \nScanOut719[1] , \nOut26_6[7] , \nScanOut18[6] , 
        \nOut1_3[2] , \nOut7_3[6] , \nOut11_19[3] , \nOut14_3[3] , 
        \nOut14_26[7] , \nOut18_29[2] , \nScanOut1008[3] , \nOut27_12[6] , 
        \nOut12_3[7] , \nScanOut64[0] , \nScanOut878[5] , \nScanOut67[3] , 
        \nScanOut165[3] , \nOut7_20[3] , \nScanOut405[2] , \nScanOut683[2] , 
        \nScanOut930[0] , \nScanOut804[3] , \nScanOut531[1] , \nOut20_21[0] , 
        \nScanOut166[0] , \nScanOut205[6] , \nScanOut331[5] , \nOut13_15[1] , 
        \nOut28_30[7] , \nOut29_11[1] , \nScanOut651[4] , \nScanOut765[7] , 
        \nOut13_16[2] , \nScanOut206[5] , \nScanOut332[6] , \nScanOut406[1] , 
        \nOut29_12[2] , \nOut16_29[6] , \nScanOut532[2] , \nOut20_22[3] , 
        \nOut7_23[0] , \nScanOut652[7] , \nScanOut766[4] , \nScanOut933[3] , 
        \nScanOut101[7] , \nScanOut680[1] , \nScanOut807[0] , \nOut4_15[5] , 
        \nScanOut355[1] , \nScanOut461[6] , \nScanOut555[5] , \nScanOut261[2] , 
        \nOut10_20[7] , \nOut19_10[6] , \nOut18_31[0] , \nScanOut635[0] , 
        \nScanOut701[3] , \nScanOut986[2] , \nOut23_14[6] , \nScanOut1010[1] , 
        \nOut0_8[6] , \nOut1_29[2] , \nScanOut102[4] , \nOut10_23[4] , 
        \nScanOut387[7] , \nScanOut587[3] , \nOut30_13[5] , \nScanOut584[0] , 
        \nOut26_28[1] , \nScanOut860[7] , \nScanOut954[4] , \nScanOut1013[2] , 
        \nScanOut384[4] , \nOut19_13[5] , \nOut23_17[5] , \nScanOut863[4] , 
        \nScanOut957[7] , \nScanOut462[5] , \nOut30_10[6] , \nScanOut556[6] , 
        \nOut31_8[7] , \nScanOut702[0] , \nScanOut985[1] , \nOut4_16[6] , 
        \nOut8_19[3] , \nScanOut636[3] , \nScanOut356[2] , \nScanOut262[1] , 
        \nScanOut294[1] , \nOut31_15[6] , \nScanOut27[1] , \nScanOut973[1] , 
        \nOut6_8[2] , \nOut13_8[3] , \nScanOut847[2] , \nOut14_19[0] , 
        \nOut15_8[7] , \nOut18_16[5] , \nScanOut494[5] , \nOut22_12[5] , 
        \nOut11_26[4] , \nScanOut24[2] , \nScanOut125[1] , \nScanOut126[2] , 
        \nOut5_13[6] , \nScanOut246[7] , \nScanOut372[4] , \nOut19_9[6] , 
        \nScanOut612[5] , \nScanOut726[6] , \nScanOut895[4] , \nOut5_10[5] , 
        \nOut4_31[3] , \nScanOut446[3] , \nScanOut572[0] , \nScanOut611[6] , 
        \nScanOut725[5] , \nScanOut896[7] , \nScanOut245[4] , \nScanOut371[7] , 
        \nScanOut445[0] , \nScanOut571[3] , \nScanOut43[5] , \nScanOut91[3] , 
        \nScanOut297[2] , \nScanOut844[1] , \nScanOut970[2] , \nOut31_16[5] , 
        \nOut11_25[7] , \nScanOut497[6] , \nOut18_15[6] , \nOut22_11[6] , 
        \nOut23_30[0] , \nScanOut142[6] , \nScanOut222[3] , \nScanOut316[0] , 
        \nScanOut676[1] , \nScanOut742[2] , \nOut22_9[6] , \nScanOut422[7] , 
        \nScanOut516[4] , \nOut21_27[3] , \nOut24_9[2] , \nOut28_17[2] , 
        \nOut12_13[2] , \nOut24_18[7] , \nOut28_8[3] , \nOut6_26[0] , 
        \nScanOut790[4] , \nScanOut823[6] , \nScanOut917[5] , \nOut0_15[2] , 
        \nOut0_16[1] , \nOut1_6[6] , \nScanOut40[6] , \nOut3_19[4] , 
        \nOut6_25[3] , \nScanOut190[0] , \nScanOut914[6] , \nOut1_15[6] , 
        \nOut1_16[5] , \nScanOut92[0] , \nScanOut193[3] , \nScanOut793[7] , 
        \nScanOut820[5] , \nScanOut221[0] , \nScanOut315[3] , \nScanOut141[5] , 
        \nOut12_10[1] , \nOut13_31[7] , \nScanOut675[2] , \nScanOut741[1] , 
        \nOut28_14[1] , \nScanOut421[4] , \nScanOut515[7] , \nOut21_24[0] , 
        \nScanOut609[4] , \nOut4_29[1] , \nOut8_25[7] , \nOut8_26[4] , 
        \nScanOut369[5] , \nOut15_20[4] , \nOut15_23[7] , \nScanOut569[1] , 
        \nOut23_28[2] , \nOut26_17[6] , \nOut30_3[3] , \nScanOut968[0] , 
        \nOut26_14[5] , \nOut2_20[0] , \nOut2_23[3] , \nOut30_0[0] , 
        \nScanOut58[4] , \nScanOut89[1] , \nScanOut159[7] , \nScanOut239[2] , 
        \nScanOut838[7] , \nScanOut759[3] , \nOut13_29[5] , \nScanOut439[6] , 
        \nOut16_16[1] , \nOut25_22[0] , \nOut16_15[2] , \nScanOut788[6] , 
        \nOut25_21[3] , \nScanOut188[2] , \nOut5_29[5] , \nOut7_6[2] , 
        \nOut12_6[3] , \nScanOut949[2] , \nOut14_6[7] , \nOut14_23[3] , 
        \nOut22_28[6] , \nOut27_17[2] , \nOut9_26[0] , \nScanOut348[7] , 
        \nOut18_7[6] , \nScanOut628[6] , \nOut26_3[3] , \nScanOut548[3] , 
        \nOut20_3[7] , \nOut26_0[0] , \nScanOut998[7] , \nScanOut21[6] , 
        \nOut2_1[4] , \nOut2_2[7] , \nOut1_5[5] , \nOut9_25[3] , \nOut18_4[5] , 
        \nOut12_5[0] , \nOut20_0[4] , \nScanOut399[2] , \nScanOut79[6] , 
        \nScanOut178[5] , \nOut7_5[1] , \nScanOut599[6] , \nScanOut218[0] , 
        \nOut14_5[4] , \nOut14_20[0] , \nOut27_14[1] , \nOut23_7[6] , 
        \nScanOut778[1] , \nOut8_3[2] , \nScanOut418[4] , \nOut17_16[5] , 
        \nOut25_7[2] , \nOut12_29[1] , \nOut24_22[4] , \nOut3_23[7] , 
        \nOut4_2[3] , \nOut17_2[6] , \nScanOut819[5] , \nOut29_6[3] , 
        \nOut11_2[2] , \nOut3_20[4] , \nOut4_1[0] , \nOut17_1[5] , 
        \nOut29_5[0] , \nScanOut45[2] , \nOut2_19[0] , \nScanOut104[3] , 
        \nOut4_10[1] , \nScanOut107[0] , \nOut4_13[2] , \nOut8_0[1] , 
        \nOut11_1[1] , \nOut23_4[5] , \nOut24_21[7] , \nOut25_4[1] , 
        \nScanOut353[6] , \nOut17_15[6] , \nScanOut633[7] , \nScanOut707[4] , 
        \nScanOut980[5] , \nScanOut267[5] , \nScanOut467[1] , \nScanOut553[2] , 
        \nOut5_31[7] , \nOut10_25[3] , \nOut10_26[0] , \nScanOut381[0] , 
        \nScanOut866[0] , \nScanOut952[3] , \nOut30_15[2] , \nScanOut1016[6] , 
        \nScanOut382[3] , \nOut15_19[4] , \nScanOut581[4] , \nOut19_16[1] , 
        \nOut23_12[1] , \nScanOut582[7] , \nOut19_15[2] , \nOut22_30[4] , 
        \nOut23_11[2] , \nScanOut865[3] , \nOut30_16[1] , \nScanOut951[0] , 
        \nScanOut1015[5] , \nScanOut350[5] , \nScanOut264[6] , 
        \nScanOut630[4] , \nScanOut704[7] , \nScanOut983[6] , \nScanOut464[2] , 
        \nScanOut550[1] , \nScanOut61[4] , \nScanOut62[7] , \nScanOut160[7] , 
        \nScanOut163[4] , \nScanOut203[1] , \nOut7_26[4] , \nScanOut337[2] , 
        \nScanOut685[5] , \nScanOut936[7] , \nScanOut802[4] , \nScanOut657[3] , 
        \nScanOut763[0] , \nScanOut200[2] , \nScanOut334[1] , \nOut13_13[6] , 
        \nOut29_17[6] , \nScanOut403[5] , \nOut25_18[3] , \nScanOut537[6] , 
        \nOut20_27[7] , \nScanOut654[0] , \nScanOut760[3] , \nOut13_10[5] , 
        \nScanOut400[6] , \nOut12_31[3] , \nScanOut534[5] , \nOut20_24[4] , 
        \nOut7_25[7] , \nOut29_14[5] , \nScanOut935[4] , \nScanOut97[4] , 
        \nScanOut144[1] , \nScanOut686[6] , \nScanOut801[7] , \nOut28_11[5] , 
        \nScanOut224[4] , \nScanOut310[7] , \nOut12_15[5] , \nOut29_30[3] , 
        \nScanOut424[0] , \nScanOut510[3] , \nOut21_21[4] , \nScanOut196[7] , 
        \nScanOut670[6] , \nScanOut744[5] , \nScanOut46[1] , \nOut3_9[3] , 
        \nOut6_20[7] , \nScanOut796[3] , \nOut10_9[6] , \nScanOut825[1] , 
        \nScanOut911[2] , \nOut5_9[7] , \nOut6_23[4] , \nScanOut195[4] , 
        \nScanOut912[1] , \nScanOut94[7] , \nScanOut147[2] , \nOut9_8[6] , 
        \nScanOut427[3] , \nOut16_9[2] , \nScanOut795[0] , \nScanOut826[2] , 
        \nOut17_29[2] , \nOut21_22[7] , \nOut12_16[6] , \nScanOut513[0] , 
        \nOut28_12[6] , \nScanOut227[7] , \nScanOut313[4] , \nScanOut673[5] , 
        \nScanOut747[6] , \nOut11_20[3] , \nScanOut492[2] , \nOut18_10[2] , 
        \nOut19_31[4] , \nOut22_14[2] , \nScanOut975[6] , \nScanOut22[5] , 
        \nOut0_29[6] , \nScanOut120[5] , \nScanOut292[6] , \nScanOut841[5] , 
        \nOut31_13[1] , \nScanOut440[4] , \nScanOut574[7] , \nScanOut123[6] , 
        \nOut5_15[1] , \nScanOut614[2] , \nScanOut720[1] , \nScanOut893[3] , 
        \nScanOut240[0] , \nScanOut374[3] , \nOut21_8[3] , \nOut5_16[2] , 
        \nOut9_19[7] , \nScanOut443[7] , \nScanOut577[4] , \nScanOut243[3] , 
        \nScanOut377[0] , \nScanOut723[2] , \nScanOut890[0] , \nScanOut291[5] , 
        \nOut11_23[0] , \nScanOut491[1] , \nOut18_13[1] , \nScanOut617[1] , 
        \nOut27_8[7] , \nOut22_17[1] , \nOut27_28[5] , \nOut31_10[2] , 
        \nOut30_31[4] , \nOut2_25[4] , \nScanOut842[6] , \nScanOut976[5] , 
        \nOut16_10[6] , \nOut17_31[0] , \nOut25_24[7] , \nScanOut8[2] , 
        \nOut25_27[4] , \nOut29_28[1] , \nOut1_10[2] , \nOut2_26[7] , 
        \nScanOut308[5] , \nOut16_13[5] , \nScanOut508[1] , \nOut20_18[0] , 
        \nScanOut668[4] , \nOut7_19[3] , \nScanOut909[0] , \nOut8_20[3] , 
        \nOut30_5[4] , \nScanOut888[2] , \nScanOut289[7] , \nOut15_25[0] , 
        \nScanOut489[3] , \nOut26_11[1] , \nOut27_30[7] , \nOut30_29[6] , 
        \nOut10_19[7] , \nOut26_12[2] , \nOut0_24[3] , \nScanOut39[4] , 
        \nOut15_26[3] , \nOut19_29[6] , \nOut1_13[1] , \nScanOut138[7] , 
        \nScanOut458[6] , \nScanOut859[7] , \nScanOut738[3] , \nOut30_6[7] , 
        \nOut8_23[0] , \nScanOut258[2] , \nOut21_5[6] , \nOut27_5[2] , 
        \nOut6_0[3] , \nOut9_14[2] , \nOut19_1[7] , \nOut13_0[2] , 
        \nOut14_11[1] , \nOut27_25[0] , \nOut15_30[7] , \nOut15_0[6] , 
        \nOut0_3[4] , \nOut6_3[0] , \nOut14_12[2] , \nOut15_3[5] , 
        \nOut22_19[7] , \nOut27_26[3] , \nScanOut5[7] , \nOut0_27[0] , 
        \nOut5_18[4] , \nOut13_3[1] , \nScanOut978[3] , \nScanOut579[2] , 
        \nOut21_6[5] , \nOut9_17[1] , \nScanOut379[6] , \nOut19_2[4] , 
        \nScanOut619[7] , \nScanOut34[1] , \nScanOut48[7] , \nOut2_30[3] , 
        \nOut3_4[6] , \nOut27_6[1] , \nOut3_11[5] , \nScanOut198[1] , 
        \nOut10_4[3] , \nOut16_4[7] , \nOut3_7[5] , \nScanOut99[2] , 
        \nOut5_4[2] , \nOut9_5[3] , \nOut17_24[7] , \nOut24_10[6] , 
        \nScanOut798[5] , \nOut28_0[2] , \nOut25_31[0] , \nOut24_1[3] , 
        \nOut22_1[7] , \nScanOut149[4] , \nOut9_6[0] , \nScanOut429[5] , 
        \nOut17_27[4] , \nOut24_2[0] , \nScanOut229[1] , \nOut12_18[0] , 
        \nOut22_2[4] , \nScanOut749[0] , \nOut24_13[5] , \nOut10_7[0] , 
        \nOut5_7[1] , \nOut3_12[6] , \nOut16_7[4] , \nScanOut828[4] , 
        \nOut28_3[1] , \nScanOut287[1] , \nOut10_14[2] , \nScanOut487[5] , 
        \nOut19_24[3] , \nOut23_20[3] , \nScanOut1024[4] , \nOut30_27[0] , 
        \nScanOut37[2] , \nOut4_21[0] , \nScanOut135[2] , \nScanOut854[2] , 
        \nScanOut960[1] , \nScanOut455[3] , \nScanOut561[0] , \nOut4_22[3] , 
        \nScanOut136[1] , \nScanOut255[7] , \nScanOut361[4] , \nScanOut456[0] , 
        \nScanOut601[5] , \nScanOut735[6] , \nScanOut886[4] , \nScanOut562[3] , 
        \nOut30_8[1] , \nScanOut602[6] , \nScanOut736[5] , \nScanOut885[7] , 
        \nScanOut256[4] , \nScanOut362[7] , \nOut10_17[1] , \nScanOut484[6] , 
        \nOut15_28[5] , \nOut19_27[0] , \nOut23_23[0] , \nScanOut963[2] , 
        \nScanOut151[6] , \nScanOut284[2] , \nScanOut857[1] , \nOut30_24[3] , 
        \nOut13_21[4] , \nScanOut431[7] , \nOut20_15[5] , \nScanOut505[4] , 
        \nScanOut6[4] , \nScanOut50[5] , \nScanOut82[3] , \nOut29_25[4] , 
        \nScanOut183[0] , \nScanOut231[3] , \nScanOut305[0] , \nScanOut665[1] , 
        \nScanOut751[2] , \nOut7_14[6] , \nScanOut904[5] , \nScanOut53[6] , 
        \nOut2_28[1] , \nScanOut180[3] , \nScanOut783[4] , \nScanOut830[6] , 
        \nScanOut152[5] , \nOut7_17[5] , \nScanOut780[7] , \nScanOut907[6] , 
        \nScanOut833[5] , \nOut29_26[7] , \nScanOut10[7] , \nScanOut13[4] , 
        \nOut0_18[7] , \nScanOut74[3] , \nScanOut77[0] , \nScanOut81[0] , 
        \nScanOut232[0] , \nScanOut306[3] , \nOut13_22[7] , \nOut25_29[2] , 
        \nScanOut432[4] , \nOut20_16[6] , \nScanOut506[7] , \nOut6_12[5] , 
        \nScanOut666[2] , \nScanOut752[1] , \nScanOut923[0] , \nScanOut175[0] , 
        \nScanOut176[3] , \nScanOut216[6] , \nScanOut322[5] , \nScanOut642[4] , 
        \nScanOut690[2] , \nScanOut817[3] , \nOut29_8[5] , \nScanOut776[7] , 
        \nOut12_27[7] , \nScanOut416[2] , \nOut17_18[3] , \nOut23_9[0] , 
        \nOut25_9[4] , \nScanOut522[1] , \nOut21_13[6] , \nScanOut215[5] , 
        \nScanOut321[6] , \nOut28_23[7] , \nScanOut641[7] , \nScanOut775[4] , 
        \nOut12_24[4] , \nOut28_20[4] , \nScanOut415[1] , \nScanOut521[2] , 
        \nOut21_10[5] , \nOut20_31[3] , \nOut5_27[3] , \nOut6_11[6] , 
        \nOut7_30[0] , \nOut9_28[6] , \nOut18_9[0] , \nScanOut693[1] , 
        \nScanOut920[3] , \nScanOut814[0] , \nScanOut272[2] , \nScanOut346[1] , 
        \nScanOut712[3] , \nScanOut995[2] , \nOut1_8[0] , \nScanOut112[7] , 
        \nScanOut626[0] , \nScanOut394[7] , \nScanOut472[6] , \nScanOut546[5] , 
        \nOut31_21[3] , \nOut7_8[4] , \nOut11_12[1] , \nOut12_8[5] , 
        \nOut14_8[1] , \nOut18_22[0] , \nOut22_26[0] , \nScanOut873[7] , 
        \nScanOut947[4] , \nScanOut594[3] , \nScanOut1003[1] , \nOut27_19[4] , 
        \nScanOut944[7] , \nScanOut24[6] , \nOut1_15[2] , \nOut2_14[5] , 
        \nOut2_17[6] , \nScanOut111[4] , \nOut5_24[0] , \nOut10_30[4] , 
        \nScanOut397[4] , \nScanOut870[4] , \nOut31_22[0] , \nScanOut1000[2] , 
        \nOut11_11[2] , \nScanOut597[0] , \nOut18_21[3] , \nScanOut625[3] , 
        \nOut22_25[3] , \nScanOut711[0] , \nScanOut996[1] , \nScanOut271[1] , 
        \nScanOut345[2] , \nScanOut471[5] , \nScanOut545[6] , \nScanOut339[4] , 
        \nOut16_22[4] , \nOut20_29[1] , \nScanOut659[5] , \nOut25_16[5] , 
        \nOut29_19[0] , \nScanOut539[0] , \nOut7_28[2] , \nScanOut688[0] , 
        \nScanOut938[1] , \nOut1_21[3] , \nOut1_22[0] , \nOut10_28[6] , 
        \nOut16_21[7] , \nOut25_15[6] , \nScanOut868[6] , \nScanOut1018[0] , 
        \nOut15_17[2] , \nOut26_23[3] , \nOut19_18[7] , \nScanOut709[2] , 
        \nScanOut109[6] , \nOut8_12[1] , \nScanOut269[3] , \nScanOut469[7] , 
        \nOut31_3[5] , \nOut8_11[2] , \nOut9_30[4] , \nOut15_14[1] , 
        \nOut30_18[7] , \nOut26_20[0] , \nOut30_0[4] , \nOut1_16[1] , 
        \nOut4_29[5] , \nOut8_25[3] , \nOut15_20[0] , \nOut26_14[1] , 
        \nOut15_23[3] , \nScanOut569[5] , \nOut23_28[6] , \nOut26_17[2] , 
        \nOut30_3[7] , \nScanOut968[4] , \nOut8_26[0] , \nScanOut369[1] , 
        \nScanOut609[0] , \nOut2_20[4] , \nScanOut188[6] , \nOut2_23[7] , 
        \nScanOut58[0] , \nScanOut89[5] , \nOut16_15[6] , \nScanOut788[2] , 
        \nOut25_21[7] , \nScanOut159[3] , \nScanOut439[2] , \nOut16_16[5] , 
        \nScanOut239[6] , \nOut13_29[1] , \nOut25_22[4] , \nScanOut759[7] , 
        \nScanOut838[3] , \nScanOut297[6] , \nOut11_25[3] , \nScanOut497[2] , 
        \nOut18_15[2] , \nOut22_11[2] , \nOut23_30[4] , \nOut31_16[1] , 
        \nScanOut125[5] , \nScanOut844[5] , \nScanOut970[6] , \nScanOut126[6] , 
        \nOut5_10[1] , \nOut4_31[7] , \nScanOut445[4] , \nScanOut571[7] , 
        \nScanOut245[0] , \nScanOut371[3] , \nScanOut446[7] , \nScanOut611[2] , 
        \nScanOut725[1] , \nScanOut896[3] , \nScanOut572[4] , \nOut5_13[2] , 
        \nScanOut612[1] , \nScanOut726[2] , \nScanOut895[0] , \nOut6_8[6] , 
        \nScanOut246[3] , \nScanOut372[0] , \nScanOut494[1] , \nOut19_9[2] , 
        \nOut11_26[0] , \nOut0_8[2] , \nScanOut27[5] , \nOut14_19[4] , 
        \nOut15_8[3] , \nOut18_16[1] , \nOut22_12[1] , \nScanOut973[5] , 
        \nScanOut294[5] , \nOut13_8[7] , \nScanOut847[6] , \nOut31_15[2] , 
        \nScanOut40[2] , \nScanOut92[4] , \nScanOut141[1] , \nOut12_10[5] , 
        \nScanOut421[0] , \nOut13_31[3] , \nScanOut515[3] , \nOut21_24[4] , 
        \nOut28_14[5] , \nOut6_25[7] , \nScanOut193[7] , \nScanOut221[4] , 
        \nScanOut315[7] , \nScanOut675[6] , \nScanOut741[5] , \nScanOut914[2] , 
        \nScanOut190[4] , \nScanOut793[3] , \nScanOut820[1] , \nOut0_10[2] , 
        \nOut0_13[1] , \nScanOut18[2] , \nOut2_4[4] , \nOut2_7[7] , 
        \nScanOut43[1] , \nOut3_19[0] , \nOut1_29[6] , \nScanOut64[4] , 
        \nScanOut67[7] , \nScanOut91[7] , \nScanOut142[2] , \nOut6_26[4] , 
        \nScanOut790[0] , \nOut28_8[7] , \nScanOut823[2] , \nScanOut917[1] , 
        \nOut28_17[6] , \nScanOut222[7] , \nScanOut316[4] , \nOut12_13[6] , 
        \nScanOut422[3] , \nOut24_18[3] , \nScanOut516[0] , \nOut21_27[7] , 
        \nOut22_9[2] , \nOut24_9[6] , \nOut7_23[4] , \nScanOut676[5] , 
        \nScanOut742[6] , \nScanOut933[7] , \nScanOut165[7] , \nScanOut166[4] , 
        \nScanOut206[1] , \nScanOut332[2] , \nScanOut652[3] , \nScanOut680[5] , 
        \nScanOut807[4] , \nScanOut766[0] , \nOut13_16[6] , \nScanOut406[5] , 
        \nOut16_29[2] , \nOut20_22[7] , \nScanOut532[6] , \nScanOut205[2] , 
        \nScanOut331[1] , \nOut29_12[6] , \nScanOut651[0] , \nScanOut765[3] , 
        \nOut13_15[5] , \nOut28_30[3] , \nOut29_11[5] , \nScanOut405[6] , 
        \nScanOut531[5] , \nOut20_21[4] , \nOut4_16[2] , \nOut7_20[7] , 
        \nOut8_19[7] , \nScanOut683[6] , \nScanOut930[4] , \nScanOut804[7] , 
        \nScanOut356[6] , \nScanOut262[5] , \nScanOut702[4] , \nScanOut985[5] , 
        \nOut3_26[7] , \nScanOut101[3] , \nScanOut102[0] , \nScanOut636[7] , 
        \nOut31_8[3] , \nOut4_15[1] , \nOut10_20[3] , \nOut10_23[0] , 
        \nScanOut384[0] , \nScanOut462[1] , \nScanOut556[2] , \nOut19_13[1] , 
        \nOut23_17[1] , \nScanOut863[0] , \nOut30_10[2] , \nScanOut957[3] , 
        \nScanOut1013[6] , \nScanOut387[3] , \nScanOut584[4] , \nOut26_28[5] , 
        \nScanOut860[3] , \nScanOut954[0] , \nOut30_13[1] , \nScanOut587[7] , 
        \nScanOut1010[5] , \nScanOut355[5] , \nOut19_10[2] , \nOut18_31[4] , 
        \nScanOut635[4] , \nScanOut701[7] , \nOut23_14[2] , \nScanOut986[6] , 
        \nScanOut261[6] , \nScanOut461[2] , \nScanOut555[1] , \nOut8_6[2] , 
        \nScanOut329[3] , \nScanOut649[2] , \nOut23_2[6] , \nOut24_27[4] , 
        \nOut25_2[2] , \nOut28_28[1] , \nOut17_7[6] , \nOut17_13[5] , 
        \nScanOut529[7] , \nOut21_18[0] , \nOut4_7[3] , \nOut6_19[3] , 
        \nScanOut928[6] , \nOut29_3[3] , \nOut3_25[4] , \nOut4_4[0] , 
        \nOut11_7[2] , \nScanOut698[7] , \nOut29_0[0] , \nOut11_4[1] , 
        \nOut17_4[5] , \nOut8_5[1] , \nOut17_10[6] , \nOut23_1[5] , 
        \nOut16_31[0] , \nOut25_1[1] , \nOut24_24[7] , \nOut1_3[6] , 
        \nOut12_3[3] , \nScanOut878[1] , \nOut7_3[2] , \nOut11_19[7] , 
        \nOut27_12[2] , \nScanOut1008[7] , \nOut14_3[7] , \nOut14_26[3] , 
        \nOut18_29[6] , \nScanOut719[5] , \nOut26_6[3] , \nScanOut119[1] , 
        \nScanOut279[4] , \nOut9_23[0] , \nOut18_2[6] , \nScanOut479[0] , 
        \nOut9_20[3] , \nOut18_1[5] , \nOut20_6[7] , \nOut26_5[0] , 
        \nOut1_0[5] , \nOut1_31[4] , \nOut20_5[4] , \nOut31_29[6] , 
        \nOut2_12[6] , \nOut1_24[3] , \nOut1_27[0] , \nOut4_18[4] , 
        \nOut7_0[1] , \nOut12_0[0] , \nOut14_25[0] , \nOut14_0[4] , 
        \nOut26_30[7] , \nScanOut358[0] , \nOut15_12[2] , \nOut23_19[7] , 
        \nOut27_11[1] , \nScanOut959[5] , \nOut26_26[3] , \nOut8_17[1] , 
        \nScanOut638[1] , \nScanOut558[4] , \nOut31_6[5] , \nScanOut988[0] , 
        \nScanOut69[1] , \nScanOut168[2] , \nScanOut208[7] , \nOut8_14[2] , 
        \nScanOut389[5] , \nOut31_5[6] , \nOut14_30[7] , \nOut15_11[1] , 
        \nScanOut589[1] , \nOut26_25[0] , \nScanOut768[6] , \nScanOut408[3] , 
        \nOut16_27[4] , \nOut13_18[0] , \nOut25_13[5] , \nScanOut809[2] , 
        \nScanOut0[7] , \nScanOut15[7] , \nScanOut16[4] , \nOut2_11[5] , 
        \nOut3_30[3] , \nScanOut117[7] , \nOut5_22[3] , \nOut16_24[7] , 
        \nOut25_10[6] , \nOut24_31[0] , \nScanOut623[0] , \nScanOut717[3] , 
        \nOut26_8[5] , \nScanOut990[2] , \nScanOut277[2] , \nScanOut343[1] , 
        \nScanOut477[6] , \nScanOut543[5] , \nOut20_8[1] , \nScanOut942[4] , 
        \nOut11_17[1] , \nScanOut391[7] , \nScanOut876[7] , \nOut31_24[3] , 
        \nScanOut591[3] , \nScanOut1006[1] , \nScanOut392[4] , \nOut14_28[5] , 
        \nOut18_27[0] , \nOut22_23[0] , \nOut31_27[0] , \nOut2_9[1] , 
        \nScanOut72[0] , \nOut3_28[1] , \nScanOut114[4] , \nOut5_21[0] , 
        \nOut11_14[2] , \nOut18_24[3] , \nOut22_20[3] , \nScanOut875[4] , 
        \nScanOut941[7] , \nScanOut592[0] , \nScanOut1005[2] , 
        \nScanOut274[1] , \nScanOut340[2] , \nScanOut620[3] , \nScanOut714[0] , 
        \nScanOut993[1] , \nScanOut474[5] , \nOut17_9[0] , \nScanOut540[6] , 
        \nOut4_9[5] , \nOut6_17[5] , \nScanOut926[0] , \nScanOut695[2] , 
        \nScanOut812[3] , \nScanOut71[3] , \nScanOut170[0] , \nScanOut173[3] , 
        \nScanOut213[6] , \nScanOut327[5] , \nOut11_9[4] , \nScanOut647[4] , 
        \nScanOut773[7] , \nScanOut210[5] , \nOut8_8[4] , \nOut12_22[7] , 
        \nOut24_29[2] , \nOut28_26[7] , \nScanOut413[2] , \nOut21_16[6] , 
        \nScanOut324[6] , \nScanOut527[1] , \nScanOut644[7] , \nScanOut770[4] , 
        \nOut12_21[4] , \nScanOut410[1] , \nScanOut524[2] , \nOut21_15[5] , 
        \nOut6_14[6] , \nOut28_25[4] , \nScanOut925[3] , \nScanOut154[6] , 
        \nScanOut696[1] , \nScanOut811[0] , \nScanOut3[4] , \nScanOut55[5] , 
        \nScanOut87[3] , \nScanOut234[3] , \nScanOut300[0] , \nOut13_24[4] , 
        \nOut29_20[4] , \nScanOut434[7] , \nOut20_10[5] , \nScanOut500[4] , 
        \nOut21_31[3] , \nScanOut186[0] , \nScanOut660[1] , \nScanOut754[2] , 
        \nScanOut56[6] , \nScanOut185[3] , \nOut6_30[0] , \nScanOut786[4] , 
        \nOut7_11[6] , \nScanOut901[5] , \nScanOut835[6] , \nOut7_12[5] , 
        \nScanOut902[6] , \nScanOut157[5] , \nOut13_27[7] , \nScanOut437[4] , 
        \nOut16_18[3] , \nScanOut785[7] , \nScanOut836[5] , \nOut20_13[6] , 
        \nScanOut503[7] , \nOut29_23[7] , \nOut0_3[0] , \nScanOut5[3] , 
        \nOut0_5[7] , \nOut0_21[3] , \nScanOut31[1] , \nScanOut84[0] , 
        \nScanOut237[0] , \nScanOut303[3] , \nScanOut663[2] , \nScanOut757[1] , 
        \nOut10_11[2] , \nOut11_30[4] , \nScanOut482[5] , \nScanOut1021[4] , 
        \nOut19_21[3] , \nOut23_25[3] , \nScanOut965[1] , \nScanOut32[2] , 
        \nOut1_18[7] , \nOut4_24[0] , \nScanOut130[2] , \nScanOut282[1] , 
        \nScanOut851[2] , \nOut30_22[0] , \nScanOut450[3] , \nScanOut564[0] , 
        \nScanOut604[5] , \nScanOut730[6] , \nScanOut883[4] , \nOut4_27[3] , 
        \nScanOut133[1] , \nScanOut250[7] , \nScanOut364[4] , \nOut8_28[6] , 
        \nScanOut453[0] , \nScanOut567[3] , \nScanOut253[4] , \nScanOut367[7] , 
        \nScanOut733[5] , \nScanOut880[7] , \nScanOut281[2] , \nOut10_12[1] , 
        \nScanOut481[6] , \nOut19_22[0] , \nScanOut607[6] , \nOut23_26[0] , 
        \nScanOut1022[7] , \nOut26_19[4] , \nOut30_21[3] , \nOut3_1[6] , 
        \nOut10_1[3] , \nScanOut852[1] , \nScanOut966[2] , \nOut3_2[5] , 
        \nOut3_14[5] , \nOut5_1[2] , \nOut16_1[7] , \nOut28_5[2] , 
        \nOut9_3[0] , \nOut9_0[3] , \nOut17_21[7] , \nOut24_4[3] , 
        \nOut17_22[4] , \nOut21_29[1] , \nOut22_4[7] , \nOut24_15[6] , 
        \nOut24_16[5] , \nOut28_19[0] , \nOut24_7[0] , \nScanOut318[2] , 
        \nScanOut518[6] , \nScanOut678[3] , \nOut22_7[4] , \nOut3_17[6] , 
        \nOut10_2[0] , \nOut16_2[4] , \nOut5_2[1] , \nOut6_28[2] , 
        \nScanOut919[7] , \nOut8_30[4] , \nOut9_11[2] , \nOut21_0[6] , 
        \nOut28_6[1] , \nOut19_4[7] , \nOut27_0[2] , \nScanOut898[5] , 
        \nOut6_5[3] , \nOut14_14[1] , \nOut15_5[6] , \nScanOut499[4] , 
        \nScanOut299[0] , \nOut27_20[0] , \nOut31_18[7] , \nScanOut6[0] , 
        \nOut0_6[4] , \nScanOut29[3] , \nOut6_6[0] , \nOut13_5[2] , 
        \nOut11_28[6] , \nOut14_17[2] , \nOut27_23[3] , \nOut15_6[5] , 
        \nOut18_18[7] , \nOut13_6[1] , \nScanOut849[0] , \nScanOut10[3] , 
        \nOut0_22[0] , \nScanOut128[0] , \nScanOut448[1] , \nOut21_3[5] , 
        \nScanOut728[4] , \nOut2_14[1] , \nScanOut248[5] , \nOut9_12[1] , 
        \nOut27_3[1] , \nOut19_7[4] , \nOut16_21[3] , \nOut25_15[2] , 
        \nOut2_17[2] , \nOut7_28[6] , \nScanOut688[4] , \nScanOut938[5] , 
        \nOut1_21[7] , \nScanOut339[0] , \nOut16_22[0] , \nScanOut539[4] , 
        \nOut20_29[5] , \nScanOut659[1] , \nOut25_16[1] , \nOut29_19[4] , 
        \nOut15_14[5] , \nOut26_20[4] , \nOut30_18[3] , \nOut1_22[4] , 
        \nScanOut109[2] , \nOut8_11[6] , \nOut9_30[0] , \nOut31_3[1] , 
        \nOut8_12[5] , \nScanOut469[3] , \nScanOut269[7] , \nScanOut709[6] , 
        \nScanOut74[7] , \nOut10_28[2] , \nOut15_17[6] , \nOut19_18[3] , 
        \nOut26_23[7] , \nScanOut1018[4] , \nScanOut868[2] , \nScanOut77[4] , 
        \nOut6_11[2] , \nOut7_30[4] , \nOut6_12[1] , \nScanOut175[4] , 
        \nScanOut415[5] , \nScanOut693[5] , \nScanOut920[7] , \nScanOut814[4] , 
        \nScanOut521[6] , \nOut21_10[1] , \nOut20_31[7] , \nScanOut176[7] , 
        \nScanOut215[1] , \nScanOut321[2] , \nOut12_24[0] , \nOut28_20[0] , 
        \nScanOut641[3] , \nScanOut775[0] , \nOut12_27[3] , \nScanOut216[2] , 
        \nScanOut322[1] , \nScanOut416[6] , \nOut25_9[0] , \nOut28_23[3] , 
        \nScanOut522[5] , \nOut17_18[7] , \nOut21_13[2] , \nScanOut642[0] , 
        \nOut23_9[4] , \nScanOut776[3] , \nScanOut923[4] , \nScanOut111[0] , 
        \nScanOut690[6] , \nScanOut817[7] , \nOut29_8[1] , \nOut5_24[4] , 
        \nScanOut471[1] , \nScanOut545[2] , \nScanOut271[5] , \nScanOut345[6] , 
        \nOut10_30[0] , \nOut18_21[7] , \nScanOut625[7] , \nScanOut711[4] , 
        \nScanOut996[5] , \nScanOut597[4] , \nOut22_25[7] , \nScanOut1000[6] , 
        \nOut11_11[6] , \nScanOut397[0] , \nOut31_22[4] , \nScanOut944[3] , 
        \nScanOut13[0] , \nOut7_8[0] , \nOut11_12[5] , \nScanOut594[7] , 
        \nScanOut870[0] , \nScanOut1003[5] , \nOut12_8[1] , \nOut14_8[5] , 
        \nOut18_22[4] , \nOut22_26[4] , \nOut27_19[0] , \nOut0_18[3] , 
        \nOut1_8[4] , \nScanOut394[3] , \nScanOut873[3] , \nScanOut947[0] , 
        \nScanOut112[3] , \nScanOut472[2] , \nOut31_21[7] , \nScanOut546[1] , 
        \nScanOut712[7] , \nScanOut995[6] , \nScanOut34[5] , \nScanOut37[6] , 
        \nOut5_27[7] , \nOut9_28[2] , \nOut18_9[4] , \nScanOut626[4] , 
        \nScanOut272[6] , \nScanOut346[5] , \nScanOut284[6] , \nOut30_24[7] , 
        \nScanOut963[6] , \nOut4_21[4] , \nOut4_22[7] , \nOut10_17[5] , 
        \nOut15_28[1] , \nOut19_27[4] , \nScanOut857[5] , \nOut23_23[4] , 
        \nScanOut484[2] , \nScanOut136[5] , \nScanOut256[0] , \nScanOut362[3] , 
        \nScanOut602[2] , \nScanOut736[1] , \nScanOut885[3] , \nOut30_8[5] , 
        \nScanOut456[4] , \nScanOut562[7] , \nScanOut601[1] , \nScanOut735[2] , 
        \nScanOut886[0] , \nScanOut135[6] , \nScanOut255[3] , \nScanOut361[0] , 
        \nScanOut455[7] , \nScanOut561[4] , \nScanOut81[4] , \nScanOut287[5] , 
        \nScanOut854[6] , \nScanOut960[5] , \nOut30_27[4] , \nOut10_14[6] , 
        \nScanOut487[1] , \nScanOut1024[0] , \nOut19_24[7] , \nOut23_20[7] , 
        \nScanOut152[1] , \nScanOut232[4] , \nScanOut306[7] , \nScanOut666[6] , 
        \nScanOut752[5] , \nScanOut432[0] , \nOut20_16[2] , \nScanOut506[3] , 
        \nScanOut50[1] , \nScanOut53[2] , \nOut13_22[3] , \nOut29_26[3] , 
        \nOut25_29[6] , \nOut2_28[5] , \nOut7_17[1] , \nScanOut780[3] , 
        \nScanOut907[2] , \nScanOut833[1] , \nScanOut180[7] , \nOut7_14[2] , 
        \nScanOut904[1] , \nScanOut82[7] , \nScanOut183[4] , \nScanOut783[0] , 
        \nScanOut830[2] , \nScanOut231[7] , \nScanOut305[4] , \nScanOut151[2] , 
        \nOut13_21[0] , \nScanOut665[5] , \nScanOut751[6] , \nOut29_25[0] , 
        \nOut0_27[4] , \nScanOut431[3] , \nOut20_15[1] , \nScanOut505[0] , 
        \nScanOut619[3] , \nOut27_6[5] , \nOut5_18[0] , \nOut9_17[5] , 
        \nScanOut379[2] , \nOut13_3[5] , \nOut19_2[0] , \nScanOut579[6] , 
        \nOut21_6[1] , \nScanOut978[7] , \nOut6_3[4] , \nOut14_12[6] , 
        \nOut15_3[1] , \nOut27_26[7] , \nOut22_19[3] , \nScanOut8[6] , 
        \nOut0_24[7] , \nOut6_0[7] , \nOut13_0[6] , \nOut14_11[5] , 
        \nOut15_30[3] , \nOut15_0[2] , \nOut9_14[6] , \nOut27_25[4] , 
        \nOut19_1[3] , \nScanOut48[3] , \nOut3_12[2] , \nOut16_7[0] , 
        \nOut21_5[2] , \nOut27_5[6] , \nOut5_7[5] , \nOut28_3[5] , 
        \nOut2_26[3] , \nOut2_30[7] , \nOut3_7[1] , \nScanOut828[0] , 
        \nOut3_11[1] , \nScanOut99[6] , \nScanOut149[0] , \nScanOut229[5] , 
        \nOut10_7[4] , \nOut22_2[0] , \nScanOut749[4] , \nOut9_6[4] , 
        \nOut12_18[4] , \nOut24_13[1] , \nScanOut429[1] , \nOut17_27[0] , 
        \nOut24_2[4] , \nOut5_4[6] , \nOut9_5[7] , \nOut17_24[3] , 
        \nOut22_1[3] , \nOut24_1[7] , \nOut24_10[2] , \nOut25_31[4] , 
        \nOut16_4[3] , \nScanOut798[1] , \nOut28_0[6] , \nOut3_4[2] , 
        \nOut10_4[7] , \nScanOut198[5] , \nOut7_19[7] , \nScanOut909[4] , 
        \nScanOut308[1] , \nScanOut668[0] , \nOut16_13[1] , \nOut20_18[4] , 
        \nScanOut508[5] , \nOut25_27[0] , \nScanOut39[0] , \nOut1_13[5] , 
        \nOut2_25[0] , \nOut16_10[2] , \nOut25_24[3] , \nOut29_28[5] , 
        \nOut17_31[4] , \nOut8_23[4] , \nScanOut258[6] , \nScanOut738[7] , 
        \nScanOut138[3] , \nScanOut458[2] , \nOut30_6[3] , \nScanOut859[3] , 
        \nScanOut21[2] , \nScanOut22[1] , \nOut1_10[6] , \nScanOut289[3] , 
        \nOut10_19[3] , \nOut15_26[7] , \nOut19_29[2] , \nOut26_12[6] , 
        \nOut30_29[2] , \nOut15_25[4] , \nScanOut489[7] , \nOut26_11[5] , 
        \nOut27_30[3] , \nScanOut888[6] , \nScanOut45[6] , \nScanOut46[5] , 
        \nScanOut94[3] , \nScanOut227[3] , \nOut8_20[7] , \nScanOut313[0] , 
        \nOut30_5[0] , \nOut5_9[3] , \nScanOut147[6] , \nOut12_16[2] , 
        \nScanOut673[1] , \nScanOut747[2] , \nOut28_12[2] , \nOut6_23[0] , 
        \nOut9_8[2] , \nScanOut427[7] , \nOut17_29[6] , \nOut21_22[3] , 
        \nOut16_9[6] , \nScanOut513[4] , \nScanOut912[5] , \nOut3_9[7] , 
        \nScanOut795[4] , \nScanOut826[6] , \nScanOut195[0] , \nOut10_9[2] , 
        \nScanOut97[0] , \nOut6_20[3] , \nScanOut796[7] , \nScanOut196[3] , 
        \nScanOut825[5] , \nScanOut911[6] , \nScanOut144[5] , \nScanOut224[0] , 
        \nScanOut310[3] , \nScanOut670[2] , \nScanOut744[1] , \nScanOut424[4] , 
        \nScanOut510[7] , \nOut21_21[0] , \nOut28_11[1] , \nOut12_15[1] , 
        \nOut29_30[7] , \nOut0_29[2] , \nScanOut291[1] , \nScanOut842[2] , 
        \nScanOut976[1] , \nOut31_10[6] , \nOut30_31[0] , \nOut11_23[4] , 
        \nScanOut491[5] , \nOut27_28[1] , \nOut18_13[5] , \nOut22_17[5] , 
        \nScanOut723[6] , \nOut27_8[3] , \nScanOut890[4] , \nScanOut120[1] , 
        \nScanOut123[2] , \nOut5_16[6] , \nOut9_19[3] , \nScanOut617[5] , 
        \nScanOut243[7] , \nScanOut377[4] , \nScanOut443[3] , \nScanOut577[0] , 
        \nOut21_8[7] , \nOut5_15[5] , \nScanOut240[4] , \nScanOut374[7] , 
        \nScanOut614[6] , \nScanOut720[5] , \nScanOut893[7] , \nScanOut292[2] , 
        \nScanOut440[0] , \nScanOut574[3] , \nOut31_13[5] , \nScanOut975[2] , 
        \nScanOut104[7] , \nOut11_20[7] , \nScanOut492[6] , \nOut18_10[6] , 
        \nOut19_31[0] , \nScanOut841[1] , \nOut22_14[6] , \nScanOut464[6] , 
        \nScanOut550[5] , \nOut4_10[5] , \nOut5_31[3] , \nScanOut630[0] , 
        \nScanOut704[3] , \nScanOut983[2] , \nScanOut350[1] , \nScanOut264[2] , 
        \nOut10_25[7] , \nScanOut1015[1] , \nScanOut582[3] , \nOut22_30[0] , 
        \nOut23_11[6] , \nScanOut8[4] , \nOut0_15[6] , \nOut1_5[1] , 
        \nOut2_19[4] , \nScanOut61[0] , \nScanOut107[4] , \nOut10_26[4] , 
        \nScanOut382[7] , \nOut19_15[6] , \nScanOut865[7] , \nScanOut951[4] , 
        \nOut15_19[0] , \nOut19_16[5] , \nOut30_16[5] , \nScanOut581[0] , 
        \nOut23_12[5] , \nScanOut1016[2] , \nScanOut381[4] , \nOut30_15[6] , 
        \nScanOut866[4] , \nScanOut952[7] , \nOut4_13[6] , \nScanOut353[2] , 
        \nScanOut467[5] , \nScanOut553[6] , \nOut7_25[3] , \nScanOut267[1] , 
        \nScanOut633[3] , \nScanOut707[0] , \nScanOut980[1] , \nScanOut935[0] , 
        \nScanOut62[3] , \nScanOut160[3] , \nOut13_10[1] , \nOut12_31[7] , 
        \nScanOut686[2] , \nScanOut801[3] , \nScanOut163[0] , \nScanOut200[6] , 
        \nScanOut334[5] , \nScanOut400[2] , \nOut29_14[1] , \nScanOut534[1] , 
        \nOut20_24[0] , \nScanOut403[1] , \nScanOut654[4] , \nScanOut760[7] , 
        \nScanOut537[2] , \nOut20_27[3] , \nScanOut203[5] , \nScanOut337[6] , 
        \nOut13_13[2] , \nOut25_18[7] , \nOut29_17[2] , \nScanOut657[7] , 
        \nScanOut763[4] , \nOut7_26[0] , \nScanOut685[1] , \nScanOut936[3] , 
        \nScanOut802[0] , \nOut7_5[5] , \nOut14_5[0] , \nOut14_20[4] , 
        \nScanOut599[2] , \nOut27_14[5] , \nScanOut399[6] , \nOut9_25[7] , 
        \nOut12_5[4] , \nOut18_4[1] , \nOut20_0[0] , \nOut26_0[4] , 
        \nScanOut998[3] , \nOut0_16[5] , \nScanOut548[7] , \nOut20_3[3] , 
        \nScanOut628[2] , \nOut26_3[7] , \nOut2_1[0] , \nOut1_6[2] , 
        \nOut5_29[1] , \nOut7_6[6] , \nOut9_26[4] , \nScanOut348[3] , 
        \nOut18_7[2] , \nOut12_6[7] , \nOut14_6[3] , \nOut14_23[7] , 
        \nOut22_28[2] , \nOut27_17[6] , \nScanOut949[6] , \nOut8_0[5] , 
        \nOut25_4[5] , \nOut11_1[5] , \nOut17_15[2] , \nOut23_4[1] , 
        \nOut24_21[3] , \nOut2_2[3] , \nOut3_20[0] , \nOut4_1[4] , 
        \nOut17_1[1] , \nOut29_5[4] , \nOut2_25[2] , \nScanOut79[2] , 
        \nOut3_23[3] , \nOut11_2[6] , \nOut17_2[2] , \nOut4_2[7] , 
        \nScanOut178[1] , \nScanOut819[1] , \nOut29_6[7] , \nScanOut218[4] , 
        \nOut8_3[6] , \nOut12_29[5] , \nScanOut418[0] , \nOut24_22[0] , 
        \nOut17_16[1] , \nOut25_7[6] , \nOut23_7[2] , \nScanOut778[5] , 
        \nOut16_10[0] , \nOut17_31[6] , \nOut25_24[1] , \nOut16_13[3] , 
        \nScanOut508[7] , \nOut20_18[6] , \nOut25_27[2] , \nOut29_28[7] , 
        \nOut2_26[1] , \nOut7_19[5] , \nScanOut308[3] , \nScanOut668[2] , 
        \nScanOut909[6] , \nOut30_5[2] , \nOut1_10[4] , \nOut8_20[5] , 
        \nScanOut888[4] , \nScanOut289[1] , \nOut15_25[6] , \nScanOut489[5] , 
        \nOut26_11[7] , \nOut27_30[1] , \nOut15_26[5] , \nOut30_29[0] , 
        \nOut0_15[4] , \nOut0_16[7] , \nScanOut21[0] , \nScanOut39[2] , 
        \nOut10_19[1] , \nOut19_29[0] , \nOut26_12[4] , \nScanOut859[1] , 
        \nOut1_13[7] , \nScanOut138[1] , \nOut8_23[6] , \nScanOut258[4] , 
        \nScanOut458[0] , \nOut30_6[1] , \nScanOut45[4] , \nScanOut97[2] , 
        \nScanOut144[7] , \nScanOut424[6] , \nScanOut510[5] , \nScanOut738[5] , 
        \nOut21_21[2] , \nOut29_30[5] , \nOut12_15[3] , \nOut28_11[3] , 
        \nScanOut670[0] , \nScanOut744[3] , \nScanOut196[1] , \nScanOut224[2] , 
        \nScanOut310[1] , \nScanOut796[5] , \nScanOut825[7] , \nScanOut46[7] , 
        \nOut3_9[5] , \nOut6_20[1] , \nScanOut911[4] , \nScanOut195[2] , 
        \nOut6_23[2] , \nOut10_9[0] , \nOut16_9[4] , \nScanOut826[4] , 
        \nScanOut912[7] , \nScanOut795[6] , \nScanOut94[1] , \nOut5_9[1] , 
        \nScanOut147[4] , \nOut12_16[0] , \nScanOut227[1] , \nOut9_8[0] , 
        \nOut28_12[0] , \nScanOut427[5] , \nScanOut513[6] , \nOut21_22[1] , 
        \nOut17_29[4] , \nScanOut313[2] , \nScanOut673[3] , \nScanOut747[0] , 
        \nScanOut292[0] , \nOut11_20[5] , \nOut18_10[4] , \nOut19_31[2] , 
        \nOut22_14[4] , \nScanOut492[4] , \nScanOut841[3] , \nOut31_13[7] , 
        \nScanOut975[0] , \nScanOut22[3] , \nOut0_29[0] , \nScanOut120[3] , 
        \nScanOut123[0] , \nOut5_15[7] , \nScanOut240[6] , \nScanOut440[2] , 
        \nScanOut574[1] , \nScanOut374[5] , \nScanOut443[1] , \nScanOut577[2] , 
        \nScanOut614[4] , \nScanOut720[7] , \nScanOut893[5] , \nOut21_8[5] , 
        \nOut5_16[4] , \nScanOut243[5] , \nScanOut617[7] , \nOut27_8[1] , 
        \nScanOut890[6] , \nScanOut723[4] , \nOut9_19[1] , \nScanOut377[6] , 
        \nOut11_23[6] , \nScanOut491[7] , \nOut27_28[3] , \nOut18_13[7] , 
        \nOut22_17[7] , \nScanOut842[0] , \nOut1_6[0] , \nOut2_19[6] , 
        \nScanOut62[1] , \nScanOut104[5] , \nOut4_10[7] , \nScanOut107[6] , 
        \nOut4_13[4] , \nScanOut267[3] , \nScanOut291[3] , \nScanOut976[3] , 
        \nOut31_10[4] , \nOut30_31[2] , \nScanOut353[0] , \nScanOut633[1] , 
        \nScanOut707[2] , \nScanOut980[3] , \nScanOut264[0] , \nOut10_25[5] , 
        \nOut10_26[6] , \nScanOut381[6] , \nScanOut467[7] , \nScanOut553[4] , 
        \nOut30_15[4] , \nOut15_19[2] , \nOut19_16[7] , \nScanOut866[6] , 
        \nScanOut952[5] , \nOut23_12[7] , \nScanOut382[5] , \nScanOut581[2] , 
        \nScanOut865[5] , \nScanOut1016[0] , \nScanOut951[6] , 
        \nScanOut582[1] , \nOut30_16[7] , \nOut19_15[4] , \nOut22_30[2] , 
        \nScanOut1015[3] , \nOut23_11[4] , \nScanOut630[2] , \nScanOut704[1] , 
        \nScanOut983[0] , \nOut5_31[1] , \nScanOut350[3] , \nScanOut464[4] , 
        \nScanOut550[7] , \nScanOut685[3] , \nScanOut802[2] , \nOut7_26[2] , 
        \nScanOut936[1] , \nScanOut61[2] , \nScanOut160[1] , \nScanOut163[2] , 
        \nScanOut203[7] , \nScanOut657[5] , \nScanOut763[6] , \nScanOut337[4] , 
        \nScanOut403[3] , \nScanOut537[0] , \nOut20_27[1] , \nOut29_17[0] , 
        \nScanOut200[4] , \nOut13_13[0] , \nOut25_18[5] , \nScanOut334[7] , 
        \nOut13_10[3] , \nScanOut654[6] , \nScanOut760[5] , \nOut12_31[5] , 
        \nOut29_14[3] , \nOut7_25[1] , \nScanOut400[0] , \nScanOut534[3] , 
        \nOut20_24[2] , \nScanOut686[0] , \nScanOut801[1] , \nScanOut935[2] , 
        \nOut12_6[5] , \nScanOut949[4] , \nOut7_6[4] , \nOut27_17[4] , 
        \nOut14_6[1] , \nOut14_23[5] , \nScanOut628[0] , \nOut22_28[0] , 
        \nOut5_29[3] , \nScanOut348[1] , \nOut26_3[5] , \nOut9_25[5] , 
        \nOut9_26[6] , \nScanOut548[5] , \nOut18_7[0] , \nOut20_3[1] , 
        \nOut18_4[3] , \nOut2_1[2] , \nOut2_2[1] , \nOut1_5[3] , \nOut20_0[2] , 
        \nOut26_0[6] , \nScanOut998[1] , \nScanOut79[0] , \nOut3_23[1] , 
        \nScanOut178[3] , \nOut7_5[7] , \nOut12_5[6] , \nScanOut399[4] , 
        \nOut14_5[2] , \nOut14_20[6] , \nScanOut218[6] , \nScanOut599[0] , 
        \nOut27_14[7] , \nOut23_7[0] , \nScanOut778[7] , \nOut8_3[4] , 
        \nOut12_29[7] , \nOut24_22[2] , \nScanOut418[2] , \nOut17_16[3] , 
        \nOut17_2[0] , \nOut25_7[4] , \nOut4_2[5] , \nOut29_6[5] , 
        \nScanOut819[3] , \nOut3_20[2] , \nOut4_1[6] , \nOut11_2[4] , 
        \nOut29_5[6] , \nOut11_1[7] , \nOut17_1[3] , \nOut2_14[3] , 
        \nOut2_17[0] , \nOut7_28[4] , \nOut8_0[7] , \nOut23_4[3] , 
        \nScanOut339[2] , \nOut17_15[0] , \nOut25_4[7] , \nScanOut659[3] , 
        \nOut24_21[1] , \nOut16_22[2] , \nScanOut539[6] , \nOut20_29[7] , 
        \nOut25_16[3] , \nOut29_19[6] , \nScanOut938[7] , \nOut1_21[5] , 
        \nOut1_22[6] , \nOut8_12[7] , \nScanOut269[5] , \nOut10_28[0] , 
        \nOut15_17[4] , \nOut16_21[1] , \nScanOut688[6] , \nOut25_15[0] , 
        \nScanOut868[0] , \nOut19_18[1] , \nOut26_23[5] , \nScanOut1018[6] , 
        \nScanOut109[0] , \nScanOut709[4] , \nScanOut469[1] , \nOut31_3[3] , 
        \nScanOut77[6] , \nOut6_12[3] , \nOut8_11[4] , \nOut9_30[2] , 
        \nOut15_14[7] , \nOut26_20[6] , \nOut30_18[1] , \nScanOut690[4] , 
        \nScanOut817[5] , \nOut29_8[3] , \nScanOut923[6] , \nScanOut5[1] , 
        \nScanOut10[1] , \nScanOut13[2] , \nOut0_18[1] , \nScanOut74[5] , 
        \nScanOut175[6] , \nScanOut176[5] , \nScanOut216[0] , \nScanOut322[3] , 
        \nOut23_9[6] , \nOut12_27[1] , \nScanOut642[2] , \nScanOut776[1] , 
        \nOut28_23[1] , \nScanOut215[3] , \nScanOut416[4] , \nScanOut522[7] , 
        \nOut17_18[5] , \nOut25_9[2] , \nOut21_13[0] , \nScanOut641[1] , 
        \nScanOut775[2] , \nScanOut321[0] , \nScanOut415[7] , \nScanOut521[4] , 
        \nOut21_10[3] , \nOut20_31[5] , \nOut28_20[2] , \nOut12_24[2] , 
        \nScanOut693[7] , \nScanOut814[6] , \nOut6_11[0] , \nScanOut920[5] , 
        \nOut7_30[6] , \nScanOut112[1] , \nOut5_27[5] , \nScanOut272[4] , 
        \nScanOut626[6] , \nScanOut712[5] , \nScanOut995[4] , \nOut9_28[0] , 
        \nScanOut346[7] , \nOut18_9[6] , \nScanOut472[0] , \nScanOut546[3] , 
        \nScanOut873[1] , \nOut1_8[6] , \nOut12_8[3] , \nScanOut947[2] , 
        \nOut7_8[2] , \nScanOut394[1] , \nOut27_19[2] , \nOut31_21[5] , 
        \nOut11_12[7] , \nScanOut397[2] , \nOut14_8[7] , \nScanOut594[5] , 
        \nScanOut1003[7] , \nOut18_22[6] , \nOut22_26[6] , \nOut31_22[6] , 
        \nScanOut870[2] , \nScanOut944[1] , \nScanOut34[7] , \nScanOut111[2] , 
        \nOut5_24[6] , \nScanOut271[7] , \nOut10_30[2] , \nOut11_11[4] , 
        \nOut18_21[5] , \nOut22_25[5] , \nScanOut597[6] , \nScanOut1000[4] , 
        \nScanOut345[4] , \nScanOut625[5] , \nScanOut711[6] , \nScanOut996[7] , 
        \nOut10_14[4] , \nScanOut471[3] , \nScanOut545[0] , \nScanOut487[3] , 
        \nScanOut1024[2] , \nOut19_24[5] , \nOut23_20[5] , \nScanOut854[4] , 
        \nScanOut37[4] , \nOut4_21[6] , \nScanOut135[4] , \nScanOut287[7] , 
        \nScanOut960[7] , \nScanOut455[5] , \nScanOut561[6] , \nOut30_27[6] , 
        \nScanOut255[1] , \nScanOut601[3] , \nScanOut886[2] , \nScanOut735[0] , 
        \nScanOut361[2] , \nOut4_22[5] , \nScanOut136[7] , \nOut30_8[7] , 
        \nScanOut256[2] , \nScanOut456[6] , \nScanOut562[5] , \nScanOut362[1] , 
        \nScanOut284[4] , \nOut10_17[7] , \nOut15_28[3] , \nScanOut602[0] , 
        \nOut19_27[6] , \nScanOut736[3] , \nScanOut885[1] , \nOut23_23[6] , 
        \nScanOut484[0] , \nScanOut857[7] , \nOut30_24[5] , \nScanOut963[4] , 
        \nOut13_21[2] , \nScanOut6[2] , \nScanOut50[3] , \nScanOut82[5] , 
        \nScanOut151[0] , \nOut29_25[2] , \nScanOut231[5] , \nScanOut431[1] , 
        \nScanOut505[2] , \nOut20_15[3] , \nScanOut305[6] , \nScanOut665[7] , 
        \nScanOut751[4] , \nScanOut183[6] , \nOut7_14[0] , \nScanOut830[0] , 
        \nScanOut783[2] , \nScanOut904[3] , \nScanOut53[0] , \nScanOut180[5] , 
        \nScanOut780[1] , \nScanOut833[3] , \nOut2_28[7] , \nOut7_17[3] , 
        \nScanOut907[0] , \nScanOut432[2] , \nScanOut506[1] , \nOut20_16[0] , 
        \nOut29_26[1] , \nOut0_24[5] , \nScanOut81[6] , \nScanOut152[3] , 
        \nOut13_22[1] , \nOut25_29[4] , \nScanOut666[4] , \nScanOut752[7] , 
        \nScanOut232[6] , \nOut9_14[4] , \nScanOut306[5] , \nOut19_1[1] , 
        \nOut21_5[0] , \nOut27_5[4] , \nOut6_0[5] , \nOut14_11[7] , 
        \nOut15_30[1] , \nOut15_0[0] , \nOut27_25[6] , \nOut0_3[2] , 
        \nOut6_3[6] , \nOut13_0[4] , \nOut27_26[5] , \nOut13_3[7] , 
        \nOut14_12[4] , \nOut15_3[3] , \nOut22_19[1] , \nScanOut978[5] , 
        \nOut0_27[6] , \nScanOut579[4] , \nScanOut619[1] , \nOut21_6[3] , 
        \nScanOut48[1] , \nOut2_30[5] , \nOut3_4[0] , \nOut5_18[2] , 
        \nScanOut379[0] , \nOut19_2[2] , \nOut27_6[7] , \nScanOut198[7] , 
        \nOut9_17[7] , \nOut10_4[5] , \nOut5_4[4] , \nScanOut798[3] , 
        \nOut28_0[4] , \nOut3_7[3] , \nOut3_11[3] , \nScanOut99[4] , 
        \nOut9_5[5] , \nOut16_4[1] , \nOut17_24[1] , \nOut24_1[5] , 
        \nOut24_10[0] , \nOut25_31[6] , \nScanOut149[2] , \nOut22_1[1] , 
        \nScanOut229[7] , \nOut9_6[6] , \nOut12_18[6] , \nOut24_13[3] , 
        \nScanOut429[3] , \nOut24_2[6] , \nOut17_27[2] , \nOut22_2[2] , 
        \nScanOut749[6] , \nOut3_12[0] , \nOut10_7[6] , \nOut16_7[2] , 
        \nScanOut828[2] , \nOut1_24[1] , \nOut5_7[7] , \nOut28_3[7] , 
        \nScanOut389[7] , \nOut14_30[5] , \nScanOut589[3] , \nOut26_25[2] , 
        \nOut15_11[3] , \nOut31_5[4] , \nOut1_27[2] , \nOut4_18[6] , 
        \nOut8_14[0] , \nScanOut988[2] , \nScanOut558[6] , \nOut31_6[7] , 
        \nOut8_17[3] , \nScanOut358[2] , \nScanOut638[3] , \nOut15_12[0] , 
        \nOut16_24[5] , \nOut23_19[5] , \nOut25_10[4] , \nOut26_26[1] , 
        \nScanOut959[7] , \nOut24_31[2] , \nScanOut15[5] , \nOut2_11[7] , 
        \nOut3_30[1] , \nOut2_12[4] , \nScanOut69[3] , \nScanOut809[0] , 
        \nScanOut114[6] , \nScanOut168[0] , \nScanOut408[1] , \nOut16_27[6] , 
        \nScanOut208[5] , \nOut13_18[2] , \nOut25_13[7] , \nScanOut768[4] , 
        \nOut5_21[2] , \nScanOut274[3] , \nScanOut474[7] , \nScanOut540[4] , 
        \nScanOut340[0] , \nOut11_14[0] , \nOut18_24[1] , \nScanOut620[1] , 
        \nOut22_20[1] , \nScanOut714[2] , \nScanOut993[3] , \nScanOut392[6] , 
        \nScanOut592[2] , \nScanOut1005[0] , \nScanOut875[6] , \nOut31_27[2] , 
        \nScanOut16[6] , \nOut11_17[3] , \nScanOut941[5] , \nOut14_28[7] , 
        \nOut18_27[2] , \nScanOut591[1] , \nScanOut1006[3] , \nOut22_23[2] , 
        \nScanOut876[5] , \nScanOut942[6] , \nScanOut117[5] , \nScanOut391[5] , 
        \nOut31_24[1] , \nScanOut477[4] , \nScanOut543[7] , \nOut20_8[3] , 
        \nOut5_22[1] , \nScanOut277[0] , \nScanOut623[2] , \nScanOut717[1] , 
        \nOut26_8[7] , \nScanOut990[0] , \nScanOut343[3] , \nScanOut811[2] , 
        \nScanOut0[5] , \nScanOut3[6] , \nOut2_9[3] , \nScanOut71[1] , 
        \nOut6_14[4] , \nScanOut696[3] , \nScanOut925[1] , \nScanOut170[2] , 
        \nOut12_21[6] , \nScanOut410[3] , \nScanOut524[0] , \nOut21_15[7] , 
        \nOut28_25[6] , \nScanOut173[1] , \nScanOut210[7] , \nScanOut644[5] , 
        \nScanOut770[6] , \nScanOut324[4] , \nOut28_26[5] , \nScanOut213[4] , 
        \nOut8_8[6] , \nOut12_22[5] , \nScanOut413[0] , \nScanOut527[3] , 
        \nOut24_29[0] , \nOut21_16[4] , \nScanOut327[7] , \nScanOut647[6] , 
        \nScanOut773[5] , \nScanOut72[2] , \nOut3_28[3] , \nOut11_9[6] , 
        \nOut4_9[7] , \nOut17_9[2] , \nScanOut695[0] , \nScanOut812[1] , 
        \nScanOut84[2] , \nOut6_17[7] , \nScanOut926[2] , \nScanOut663[0] , 
        \nScanOut757[3] , \nScanOut237[2] , \nScanOut303[1] , \nOut13_27[5] , 
        \nScanOut437[6] , \nScanOut503[5] , \nOut16_18[1] , \nOut20_13[4] , 
        \nScanOut55[7] , \nScanOut56[4] , \nScanOut157[7] , \nOut29_23[5] , 
        \nOut7_12[7] , \nScanOut836[7] , \nScanOut785[5] , \nScanOut902[4] , 
        \nScanOut185[1] , \nScanOut786[6] , \nScanOut835[4] , \nScanOut87[1] , 
        \nScanOut186[2] , \nOut6_30[2] , \nOut7_11[4] , \nScanOut901[7] , 
        \nScanOut234[1] , \nScanOut300[2] , \nScanOut660[3] , \nScanOut754[0] , 
        \nOut29_20[6] , \nOut0_5[5] , \nOut0_6[6] , \nOut0_22[2] , 
        \nScanOut31[3] , \nScanOut32[0] , \nScanOut154[4] , \nScanOut281[0] , 
        \nOut13_24[6] , \nScanOut434[5] , \nScanOut500[6] , \nOut21_31[1] , 
        \nOut20_10[7] , \nScanOut852[3] , \nOut30_21[1] , \nOut1_18[5] , 
        \nOut4_27[1] , \nOut8_28[4] , \nScanOut253[6] , \nOut10_12[3] , 
        \nOut19_22[2] , \nOut23_26[2] , \nScanOut966[0] , \nScanOut481[4] , 
        \nOut26_19[6] , \nScanOut1022[5] , \nScanOut367[5] , \nOut4_24[2] , 
        \nScanOut133[3] , \nScanOut607[4] , \nScanOut880[5] , \nScanOut733[7] , 
        \nScanOut250[5] , \nScanOut453[2] , \nScanOut567[1] , \nScanOut604[7] , 
        \nScanOut730[4] , \nScanOut883[6] , \nScanOut364[6] , \nScanOut130[0] , 
        \nScanOut450[1] , \nScanOut564[2] , \nScanOut851[0] , \nScanOut965[3] , 
        \nOut3_1[4] , \nOut3_2[7] , \nOut3_17[4] , \nScanOut282[3] , 
        \nOut10_11[0] , \nOut30_22[2] , \nOut11_30[6] , \nScanOut482[7] , 
        \nOut19_21[1] , \nScanOut1021[6] , \nOut23_25[1] , \nOut5_2[3] , 
        \nOut6_28[0] , \nOut16_2[6] , \nScanOut919[5] , \nOut28_6[3] , 
        \nOut3_14[7] , \nOut5_1[0] , \nOut9_3[2] , \nOut10_2[2] , 
        \nScanOut318[0] , \nScanOut678[1] , \nOut22_7[6] , \nOut24_16[7] , 
        \nOut28_19[2] , \nOut9_0[1] , \nScanOut518[4] , \nOut24_7[2] , 
        \nOut17_22[6] , \nOut21_29[3] , \nOut22_4[5] , \nOut17_21[5] , 
        \nOut24_4[1] , \nOut24_15[4] , \nOut28_5[0] , \nOut10_1[1] , 
        \nOut16_1[5] , \nOut27_3[3] , \nScanOut29[1] , \nScanOut128[2] , 
        \nScanOut248[7] , \nOut19_7[6] , \nScanOut728[6] , \nOut9_12[3] , 
        \nScanOut448[3] , \nOut13_6[3] , \nOut21_3[7] , \nScanOut849[2] , 
        \nOut6_6[2] , \nOut11_28[4] , \nOut27_23[1] , \nOut14_17[0] , 
        \nOut15_6[7] , \nOut18_18[5] , \nOut0_8[0] , \nOut0_21[1] , 
        \nOut6_5[1] , \nScanOut299[2] , \nOut13_5[0] , \nOut31_18[5] , 
        \nOut14_14[3] , \nOut15_5[4] , \nOut27_20[2] , \nOut8_30[6] , 
        \nScanOut499[6] , \nOut19_4[5] , \nOut9_11[0] , \nScanOut27[7] , 
        \nOut1_15[0] , \nOut1_16[3] , \nOut4_29[7] , \nScanOut369[3] , 
        \nOut21_0[4] , \nOut27_0[0] , \nScanOut898[7] , \nOut8_26[2] , 
        \nScanOut609[2] , \nOut15_20[2] , \nOut15_23[1] , \nScanOut569[7] , 
        \nOut30_3[5] , \nOut23_28[4] , \nScanOut968[6] , \nOut26_14[3] , 
        \nOut26_17[0] , \nOut2_20[6] , \nOut2_23[5] , \nScanOut58[2] , 
        \nOut8_25[1] , \nScanOut838[1] , \nOut30_0[6] , \nScanOut89[7] , 
        \nScanOut159[1] , \nScanOut239[4] , \nScanOut759[5] , \nScanOut439[0] , 
        \nOut16_16[7] , \nOut13_29[3] , \nOut25_22[6] , \nOut16_15[4] , 
        \nOut25_21[5] , \nScanOut188[4] , \nScanOut788[0] , \nOut13_8[5] , 
        \nScanOut847[4] , \nScanOut973[7] , \nScanOut294[7] , \nOut11_26[2] , 
        \nOut31_15[0] , \nScanOut24[4] , \nScanOut125[7] , \nScanOut126[4] , 
        \nOut5_13[0] , \nOut6_8[4] , \nScanOut246[1] , \nOut14_19[6] , 
        \nOut15_8[1] , \nScanOut494[3] , \nOut18_16[3] , \nScanOut612[3] , 
        \nOut22_12[3] , \nScanOut726[0] , \nScanOut895[2] , \nScanOut372[2] , 
        \nOut19_9[0] , \nScanOut446[5] , \nScanOut572[6] , \nOut5_10[3] , 
        \nScanOut245[2] , \nScanOut371[1] , \nOut4_31[5] , \nScanOut611[0] , 
        \nScanOut896[1] , \nScanOut725[3] , \nScanOut297[4] , \nScanOut445[6] , 
        \nScanOut571[5] , \nScanOut844[7] , \nOut31_16[3] , \nOut3_19[2] , 
        \nScanOut91[5] , \nScanOut222[5] , \nOut11_25[1] , \nOut18_15[0] , 
        \nOut22_11[0] , \nOut23_30[6] , \nScanOut970[4] , \nScanOut497[0] , 
        \nScanOut316[6] , \nOut22_9[0] , \nScanOut676[7] , \nScanOut742[4] , 
        \nScanOut142[0] , \nOut12_13[4] , \nOut24_18[1] , \nOut28_17[4] , 
        \nScanOut422[1] , \nScanOut516[2] , \nOut21_27[5] , \nOut24_9[4] , 
        \nOut0_3[6] , \nOut0_10[0] , \nOut1_0[7] , \nOut2_4[6] , 
        \nScanOut40[0] , \nScanOut43[3] , \nScanOut790[2] , \nScanOut823[0] , 
        \nOut28_8[5] , \nOut6_25[5] , \nOut6_26[6] , \nScanOut917[3] , 
        \nScanOut190[6] , \nScanOut820[3] , \nScanOut914[0] , \nScanOut793[1] , 
        \nOut1_29[4] , \nScanOut64[6] , \nScanOut92[6] , \nScanOut193[5] , 
        \nScanOut675[4] , \nScanOut741[7] , \nScanOut141[3] , \nScanOut221[6] , 
        \nScanOut315[5] , \nOut12_10[7] , \nScanOut421[2] , \nScanOut515[1] , 
        \nOut21_24[6] , \nOut13_31[1] , \nScanOut683[4] , \nOut28_14[7] , 
        \nScanOut804[5] , \nScanOut67[5] , \nScanOut165[5] , \nOut7_20[5] , 
        \nScanOut930[6] , \nOut28_30[1] , \nOut29_11[7] , \nScanOut166[6] , 
        \nScanOut205[0] , \nOut13_15[7] , \nScanOut405[4] , \nScanOut531[7] , 
        \nOut20_21[6] , \nScanOut331[3] , \nOut13_16[4] , \nScanOut406[7] , 
        \nOut16_29[0] , \nScanOut532[4] , \nScanOut651[2] , \nScanOut765[1] , 
        \nOut20_22[5] , \nOut29_12[4] , \nScanOut206[3] , \nScanOut652[1] , 
        \nScanOut766[2] , \nOut7_23[6] , \nScanOut332[0] , \nScanOut680[7] , 
        \nScanOut807[6] , \nScanOut933[5] , \nScanOut101[1] , \nScanOut461[0] , 
        \nScanOut555[3] , \nScanOut102[2] , \nOut4_15[3] , \nScanOut261[4] , 
        \nScanOut635[6] , \nScanOut701[5] , \nScanOut986[4] , \nOut10_20[1] , 
        \nScanOut355[7] , \nOut10_23[2] , \nScanOut387[1] , \nOut19_10[0] , 
        \nScanOut587[5] , \nScanOut1010[7] , \nOut18_31[6] , \nOut23_14[0] , 
        \nScanOut860[1] , \nOut30_13[3] , \nScanOut954[2] , \nScanOut584[6] , 
        \nOut19_13[3] , \nOut23_17[3] , \nOut26_28[7] , \nScanOut384[2] , 
        \nScanOut1013[4] , \nScanOut863[2] , \nOut30_10[0] , \nScanOut957[1] , 
        \nOut4_16[0] , \nOut8_19[5] , \nScanOut262[7] , \nScanOut462[3] , 
        \nScanOut556[0] , \nOut31_8[1] , \nScanOut356[4] , \nOut8_5[3] , 
        \nOut17_10[4] , \nOut16_31[2] , \nScanOut636[5] , \nScanOut702[6] , 
        \nScanOut985[7] , \nOut11_4[3] , \nOut23_1[7] , \nOut24_24[5] , 
        \nOut25_1[3] , \nOut2_7[5] , \nOut3_25[6] , \nOut4_4[2] , 
        \nScanOut698[5] , \nOut29_0[2] , \nOut17_4[7] , \nOut3_26[5] , 
        \nOut11_7[0] , \nOut4_7[1] , \nOut17_7[4] , \nOut29_3[1] , 
        \nOut6_19[1] , \nScanOut928[4] , \nOut7_0[3] , \nOut8_6[0] , 
        \nScanOut529[5] , \nOut24_27[6] , \nOut28_28[3] , \nScanOut329[1] , 
        \nOut17_13[7] , \nOut21_18[2] , \nOut25_2[0] , \nOut23_2[4] , 
        \nOut14_25[2] , \nOut14_0[6] , \nScanOut649[0] , \nOut27_11[3] , 
        \nOut26_30[5] , \nOut31_29[4] , \nOut1_31[6] , \nOut9_20[1] , 
        \nOut12_0[2] , \nOut20_5[6] , \nOut18_1[7] , \nOut0_13[3] , 
        \nScanOut119[3] , \nScanOut479[2] , \nOut26_5[2] , \nOut20_6[5] , 
        \nScanOut18[0] , \nOut7_3[0] , \nScanOut279[6] , \nScanOut719[7] , 
        \nOut26_6[1] , \nOut9_23[2] , \nOut18_2[4] , \nOut11_19[5] , 
        \nOut12_3[1] , \nOut14_3[5] , \nOut27_12[0] , \nScanOut1008[5] , 
        \nOut14_26[1] , \nOut18_29[4] , \nScanOut878[3] , \nOut0_27[2] , 
        \nOut1_3[4] , \nOut5_18[6] , \nScanOut379[4] , \nOut19_2[6] , 
        \nOut9_17[3] , \nScanOut619[5] , \nOut27_6[3] , \nScanOut579[0] , 
        \nOut21_6[7] , \nOut6_3[2] , \nOut13_3[3] , \nOut14_12[0] , 
        \nOut15_3[7] , \nScanOut978[1] , \nOut22_19[5] , \nOut27_26[1] , 
        \nOut13_0[0] , \nScanOut5[5] , \nScanOut6[6] , \nOut0_24[1] , 
        \nOut6_0[1] , \nOut27_25[2] , \nOut14_11[3] , \nOut15_30[5] , 
        \nOut15_0[4] , \nScanOut34[3] , \nScanOut37[0] , \nScanOut48[5] , 
        \nOut9_14[0] , \nOut19_1[5] , \nOut27_5[0] , \nOut21_5[4] , 
        \nScanOut828[6] , \nOut28_3[3] , \nOut2_30[1] , \nOut3_7[7] , 
        \nOut3_12[4] , \nOut5_7[3] , \nOut10_7[2] , \nOut16_7[6] , 
        \nScanOut99[0] , \nScanOut149[6] , \nScanOut229[3] , \nScanOut749[2] , 
        \nOut9_6[2] , \nOut22_2[6] , \nScanOut429[7] , \nOut17_27[6] , 
        \nOut24_2[2] , \nOut12_18[2] , \nOut24_13[7] , \nOut22_1[5] , 
        \nOut9_5[1] , \nOut24_10[4] , \nOut25_31[2] , \nOut17_24[5] , 
        \nOut24_1[1] , \nOut3_4[4] , \nOut3_11[7] , \nOut5_4[0] , 
        \nOut16_4[5] , \nScanOut798[7] , \nOut28_0[0] , \nScanOut198[3] , 
        \nOut10_4[1] , \nScanOut857[3] , \nScanOut963[0] , \nOut4_21[2] , 
        \nOut4_22[1] , \nScanOut256[6] , \nScanOut284[0] , \nOut10_17[3] , 
        \nOut30_24[1] , \nOut15_28[7] , \nScanOut484[4] , \nOut19_27[2] , 
        \nOut23_23[2] , \nScanOut602[4] , \nScanOut736[7] , \nScanOut885[5] , 
        \nScanOut362[5] , \nScanOut136[3] , \nScanOut456[2] , \nScanOut562[1] , 
        \nOut30_8[3] , \nScanOut255[5] , \nScanOut361[6] , \nScanOut135[0] , 
        \nScanOut601[7] , \nScanOut886[6] , \nScanOut735[4] , \nScanOut287[3] , 
        \nScanOut455[1] , \nScanOut561[2] , \nScanOut854[0] , \nOut30_27[2] , 
        \nScanOut81[2] , \nScanOut232[2] , \nOut10_14[0] , \nOut19_24[1] , 
        \nOut23_20[1] , \nScanOut960[3] , \nScanOut487[7] , \nScanOut1024[6] , 
        \nScanOut306[1] , \nScanOut666[0] , \nScanOut752[3] , \nScanOut50[7] , 
        \nScanOut53[4] , \nOut2_28[3] , \nScanOut152[7] , \nOut29_26[5] , 
        \nOut13_22[5] , \nScanOut432[6] , \nScanOut506[5] , \nOut25_29[0] , 
        \nOut20_16[4] , \nScanOut780[5] , \nScanOut833[7] , \nScanOut180[1] , 
        \nOut7_17[7] , \nScanOut907[4] , \nOut7_14[4] , \nScanOut830[4] , 
        \nScanOut783[6] , \nScanOut904[7] , \nScanOut82[1] , \nScanOut183[2] , 
        \nScanOut665[3] , \nScanOut751[0] , \nScanOut231[1] , \nScanOut305[2] , 
        \nOut13_21[6] , \nScanOut431[5] , \nScanOut505[6] , \nOut20_15[7] , 
        \nOut29_25[6] , \nScanOut8[0] , \nScanOut10[5] , \nScanOut74[1] , 
        \nScanOut151[4] , \nScanOut693[3] , \nScanOut814[2] , \nScanOut77[2] , 
        \nOut6_11[4] , \nScanOut920[1] , \nOut6_12[7] , \nScanOut175[2] , 
        \nOut7_30[2] , \nOut28_20[6] , \nScanOut176[1] , \nScanOut215[7] , 
        \nOut12_24[6] , \nScanOut415[3] , \nScanOut521[0] , \nOut21_10[7] , 
        \nOut20_31[1] , \nScanOut321[4] , \nOut12_27[5] , \nScanOut416[0] , 
        \nScanOut522[3] , \nScanOut641[5] , \nScanOut775[6] , \nOut21_13[4] , 
        \nOut25_9[6] , \nOut17_18[1] , \nOut28_23[5] , \nScanOut216[4] , 
        \nScanOut642[6] , \nScanOut776[5] , \nScanOut322[7] , \nOut23_9[2] , 
        \nScanOut690[0] , \nScanOut817[1] , \nOut29_8[7] , \nScanOut923[2] , 
        \nScanOut111[6] , \nScanOut471[7] , \nScanOut545[4] , \nOut5_24[2] , 
        \nScanOut271[3] , \nScanOut625[1] , \nScanOut711[2] , \nScanOut996[3] , 
        \nScanOut345[0] , \nOut10_30[6] , \nOut11_11[0] , \nScanOut597[2] , 
        \nOut18_21[1] , \nScanOut1000[0] , \nOut22_25[1] , \nScanOut870[6] , 
        \nScanOut944[5] , \nScanOut13[6] , \nOut1_8[2] , \nOut7_8[6] , 
        \nScanOut397[6] , \nOut31_22[2] , \nOut14_8[3] , \nOut18_22[2] , 
        \nOut22_26[2] , \nOut11_12[3] , \nScanOut594[1] , \nOut27_19[6] , 
        \nScanOut1003[3] , \nOut12_8[7] , \nScanOut394[5] , \nScanOut873[5] , 
        \nOut31_21[1] , \nOut0_15[0] , \nOut0_18[5] , \nScanOut112[5] , 
        \nScanOut947[6] , \nOut5_27[1] , \nScanOut272[0] , \nScanOut472[4] , 
        \nScanOut546[7] , \nOut9_28[4] , \nScanOut346[3] , \nOut18_9[2] , 
        \nOut1_5[7] , \nOut2_14[7] , \nOut16_21[5] , \nScanOut626[2] , 
        \nScanOut712[1] , \nScanOut995[0] , \nScanOut688[2] , \nOut25_15[4] , 
        \nOut2_17[4] , \nOut1_21[1] , \nOut7_28[0] , \nScanOut938[3] , 
        \nOut8_11[0] , \nOut9_30[6] , \nScanOut339[6] , \nOut16_22[6] , 
        \nScanOut539[2] , \nOut25_16[7] , \nOut29_19[2] , \nOut20_29[3] , 
        \nOut15_14[3] , \nScanOut659[7] , \nOut26_20[2] , \nOut30_18[5] , 
        \nOut1_22[2] , \nScanOut109[4] , \nScanOut469[5] , \nOut31_3[7] , 
        \nOut7_5[3] , \nOut8_12[3] , \nScanOut269[1] , \nScanOut709[0] , 
        \nOut10_28[4] , \nOut26_23[1] , \nOut15_17[0] , \nScanOut1018[2] , 
        \nOut19_18[5] , \nOut27_14[3] , \nScanOut868[4] , \nOut12_5[2] , 
        \nOut14_5[6] , \nScanOut599[4] , \nOut14_20[2] , \nScanOut399[0] , 
        \nOut20_0[6] , \nOut0_16[3] , \nOut5_29[7] , \nOut9_25[1] , 
        \nOut26_0[2] , \nScanOut998[5] , \nScanOut348[5] , \nScanOut548[1] , 
        \nOut18_4[7] , \nOut20_3[5] , \nOut9_26[2] , \nOut18_7[4] , 
        \nScanOut628[4] , \nScanOut21[4] , \nScanOut22[7] , \nOut2_1[6] , 
        \nOut1_6[4] , \nOut7_6[0] , \nOut14_6[5] , \nOut26_3[1] , 
        \nOut14_23[1] , \nOut22_28[4] , \nOut27_17[0] , \nOut8_0[3] , 
        \nOut12_6[1] , \nScanOut949[0] , \nOut24_21[5] , \nOut17_15[4] , 
        \nOut25_4[3] , \nOut23_4[7] , \nOut2_2[5] , \nOut3_20[6] , 
        \nOut11_1[3] , \nOut17_1[7] , \nOut4_1[2] , \nOut29_5[2] , 
        \nOut11_2[0] , \nScanOut45[0] , \nScanOut46[3] , \nOut2_19[2] , 
        \nScanOut61[6] , \nScanOut79[4] , \nOut4_2[1] , \nOut29_6[1] , 
        \nScanOut819[7] , \nOut3_23[5] , \nScanOut104[1] , \nScanOut178[7] , 
        \nOut8_3[0] , \nScanOut418[6] , \nOut17_2[4] , \nOut17_16[7] , 
        \nOut25_7[0] , \nScanOut218[2] , \nOut12_29[3] , \nOut23_7[4] , 
        \nOut24_22[6] , \nScanOut778[3] , \nOut4_10[3] , \nScanOut264[4] , 
        \nScanOut464[0] , \nScanOut550[3] , \nScanOut107[2] , \nOut5_31[5] , 
        \nScanOut350[7] , \nOut10_25[1] , \nOut19_15[0] , \nScanOut630[6] , 
        \nOut22_30[6] , \nScanOut704[5] , \nScanOut983[4] , \nOut23_11[0] , 
        \nOut10_26[2] , \nScanOut382[1] , \nScanOut582[5] , \nScanOut1015[7] , 
        \nScanOut581[6] , \nScanOut865[1] , \nOut30_16[3] , \nScanOut951[2] , 
        \nScanOut381[2] , \nOut15_19[6] , \nOut19_16[3] , \nScanOut1016[4] , 
        \nOut23_12[3] , \nScanOut866[2] , \nOut30_15[0] , \nScanOut952[1] , 
        \nScanOut467[3] , \nScanOut553[0] , \nOut4_13[0] , \nScanOut267[7] , 
        \nScanOut633[5] , \nScanOut707[6] , \nScanOut980[7] , \nOut7_25[5] , 
        \nScanOut353[4] , \nScanOut686[4] , \nScanOut801[5] , \nScanOut935[6] , 
        \nScanOut160[5] , \nOut13_10[7] , \nScanOut400[4] , \nScanOut534[7] , 
        \nOut20_24[6] , \nOut12_31[1] , \nOut29_14[7] , \nScanOut163[6] , 
        \nScanOut200[0] , \nScanOut654[2] , \nScanOut760[1] , \nScanOut334[3] , 
        \nOut29_17[4] , \nScanOut203[3] , \nOut13_13[4] , \nOut25_18[1] , 
        \nScanOut403[7] , \nScanOut537[4] , \nOut20_27[5] , \nScanOut337[0] , 
        \nScanOut657[1] , \nScanOut763[2] , \nScanOut62[5] , \nScanOut685[7] , 
        \nScanOut802[6] , \nScanOut94[5] , \nOut7_26[6] , \nScanOut936[5] , 
        \nScanOut673[7] , \nScanOut747[4] , \nScanOut147[0] , \nScanOut227[5] , 
        \nOut9_8[4] , \nScanOut313[6] , \nOut12_16[4] , \nScanOut427[1] , 
        \nScanOut513[2] , \nOut17_29[0] , \nOut21_22[5] , \nOut6_23[6] , 
        \nScanOut826[0] , \nOut28_12[4] , \nScanOut912[3] , \nScanOut795[2] , 
        \nOut3_9[1] , \nOut5_9[5] , \nScanOut195[6] , \nOut10_9[4] , 
        \nOut16_9[0] , \nScanOut796[1] , \nScanOut825[3] , \nScanOut97[6] , 
        \nOut6_20[5] , \nScanOut911[0] , \nScanOut196[5] , \nScanOut224[6] , 
        \nScanOut310[5] , \nScanOut670[4] , \nScanOut744[7] , \nScanOut144[3] , 
        \nOut29_30[1] , \nScanOut291[7] , \nOut12_15[7] , \nOut28_11[7] , 
        \nScanOut424[2] , \nScanOut510[1] , \nOut21_21[6] , \nScanOut842[4] , 
        \nOut31_10[0] , \nOut30_31[6] , \nOut0_29[4] , \nOut5_16[0] , 
        \nScanOut243[1] , \nOut11_23[2] , \nOut18_13[3] , \nOut22_17[3] , 
        \nScanOut976[7] , \nOut27_28[7] , \nScanOut491[3] , \nOut9_19[5] , 
        \nScanOut377[2] , \nOut27_8[5] , \nScanOut120[7] , \nScanOut123[4] , 
        \nScanOut617[3] , \nScanOut890[2] , \nScanOut723[0] , \nOut5_15[3] , 
        \nScanOut240[2] , \nScanOut443[5] , \nScanOut577[6] , \nOut21_8[1] , 
        \nScanOut614[0] , \nScanOut720[3] , \nScanOut893[1] , \nScanOut374[1] , 
        \nScanOut440[6] , \nScanOut574[5] , \nScanOut841[7] , \nScanOut975[4] , 
        \nOut2_26[5] , \nScanOut292[4] , \nOut11_20[1] , \nOut31_13[3] , 
        \nScanOut492[0] , \nOut18_10[0] , \nOut19_31[6] , \nOut22_14[0] , 
        \nOut7_19[1] , \nScanOut308[7] , \nScanOut909[2] , \nScanOut668[6] , 
        \nOut25_27[6] , \nScanOut39[6] , \nOut1_13[3] , \nOut2_25[6] , 
        \nOut16_10[4] , \nOut16_13[7] , \nScanOut508[3] , \nOut29_28[3] , 
        \nOut20_18[2] , \nOut17_31[2] , \nOut25_24[5] , \nScanOut138[5] , 
        \nOut8_23[2] , \nScanOut258[0] , \nScanOut738[1] , \nScanOut458[4] , 
        \nScanOut859[5] , \nOut30_6[5] , \nOut10_19[5] , \nOut15_26[1] , 
        \nOut26_12[0] , \nOut8_20[1] , \nScanOut289[5] , \nOut19_29[4] , 
        \nOut15_25[2] , \nOut30_29[4] , \nScanOut489[1] , \nOut26_11[3] , 
        \nOut27_30[5] , \nOut1_10[0] , \nScanOut888[0] , \nOut30_5[6] , 
        \nOut0_10[4] , \nOut0_13[7] , \nScanOut18[4] , \nOut1_3[0] , 
        \nOut2_4[2] , \nOut2_7[1] , \nOut3_26[1] , \nOut4_7[5] , \nOut8_6[4] , 
        \nScanOut329[5] , \nScanOut649[4] , \nOut23_2[0] , \nScanOut529[1] , 
        \nOut17_13[3] , \nOut25_2[4] , \nOut21_18[6] , \nOut24_27[2] , 
        \nOut28_28[7] , \nOut29_3[5] , \nOut6_19[5] , \nScanOut928[0] , 
        \nOut17_7[0] , \nOut11_7[4] , \nOut3_25[2] , \nOut4_4[6] , 
        \nOut17_4[3] , \nScanOut698[1] , \nOut29_0[6] , \nOut8_5[7] , 
        \nOut11_4[7] , \nOut17_10[0] , \nOut16_31[6] , \nOut23_1[3] , 
        \nOut24_24[1] , \nOut25_1[7] , \nScanOut878[7] , \nOut7_3[4] , 
        \nOut12_3[5] , \nOut14_3[1] , \nOut14_26[5] , \nOut18_29[0] , 
        \nOut27_12[4] , \nScanOut279[2] , \nOut11_19[1] , \nScanOut1008[1] , 
        \nOut9_23[6] , \nOut18_2[0] , \nOut1_31[2] , \nScanOut119[7] , 
        \nScanOut719[3] , \nOut26_6[5] , \nScanOut479[6] , \nOut20_6[1] , 
        \nScanOut24[0] , \nOut1_0[3] , \nOut9_20[5] , \nOut26_5[6] , 
        \nOut12_0[6] , \nOut18_1[3] , \nOut20_5[2] , \nOut31_29[0] , 
        \nOut1_29[0] , \nScanOut64[2] , \nScanOut67[1] , \nOut7_23[2] , 
        \nOut7_0[7] , \nOut14_25[6] , \nOut14_0[2] , \nOut26_30[1] , 
        \nOut27_11[7] , \nScanOut680[3] , \nScanOut807[2] , \nScanOut933[1] , 
        \nScanOut165[1] , \nScanOut166[2] , \nScanOut206[7] , \nScanOut332[4] , 
        \nOut13_16[0] , \nScanOut652[5] , \nScanOut766[6] , \nOut29_12[0] , 
        \nScanOut205[4] , \nScanOut406[3] , \nOut16_29[4] , \nScanOut532[0] , 
        \nOut20_22[1] , \nScanOut651[6] , \nScanOut765[5] , \nScanOut331[7] , 
        \nScanOut405[0] , \nScanOut531[3] , \nOut20_21[2] , \nOut28_30[5] , 
        \nOut29_11[3] , \nOut13_15[3] , \nScanOut683[0] , \nScanOut804[1] , 
        \nOut7_20[1] , \nScanOut930[2] , \nScanOut101[5] , \nScanOut102[6] , 
        \nOut4_16[4] , \nOut8_19[1] , \nScanOut262[3] , \nScanOut636[1] , 
        \nScanOut702[2] , \nScanOut985[3] , \nScanOut356[0] , \nScanOut462[7] , 
        \nScanOut556[4] , \nOut4_15[7] , \nScanOut261[0] , \nOut10_20[5] , 
        \nOut10_23[6] , \nScanOut384[6] , \nScanOut863[6] , \nOut31_8[5] , 
        \nScanOut957[5] , \nOut30_10[4] , \nScanOut387[5] , \nScanOut584[2] , 
        \nOut19_13[7] , \nOut23_17[7] , \nOut26_28[3] , \nScanOut1013[0] , 
        \nOut30_13[7] , \nOut19_10[4] , \nScanOut860[5] , \nScanOut954[6] , 
        \nScanOut587[1] , \nOut18_31[2] , \nOut23_14[4] , \nScanOut1010[3] , 
        \nScanOut355[3] , \nScanOut635[2] , \nScanOut701[1] , \nScanOut986[0] , 
        \nOut11_25[5] , \nScanOut461[4] , \nScanOut555[7] , \nScanOut497[4] , 
        \nOut18_15[4] , \nOut22_11[4] , \nOut23_30[2] , \nScanOut844[3] , 
        \nScanOut125[3] , \nScanOut297[0] , \nScanOut970[0] , \nScanOut445[2] , 
        \nScanOut571[1] , \nOut31_16[7] , \nScanOut126[0] , \nOut5_10[7] , 
        \nScanOut245[6] , \nScanOut611[4] , \nScanOut896[5] , \nScanOut725[7] , 
        \nScanOut371[5] , \nOut4_31[1] , \nOut5_13[4] , \nScanOut246[5] , 
        \nScanOut446[1] , \nScanOut572[2] , \nScanOut372[6] , \nOut19_9[4] , 
        \nOut11_26[6] , \nOut14_19[2] , \nOut15_8[5] , \nOut18_16[7] , 
        \nScanOut612[7] , \nScanOut726[4] , \nScanOut895[6] , \nOut22_12[7] , 
        \nOut0_8[4] , \nOut6_8[0] , \nScanOut494[7] , \nScanOut27[3] , 
        \nScanOut294[3] , \nOut13_8[1] , \nScanOut847[0] , \nOut31_15[4] , 
        \nScanOut973[3] , \nScanOut40[4] , \nScanOut92[2] , \nScanOut141[7] , 
        \nOut12_10[3] , \nOut13_31[5] , \nScanOut221[2] , \nScanOut421[6] , 
        \nScanOut515[5] , \nOut28_14[3] , \nOut21_24[2] , \nScanOut315[1] , 
        \nScanOut675[0] , \nScanOut741[3] , \nOut6_25[1] , \nScanOut193[1] , 
        \nScanOut820[7] , \nScanOut914[4] , \nScanOut793[5] , \nScanOut43[7] , 
        \nScanOut190[2] , \nScanOut790[6] , \nScanOut823[4] , \nOut3_19[6] , 
        \nOut6_26[2] , \nOut28_8[1] , \nScanOut917[7] , \nScanOut0[1] , 
        \nOut0_5[1] , \nOut0_21[5] , \nOut1_15[4] , \nScanOut91[1] , 
        \nScanOut142[4] , \nScanOut422[5] , \nScanOut516[6] , \nOut21_27[1] , 
        \nOut24_9[0] , \nOut12_13[0] , \nOut28_17[0] , \nScanOut676[3] , 
        \nOut24_18[5] , \nScanOut742[0] , \nScanOut222[1] , \nOut8_25[5] , 
        \nScanOut316[2] , \nOut22_9[4] , \nOut30_0[2] , \nOut1_16[7] , 
        \nOut15_20[6] , \nOut15_23[5] , \nOut26_14[7] , \nOut26_17[4] , 
        \nScanOut569[3] , \nOut23_28[0] , \nScanOut968[2] , \nScanOut609[6] , 
        \nOut30_3[1] , \nOut2_20[2] , \nOut4_29[3] , \nScanOut369[7] , 
        \nScanOut188[0] , \nOut8_26[6] , \nScanOut788[4] , \nOut2_23[1] , 
        \nScanOut89[3] , \nOut16_15[0] , \nOut25_21[1] , \nScanOut159[5] , 
        \nScanOut239[0] , \nOut13_29[7] , \nOut25_22[2] , \nScanOut439[4] , 
        \nOut16_16[3] , \nScanOut759[1] , \nScanOut58[6] , \nScanOut838[5] , 
        \nOut3_1[0] , \nOut3_2[3] , \nOut3_14[3] , \nOut10_1[5] , \nOut5_1[4] , 
        \nOut16_1[1] , \nOut28_5[4] , \nOut9_3[6] , \nOut9_0[5] , 
        \nOut24_15[0] , \nOut17_21[1] , \nOut24_4[5] , \nOut22_4[1] , 
        \nOut10_2[6] , \nScanOut318[4] , \nScanOut518[0] , \nOut24_7[6] , 
        \nOut17_22[2] , \nOut21_29[7] , \nScanOut678[5] , \nOut24_16[3] , 
        \nOut28_19[6] , \nOut22_7[2] , \nOut3_17[0] , \nOut5_2[7] , 
        \nOut6_28[4] , \nScanOut919[1] , \nOut28_6[7] , \nOut16_2[2] , 
        \nOut21_0[0] , \nOut27_0[4] , \nOut6_5[5] , \nOut8_30[2] , 
        \nOut19_4[1] , \nScanOut898[3] , \nOut9_11[4] , \nOut27_20[6] , 
        \nOut13_5[4] , \nOut14_14[7] , \nOut15_5[0] , \nScanOut499[2] , 
        \nOut0_6[2] , \nOut6_6[6] , \nScanOut299[6] , \nOut11_28[0] , 
        \nOut14_17[4] , \nOut31_18[1] , \nOut15_6[3] , \nOut18_18[1] , 
        \nOut27_23[5] , \nOut0_22[6] , \nScanOut29[5] , \nOut13_6[7] , 
        \nScanOut849[6] , \nScanOut128[6] , \nScanOut248[3] , \nScanOut448[7] , 
        \nOut21_3[3] , \nOut19_7[2] , \nOut9_12[7] , \nScanOut434[1] , 
        \nScanOut500[2] , \nScanOut728[2] , \nOut27_3[7] , \nOut21_31[5] , 
        \nOut20_10[3] , \nScanOut3[2] , \nScanOut55[3] , \nScanOut87[5] , 
        \nScanOut154[0] , \nOut29_20[2] , \nOut13_24[2] , \nScanOut660[7] , 
        \nScanOut754[4] , \nScanOut186[6] , \nScanOut234[5] , \nScanOut300[6] , 
        \nScanOut786[2] , \nScanOut835[0] , \nScanOut56[0] , \nScanOut185[5] , 
        \nOut6_30[6] , \nOut7_11[0] , \nScanOut901[3] , \nOut7_12[3] , 
        \nScanOut836[3] , \nScanOut785[1] , \nScanOut902[0] , \nOut13_27[1] , 
        \nOut29_23[1] , \nScanOut15[1] , \nScanOut16[2] , \nScanOut31[7] , 
        \nScanOut84[6] , \nScanOut157[3] , \nScanOut237[6] , \nScanOut437[2] , 
        \nScanOut503[1] , \nOut16_18[5] , \nOut20_13[0] , \nScanOut303[5] , 
        \nScanOut663[4] , \nScanOut757[7] , \nScanOut282[7] , \nOut10_11[4] , 
        \nOut19_21[5] , \nOut23_25[5] , \nOut11_30[2] , \nScanOut482[3] , 
        \nScanOut1021[2] , \nScanOut851[4] , \nOut30_22[6] , \nScanOut965[7] , 
        \nScanOut32[4] , \nOut1_18[1] , \nOut4_24[6] , \nScanOut130[4] , 
        \nScanOut250[1] , \nScanOut450[5] , \nScanOut564[6] , \nScanOut364[2] , 
        \nScanOut133[7] , \nScanOut453[6] , \nScanOut567[5] , \nScanOut604[3] , 
        \nScanOut730[0] , \nScanOut883[2] , \nOut4_27[5] , \nOut8_28[0] , 
        \nScanOut253[2] , \nScanOut607[0] , \nScanOut880[1] , \nScanOut733[3] , 
        \nScanOut367[1] , \nOut10_12[7] , \nOut26_19[2] , \nScanOut481[0] , 
        \nScanOut1022[1] , \nOut19_22[6] , \nOut23_26[6] , \nScanOut852[7] , 
        \nScanOut117[1] , \nOut5_22[5] , \nScanOut277[4] , \nScanOut281[4] , 
        \nScanOut966[4] , \nOut30_21[5] , \nScanOut343[7] , \nOut20_8[7] , 
        \nScanOut623[6] , \nScanOut717[5] , \nOut26_8[3] , \nScanOut990[4] , 
        \nScanOut391[1] , \nScanOut477[0] , \nScanOut543[3] , \nOut31_24[5] , 
        \nScanOut876[1] , \nScanOut942[2] , \nOut11_17[7] , \nOut14_28[3] , 
        \nOut18_27[6] , \nOut22_23[6] , \nScanOut591[5] , \nScanOut875[2] , 
        \nScanOut1006[7] , \nOut2_9[7] , \nScanOut72[6] , \nOut4_9[3] , 
        \nScanOut114[2] , \nOut5_21[6] , \nScanOut274[7] , \nOut11_14[4] , 
        \nScanOut392[2] , \nScanOut941[1] , \nOut31_27[6] , \nOut18_24[5] , 
        \nScanOut592[6] , \nOut22_20[5] , \nScanOut1005[4] , \nScanOut620[5] , 
        \nScanOut714[6] , \nScanOut993[7] , \nScanOut340[4] , \nScanOut474[3] , 
        \nScanOut540[0] , \nScanOut695[4] , \nScanOut812[5] , \nOut3_28[7] , 
        \nOut6_17[3] , \nScanOut926[6] , \nOut17_9[6] , \nOut11_9[2] , 
        \nOut2_12[0] , \nOut1_24[5] , \nOut1_27[6] , \nScanOut71[5] , 
        \nScanOut170[6] , \nScanOut173[5] , \nScanOut213[0] , \nScanOut647[2] , 
        \nScanOut773[1] , \nOut8_8[2] , \nScanOut327[3] , \nScanOut413[4] , 
        \nScanOut527[7] , \nOut21_16[0] , \nOut28_26[1] , \nScanOut210[3] , 
        \nOut12_22[1] , \nOut24_29[4] , \nScanOut324[0] , \nOut12_21[2] , 
        \nScanOut644[1] , \nScanOut770[2] , \nOut28_25[2] , \nOut6_14[0] , 
        \nScanOut410[7] , \nScanOut524[4] , \nOut21_15[3] , \nScanOut696[7] , 
        \nScanOut811[6] , \nScanOut925[5] , \nOut15_12[4] , \nOut23_19[1] , 
        \nOut26_26[5] , \nScanOut959[3] , \nScanOut638[7] , \nOut4_18[2] , 
        \nOut8_14[4] , \nOut8_17[7] , \nScanOut358[6] , \nScanOut558[2] , 
        \nOut31_6[3] , \nScanOut168[4] , \nScanOut208[1] , \nScanOut389[3] , 
        \nOut31_5[0] , \nScanOut988[6] , \nOut14_30[1] , \nOut15_11[7] , 
        \nScanOut589[7] , \nOut26_25[6] , \nScanOut768[0] , \nOut13_18[6] , 
        \nScanOut408[5] , \nOut16_27[2] , \nOut25_13[3] , \nScanOut69[7] , 
        \nScanOut809[4] , \nScanOut5[4] , \nScanOut34[2] , \nOut2_11[3] , 
        \nOut3_30[5] , \nOut4_21[3] , \nScanOut135[1] , \nScanOut455[0] , 
        \nOut16_24[1] , \nScanOut561[3] , \nOut25_10[0] , \nOut24_31[6] , 
        \nScanOut255[4] , \nScanOut601[6] , \nScanOut735[5] , \nScanOut886[7] , 
        \nScanOut361[7] , \nOut10_14[1] , \nScanOut487[6] , \nOut19_24[0] , 
        \nScanOut1024[7] , \nOut23_20[0] , \nScanOut854[1] , \nScanOut960[2] , 
        \nScanOut37[1] , \nScanOut284[1] , \nScanOut287[2] , \nOut10_17[2] , 
        \nOut15_28[6] , \nOut30_27[3] , \nOut19_27[3] , \nOut23_23[3] , 
        \nScanOut484[5] , \nScanOut857[2] , \nOut30_24[0] , \nScanOut50[6] , 
        \nOut4_22[0] , \nScanOut136[2] , \nScanOut963[1] , \nScanOut256[7] , 
        \nScanOut456[3] , \nScanOut562[0] , \nOut30_8[2] , \nScanOut362[4] , 
        \nScanOut183[3] , \nScanOut602[5] , \nScanOut885[4] , \nScanOut736[6] , 
        \nScanOut783[7] , \nScanOut830[5] , \nScanOut151[5] , \nOut7_14[5] , 
        \nScanOut904[6] , \nScanOut6[7] , \nScanOut82[0] , \nScanOut231[0] , 
        \nOut13_21[7] , \nOut29_25[7] , \nScanOut431[4] , \nScanOut505[7] , 
        \nOut20_15[6] , \nScanOut305[3] , \nScanOut665[2] , \nScanOut751[1] , 
        \nScanOut152[6] , \nOut13_22[4] , \nScanOut432[7] , \nScanOut506[4] , 
        \nOut20_16[5] , \nOut25_29[1] , \nOut29_26[4] , \nScanOut53[5] , 
        \nScanOut81[3] , \nScanOut666[1] , \nScanOut752[2] , \nScanOut180[0] , 
        \nScanOut232[3] , \nScanOut306[0] , \nOut7_17[6] , \nScanOut833[6] , 
        \nScanOut780[4] , \nScanOut907[5] , \nOut2_28[2] , \nOut6_0[0] , 
        \nOut14_11[2] , \nOut15_30[4] , \nOut15_0[5] , \nOut27_25[3] , 
        \nOut0_3[7] , \nOut0_24[0] , \nOut9_14[1] , \nOut13_0[1] , 
        \nOut19_1[4] , \nOut21_5[5] , \nOut27_5[1] , \nOut0_27[3] , 
        \nScanOut579[1] , \nOut21_6[6] , \nOut5_18[7] , \nOut9_17[2] , 
        \nOut19_2[7] , \nScanOut619[4] , \nOut27_6[2] , \nOut6_3[3] , 
        \nScanOut379[5] , \nOut27_26[0] , \nOut13_3[2] , \nOut14_12[1] , 
        \nOut22_19[4] , \nOut15_3[6] , \nScanOut978[0] , \nScanOut8[1] , 
        \nScanOut10[4] , \nScanOut13[7] , \nOut2_14[6] , \nScanOut48[4] , 
        \nOut2_30[0] , \nOut3_4[5] , \nScanOut99[1] , \nOut9_5[0] , 
        \nOut24_1[0] , \nOut17_24[4] , \nOut24_10[5] , \nOut25_31[3] , 
        \nScanOut198[2] , \nOut10_4[0] , \nOut22_1[4] , \nOut5_4[1] , 
        \nScanOut798[6] , \nOut28_0[1] , \nOut3_7[6] , \nOut3_11[6] , 
        \nOut16_4[4] , \nOut3_12[5] , \nOut10_7[3] , \nOut5_7[2] , 
        \nOut16_7[7] , \nScanOut828[7] , \nOut2_17[5] , \nScanOut149[7] , 
        \nOut12_18[3] , \nOut28_3[2] , \nOut24_13[6] , \nOut7_28[1] , 
        \nScanOut229[2] , \nOut9_6[3] , \nOut24_2[3] , \nScanOut429[6] , 
        \nOut17_27[7] , \nOut22_2[7] , \nScanOut749[3] , \nScanOut938[2] , 
        \nScanOut339[7] , \nScanOut659[6] , \nOut16_21[4] , \nOut16_22[7] , 
        \nScanOut539[3] , \nOut20_29[2] , \nOut25_15[5] , \nOut25_16[6] , 
        \nOut29_19[3] , \nOut1_21[0] , \nOut1_22[3] , \nOut8_12[2] , 
        \nScanOut269[0] , \nScanOut688[3] , \nScanOut109[5] , \nScanOut709[1] , 
        \nOut10_28[5] , \nOut15_17[1] , \nScanOut469[4] , \nOut31_3[6] , 
        \nOut19_18[4] , \nScanOut868[5] , \nOut15_14[2] , \nOut26_20[3] , 
        \nOut26_23[0] , \nOut30_18[4] , \nScanOut1018[3] , \nScanOut74[0] , 
        \nScanOut77[3] , \nScanOut176[0] , \nScanOut216[5] , \nOut8_11[1] , 
        \nOut9_30[7] , \nOut23_9[3] , \nScanOut322[6] , \nScanOut642[7] , 
        \nScanOut776[4] , \nOut28_23[4] , \nOut12_27[4] , \nScanOut416[1] , 
        \nScanOut522[2] , \nOut17_18[0] , \nOut21_13[5] , \nScanOut690[1] , 
        \nOut25_9[7] , \nScanOut817[0] , \nOut29_8[6] , \nOut6_11[5] , 
        \nOut6_12[6] , \nScanOut693[2] , \nScanOut814[3] , \nScanOut923[3] , 
        \nOut7_30[3] , \nScanOut920[0] , \nScanOut175[3] , \nScanOut215[6] , 
        \nScanOut641[4] , \nScanOut775[7] , \nScanOut321[5] , \nOut12_24[7] , 
        \nScanOut415[2] , \nScanOut521[1] , \nOut20_31[0] , \nOut21_10[6] , 
        \nOut28_20[7] , \nScanOut873[4] , \nScanOut947[7] , \nOut0_18[4] , 
        \nOut1_8[3] , \nOut12_8[6] , \nOut31_21[0] , \nOut7_8[7] , 
        \nOut11_12[2] , \nScanOut394[4] , \nOut27_19[7] , \nOut14_8[2] , 
        \nScanOut594[0] , \nScanOut1003[2] , \nOut18_22[3] , \nScanOut626[3] , 
        \nOut22_26[3] , \nScanOut111[7] , \nScanOut112[4] , \nOut5_27[0] , 
        \nScanOut272[1] , \nScanOut712[0] , \nScanOut995[1] , \nOut9_28[5] , 
        \nScanOut346[2] , \nScanOut472[5] , \nScanOut546[6] , \nOut18_9[3] , 
        \nOut5_24[3] , \nScanOut271[2] , \nScanOut345[1] , \nScanOut625[0] , 
        \nScanOut711[3] , \nScanOut996[2] , \nScanOut397[7] , \nScanOut471[6] , 
        \nScanOut545[5] , \nScanOut870[7] , \nOut31_22[3] , \nOut0_15[1] , 
        \nOut0_16[2] , \nOut2_19[3] , \nScanOut62[4] , \nScanOut104[0] , 
        \nOut4_10[2] , \nScanOut107[3] , \nOut4_13[1] , \nScanOut267[6] , 
        \nOut10_26[3] , \nOut10_30[7] , \nOut11_11[1] , \nOut18_21[0] , 
        \nOut22_25[0] , \nScanOut944[4] , \nScanOut381[3] , \nScanOut597[3] , 
        \nScanOut1000[1] , \nOut15_19[7] , \nOut23_12[2] , \nScanOut866[3] , 
        \nOut30_15[1] , \nScanOut952[0] , \nOut19_16[2] , \nScanOut581[7] , 
        \nScanOut1016[5] , \nScanOut353[5] , \nScanOut633[4] , 
        \nScanOut707[7] , \nScanOut980[6] , \nScanOut264[5] , \nScanOut467[2] , 
        \nScanOut553[1] , \nScanOut630[7] , \nScanOut704[4] , \nScanOut983[5] , 
        \nOut5_31[4] , \nScanOut350[6] , \nScanOut464[1] , \nScanOut550[2] , 
        \nScanOut163[7] , \nScanOut203[2] , \nOut10_25[0] , \nScanOut382[0] , 
        \nScanOut865[0] , \nOut30_16[2] , \nScanOut951[3] , \nScanOut582[4] , 
        \nOut19_15[1] , \nScanOut1015[6] , \nScanOut657[0] , \nOut22_30[7] , 
        \nOut23_11[1] , \nScanOut763[3] , \nScanOut337[1] , \nOut13_13[5] , 
        \nScanOut403[6] , \nScanOut537[5] , \nOut20_27[4] , \nOut25_18[0] , 
        \nOut7_26[7] , \nScanOut685[6] , \nScanOut802[7] , \nOut29_17[5] , 
        \nScanOut936[4] , \nScanOut61[7] , \nScanOut686[5] , \nScanOut801[4] , 
        \nScanOut160[4] , \nScanOut200[1] , \nOut7_25[4] , \nScanOut935[7] , 
        \nScanOut334[2] , \nScanOut654[3] , \nScanOut760[0] , \nOut13_10[6] , 
        \nOut29_14[6] , \nScanOut400[5] , \nOut12_31[0] , \nScanOut534[6] , 
        \nOut20_24[7] , \nOut1_5[6] , \nOut1_6[5] , \nOut5_29[6] , 
        \nOut9_26[3] , \nScanOut628[5] , \nOut26_3[0] , \nOut18_7[5] , 
        \nScanOut348[4] , \nOut12_6[0] , \nScanOut548[0] , \nOut20_3[4] , 
        \nScanOut949[1] , \nOut7_6[1] , \nOut27_17[1] , \nOut14_6[4] , 
        \nOut14_23[0] , \nOut22_28[5] , \nOut7_5[2] , \nOut12_5[3] , 
        \nScanOut399[1] , \nOut14_5[7] , \nOut14_20[3] , \nOut9_25[0] , 
        \nScanOut599[5] , \nOut27_14[2] , \nOut18_4[6] , \nOut2_1[7] , 
        \nOut2_2[4] , \nScanOut79[5] , \nOut3_23[4] , \nOut17_2[5] , 
        \nOut20_0[7] , \nOut26_0[3] , \nScanOut998[4] , \nOut4_2[0] , 
        \nScanOut819[6] , \nOut29_6[0] , \nOut3_20[7] , \nOut4_1[3] , 
        \nScanOut178[6] , \nScanOut218[3] , \nOut11_2[1] , \nOut12_29[2] , 
        \nOut23_7[5] , \nOut24_22[7] , \nScanOut778[2] , \nOut8_3[1] , 
        \nOut25_7[1] , \nOut8_0[2] , \nScanOut418[7] , \nOut17_16[6] , 
        \nOut17_15[5] , \nOut23_4[6] , \nOut25_4[2] , \nOut24_21[4] , 
        \nOut29_5[3] , \nOut11_1[2] , \nOut17_1[6] , \nOut2_25[7] , 
        \nOut16_10[5] , \nOut17_31[3] , \nOut25_24[4] , \nOut2_26[4] , 
        \nOut7_19[0] , \nScanOut909[3] , \nOut16_13[6] , \nScanOut508[2] , 
        \nOut20_18[3] , \nOut29_28[2] , \nScanOut289[4] , \nScanOut308[6] , 
        \nScanOut668[7] , \nOut25_27[7] , \nOut15_25[3] , \nScanOut489[0] , 
        \nOut26_11[2] , \nOut27_30[4] , \nOut30_29[5] , \nOut30_5[7] , 
        \nOut1_10[1] , \nScanOut888[1] , \nOut1_13[2] , \nScanOut138[4] , 
        \nOut8_20[0] , \nOut30_6[4] , \nOut8_23[3] , \nScanOut258[1] , 
        \nScanOut458[5] , \nOut15_26[0] , \nOut19_29[5] , \nScanOut738[0] , 
        \nOut0_8[5] , \nOut0_10[5] , \nScanOut21[5] , \nScanOut39[7] , 
        \nOut10_19[4] , \nOut26_12[1] , \nScanOut859[4] , \nScanOut45[1] , 
        \nOut6_20[4] , \nScanOut196[4] , \nScanOut825[2] , \nScanOut796[0] , 
        \nScanOut911[1] , \nScanOut46[2] , \nOut3_9[0] , \nScanOut94[4] , 
        \nScanOut97[7] , \nScanOut144[2] , \nOut12_15[6] , \nScanOut424[3] , 
        \nScanOut510[0] , \nOut21_21[7] , \nScanOut670[5] , \nOut28_11[6] , 
        \nOut29_30[0] , \nScanOut744[6] , \nScanOut147[1] , \nScanOut224[7] , 
        \nScanOut310[4] , \nScanOut227[4] , \nOut9_8[5] , \nOut12_16[5] , 
        \nOut28_12[5] , \nScanOut513[3] , \nScanOut427[0] , \nOut17_29[1] , 
        \nOut21_22[4] , \nScanOut313[7] , \nScanOut673[6] , \nScanOut747[5] , 
        \nScanOut195[7] , \nOut5_9[4] , \nOut10_9[5] , \nOut16_9[1] , 
        \nScanOut795[3] , \nScanOut826[1] , \nScanOut120[6] , \nOut6_23[7] , 
        \nScanOut912[2] , \nOut5_15[2] , \nScanOut240[3] , \nScanOut440[7] , 
        \nScanOut574[4] , \nScanOut292[5] , \nOut11_20[0] , \nScanOut374[0] , 
        \nOut18_10[1] , \nScanOut614[1] , \nScanOut893[0] , \nOut22_14[1] , 
        \nScanOut720[2] , \nOut19_31[7] , \nScanOut492[1] , \nScanOut841[6] , 
        \nOut31_13[2] , \nScanOut22[6] , \nOut11_23[3] , \nScanOut975[5] , 
        \nScanOut491[2] , \nOut27_28[6] , \nOut18_13[2] , \nOut22_17[2] , 
        \nScanOut842[5] , \nScanOut976[6] , \nOut0_29[5] , \nScanOut123[5] , 
        \nScanOut291[6] , \nScanOut443[4] , \nScanOut577[7] , \nOut31_10[1] , 
        \nOut30_31[7] , \nScanOut617[2] , \nOut21_8[0] , \nOut2_4[3] , 
        \nOut1_29[1] , \nScanOut64[3] , \nOut5_16[1] , \nScanOut243[0] , 
        \nScanOut723[1] , \nOut27_8[4] , \nScanOut890[3] , \nScanOut165[0] , 
        \nOut9_19[4] , \nScanOut377[3] , \nOut13_15[2] , \nOut28_30[4] , 
        \nScanOut205[5] , \nScanOut405[1] , \nScanOut531[2] , \nOut29_11[2] , 
        \nOut20_21[3] , \nOut7_20[0] , \nScanOut331[6] , \nScanOut651[7] , 
        \nScanOut683[1] , \nScanOut765[4] , \nScanOut804[0] , \nScanOut930[3] , 
        \nScanOut67[0] , \nScanOut680[2] , \nScanOut807[3] , \nScanOut101[4] , 
        \nScanOut166[3] , \nOut7_23[3] , \nScanOut933[0] , \nScanOut406[2] , 
        \nOut16_29[5] , \nScanOut532[1] , \nOut20_22[0] , \nScanOut206[6] , 
        \nOut13_16[1] , \nOut29_12[1] , \nScanOut652[4] , \nScanOut766[7] , 
        \nOut10_20[4] , \nScanOut332[5] , \nScanOut387[4] , \nOut19_10[5] , 
        \nScanOut587[0] , \nOut23_14[5] , \nScanOut1010[2] , \nOut18_31[3] , 
        \nScanOut860[4] , \nScanOut954[7] , \nScanOut461[5] , \nScanOut555[6] , 
        \nOut30_13[6] , \nScanOut102[7] , \nOut4_15[6] , \nScanOut261[1] , 
        \nScanOut635[3] , \nScanOut701[0] , \nScanOut986[1] , \nScanOut355[2] , 
        \nOut4_16[5] , \nScanOut262[2] , \nScanOut462[6] , \nScanOut556[5] , 
        \nOut31_8[4] , \nOut8_19[0] , \nScanOut356[1] , \nScanOut636[0] , 
        \nOut10_23[7] , \nScanOut584[3] , \nOut19_13[6] , \nScanOut702[3] , 
        \nScanOut985[2] , \nOut23_17[6] , \nOut26_28[2] , \nOut11_4[6] , 
        \nScanOut384[7] , \nOut30_10[5] , \nScanOut1013[1] , \nScanOut863[7] , 
        \nScanOut957[4] , \nOut2_7[0] , \nOut3_25[3] , \nOut4_4[7] , 
        \nScanOut698[0] , \nOut17_4[2] , \nOut29_0[7] , \nOut8_5[6] , 
        \nOut25_1[6] , \nOut8_6[5] , \nOut17_10[1] , \nOut16_31[7] , 
        \nOut17_13[2] , \nScanOut529[0] , \nOut23_1[2] , \nOut24_24[0] , 
        \nOut24_27[3] , \nOut28_28[6] , \nOut21_18[7] , \nOut25_2[5] , 
        \nScanOut329[4] , \nOut23_2[1] , \nScanOut649[5] , \nOut1_31[3] , 
        \nOut3_26[0] , \nOut11_7[5] , \nOut4_7[4] , \nOut17_7[1] , 
        \nOut6_19[4] , \nOut29_3[4] , \nOut9_20[4] , \nOut20_5[3] , 
        \nScanOut928[1] , \nOut18_1[2] , \nOut0_13[6] , \nScanOut18[5] , 
        \nOut1_0[2] , \nOut7_0[6] , \nOut14_25[7] , \nOut14_0[3] , 
        \nOut26_5[7] , \nOut27_11[6] , \nOut26_30[0] , \nOut7_3[5] , 
        \nOut11_19[0] , \nOut12_0[7] , \nOut31_29[1] , \nOut12_3[4] , 
        \nOut14_3[0] , \nOut27_12[5] , \nScanOut1008[0] , \nOut14_26[4] , 
        \nOut18_29[1] , \nScanOut878[6] , \nOut1_3[1] , \nScanOut119[6] , 
        \nScanOut479[7] , \nOut20_6[0] , \nScanOut27[2] , \nOut1_15[5] , 
        \nOut1_16[6] , \nOut4_29[2] , \nOut8_26[7] , \nScanOut279[3] , 
        \nScanOut719[2] , \nOut26_6[4] , \nOut9_23[7] , \nOut15_23[4] , 
        \nOut18_2[1] , \nOut23_28[1] , \nScanOut968[3] , \nOut26_17[5] , 
        \nScanOut369[6] , \nScanOut569[2] , \nScanOut609[7] , \nOut30_3[0] , 
        \nOut2_20[3] , \nOut2_23[0] , \nScanOut58[7] , \nScanOut159[4] , 
        \nScanOut239[1] , \nOut8_25[4] , \nOut15_20[7] , \nOut26_14[6] , 
        \nOut30_0[3] , \nScanOut759[0] , \nOut13_29[6] , \nScanOut439[5] , 
        \nOut16_16[2] , \nOut25_22[3] , \nScanOut838[4] , \nScanOut89[2] , 
        \nScanOut188[1] , \nScanOut788[5] , \nScanOut126[1] , \nOut5_13[5] , 
        \nScanOut246[4] , \nOut16_15[1] , \nOut25_21[0] , \nOut19_9[5] , 
        \nScanOut612[6] , \nScanOut895[7] , \nScanOut726[5] , \nScanOut372[7] , 
        \nScanOut446[0] , \nScanOut572[3] , \nOut13_8[0] , \nScanOut847[1] , 
        \nScanOut973[2] , \nScanOut294[2] , \nOut31_15[5] , \nScanOut24[1] , 
        \nOut6_8[1] , \nOut11_26[7] , \nScanOut297[1] , \nOut14_19[3] , 
        \nScanOut494[6] , \nOut15_8[4] , \nOut18_16[6] , \nOut22_12[6] , 
        \nScanOut844[2] , \nOut31_16[6] , \nScanOut970[1] , \nScanOut125[2] , 
        \nOut5_10[6] , \nScanOut245[7] , \nOut11_25[4] , \nOut18_15[5] , 
        \nOut22_11[5] , \nOut23_30[3] , \nScanOut497[5] , \nOut4_31[0] , 
        \nScanOut371[4] , \nScanOut611[5] , \nScanOut725[6] , \nScanOut896[4] , 
        \nOut3_19[7] , \nScanOut445[3] , \nScanOut571[0] , \nScanOut0[0] , 
        \nScanOut3[3] , \nScanOut40[5] , \nScanOut43[6] , \nOut6_26[3] , 
        \nScanOut823[5] , \nScanOut790[7] , \nScanOut917[6] , \nOut28_8[0] , 
        \nScanOut91[0] , \nScanOut190[3] , \nScanOut222[0] , \nScanOut316[3] , 
        \nScanOut676[2] , \nOut22_9[5] , \nScanOut742[1] , \nScanOut92[3] , 
        \nScanOut142[5] , \nOut12_13[1] , \nOut24_18[4] , \nScanOut422[4] , 
        \nScanOut516[7] , \nOut24_9[1] , \nOut28_17[1] , \nOut21_27[0] , 
        \nScanOut675[1] , \nScanOut741[2] , \nScanOut141[6] , \nScanOut221[3] , 
        \nScanOut315[0] , \nScanOut421[7] , \nScanOut515[4] , \nOut21_24[3] , 
        \nOut12_10[2] , \nOut28_14[2] , \nOut13_31[4] , \nScanOut793[4] , 
        \nScanOut820[6] , \nScanOut56[1] , \nOut6_25[0] , \nScanOut193[0] , 
        \nScanOut914[5] , \nScanOut785[0] , \nScanOut836[2] , \nScanOut84[7] , 
        \nScanOut185[4] , \nOut7_12[2] , \nScanOut902[1] , \nScanOut663[5] , 
        \nScanOut757[6] , \nScanOut157[2] , \nScanOut237[7] , \nScanOut303[4] , 
        \nScanOut437[3] , \nScanOut503[0] , \nOut16_18[4] , \nOut20_13[1] , 
        \nScanOut87[4] , \nScanOut234[4] , \nOut13_27[0] , \nOut29_23[0] , 
        \nScanOut300[7] , \nScanOut660[6] , \nScanOut754[5] , \nScanOut154[1] , 
        \nOut13_24[3] , \nOut29_20[3] , \nOut0_5[0] , \nOut0_6[3] , 
        \nScanOut29[4] , \nScanOut31[6] , \nScanOut32[5] , \nOut1_18[0] , 
        \nScanOut55[2] , \nOut6_30[7] , \nOut7_11[1] , \nScanOut434[0] , 
        \nScanOut500[3] , \nOut20_10[2] , \nOut21_31[4] , \nScanOut835[1] , 
        \nScanOut786[3] , \nScanOut901[2] , \nOut4_27[4] , \nScanOut186[7] , 
        \nScanOut253[3] , \nScanOut367[0] , \nOut8_28[1] , \nScanOut607[1] , 
        \nScanOut880[0] , \nScanOut133[6] , \nScanOut733[2] , \nScanOut281[5] , 
        \nScanOut453[7] , \nScanOut567[4] , \nScanOut852[6] , \nOut30_21[4] , 
        \nScanOut966[5] , \nOut10_12[6] , \nOut19_22[7] , \nOut23_26[7] , 
        \nScanOut481[1] , \nOut26_19[3] , \nScanOut851[5] , \nScanOut1022[0] , 
        \nOut3_1[1] , \nOut3_2[2] , \nOut3_17[1] , \nOut4_24[7] , 
        \nScanOut250[0] , \nScanOut282[6] , \nScanOut965[6] , \nOut10_11[5] , 
        \nOut30_22[7] , \nOut11_30[3] , \nScanOut482[2] , \nScanOut1021[3] , 
        \nOut19_21[4] , \nOut23_25[4] , \nScanOut604[2] , \nScanOut883[3] , 
        \nScanOut730[1] , \nScanOut364[3] , \nScanOut130[5] , \nScanOut450[4] , 
        \nScanOut564[7] , \nOut9_3[7] , \nScanOut318[5] , \nOut22_7[3] , 
        \nScanOut518[1] , \nScanOut678[4] , \nOut24_16[2] , \nOut28_19[7] , 
        \nOut24_7[7] , \nOut17_22[3] , \nOut21_29[6] , \nOut5_2[6] , 
        \nOut16_2[3] , \nOut6_28[5] , \nOut28_6[6] , \nScanOut919[0] , 
        \nOut3_14[2] , \nOut5_1[5] , \nOut10_2[7] , \nOut28_5[5] , 
        \nOut10_1[4] , \nOut16_1[0] , \nOut9_0[4] , \nOut22_4[0] , 
        \nOut24_4[4] , \nOut13_6[6] , \nOut17_21[0] , \nOut24_15[1] , 
        \nScanOut849[7] , \nOut0_21[4] , \nOut0_22[7] , \nOut6_6[7] , 
        \nOut11_28[1] , \nOut27_23[4] , \nOut14_17[5] , \nOut15_6[2] , 
        \nOut18_18[0] , \nOut27_3[6] , \nScanOut128[7] , \nScanOut248[2] , 
        \nScanOut728[3] , \nOut9_12[6] , \nOut19_7[3] , \nScanOut448[6] , 
        \nOut8_30[3] , \nOut19_4[0] , \nOut21_3[2] , \nOut9_11[5] , 
        \nOut21_0[1] , \nOut27_0[5] , \nScanOut898[2] , \nOut2_11[2] , 
        \nOut1_24[4] , \nOut6_5[4] , \nScanOut299[7] , \nOut13_5[5] , 
        \nOut31_18[0] , \nOut14_14[6] , \nOut15_5[1] , \nOut27_20[7] , 
        \nScanOut499[3] , \nOut31_5[1] , \nOut1_27[7] , \nOut4_18[3] , 
        \nOut8_14[5] , \nScanOut988[7] , \nOut8_17[6] , \nScanOut389[2] , 
        \nOut14_30[0] , \nScanOut589[6] , \nOut26_25[7] , \nOut15_11[6] , 
        \nOut15_12[5] , \nScanOut558[3] , \nOut23_19[0] , \nOut26_26[4] , 
        \nScanOut959[2] , \nOut31_6[2] , \nScanOut358[7] , \nOut3_30[4] , 
        \nScanOut638[6] , \nScanOut8[5] , \nScanOut15[0] , \nOut2_12[1] , 
        \nScanOut69[6] , \nScanOut168[5] , \nOut13_18[7] , \nScanOut408[4] , 
        \nOut16_24[0] , \nOut25_10[1] , \nOut24_31[7] , \nOut16_27[3] , 
        \nOut25_13[2] , \nScanOut208[0] , \nScanOut768[1] , \nScanOut809[5] , 
        \nOut11_14[5] , \nOut18_24[4] , \nOut22_20[4] , \nScanOut392[3] , 
        \nScanOut592[7] , \nOut31_27[7] , \nScanOut1005[5] , \nScanOut875[3] , 
        \nScanOut941[0] , \nScanOut16[3] , \nScanOut114[3] , \nScanOut117[0] , 
        \nOut5_21[7] , \nScanOut274[6] , \nScanOut474[2] , \nScanOut540[1] , 
        \nScanOut340[5] , \nScanOut477[1] , \nScanOut543[2] , \nScanOut620[4] , 
        \nScanOut714[7] , \nScanOut993[6] , \nOut5_22[4] , \nScanOut277[5] , 
        \nOut20_8[6] , \nScanOut623[7] , \nScanOut717[4] , \nOut26_8[2] , 
        \nScanOut990[5] , \nOut11_17[6] , \nScanOut343[6] , \nOut14_28[2] , 
        \nScanOut591[4] , \nOut22_23[7] , \nScanOut1006[6] , \nOut18_27[7] , 
        \nScanOut876[0] , \nScanOut21[1] , \nScanOut22[2] , \nOut0_29[1] , 
        \nOut2_9[6] , \nScanOut71[4] , \nScanOut170[7] , \nScanOut391[0] , 
        \nScanOut942[3] , \nScanOut410[6] , \nScanOut524[5] , \nOut31_24[4] , 
        \nOut21_15[2] , \nOut28_25[3] , \nScanOut210[2] , \nOut12_21[3] , 
        \nScanOut644[0] , \nScanOut770[3] , \nScanOut324[1] , \nScanOut696[6] , 
        \nScanOut811[7] , \nOut6_14[1] , \nScanOut925[4] , \nScanOut45[5] , 
        \nScanOut46[6] , \nScanOut72[7] , \nOut3_28[6] , \nOut11_9[3] , 
        \nOut4_9[2] , \nOut17_9[7] , \nScanOut695[5] , \nScanOut812[4] , 
        \nOut6_17[2] , \nScanOut926[7] , \nOut5_9[0] , \nScanOut173[4] , 
        \nOut12_22[0] , \nOut24_29[5] , \nOut28_26[0] , \nScanOut213[1] , 
        \nOut8_8[3] , \nScanOut527[6] , \nScanOut413[5] , \nOut21_16[1] , 
        \nScanOut327[2] , \nScanOut647[3] , \nScanOut773[0] , \nScanOut795[7] , 
        \nScanOut826[5] , \nOut3_9[4] , \nOut6_23[3] , \nScanOut195[3] , 
        \nOut10_9[1] , \nOut16_9[5] , \nScanOut912[6] , \nScanOut94[0] , 
        \nScanOut673[2] , \nScanOut747[1] , \nScanOut97[3] , \nScanOut147[5] , 
        \nScanOut227[0] , \nOut9_8[1] , \nScanOut313[3] , \nScanOut513[7] , 
        \nScanOut427[4] , \nOut17_29[5] , \nOut21_22[0] , \nScanOut224[3] , 
        \nOut12_16[1] , \nOut28_12[1] , \nScanOut310[0] , \nScanOut670[1] , 
        \nScanOut744[2] , \nScanOut144[6] , \nOut12_15[2] , \nOut6_20[0] , 
        \nScanOut424[7] , \nScanOut510[4] , \nOut28_11[2] , \nOut29_30[4] , 
        \nOut21_21[3] , \nScanOut825[6] , \nScanOut796[4] , \nScanOut911[5] , 
        \nOut5_16[5] , \nScanOut196[0] , \nScanOut243[4] , \nOut9_19[0] , 
        \nScanOut377[7] , \nScanOut617[6] , \nOut27_8[0] , \nScanOut123[1] , 
        \nScanOut723[5] , \nScanOut890[7] , \nScanOut291[2] , \nScanOut443[0] , 
        \nScanOut577[3] , \nOut21_8[4] , \nScanOut842[1] , \nOut31_10[5] , 
        \nOut30_31[3] , \nScanOut976[2] , \nOut11_23[7] , \nOut18_13[6] , 
        \nOut22_17[6] , \nOut27_28[2] , \nScanOut491[6] , \nScanOut841[2] , 
        \nScanOut120[2] , \nOut5_15[6] , \nScanOut240[7] , \nScanOut292[1] , 
        \nScanOut975[1] , \nOut11_20[4] , \nOut31_13[6] , \nScanOut492[5] , 
        \nOut18_10[5] , \nOut22_14[5] , \nScanOut614[5] , \nOut19_31[3] , 
        \nScanOut893[4] , \nScanOut720[6] , \nScanOut374[4] , \nScanOut440[3] , 
        \nScanOut574[0] , \nScanOut308[2] , \nScanOut668[3] , \nScanOut39[3] , 
        \nOut2_25[3] , \nOut2_26[0] , \nOut16_13[2] , \nScanOut508[6] , 
        \nOut25_27[3] , \nOut29_28[6] , \nOut20_18[7] , \nOut7_19[4] , 
        \nScanOut909[7] , \nOut16_10[1] , \nOut17_31[7] , \nOut25_24[0] , 
        \nScanOut859[0] , \nOut10_19[0] , \nOut15_26[4] , \nOut19_29[1] , 
        \nOut26_12[5] , \nOut0_15[5] , \nOut1_13[6] , \nScanOut138[0] , 
        \nOut8_23[7] , \nScanOut258[5] , \nScanOut738[4] , \nScanOut458[1] , 
        \nOut30_6[0] , \nOut8_20[4] , \nOut1_10[5] , \nScanOut888[5] , 
        \nScanOut289[0] , \nOut30_5[3] , \nOut15_25[7] , \nOut30_29[1] , 
        \nScanOut489[4] , \nOut26_11[6] , \nOut27_30[0] , \nOut20_0[3] , 
        \nOut0_16[6] , \nOut1_5[2] , \nOut7_5[6] , \nOut9_25[4] , 
        \nOut26_0[7] , \nScanOut998[0] , \nOut18_4[2] , \nOut27_14[6] , 
        \nOut12_5[7] , \nOut14_5[3] , \nScanOut599[1] , \nOut14_20[7] , 
        \nOut1_6[1] , \nOut7_6[5] , \nScanOut399[5] , \nOut14_6[0] , 
        \nOut14_23[4] , \nOut22_28[1] , \nOut27_17[5] , \nOut5_29[2] , 
        \nOut9_26[7] , \nOut12_6[4] , \nScanOut548[4] , \nOut20_3[0] , 
        \nScanOut949[5] , \nOut18_7[1] , \nScanOut348[0] , \nOut2_1[3] , 
        \nScanOut628[1] , \nOut26_3[4] , \nOut2_2[0] , \nOut3_20[3] , 
        \nOut11_1[6] , \nOut17_1[2] , \nOut4_1[7] , \nScanOut178[2] , 
        \nOut8_3[5] , \nOut8_0[6] , \nOut17_15[1] , \nOut24_21[0] , 
        \nOut29_5[7] , \nOut25_4[6] , \nOut23_4[2] , \nOut25_7[5] , 
        \nOut12_29[6] , \nScanOut418[3] , \nOut17_16[2] , \nOut24_22[3] , 
        \nScanOut218[7] , \nScanOut778[6] , \nOut11_2[5] , \nOut23_7[1] , 
        \nOut2_19[7] , \nScanOut61[3] , \nScanOut79[1] , \nOut4_2[4] , 
        \nScanOut819[2] , \nOut29_6[4] , \nOut3_23[0] , \nScanOut104[4] , 
        \nOut10_25[4] , \nOut17_2[1] , \nOut19_15[5] , \nOut22_30[3] , 
        \nOut23_11[5] , \nScanOut382[4] , \nScanOut582[0] , \nOut30_16[6] , 
        \nScanOut1015[2] , \nScanOut865[4] , \nScanOut951[7] , \nOut4_10[6] , 
        \nScanOut264[1] , \nScanOut464[5] , \nScanOut550[6] , \nScanOut107[7] , 
        \nOut5_31[0] , \nScanOut350[2] , \nScanOut467[6] , \nScanOut553[5] , 
        \nScanOut630[3] , \nScanOut704[0] , \nScanOut983[1] , \nOut4_13[5] , 
        \nScanOut267[2] , \nScanOut633[0] , \nScanOut707[3] , \nScanOut980[2] , 
        \nScanOut160[0] , \nOut10_26[7] , \nScanOut353[1] , \nScanOut581[3] , 
        \nScanOut381[7] , \nOut15_19[3] , \nScanOut1016[1] , \nOut19_16[6] , 
        \nOut23_12[6] , \nScanOut866[7] , \nScanOut952[4] , \nScanOut400[1] , 
        \nScanOut534[2] , \nOut30_15[5] , \nOut20_24[3] , \nScanOut200[5] , 
        \nOut13_10[2] , \nOut29_14[2] , \nOut12_31[4] , \nScanOut654[7] , 
        \nScanOut760[4] , \nScanOut334[6] , \nScanOut686[1] , \nScanOut801[0] , 
        \nOut7_25[0] , \nScanOut935[3] , \nScanOut62[0] , \nOut7_26[3] , 
        \nScanOut685[2] , \nScanOut802[3] , \nScanOut936[0] , \nScanOut74[4] , 
        \nScanOut163[3] , \nOut13_13[1] , \nOut25_18[4] , \nOut6_11[1] , 
        \nScanOut175[7] , \nScanOut203[6] , \nScanOut403[2] , \nScanOut537[1] , 
        \nOut29_17[1] , \nOut20_27[0] , \nScanOut337[5] , \nOut12_24[3] , 
        \nScanOut657[4] , \nScanOut763[7] , \nOut28_20[3] , \nScanOut215[2] , 
        \nScanOut415[6] , \nScanOut521[5] , \nOut20_31[4] , \nOut21_10[2] , 
        \nScanOut321[1] , \nScanOut641[0] , \nScanOut693[6] , \nScanOut775[3] , 
        \nScanOut814[7] , \nOut7_30[7] , \nScanOut920[4] , \nScanOut77[7] , 
        \nScanOut690[5] , \nScanOut817[4] , \nOut29_8[2] , \nOut6_12[2] , 
        \nScanOut176[4] , \nScanOut416[5] , \nScanOut522[6] , \nScanOut923[7] , 
        \nOut17_18[4] , \nOut21_13[1] , \nOut25_9[3] , \nOut28_23[0] , 
        \nOut12_27[0] , \nScanOut642[3] , \nOut23_9[7] , \nScanOut776[0] , 
        \nOut0_3[3] , \nScanOut10[0] , \nScanOut216[1] , \nOut10_30[3] , 
        \nScanOut322[2] , \nOut11_11[5] , \nScanOut597[7] , \nOut18_21[4] , 
        \nOut22_25[4] , \nScanOut1000[5] , \nScanOut870[3] , \nScanOut13[3] , 
        \nOut0_18[0] , \nScanOut111[3] , \nScanOut397[3] , \nScanOut944[0] , 
        \nScanOut471[2] , \nScanOut545[1] , \nOut31_22[7] , \nScanOut112[0] , 
        \nOut5_24[7] , \nScanOut271[6] , \nScanOut625[4] , \nScanOut711[7] , 
        \nScanOut996[6] , \nScanOut345[5] , \nOut5_27[4] , \nScanOut272[5] , 
        \nScanOut472[1] , \nScanOut546[2] , \nOut9_28[1] , \nScanOut346[6] , 
        \nOut18_9[7] , \nScanOut626[7] , \nOut1_8[7] , \nOut7_8[3] , 
        \nOut11_12[6] , \nOut14_8[6] , \nScanOut712[4] , \nScanOut995[5] , 
        \nOut18_22[7] , \nOut22_26[7] , \nScanOut594[4] , \nOut27_19[3] , 
        \nOut31_21[4] , \nScanOut1003[6] , \nOut12_8[2] , \nScanOut394[0] , 
        \nScanOut873[0] , \nScanOut947[3] , \nOut2_14[2] , \nScanOut688[7] , 
        \nOut2_17[1] , \nScanOut339[3] , \nOut16_21[0] , \nOut16_22[3] , 
        \nScanOut539[7] , \nOut25_15[1] , \nOut25_16[2] , \nOut29_19[7] , 
        \nOut20_29[6] , \nScanOut659[2] , \nOut1_21[4] , \nOut7_28[5] , 
        \nScanOut938[6] , \nOut8_11[5] , \nOut9_30[3] , \nOut1_22[7] , 
        \nScanOut109[1] , \nOut10_28[1] , \nOut15_14[6] , \nOut26_20[7] , 
        \nOut26_23[4] , \nOut30_18[0] , \nOut15_17[5] , \nOut19_18[0] , 
        \nScanOut1018[7] , \nScanOut469[0] , \nScanOut868[1] , \nOut31_3[2] , 
        \nOut8_12[6] , \nScanOut269[4] , \nScanOut709[5] , \nOut0_24[4] , 
        \nOut0_27[7] , \nOut5_18[3] , \nOut6_3[7] , \nOut13_3[6] , 
        \nOut14_12[5] , \nScanOut978[4] , \nOut15_3[2] , \nOut22_19[0] , 
        \nOut27_26[4] , \nOut9_17[6] , \nOut19_2[3] , \nScanOut379[1] , 
        \nOut27_6[6] , \nScanOut579[5] , \nScanOut619[0] , \nOut21_6[2] , 
        \nOut9_14[5] , \nOut19_1[0] , \nOut27_5[5] , \nOut13_0[5] , 
        \nOut21_5[1] , \nScanOut5[0] , \nScanOut6[3] , \nScanOut34[6] , 
        \nScanOut37[5] , \nScanOut48[0] , \nOut5_7[6] , \nScanOut149[3] , 
        \nOut6_0[4] , \nOut27_25[7] , \nScanOut229[6] , \nOut14_11[6] , 
        \nOut15_30[0] , \nOut15_0[1] , \nScanOut749[7] , \nOut9_6[7] , 
        \nOut22_2[3] , \nOut24_2[7] , \nOut12_18[7] , \nScanOut429[2] , 
        \nOut17_27[3] , \nOut24_13[2] , \nScanOut828[3] , \nOut28_3[6] , 
        \nOut2_30[4] , \nOut3_7[2] , \nOut3_12[1] , \nOut10_7[7] , 
        \nOut16_7[3] , \nOut3_4[1] , \nOut3_11[2] , \nOut5_4[5] , 
        \nOut16_4[0] , \nScanOut798[2] , \nScanOut198[6] , \nOut28_0[5] , 
        \nScanOut99[5] , \nOut10_4[4] , \nOut22_1[0] , \nOut4_22[4] , 
        \nScanOut256[3] , \nOut9_5[4] , \nOut24_1[4] , \nOut24_10[1] , 
        \nOut25_31[7] , \nOut17_24[0] , \nScanOut602[1] , \nScanOut885[0] , 
        \nScanOut736[2] , \nScanOut362[0] , \nScanOut136[6] , \nScanOut456[7] , 
        \nScanOut562[4] , \nScanOut857[6] , \nOut30_8[6] , \nScanOut284[5] , 
        \nScanOut963[5] , \nScanOut287[6] , \nOut10_17[6] , \nOut30_24[4] , 
        \nOut15_28[2] , \nScanOut484[1] , \nOut23_23[7] , \nOut19_27[7] , 
        \nScanOut854[5] , \nOut30_27[7] , \nScanOut960[6] , \nScanOut53[1] , 
        \nOut2_28[6] , \nOut4_21[7] , \nScanOut255[0] , \nOut10_14[5] , 
        \nOut19_24[4] , \nOut23_20[4] , \nScanOut487[2] , \nScanOut1024[3] , 
        \nScanOut361[3] , \nScanOut135[5] , \nScanOut601[2] , \nScanOut735[1] , 
        \nScanOut886[3] , \nScanOut455[4] , \nScanOut561[7] , \nOut7_17[2] , 
        \nScanOut833[2] , \nScanOut780[0] , \nScanOut907[1] , \nScanOut81[7] , 
        \nScanOut180[4] , \nScanOut232[7] , \nScanOut306[4] , \nScanOut666[5] , 
        \nScanOut752[6] , \nScanOut152[2] , \nOut13_22[0] , \nOut25_29[5] , 
        \nScanOut82[4] , \nScanOut432[3] , \nScanOut506[0] , \nOut29_26[0] , 
        \nOut20_16[1] , \nScanOut665[6] , \nScanOut751[5] , \nScanOut151[1] , 
        \nScanOut231[4] , \nScanOut305[7] , \nScanOut431[0] , \nScanOut505[3] , 
        \nOut20_15[2] , \nOut29_25[3] , \nScanOut15[4] , \nScanOut16[7] , 
        \nScanOut50[2] , \nOut13_21[3] , \nScanOut783[3] , \nScanOut830[1] , 
        \nScanOut183[7] , \nOut7_14[1] , \nScanOut904[2] , \nScanOut391[4] , 
        \nScanOut876[4] , \nOut31_24[0] , \nScanOut114[7] , \nScanOut117[4] , 
        \nOut5_22[0] , \nScanOut277[1] , \nOut11_17[2] , \nOut14_28[6] , 
        \nScanOut942[7] , \nOut18_27[3] , \nOut22_23[3] , \nScanOut591[0] , 
        \nScanOut1006[2] , \nScanOut343[2] , \nScanOut623[3] , 
        \nScanOut717[0] , \nOut26_8[6] , \nScanOut990[1] , \nOut5_21[3] , 
        \nScanOut274[2] , \nScanOut477[5] , \nScanOut543[6] , \nOut20_8[2] , 
        \nScanOut620[0] , \nScanOut714[3] , \nScanOut993[2] , \nScanOut340[1] , 
        \nScanOut474[6] , \nScanOut540[5] , \nScanOut875[7] , \nScanOut941[4] , 
        \nOut2_9[2] , \nScanOut72[3] , \nOut4_9[6] , \nScanOut173[0] , 
        \nScanOut213[5] , \nOut11_14[1] , \nScanOut392[7] , \nOut31_27[3] , 
        \nOut18_24[0] , \nScanOut592[3] , \nScanOut1005[1] , \nScanOut647[7] , 
        \nOut22_20[0] , \nScanOut773[4] , \nOut8_8[7] , \nScanOut327[6] , 
        \nScanOut527[2] , \nOut12_22[4] , \nScanOut413[1] , \nOut21_16[5] , 
        \nOut24_29[1] , \nOut28_26[4] , \nScanOut695[1] , \nScanOut812[0] , 
        \nOut6_17[6] , \nScanOut926[3] , \nOut3_28[2] , \nOut17_9[3] , 
        \nOut11_9[7] , \nOut2_11[6] , \nOut2_12[5] , \nOut1_24[0] , 
        \nOut1_27[3] , \nScanOut71[0] , \nScanOut696[2] , \nScanOut811[3] , 
        \nScanOut170[3] , \nOut6_14[5] , \nScanOut210[6] , \nScanOut925[0] , 
        \nScanOut324[5] , \nScanOut644[4] , \nScanOut770[7] , \nOut28_25[7] , 
        \nOut12_21[7] , \nScanOut410[2] , \nScanOut524[1] , \nOut21_15[6] , 
        \nOut4_18[7] , \nOut8_17[2] , \nScanOut638[2] , \nOut8_14[1] , 
        \nScanOut358[3] , \nScanOut389[6] , \nOut15_12[1] , \nScanOut558[7] , 
        \nOut23_19[4] , \nOut26_26[0] , \nScanOut959[6] , \nOut31_6[6] , 
        \nOut14_30[4] , \nOut15_11[2] , \nScanOut589[2] , \nOut26_25[3] , 
        \nOut31_5[5] , \nScanOut988[3] , \nScanOut69[2] , \nScanOut809[1] , 
        \nOut3_30[0] , \nScanOut168[1] , \nScanOut208[4] , \nOut13_18[3] , 
        \nScanOut768[5] , \nOut25_13[6] , \nScanOut408[0] , \nOut16_27[7] , 
        \nOut16_24[4] , \nOut25_10[5] , \nOut24_31[3] , \nScanOut0[4] , 
        \nOut0_5[4] , \nOut3_1[5] , \nOut9_0[0] , \nOut24_4[0] , 
        \nOut24_15[5] , \nOut17_21[4] , \nOut22_4[4] , \nOut3_2[6] , 
        \nOut3_14[6] , \nOut10_1[0] , \nOut5_1[1] , \nOut16_1[4] , 
        \nOut10_2[3] , \nOut28_5[1] , \nOut3_17[5] , \nOut5_2[2] , 
        \nOut6_28[1] , \nOut28_6[2] , \nScanOut919[4] , \nOut6_5[0] , 
        \nOut9_3[3] , \nOut16_2[7] , \nScanOut518[5] , \nOut24_7[3] , 
        \nScanOut318[1] , \nOut17_22[7] , \nOut21_29[2] , \nScanOut678[0] , 
        \nOut24_16[6] , \nOut28_19[3] , \nOut22_7[7] , \nOut27_20[3] , 
        \nOut13_5[1] , \nOut14_14[2] , \nScanOut499[7] , \nOut15_5[5] , 
        \nOut0_6[7] , \nOut0_21[0] , \nScanOut299[3] , \nOut21_0[5] , 
        \nOut31_18[4] , \nOut27_0[1] , \nOut0_22[3] , \nScanOut128[3] , 
        \nOut8_30[7] , \nOut19_4[4] , \nScanOut898[6] , \nOut9_11[1] , 
        \nScanOut248[6] , \nScanOut448[2] , \nOut21_3[6] , \nOut9_12[2] , 
        \nOut19_7[7] , \nOut6_6[3] , \nOut11_28[5] , \nOut14_17[1] , 
        \nOut15_6[6] , \nOut18_18[4] , \nScanOut728[7] , \nOut27_3[2] , 
        \nOut27_23[0] , \nScanOut29[0] , \nOut13_6[2] , \nScanOut849[3] , 
        \nScanOut55[6] , \nScanOut186[3] , \nOut6_30[3] , \nOut7_11[5] , 
        \nScanOut835[5] , \nScanOut786[7] , \nScanOut901[6] , \nScanOut154[5] , 
        \nOut13_24[7] , \nScanOut434[4] , \nScanOut500[7] , \nOut20_10[6] , 
        \nOut21_31[0] , \nScanOut3[7] , \nScanOut87[0] , \nScanOut660[2] , 
        \nOut29_20[7] , \nScanOut754[1] , \nScanOut157[6] , \nScanOut234[0] , 
        \nScanOut300[3] , \nOut29_23[4] , \nScanOut24[5] , \nScanOut31[2] , 
        \nScanOut56[5] , \nScanOut84[3] , \nScanOut237[3] , \nOut13_27[4] , 
        \nScanOut437[7] , \nScanOut503[4] , \nOut16_18[0] , \nOut20_13[5] , 
        \nScanOut303[0] , \nScanOut663[1] , \nScanOut757[2] , \nScanOut185[0] , 
        \nScanOut785[4] , \nScanOut836[6] , \nOut4_24[3] , \nScanOut130[1] , 
        \nOut7_12[6] , \nScanOut902[5] , \nScanOut250[4] , \nScanOut450[0] , 
        \nScanOut564[3] , \nScanOut364[7] , \nScanOut282[2] , \nOut10_11[1] , 
        \nOut19_21[0] , \nScanOut604[6] , \nScanOut883[7] , \nOut23_25[0] , 
        \nScanOut730[5] , \nOut11_30[7] , \nScanOut482[6] , \nScanOut1021[7] , 
        \nScanOut851[1] , \nOut30_22[3] , \nScanOut32[1] , \nOut10_12[2] , 
        \nOut26_19[7] , \nScanOut965[2] , \nScanOut481[5] , \nOut19_22[3] , 
        \nScanOut1022[4] , \nOut23_26[3] , \nScanOut852[2] , \nScanOut966[1] , 
        \nOut1_18[4] , \nScanOut133[2] , \nScanOut281[1] , \nScanOut453[3] , 
        \nScanOut567[0] , \nOut30_21[0] , \nScanOut607[5] , \nScanOut880[4] , 
        \nOut4_27[0] , \nScanOut253[7] , \nScanOut733[6] , \nScanOut367[4] , 
        \nScanOut125[6] , \nOut8_28[5] , \nScanOut445[7] , \nScanOut571[4] , 
        \nOut5_10[2] , \nScanOut245[3] , \nScanOut611[1] , \nScanOut725[2] , 
        \nScanOut896[0] , \nOut4_31[4] , \nScanOut371[0] , \nOut11_25[0] , 
        \nScanOut497[1] , \nOut18_15[1] , \nOut22_11[1] , \nOut23_30[7] , 
        \nScanOut844[6] , \nScanOut970[5] , \nScanOut297[5] , \nOut14_19[7] , 
        \nOut22_12[2] , \nOut31_16[2] , \nOut15_8[0] , \nOut18_16[2] , 
        \nOut0_8[1] , \nOut6_8[5] , \nOut11_26[3] , \nScanOut494[2] , 
        \nScanOut27[6] , \nScanOut294[6] , \nOut13_8[4] , \nOut31_15[1] , 
        \nScanOut847[5] , \nScanOut40[1] , \nScanOut126[5] , \nScanOut973[6] , 
        \nOut5_13[1] , \nScanOut246[0] , \nScanOut446[4] , \nScanOut572[7] , 
        \nOut19_9[1] , \nScanOut193[4] , \nScanOut372[3] , \nScanOut612[2] , 
        \nScanOut895[3] , \nScanOut726[1] , \nScanOut793[0] , \nScanOut820[2] , 
        \nScanOut43[2] , \nScanOut91[4] , \nScanOut92[7] , \nScanOut141[2] , 
        \nOut6_25[4] , \nScanOut914[1] , \nScanOut221[7] , \nOut12_10[6] , 
        \nOut28_14[6] , \nScanOut421[3] , \nOut13_31[0] , \nScanOut515[0] , 
        \nOut21_24[7] , \nScanOut315[4] , \nScanOut675[5] , \nScanOut741[6] , 
        \nScanOut142[1] , \nOut12_13[5] , \nScanOut422[0] , \nScanOut516[3] , 
        \nOut24_9[5] , \nOut21_27[4] , \nOut24_18[0] , \nScanOut676[6] , 
        \nOut28_17[5] , \nScanOut742[5] , \nOut6_26[7] , \nScanOut190[7] , 
        \nScanOut222[4] , \nScanOut316[7] , \nOut22_9[1] , \nScanOut823[1] , 
        \nScanOut790[3] , \nScanOut917[2] , \nOut3_19[3] , \nOut28_8[4] , 
        \nOut0_8[3] , \nOut0_10[1] , \nOut0_13[2] , \nOut2_4[7] , \nOut2_7[4] , 
        \nOut1_15[1] , \nOut8_25[0] , \nOut15_20[3] , \nOut26_14[2] , 
        \nOut30_0[7] , \nOut1_16[2] , \nScanOut569[6] , \nOut30_3[4] , 
        \nOut2_20[7] , \nScanOut89[6] , \nOut4_29[6] , \nOut8_26[3] , 
        \nScanOut609[3] , \nScanOut369[2] , \nOut15_23[0] , \nOut26_17[1] , 
        \nOut16_15[5] , \nOut23_28[5] , \nScanOut968[7] , \nOut25_21[4] , 
        \nScanOut188[5] , \nScanOut788[1] , \nOut2_23[4] , \nScanOut58[3] , 
        \nScanOut838[0] , \nOut3_26[4] , \nOut4_7[0] , \nScanOut159[0] , 
        \nOut13_29[2] , \nOut25_22[7] , \nScanOut239[5] , \nScanOut439[1] , 
        \nOut16_16[6] , \nScanOut759[4] , \nOut6_19[0] , \nOut29_3[0] , 
        \nOut17_7[5] , \nScanOut928[5] , \nOut11_7[1] , \nOut3_25[7] , 
        \nOut8_5[2] , \nOut8_6[1] , \nScanOut329[0] , \nScanOut649[1] , 
        \nOut23_2[5] , \nOut17_13[6] , \nScanOut529[4] , \nOut21_18[3] , 
        \nOut25_2[1] , \nOut23_1[6] , \nOut24_27[7] , \nOut28_28[2] , 
        \nOut24_24[4] , \nOut25_1[2] , \nOut17_10[5] , \nOut16_31[3] , 
        \nOut4_4[3] , \nOut17_4[6] , \nScanOut698[4] , \nOut29_0[3] , 
        \nScanOut279[7] , \nOut11_4[2] , \nOut9_23[3] , \nOut18_2[5] , 
        \nScanOut18[1] , \nOut1_3[5] , \nScanOut119[2] , \nOut20_6[4] , 
        \nScanOut719[6] , \nOut26_6[0] , \nScanOut479[3] , \nScanOut878[2] , 
        \nOut1_0[6] , \nOut7_3[1] , \nOut11_19[4] , \nOut12_3[0] , 
        \nOut14_3[4] , \nOut14_26[0] , \nOut18_29[5] , \nOut27_12[1] , 
        \nOut12_0[3] , \nScanOut1008[4] , \nOut1_31[7] , \nOut7_0[2] , 
        \nOut31_29[5] , \nOut14_25[3] , \nOut14_0[7] , \nOut26_30[4] , 
        \nOut27_11[2] , \nOut1_29[5] , \nScanOut64[7] , \nScanOut67[4] , 
        \nScanOut166[7] , \nScanOut206[2] , \nOut9_20[0] , \nOut26_5[3] , 
        \nOut18_1[6] , \nOut20_5[7] , \nScanOut332[1] , \nScanOut652[0] , 
        \nScanOut766[3] , \nOut13_16[5] , \nOut29_12[5] , \nScanOut406[6] , 
        \nOut16_29[1] , \nScanOut532[5] , \nOut20_22[4] , \nScanOut680[6] , 
        \nScanOut807[7] , \nOut7_20[4] , \nOut7_23[7] , \nScanOut933[4] , 
        \nScanOut683[5] , \nScanOut804[4] , \nScanOut930[7] , \nScanOut165[4] , 
        \nScanOut205[1] , \nScanOut651[3] , \nScanOut765[0] , \nScanOut331[2] , 
        \nOut13_15[6] , \nScanOut405[5] , \nScanOut531[6] , \nOut20_21[7] , 
        \nOut28_30[0] , \nOut10_23[3] , \nScanOut384[3] , \nScanOut863[3] , 
        \nOut29_11[6] , \nOut30_10[1] , \nScanOut957[0] , \nScanOut584[7] , 
        \nOut26_28[6] , \nOut19_13[2] , \nScanOut1013[5] , \nScanOut636[4] , 
        \nOut23_17[2] , \nScanOut101[0] , \nScanOut102[3] , \nOut4_16[1] , 
        \nScanOut262[6] , \nScanOut702[7] , \nScanOut985[6] , \nOut8_19[4] , 
        \nScanOut356[5] , \nScanOut462[2] , \nScanOut556[1] , \nOut4_15[2] , 
        \nScanOut261[5] , \nOut31_8[0] , \nScanOut355[6] , \nScanOut635[7] , 
        \nScanOut701[4] , \nScanOut986[5] , \nScanOut126[7] , \nOut5_13[3] , 
        \nOut10_20[0] , \nScanOut387[0] , \nScanOut461[1] , \nScanOut555[2] , 
        \nOut19_10[1] , \nOut23_14[1] , \nScanOut860[0] , \nOut30_13[2] , 
        \nScanOut954[3] , \nScanOut587[4] , \nOut18_31[7] , \nScanOut372[1] , 
        \nScanOut1010[6] , \nScanOut246[2] , \nOut19_9[3] , \nScanOut612[0] , 
        \nScanOut726[3] , \nScanOut895[1] , \nScanOut294[4] , \nScanOut446[6] , 
        \nScanOut572[5] , \nOut31_15[3] , \nScanOut27[4] , \nOut6_8[7] , 
        \nOut13_8[6] , \nScanOut973[4] , \nOut14_19[5] , \nScanOut847[7] , 
        \nOut15_8[2] , \nOut22_12[0] , \nScanOut494[0] , \nOut18_16[0] , 
        \nScanOut24[7] , \nOut11_26[1] , \nScanOut970[7] , \nScanOut43[0] , 
        \nScanOut125[4] , \nOut5_10[0] , \nOut4_31[6] , \nScanOut297[7] , 
        \nScanOut844[4] , \nOut31_16[0] , \nOut11_25[2] , \nScanOut497[3] , 
        \nOut18_15[3] , \nScanOut611[3] , \nOut22_11[3] , \nScanOut725[0] , 
        \nOut23_30[5] , \nScanOut896[2] , \nScanOut371[2] , \nScanOut245[1] , 
        \nScanOut445[5] , \nScanOut571[6] , \nOut6_26[5] , \nScanOut917[0] , 
        \nOut28_8[6] , \nScanOut790[1] , \nScanOut823[3] , \nOut0_10[3] , 
        \nOut2_4[5] , \nScanOut40[3] , \nOut3_19[1] , \nScanOut91[6] , 
        \nScanOut190[5] , \nScanOut92[5] , \nScanOut142[3] , \nScanOut222[6] , 
        \nScanOut316[5] , \nScanOut676[4] , \nScanOut742[7] , \nOut22_9[3] , 
        \nOut12_13[7] , \nScanOut422[2] , \nOut21_27[6] , \nScanOut516[1] , 
        \nOut24_9[7] , \nOut24_18[2] , \nOut28_17[7] , \nScanOut221[5] , 
        \nScanOut315[6] , \nScanOut141[0] , \nScanOut675[7] , \nScanOut741[4] , 
        \nOut28_14[4] , \nOut12_10[4] , \nOut13_31[2] , \nScanOut421[1] , 
        \nOut21_24[5] , \nScanOut515[2] , \nOut1_15[3] , \nOut1_16[0] , 
        \nOut6_25[6] , \nScanOut793[2] , \nScanOut914[3] , \nScanOut193[6] , 
        \nScanOut820[0] , \nOut15_23[2] , \nOut23_28[7] , \nOut26_17[3] , 
        \nScanOut968[5] , \nOut4_29[4] , \nOut8_26[1] , \nScanOut609[1] , 
        \nOut8_25[2] , \nScanOut369[0] , \nScanOut569[4] , \nOut30_3[6] , 
        \nOut2_20[5] , \nOut2_23[6] , \nScanOut159[2] , \nScanOut239[7] , 
        \nOut15_20[1] , \nOut30_0[5] , \nOut26_14[0] , \nOut13_29[0] , 
        \nScanOut759[6] , \nOut25_22[5] , \nScanOut439[3] , \nOut16_16[4] , 
        \nScanOut58[1] , \nScanOut788[3] , \nScanOut838[2] , \nScanOut89[4] , 
        \nScanOut188[7] , \nOut16_15[7] , \nOut25_21[6] , \nOut2_7[6] , 
        \nOut3_25[5] , \nOut11_4[0] , \nOut17_4[4] , \nOut4_4[1] , 
        \nOut29_0[1] , \nOut8_5[0] , \nScanOut698[6] , \nOut24_24[6] , 
        \nOut8_6[3] , \nOut17_10[7] , \nOut25_1[0] , \nOut17_13[4] , 
        \nOut16_31[1] , \nOut21_18[1] , \nOut23_1[4] , \nOut11_7[3] , 
        \nScanOut329[2] , \nScanOut529[6] , \nOut25_2[3] , \nScanOut649[3] , 
        \nOut24_27[5] , \nOut28_28[0] , \nOut23_2[7] , \nOut3_26[6] , 
        \nOut4_7[2] , \nOut6_19[2] , \nScanOut928[7] , \nOut29_3[2] , 
        \nOut17_7[7] , \nOut20_5[5] , \nOut26_5[1] , \nOut0_13[0] , 
        \nScanOut18[3] , \nOut1_0[4] , \nOut1_31[5] , \nOut7_0[0] , 
        \nOut9_20[2] , \nOut18_1[4] , \nOut26_30[6] , \nOut27_11[0] , 
        \nOut12_0[1] , \nOut14_25[1] , \nOut14_0[5] , \nOut1_3[7] , 
        \nOut7_3[3] , \nOut14_3[6] , \nOut14_26[2] , \nOut18_29[7] , 
        \nOut31_29[7] , \nScanOut1008[6] , \nOut11_19[6] , \nOut27_12[3] , 
        \nOut12_3[2] , \nScanOut119[0] , \nOut20_6[6] , \nScanOut878[0] , 
        \nScanOut279[5] , \nOut9_23[1] , \nScanOut479[1] , \nOut18_2[7] , 
        \nScanOut719[4] , \nOut26_6[2] , \nScanOut15[6] , \nOut1_29[7] , 
        \nScanOut64[5] , \nScanOut165[6] , \nOut13_15[4] , \nScanOut405[7] , 
        \nScanOut531[4] , \nOut20_21[5] , \nOut29_11[4] , \nScanOut205[3] , 
        \nScanOut331[0] , \nScanOut651[1] , \nScanOut765[2] , \nOut28_30[2] , 
        \nOut7_20[6] , \nScanOut930[5] , \nScanOut67[6] , \nScanOut683[7] , 
        \nScanOut804[6] , \nScanOut101[2] , \nScanOut166[5] , \nOut7_23[5] , 
        \nScanOut680[4] , \nScanOut933[6] , \nScanOut807[5] , \nOut29_12[7] , 
        \nScanOut206[0] , \nScanOut332[3] , \nOut13_16[7] , \nScanOut406[4] , 
        \nOut16_29[3] , \nScanOut532[7] , \nOut20_22[6] , \nOut10_20[2] , 
        \nOut19_10[3] , \nOut18_31[5] , \nScanOut652[2] , \nScanOut766[1] , 
        \nOut23_14[3] , \nScanOut1010[4] , \nScanOut387[2] , \nScanOut587[6] , 
        \nScanOut860[2] , \nOut30_13[0] , \nScanOut954[1] , \nScanOut102[1] , 
        \nOut4_15[0] , \nScanOut355[4] , \nScanOut461[3] , \nScanOut555[0] , 
        \nScanOut261[7] , \nScanOut462[0] , \nScanOut635[5] , \nScanOut701[6] , 
        \nScanOut986[7] , \nScanOut556[3] , \nOut31_8[2] , \nScanOut636[6] , 
        \nScanOut702[5] , \nScanOut985[4] , \nOut4_16[3] , \nScanOut356[7] , 
        \nOut8_19[6] , \nScanOut262[4] , \nOut10_23[1] , \nScanOut584[5] , 
        \nScanOut1013[7] , \nOut26_28[4] , \nOut11_14[3] , \nScanOut384[1] , 
        \nOut19_13[0] , \nOut23_17[0] , \nScanOut863[1] , \nScanOut957[2] , 
        \nOut30_10[3] , \nScanOut592[1] , \nScanOut1005[3] , \nOut18_24[2] , 
        \nOut22_20[2] , \nScanOut941[6] , \nScanOut16[5] , \nScanOut114[5] , 
        \nScanOut392[5] , \nScanOut875[5] , \nOut31_27[1] , \nScanOut474[4] , 
        \nScanOut540[7] , \nScanOut117[6] , \nOut5_21[1] , \nScanOut340[3] , 
        \nScanOut620[2] , \nScanOut714[1] , \nScanOut993[0] , \nScanOut274[0] , 
        \nOut5_22[2] , \nScanOut343[0] , \nScanOut477[7] , \nOut20_8[0] , 
        \nScanOut543[4] , \nScanOut277[3] , \nOut11_17[0] , \nOut14_28[4] , 
        \nScanOut623[1] , \nScanOut717[2] , \nOut26_8[4] , \nScanOut990[3] , 
        \nOut22_23[1] , \nOut18_27[1] , \nScanOut591[2] , \nScanOut1006[0] , 
        \nScanOut391[6] , \nOut31_24[2] , \nOut2_9[0] , \nScanOut71[2] , 
        \nScanOut170[1] , \nScanOut876[6] , \nScanOut942[5] , \nScanOut210[4] , 
        \nScanOut324[7] , \nOut12_21[5] , \nOut28_25[5] , \nScanOut410[0] , 
        \nOut21_15[4] , \nScanOut524[3] , \nScanOut644[6] , \nScanOut770[5] , 
        \nOut6_14[7] , \nScanOut925[2] , \nOut11_9[5] , \nScanOut696[0] , 
        \nScanOut811[1] , \nOut2_11[4] , \nOut1_24[2] , \nScanOut72[1] , 
        \nOut6_17[4] , \nScanOut926[1] , \nOut3_28[0] , \nOut4_9[4] , 
        \nScanOut812[2] , \nScanOut695[3] , \nScanOut173[2] , \nOut8_8[5] , 
        \nOut17_9[1] , \nOut12_22[6] , \nScanOut413[3] , \nOut21_16[7] , 
        \nScanOut527[0] , \nOut24_29[3] , \nScanOut213[7] , \nScanOut327[4] , 
        \nScanOut647[5] , \nScanOut773[6] , \nOut28_26[6] , \nOut8_14[3] , 
        \nOut31_5[7] , \nScanOut988[1] , \nOut1_27[1] , \nScanOut389[4] , 
        \nOut14_30[6] , \nOut15_11[0] , \nScanOut589[0] , \nOut26_25[1] , 
        \nOut15_12[3] , \nOut26_26[2] , \nScanOut558[5] , \nOut23_19[6] , 
        \nScanOut959[4] , \nOut31_6[4] , \nOut4_18[5] , \nOut8_17[0] , 
        \nScanOut638[0] , \nScanOut358[1] , \nOut3_30[2] , \nScanOut0[6] , 
        \nScanOut3[5] , \nOut0_5[6] , \nOut0_6[5] , \nOut2_12[7] , 
        \nScanOut168[3] , \nOut13_18[1] , \nOut16_24[6] , \nOut25_10[7] , 
        \nOut24_31[1] , \nOut25_13[4] , \nScanOut208[6] , \nScanOut408[2] , 
        \nOut16_27[5] , \nScanOut768[7] , \nOut3_1[7] , \nOut3_2[4] , 
        \nScanOut69[0] , \nOut3_17[7] , \nOut5_2[0] , \nOut9_3[1] , 
        \nScanOut318[3] , \nScanOut678[2] , \nScanOut809[3] , \nOut22_7[5] , 
        \nScanOut518[7] , \nOut17_22[5] , \nOut21_29[0] , \nOut24_7[1] , 
        \nOut24_16[4] , \nOut28_19[1] , \nOut28_6[0] , \nOut6_28[3] , 
        \nScanOut919[6] , \nOut16_2[5] , \nOut10_2[1] , \nOut3_14[4] , 
        \nOut16_1[6] , \nOut5_1[3] , \nOut28_5[3] , \nOut9_0[2] , 
        \nOut10_1[2] , \nOut17_21[6] , \nOut22_4[6] , \nOut24_15[7] , 
        \nOut24_4[2] , \nOut0_21[2] , \nOut0_22[1] , \nScanOut29[2] , 
        \nOut6_6[1] , \nOut13_6[0] , \nScanOut849[1] , \nOut14_17[3] , 
        \nOut15_6[4] , \nOut18_18[6] , \nScanOut248[4] , \nOut9_12[0] , 
        \nOut11_28[7] , \nOut27_23[2] , \nOut19_7[5] , \nScanOut728[5] , 
        \nOut27_3[0] , \nScanOut128[1] , \nOut21_3[4] , \nScanOut448[0] , 
        \nScanOut898[4] , \nOut8_30[5] , \nOut9_11[3] , \nOut27_0[3] , 
        \nScanOut299[1] , \nOut13_5[3] , \nOut19_4[6] , \nOut21_0[7] , 
        \nOut31_18[6] , \nScanOut56[7] , \nOut6_5[2] , \nScanOut499[5] , 
        \nOut14_14[0] , \nOut27_20[1] , \nOut15_5[7] , \nScanOut84[1] , 
        \nScanOut185[2] , \nOut7_12[4] , \nScanOut785[6] , \nScanOut902[7] , 
        \nScanOut836[4] , \nScanOut237[1] , \nScanOut303[2] , \nScanOut663[3] , 
        \nScanOut757[0] , \nScanOut87[2] , \nScanOut157[4] , \nOut29_23[6] , 
        \nOut13_27[6] , \nScanOut437[5] , \nOut16_18[2] , \nOut20_13[7] , 
        \nScanOut503[6] , \nScanOut234[2] , \nScanOut300[1] , \nScanOut660[0] , 
        \nScanOut754[3] , \nOut13_24[5] , \nScanOut434[6] , \nOut20_10[4] , 
        \nOut21_31[2] , \nScanOut500[5] , \nOut29_20[5] , \nScanOut10[2] , 
        \nScanOut13[1] , \nScanOut31[0] , \nScanOut32[3] , \nOut1_18[6] , 
        \nScanOut55[4] , \nScanOut154[7] , \nOut6_30[1] , \nScanOut901[4] , 
        \nOut7_11[7] , \nScanOut186[1] , \nScanOut786[5] , \nScanOut835[7] , 
        \nScanOut607[7] , \nScanOut733[4] , \nOut4_27[2] , \nScanOut880[6] , 
        \nScanOut133[0] , \nOut8_28[7] , \nScanOut367[6] , \nScanOut253[5] , 
        \nScanOut453[1] , \nScanOut567[2] , \nScanOut966[3] , \nScanOut281[3] , 
        \nScanOut852[0] , \nOut30_21[2] , \nScanOut282[0] , \nOut10_12[0] , 
        \nScanOut481[7] , \nScanOut1022[6] , \nOut19_22[1] , \nOut26_19[5] , 
        \nOut23_26[1] , \nOut30_22[1] , \nOut1_8[5] , \nScanOut74[6] , 
        \nScanOut77[5] , \nOut4_24[1] , \nOut10_11[3] , \nOut11_30[5] , 
        \nScanOut482[4] , \nOut19_21[2] , \nOut23_25[2] , \nScanOut851[3] , 
        \nScanOut965[0] , \nScanOut1021[5] , \nScanOut130[3] , 
        \nScanOut250[6] , \nScanOut364[5] , \nScanOut604[4] , \nScanOut730[7] , 
        \nScanOut883[5] , \nScanOut176[6] , \nScanOut216[3] , \nScanOut322[0] , 
        \nScanOut450[2] , \nScanOut564[1] , \nScanOut642[1] , \nScanOut776[2] , 
        \nOut23_9[5] , \nScanOut416[7] , \nOut17_18[6] , \nOut21_13[3] , 
        \nScanOut522[4] , \nOut25_9[1] , \nOut12_27[2] , \nOut28_23[2] , 
        \nOut6_11[3] , \nOut6_12[0] , \nScanOut923[5] , \nOut7_30[5] , 
        \nScanOut690[7] , \nOut29_8[0] , \nScanOut817[6] , \nScanOut920[6] , 
        \nScanOut175[5] , \nScanOut215[0] , \nScanOut321[3] , \nScanOut693[4] , 
        \nScanOut814[5] , \nOut12_24[1] , \nScanOut641[2] , \nScanOut775[1] , 
        \nScanOut394[2] , \nScanOut415[4] , \nOut21_10[0] , \nOut28_20[1] , 
        \nScanOut521[7] , \nOut20_31[6] , \nOut31_21[6] , \nScanOut947[1] , 
        \nOut0_18[2] , \nOut5_27[6] , \nOut7_8[1] , \nOut12_8[0] , 
        \nOut14_8[4] , \nOut18_22[5] , \nScanOut873[2] , \nOut22_26[5] , 
        \nScanOut594[6] , \nScanOut1003[4] , \nOut27_19[1] , \nOut11_12[4] , 
        \nScanOut346[4] , \nScanOut272[7] , \nOut9_28[3] , \nOut18_9[5] , 
        \nScanOut626[5] , \nScanOut712[6] , \nScanOut995[7] , \nScanOut111[1] , 
        \nScanOut112[2] , \nOut5_24[5] , \nScanOut345[7] , \nScanOut472[3] , 
        \nScanOut546[0] , \nScanOut625[6] , \nScanOut711[5] , \nScanOut996[4] , 
        \nScanOut271[4] , \nScanOut471[0] , \nScanOut545[3] , \nOut2_14[0] , 
        \nOut2_17[3] , \nOut10_30[1] , \nScanOut397[1] , \nScanOut870[1] , 
        \nScanOut944[2] , \nOut31_22[5] , \nScanOut1000[7] , \nOut11_11[7] , 
        \nScanOut597[5] , \nOut18_21[6] , \nOut22_25[6] , \nOut7_28[7] , 
        \nScanOut339[1] , \nScanOut938[4] , \nOut16_21[2] , \nOut16_22[1] , 
        \nOut20_29[4] , \nScanOut659[0] , \nOut25_16[0] , \nOut29_19[5] , 
        \nScanOut539[5] , \nScanOut688[5] , \nOut25_15[3] , \nOut1_21[6] , 
        \nOut1_22[5] , \nScanOut709[7] , \nScanOut109[3] , \nOut8_12[4] , 
        \nScanOut269[6] , \nScanOut469[2] , \nOut31_3[0] , \nOut8_11[7] , 
        \nOut10_28[3] , \nScanOut868[3] , \nScanOut1018[5] , \nOut15_14[4] , 
        \nOut15_17[7] , \nOut19_18[2] , \nOut26_23[6] , \nOut30_18[2] , 
        \nOut26_20[5] , \nOut9_30[1] , \nOut6_0[6] , \nOut13_0[7] , 
        \nOut14_11[4] , \nOut15_0[3] , \nOut27_25[5] , \nOut15_30[2] , 
        \nOut0_3[1] , \nOut0_24[6] , \nOut21_5[3] , \nOut27_5[7] , 
        \nOut0_27[5] , \nOut5_18[1] , \nOut9_14[7] , \nOut9_17[4] , 
        \nOut19_1[2] , \nScanOut579[7] , \nOut21_6[0] , \nScanOut379[3] , 
        \nOut19_2[1] , \nOut6_3[5] , \nOut14_12[7] , \nScanOut619[2] , 
        \nOut27_6[4] , \nOut22_19[2] , \nOut15_3[0] , \nOut27_26[6] , 
        \nScanOut5[2] , \nScanOut34[4] , \nScanOut48[2] , \nOut2_30[6] , 
        \nOut3_4[3] , \nScanOut99[7] , \nOut9_5[6] , \nOut13_3[4] , 
        \nScanOut978[6] , \nOut17_24[2] , \nOut24_10[3] , \nOut25_31[5] , 
        \nOut22_1[2] , \nOut24_1[6] , \nOut3_11[0] , \nScanOut198[4] , 
        \nOut10_4[6] , \nOut16_4[2] , \nOut3_7[0] , \nOut5_4[7] , 
        \nOut28_0[7] , \nOut10_7[5] , \nScanOut798[0] , \nOut3_12[3] , 
        \nOut5_7[4] , \nOut28_3[4] , \nOut16_7[1] , \nScanOut828[1] , 
        \nOut4_21[5] , \nScanOut135[7] , \nScanOut149[1] , \nOut9_6[5] , 
        \nScanOut429[0] , \nOut17_27[1] , \nOut12_18[5] , \nOut24_2[5] , 
        \nOut24_13[0] , \nScanOut229[4] , \nOut22_2[1] , \nScanOut749[5] , 
        \nScanOut455[6] , \nScanOut561[5] , \nScanOut255[2] , \nScanOut361[1] , 
        \nScanOut287[4] , \nOut10_14[7] , \nScanOut487[0] , \nOut19_24[6] , 
        \nScanOut601[0] , \nScanOut735[3] , \nScanOut886[1] , \nOut23_20[6] , 
        \nScanOut1024[1] , \nOut30_27[5] , \nScanOut960[4] , \nScanOut37[7] , 
        \nOut10_17[4] , \nScanOut484[3] , \nScanOut854[7] , \nOut15_28[0] , 
        \nOut19_27[5] , \nOut23_23[5] , \nScanOut50[0] , \nOut4_22[6] , 
        \nScanOut136[4] , \nScanOut284[7] , \nScanOut857[4] , \nScanOut963[7] , 
        \nOut30_24[6] , \nScanOut456[5] , \nScanOut562[6] , \nScanOut602[3] , 
        \nScanOut736[0] , \nOut30_8[4] , \nScanOut885[2] , \nScanOut183[5] , 
        \nScanOut256[1] , \nScanOut362[2] , \nOut7_14[3] , \nScanOut783[1] , 
        \nScanOut904[0] , \nScanOut431[2] , \nOut20_15[0] , \nScanOut830[3] , 
        \nScanOut505[1] , \nScanOut6[1] , \nScanOut82[6] , \nScanOut151[3] , 
        \nOut29_25[1] , \nOut13_21[1] , \nScanOut231[6] , \nScanOut305[5] , 
        \nScanOut665[4] , \nScanOut751[7] , \nOut13_22[2] , \nOut25_29[7] , 
        \nOut29_26[2] , \nScanOut45[7] , \nScanOut53[3] , \nOut2_28[4] , 
        \nScanOut81[5] , \nScanOut152[0] , \nScanOut232[5] , \nScanOut306[6] , 
        \nScanOut432[1] , \nOut20_16[3] , \nScanOut506[2] , \nScanOut180[6] , 
        \nScanOut666[7] , \nScanOut752[4] , \nOut7_17[0] , \nScanOut907[3] , 
        \nOut6_20[2] , \nScanOut196[2] , \nScanOut780[2] , \nScanOut833[0] , 
        \nScanOut911[7] , \nScanOut94[2] , \nScanOut97[1] , \nScanOut144[4] , 
        \nOut12_15[0] , \nScanOut796[6] , \nScanOut825[4] , \nOut28_11[0] , 
        \nOut29_30[6] , \nScanOut224[1] , \nScanOut310[2] , \nScanOut424[5] , 
        \nOut21_21[1] , \nScanOut510[6] , \nScanOut147[7] , \nOut9_8[3] , 
        \nScanOut427[6] , \nOut21_22[2] , \nScanOut670[3] , \nScanOut744[0] , 
        \nScanOut513[5] , \nOut17_29[7] , \nOut28_12[3] , \nOut12_16[3] , 
        \nScanOut227[2] , \nScanOut313[1] , \nScanOut673[0] , \nScanOut747[3] , 
        \nScanOut8[7] , \nScanOut21[3] , \nScanOut46[4] , \nOut3_9[6] , 
        \nOut10_9[3] , \nScanOut195[1] , \nScanOut120[0] , \nOut5_9[2] , 
        \nOut6_23[1] , \nScanOut795[5] , \nScanOut912[4] , \nScanOut440[1] , 
        \nOut16_9[7] , \nScanOut826[7] , \nScanOut574[2] , \nOut5_15[4] , 
        \nScanOut374[6] , \nScanOut614[7] , \nScanOut720[4] , \nScanOut893[6] , 
        \nScanOut240[5] , \nOut11_20[6] , \nScanOut492[7] , \nOut18_10[7] , 
        \nOut19_31[1] , \nOut22_14[7] , \nScanOut22[0] , \nScanOut291[0] , 
        \nScanOut292[3] , \nScanOut841[0] , \nScanOut975[3] , \nOut31_13[4] , 
        \nOut11_23[5] , \nScanOut491[4] , \nOut18_13[4] , \nOut22_17[4] , 
        \nOut27_28[0] , \nOut31_10[7] , \nOut30_31[1] , \nScanOut976[0] , 
        \nOut0_29[3] , \nScanOut123[3] , \nOut21_8[6] , \nScanOut842[3] , 
        \nOut5_16[7] , \nScanOut377[5] , \nScanOut443[2] , \nScanOut577[1] , 
        \nScanOut243[6] , \nOut9_19[2] , \nScanOut617[4] , \nScanOut723[7] , 
        \nScanOut890[5] , \nOut2_25[1] , \nOut16_10[3] , \nOut27_8[2] , 
        \nOut17_31[5] , \nOut25_24[2] , \nOut2_26[2] , \nOut7_19[6] , 
        \nScanOut909[5] , \nOut29_28[4] , \nOut1_10[7] , \nOut8_20[6] , 
        \nScanOut289[2] , \nScanOut308[0] , \nOut16_13[0] , \nOut25_27[1] , 
        \nScanOut508[4] , \nOut20_18[5] , \nOut15_25[5] , \nScanOut668[1] , 
        \nScanOut489[6] , \nOut26_11[4] , \nOut27_30[2] , \nOut30_29[3] , 
        \nOut30_5[1] , \nScanOut888[7] , \nOut1_13[4] , \nScanOut138[2] , 
        \nScanOut458[3] , \nOut30_6[2] , \nScanOut738[6] , \nOut8_23[5] , 
        \nScanOut258[7] , \nOut10_19[2] , \nOut26_12[7] , \nOut19_29[3] , 
        \nScanOut0[2] , \nOut0_15[7] , \nOut0_16[4] , \nScanOut39[1] , 
        \nOut15_26[6] , \nOut5_29[0] , \nOut9_26[5] , \nOut18_7[3] , 
        \nScanOut859[2] , \nScanOut348[2] , \nOut26_3[6] , \nOut1_5[0] , 
        \nOut1_6[3] , \nScanOut548[6] , \nOut20_3[2] , \nScanOut628[3] , 
        \nOut7_6[7] , \nOut12_6[6] , \nOut14_6[2] , \nOut14_23[6] , 
        \nScanOut949[7] , \nOut22_28[3] , \nOut27_17[7] , \nOut12_5[5] , 
        \nScanOut399[7] , \nOut7_5[4] , \nScanOut599[3] , \nOut14_5[1] , 
        \nOut14_20[5] , \nOut27_14[4] , \nOut26_0[5] , \nScanOut998[2] , 
        \nOut2_1[1] , \nOut2_2[2] , \nScanOut79[3] , \nOut9_25[6] , 
        \nOut18_4[0] , \nOut20_0[1] , \nOut3_23[2] , \nOut4_2[6] , 
        \nScanOut819[0] , \nOut29_6[6] , \nOut17_2[3] , \nOut11_2[7] , 
        \nOut3_20[1] , \nScanOut178[0] , \nScanOut218[5] , \nScanOut778[4] , 
        \nOut8_3[7] , \nOut23_7[3] , \nOut12_29[4] , \nScanOut418[1] , 
        \nOut17_16[0] , \nOut25_7[7] , \nOut24_22[1] , \nOut8_0[4] , 
        \nOut17_15[3] , \nOut23_4[0] , \nOut24_21[2] , \nOut25_4[4] , 
        \nOut4_1[5] , \nOut17_1[0] , \nOut29_5[5] , \nOut2_19[5] , 
        \nScanOut104[6] , \nOut4_10[4] , \nScanOut107[5] , \nOut4_13[7] , 
        \nOut10_26[5] , \nOut11_1[4] , \nScanOut381[5] , \nScanOut866[5] , 
        \nScanOut952[6] , \nOut30_15[7] , \nScanOut1016[3] , \nScanOut353[3] , 
        \nOut15_19[1] , \nScanOut581[1] , \nOut23_12[4] , \nOut19_16[4] , 
        \nScanOut633[2] , \nScanOut707[1] , \nScanOut980[0] , \nScanOut267[0] , 
        \nScanOut467[4] , \nScanOut553[7] , \nOut5_31[2] , \nScanOut350[0] , 
        \nScanOut264[3] , \nScanOut630[1] , \nScanOut704[2] , \nScanOut983[3] , 
        \nScanOut163[1] , \nScanOut203[4] , \nOut10_25[6] , \nScanOut382[6] , 
        \nScanOut464[7] , \nScanOut550[4] , \nOut30_16[4] , \nScanOut582[2] , 
        \nOut19_15[7] , \nScanOut865[6] , \nScanOut951[5] , \nOut22_30[1] , 
        \nOut23_11[7] , \nScanOut1015[0] , \nScanOut337[7] , \nOut13_13[3] , 
        \nScanOut657[6] , \nScanOut763[5] , \nOut25_18[6] , \nOut29_17[3] , 
        \nScanOut403[0] , \nScanOut537[3] , \nOut20_27[2] , \nScanOut55[0] , 
        \nScanOut61[1] , \nScanOut62[2] , \nOut7_26[1] , \nScanOut936[2] , 
        \nScanOut685[0] , \nScanOut802[1] , \nScanOut160[2] , \nScanOut200[7] , 
        \nOut7_25[2] , \nScanOut334[4] , \nScanOut654[5] , \nScanOut686[3] , 
        \nScanOut935[1] , \nScanOut760[6] , \nScanOut801[2] , \nScanOut400[3] , 
        \nScanOut534[0] , \nOut20_24[1] , \nOut29_14[0] , \nScanOut186[5] , 
        \nOut13_10[0] , \nOut12_31[6] , \nOut6_30[5] , \nScanOut901[0] , 
        \nOut7_11[3] , \nOut13_24[1] , \nScanOut786[1] , \nScanOut835[3] , 
        \nScanOut3[1] , \nScanOut87[6] , \nScanOut154[3] , \nOut29_20[1] , 
        \nScanOut234[6] , \nScanOut300[5] , \nScanOut434[2] , \nOut20_10[0] , 
        \nOut21_31[6] , \nScanOut500[1] , \nScanOut437[1] , \nOut16_18[6] , 
        \nScanOut660[4] , \nScanOut754[7] , \nOut20_13[3] , \nScanOut503[2] , 
        \nOut29_23[2] , \nOut0_5[2] , \nScanOut31[4] , \nScanOut56[3] , 
        \nScanOut84[5] , \nScanOut157[0] , \nOut13_27[2] , \nScanOut185[6] , 
        \nScanOut237[5] , \nScanOut303[6] , \nScanOut663[7] , \nScanOut757[4] , 
        \nOut4_24[5] , \nScanOut130[7] , \nOut7_12[0] , \nScanOut785[2] , 
        \nScanOut902[3] , \nScanOut450[6] , \nScanOut836[0] , \nScanOut564[5] , 
        \nScanOut604[0] , \nScanOut730[3] , \nScanOut883[1] , \nScanOut250[2] , 
        \nScanOut364[1] , \nOut10_11[7] , \nOut11_30[1] , \nScanOut482[0] , 
        \nScanOut1021[1] , \nOut19_21[6] , \nOut23_25[6] , \nScanOut32[7] , 
        \nScanOut281[7] , \nScanOut282[4] , \nScanOut851[7] , \nScanOut965[4] , 
        \nOut30_22[5] , \nOut10_12[4] , \nScanOut481[3] , \nOut19_22[5] , 
        \nOut23_26[5] , \nOut26_19[1] , \nScanOut1022[2] , \nOut30_21[6] , 
        \nScanOut966[7] , \nOut1_18[2] , \nOut4_27[6] , \nScanOut133[4] , 
        \nScanOut852[4] , \nScanOut453[5] , \nScanOut567[6] , \nOut8_28[3] , 
        \nScanOut367[2] , \nScanOut253[1] , \nScanOut607[3] , \nScanOut733[0] , 
        \nOut3_1[3] , \nOut9_0[6] , \nOut17_21[2] , \nScanOut880[2] , 
        \nOut10_1[6] , \nOut22_4[2] , \nOut24_4[6] , \nOut24_15[3] , 
        \nOut3_2[0] , \nOut3_14[0] , \nOut5_1[7] , \nOut28_5[7] , 
        \nOut16_1[2] , \nOut3_17[3] , \nOut10_2[5] , \nOut16_2[1] , 
        \nOut5_2[4] , \nOut28_6[4] , \nOut6_5[6] , \nOut6_28[7] , 
        \nScanOut919[2] , \nOut9_3[5] , \nScanOut518[3] , \nOut17_22[1] , 
        \nOut21_29[4] , \nOut24_16[0] , \nOut28_19[5] , \nScanOut318[7] , 
        \nOut22_7[1] , \nOut24_7[5] , \nOut14_14[4] , \nScanOut678[6] , 
        \nOut15_5[3] , \nScanOut499[1] , \nScanOut299[5] , \nOut27_20[5] , 
        \nOut31_18[2] , \nOut0_6[1] , \nOut0_21[6] , \nOut8_30[1] , 
        \nOut9_11[7] , \nOut13_5[7] , \nOut21_0[3] , \nOut19_4[2] , 
        \nOut27_0[7] , \nScanOut898[0] , \nOut0_22[5] , \nScanOut128[5] , 
        \nScanOut448[4] , \nOut21_3[0] , \nScanOut728[1] , \nScanOut29[6] , 
        \nOut6_6[5] , \nScanOut248[0] , \nOut9_12[4] , \nOut27_3[4] , 
        \nOut19_7[1] , \nOut11_28[3] , \nOut14_17[7] , \nOut15_6[0] , 
        \nOut27_23[6] , \nOut18_18[2] , \nOut13_6[4] , \nScanOut849[5] , 
        \nOut2_11[0] , \nOut2_12[3] , \nOut1_24[6] , \nOut1_27[5] , 
        \nOut4_18[1] , \nOut8_17[4] , \nScanOut358[5] , \nScanOut389[0] , 
        \nOut15_12[7] , \nScanOut558[1] , \nScanOut638[4] , \nOut31_6[0] , 
        \nOut23_19[2] , \nScanOut959[0] , \nOut26_26[6] , \nOut14_30[2] , 
        \nOut15_11[4] , \nScanOut589[4] , \nOut26_25[5] , \nScanOut988[5] , 
        \nScanOut69[4] , \nOut8_14[7] , \nOut31_5[3] , \nScanOut809[7] , 
        \nScanOut168[7] , \nScanOut208[2] , \nScanOut768[3] , \nOut13_18[5] , 
        \nScanOut408[6] , \nOut16_27[1] , \nOut25_13[0] , \nOut16_24[2] , 
        \nOut25_10[3] , \nOut24_31[5] , \nOut3_30[6] , \nOut0_10[7] , 
        \nOut0_13[4] , \nScanOut15[2] , \nScanOut16[1] , \nScanOut114[1] , 
        \nScanOut117[2] , \nOut5_22[6] , \nOut11_17[4] , \nScanOut391[2] , 
        \nScanOut876[2] , \nScanOut942[1] , \nScanOut591[6] , \nOut31_24[6] , 
        \nScanOut1006[4] , \nScanOut343[4] , \nOut14_28[0] , \nOut18_27[5] , 
        \nOut22_23[5] , \nScanOut623[5] , \nScanOut717[6] , \nOut26_8[0] , 
        \nScanOut990[7] , \nScanOut277[7] , \nScanOut477[3] , \nScanOut543[0] , 
        \nOut5_21[5] , \nScanOut340[7] , \nOut20_8[4] , \nScanOut274[4] , 
        \nScanOut620[6] , \nScanOut714[5] , \nScanOut993[4] , \nScanOut392[1] , 
        \nScanOut474[0] , \nScanOut540[3] , \nOut31_27[5] , \nScanOut941[2] , 
        \nOut2_4[1] , \nOut2_7[2] , \nOut2_9[4] , \nScanOut72[5] , 
        \nOut3_28[4] , \nScanOut173[6] , \nScanOut213[3] , \nScanOut327[0] , 
        \nOut11_14[7] , \nOut18_24[6] , \nScanOut875[1] , \nScanOut592[5] , 
        \nOut22_20[6] , \nScanOut1005[7] , \nOut12_22[2] , \nScanOut647[1] , 
        \nScanOut773[2] , \nOut24_29[7] , \nOut8_8[1] , \nOut28_26[2] , 
        \nScanOut413[7] , \nOut21_16[3] , \nOut17_9[5] , \nScanOut527[4] , 
        \nOut6_17[0] , \nScanOut926[5] , \nOut4_9[0] , \nScanOut812[6] , 
        \nScanOut695[7] , \nOut1_29[3] , \nScanOut64[1] , \nScanOut67[2] , 
        \nScanOut71[6] , \nOut11_9[1] , \nScanOut166[1] , \nScanOut170[5] , 
        \nOut6_14[3] , \nScanOut925[6] , \nScanOut210[0] , \nScanOut324[3] , 
        \nScanOut644[2] , \nScanOut696[4] , \nScanOut770[1] , \nScanOut811[5] , 
        \nScanOut410[4] , \nOut21_15[0] , \nScanOut524[7] , \nScanOut206[4] , 
        \nScanOut332[7] , \nOut12_21[1] , \nOut28_25[1] , \nScanOut652[6] , 
        \nScanOut766[5] , \nScanOut406[0] , \nOut16_29[7] , \nOut20_22[2] , 
        \nScanOut532[3] , \nOut29_12[3] , \nOut13_16[3] , \nOut7_20[2] , 
        \nOut7_23[1] , \nScanOut680[0] , \nScanOut933[2] , \nScanOut807[1] , 
        \nScanOut930[1] , \nOut4_16[7] , \nScanOut165[2] , \nScanOut205[7] , 
        \nScanOut331[4] , \nScanOut683[3] , \nScanOut804[2] , \nOut13_15[0] , 
        \nScanOut651[5] , \nScanOut765[6] , \nOut29_11[0] , \nOut10_23[5] , 
        \nScanOut384[5] , \nScanOut405[3] , \nOut28_30[6] , \nScanOut531[0] , 
        \nOut20_21[1] , \nOut30_10[7] , \nOut19_13[4] , \nScanOut863[5] , 
        \nScanOut957[6] , \nOut23_17[4] , \nScanOut1013[3] , \nScanOut356[3] , 
        \nScanOut584[1] , \nOut26_28[0] , \nOut8_19[2] , \nScanOut262[0] , 
        \nScanOut636[2] , \nScanOut702[1] , \nScanOut985[0] , \nOut3_26[2] , 
        \nScanOut101[6] , \nScanOut102[5] , \nOut31_8[6] , \nOut4_15[4] , 
        \nScanOut355[0] , \nScanOut462[4] , \nScanOut556[7] , \nScanOut635[1] , 
        \nScanOut701[2] , \nScanOut986[3] , \nScanOut261[3] , \nScanOut461[7] , 
        \nScanOut555[4] , \nOut10_20[6] , \nScanOut387[6] , \nScanOut860[6] , 
        \nScanOut954[5] , \nScanOut587[2] , \nOut30_13[4] , \nScanOut1010[0] , 
        \nOut17_7[3] , \nOut19_10[7] , \nOut18_31[1] , \nOut23_14[7] , 
        \nOut4_7[6] , \nOut6_19[6] , \nScanOut928[3] , \nOut29_3[6] , 
        \nOut3_25[1] , \nOut4_4[5] , \nOut8_5[4] , \nOut8_6[7] , \nOut11_7[7] , 
        \nScanOut329[6] , \nOut17_13[0] , \nScanOut649[7] , \nOut23_2[3] , 
        \nOut24_27[1] , \nOut28_28[4] , \nOut21_18[5] , \nScanOut529[2] , 
        \nOut25_2[7] , \nOut23_1[0] , \nOut17_10[3] , \nOut25_1[4] , 
        \nOut16_31[5] , \nOut24_24[2] , \nOut29_0[5] , \nScanOut698[2] , 
        \nOut11_4[4] , \nOut17_4[0] , \nScanOut719[0] , \nOut26_6[6] , 
        \nScanOut18[7] , \nScanOut119[4] , \nScanOut279[1] , \nOut9_23[5] , 
        \nOut18_2[3] , \nScanOut479[5] , \nOut20_6[2] , \nOut1_0[0] , 
        \nOut1_3[3] , \nOut12_3[6] , \nScanOut878[4] , \nOut7_3[7] , 
        \nOut27_12[7] , \nScanOut1008[2] , \nOut11_19[2] , \nOut14_3[2] , 
        \nOut14_26[6] , \nOut18_29[3] , \nOut7_0[4] , \nOut12_0[5] , 
        \nOut31_29[3] , \nOut14_25[5] , \nOut14_0[1] , \nOut26_30[2] , 
        \nOut9_20[6] , \nOut18_1[0] , \nOut27_11[4] , \nOut26_5[5] , 
        \nScanOut24[3] , \nOut1_15[7] , \nOut1_31[1] , \nOut15_20[5] , 
        \nOut20_5[1] , \nOut26_14[4] , \nOut30_0[1] , \nOut1_16[4] , 
        \nOut4_29[0] , \nOut8_25[6] , \nOut8_26[5] , \nScanOut569[0] , 
        \nOut30_3[2] , \nScanOut369[4] , \nOut2_20[1] , \nScanOut89[0] , 
        \nOut15_23[6] , \nScanOut609[5] , \nOut16_15[3] , \nOut23_28[3] , 
        \nOut25_21[2] , \nOut26_17[7] , \nScanOut968[1] , \nScanOut188[3] , 
        \nOut2_23[2] , \nScanOut58[5] , \nScanOut788[7] , \nScanOut838[6] , 
        \nScanOut125[0] , \nScanOut159[6] , \nOut13_29[4] , \nScanOut439[7] , 
        \nOut16_16[0] , \nOut25_22[1] , \nScanOut239[3] , \nScanOut759[2] , 
        \nOut5_10[4] , \nOut4_31[2] , \nScanOut445[1] , \nScanOut571[2] , 
        \nScanOut371[6] , \nScanOut245[5] , \nScanOut297[3] , \nOut11_25[6] , 
        \nScanOut497[7] , \nOut18_15[7] , \nScanOut611[7] , \nScanOut725[4] , 
        \nScanOut896[6] , \nOut22_11[7] , \nOut23_30[1] , \nOut31_16[4] , 
        \nScanOut970[3] , \nOut6_8[3] , \nScanOut494[4] , \nScanOut844[0] , 
        \nOut0_8[7] , \nScanOut27[0] , \nOut11_26[5] , \nOut14_19[1] , 
        \nOut22_12[4] , \nOut15_8[6] , \nOut18_16[4] , \nScanOut294[0] , 
        \nOut13_8[2] , \nScanOut973[0] , \nScanOut847[3] , \nOut31_15[7] , 
        \nScanOut40[7] , \nScanOut126[3] , \nScanOut446[2] , \nScanOut572[1] , 
        \nOut5_13[7] , \nScanOut372[5] , \nScanOut612[4] , \nScanOut726[7] , 
        \nScanOut895[5] , \nScanOut193[2] , \nScanOut246[6] , \nOut19_9[7] , 
        \nScanOut91[2] , \nScanOut92[1] , \nScanOut141[4] , \nOut6_25[2] , 
        \nScanOut793[6] , \nScanOut914[7] , \nScanOut421[5] , \nOut21_24[1] , 
        \nScanOut820[4] , \nScanOut515[6] , \nOut28_14[0] , \nOut12_10[0] , 
        \nOut13_31[6] , \nScanOut142[7] , \nScanOut221[1] , \nScanOut315[2] , 
        \nScanOut675[3] , \nScanOut741[0] , \nOut12_13[3] , \nOut24_18[6] , 
        \nOut28_17[3] , \nScanOut222[2] , \nScanOut316[1] , \nScanOut422[6] , 
        \nOut21_27[2] , \nScanOut516[5] , \nOut24_9[3] , \nOut22_9[7] , 
        \nScanOut190[1] , \nScanOut676[0] , \nScanOut742[3] , \nScanOut8[3] , 
        \nOut0_15[3] , \nScanOut43[4] , \nOut3_19[5] , \nOut6_26[1] , 
        \nScanOut917[4] , \nOut2_19[1] , \nScanOut61[5] , \nScanOut104[2] , 
        \nOut10_25[2] , \nScanOut790[5] , \nOut28_8[2] , \nScanOut823[7] , 
        \nScanOut1015[4] , \nScanOut382[2] , \nScanOut582[6] , \nOut19_15[3] , 
        \nOut22_30[5] , \nOut23_11[3] , \nScanOut865[2] , \nScanOut951[1] , 
        \nOut30_16[0] , \nScanOut464[3] , \nScanOut550[0] , \nOut4_10[0] , 
        \nOut5_31[6] , \nScanOut350[4] , \nScanOut630[5] , \nScanOut704[6] , 
        \nScanOut983[7] , \nScanOut107[1] , \nScanOut264[7] , \nOut4_13[3] , 
        \nScanOut353[7] , \nScanOut467[0] , \nScanOut553[3] , \nScanOut160[6] , 
        \nScanOut267[4] , \nOut10_26[1] , \nOut15_19[5] , \nScanOut633[6] , 
        \nScanOut707[5] , \nScanOut980[4] , \nScanOut581[5] , \nOut19_16[0] , 
        \nOut23_12[0] , \nScanOut1016[7] , \nScanOut381[1] , \nScanOut866[1] , 
        \nOut30_15[3] , \nScanOut952[2] , \nOut29_14[4] , \nScanOut200[3] , 
        \nScanOut334[0] , \nOut13_10[4] , \nOut12_31[2] , \nScanOut400[7] , 
        \nScanOut534[4] , \nOut20_24[5] , \nScanOut654[1] , \nScanOut760[2] , 
        \nScanOut62[6] , \nOut7_25[6] , \nOut7_26[5] , \nScanOut686[7] , 
        \nScanOut935[5] , \nScanOut801[6] , \nScanOut936[6] , \nScanOut685[4] , 
        \nScanOut802[5] , \nScanOut163[5] , \nOut13_13[7] , \nScanOut403[4] , 
        \nScanOut537[7] , \nOut20_27[6] , \nOut25_18[2] , \nOut29_17[7] , 
        \nScanOut203[0] , \nScanOut337[3] , \nScanOut657[2] , \nScanOut763[1] , 
        \nOut9_25[2] , \nOut18_4[4] , \nOut20_0[5] , \nOut26_0[1] , 
        \nScanOut998[6] , \nOut0_16[0] , \nOut1_5[4] , \nOut7_5[0] , 
        \nOut14_5[5] , \nOut14_20[1] , \nScanOut599[7] , \nOut27_14[0] , 
        \nScanOut399[3] , \nOut1_6[7] , \nOut7_6[3] , \nOut12_5[1] , 
        \nOut12_6[2] , \nOut14_6[6] , \nOut14_23[2] , \nOut22_28[7] , 
        \nOut27_17[3] , \nScanOut949[3] , \nScanOut548[2] , \nOut20_3[6] , 
        \nOut26_3[2] , \nOut2_1[5] , \nOut5_29[4] , \nOut9_26[1] , 
        \nOut18_7[7] , \nScanOut628[7] , \nScanOut348[6] , \nOut11_1[0] , 
        \nOut2_2[6] , \nOut3_20[5] , \nOut4_1[1] , \nOut29_5[1] , 
        \nOut17_1[4] , \nScanOut178[4] , \nOut8_0[0] , \nOut17_15[7] , 
        \nOut12_29[0] , \nOut23_4[4] , \nOut24_21[6] , \nOut25_4[0] , 
        \nOut24_22[5] , \nScanOut218[1] , \nOut8_3[3] , \nScanOut418[5] , 
        \nOut25_7[3] , \nOut17_16[4] , \nOut23_7[7] , \nScanOut778[0] , 
        \nScanOut79[7] , \nOut3_23[6] , \nOut11_2[3] , \nOut17_2[7] , 
        \nOut4_2[2] , \nScanOut819[4] , \nOut29_6[2] , \nScanOut308[4] , 
        \nScanOut668[5] , \nOut16_13[4] , \nOut20_18[1] , \nScanOut508[0] , 
        \nOut2_25[5] , \nOut2_26[6] , \nOut7_19[2] , \nOut25_27[5] , 
        \nOut29_28[0] , \nScanOut909[1] , \nScanOut39[5] , \nOut16_10[7] , 
        \nOut25_24[6] , \nOut17_31[1] , \nOut19_29[7] , \nScanOut859[6] , 
        \nOut0_3[5] , \nScanOut5[6] , \nScanOut6[5] , \nScanOut21[7] , 
        \nScanOut22[4] , \nOut0_29[7] , \nOut1_10[3] , \nOut1_13[0] , 
        \nOut8_23[1] , \nOut10_19[6] , \nOut15_26[2] , \nOut26_12[3] , 
        \nScanOut258[3] , \nScanOut738[2] , \nScanOut138[6] , \nOut30_6[6] , 
        \nScanOut458[7] , \nScanOut888[3] , \nScanOut45[3] , \nScanOut46[0] , 
        \nOut8_20[2] , \nScanOut289[6] , \nOut30_5[5] , \nOut30_29[7] , 
        \nOut15_25[1] , \nScanOut489[2] , \nOut26_11[0] , \nOut27_30[6] , 
        \nOut16_9[3] , \nOut3_9[2] , \nOut5_9[6] , \nOut6_23[5] , 
        \nScanOut795[1] , \nScanOut912[0] , \nScanOut826[3] , \nScanOut94[6] , 
        \nScanOut195[5] , \nScanOut227[6] , \nOut10_9[7] , \nScanOut313[5] , 
        \nScanOut97[5] , \nScanOut147[3] , \nScanOut673[4] , \nScanOut747[7] , 
        \nOut28_12[7] , \nOut9_8[7] , \nOut12_16[7] , \nScanOut427[2] , 
        \nOut17_29[3] , \nOut21_22[6] , \nScanOut513[1] , \nScanOut144[0] , 
        \nScanOut224[5] , \nScanOut310[6] , \nScanOut670[7] , \nScanOut744[4] , 
        \nOut12_15[4] , \nScanOut424[1] , \nOut21_21[5] , \nScanOut510[2] , 
        \nOut28_11[4] , \nOut29_30[2] , \nOut6_20[6] , \nScanOut911[3] , 
        \nScanOut196[6] , \nScanOut796[2] , \nScanOut825[0] , \nScanOut617[0] , 
        \nScanOut723[3] , \nOut27_8[6] , \nScanOut890[1] , \nScanOut123[7] , 
        \nOut5_16[3] , \nScanOut377[1] , \nScanOut243[2] , \nOut9_19[6] , 
        \nScanOut443[6] , \nScanOut577[5] , \nOut21_8[2] , \nScanOut976[4] , 
        \nScanOut291[4] , \nScanOut842[7] , \nOut31_10[3] , \nOut30_31[5] , 
        \nScanOut292[7] , \nOut11_23[1] , \nScanOut491[0] , \nOut27_28[4] , 
        \nOut18_13[0] , \nOut22_17[0] , \nOut31_13[0] , \nScanOut34[0] , 
        \nScanOut37[3] , \nOut4_22[2] , \nScanOut120[4] , \nOut5_15[0] , 
        \nOut11_20[2] , \nScanOut492[3] , \nOut18_10[3] , \nOut19_31[5] , 
        \nOut22_14[3] , \nScanOut841[4] , \nScanOut975[7] , \nScanOut374[2] , 
        \nScanOut240[1] , \nScanOut614[3] , \nScanOut720[0] , \nScanOut893[2] , 
        \nScanOut440[5] , \nScanOut574[6] , \nScanOut136[0] , \nScanOut256[5] , 
        \nScanOut362[6] , \nScanOut602[7] , \nScanOut736[4] , \nScanOut885[6] , 
        \nScanOut284[3] , \nScanOut456[1] , \nOut30_8[0] , \nScanOut562[2] , 
        \nOut30_24[2] , \nOut10_17[0] , \nOut15_28[4] , \nOut23_23[1] , 
        \nScanOut857[0] , \nScanOut963[3] , \nScanOut484[7] , \nOut19_27[1] , 
        \nScanOut960[0] , \nScanOut53[7] , \nOut4_21[1] , \nScanOut287[0] , 
        \nScanOut854[3] , \nOut30_27[1] , \nOut10_14[3] , \nScanOut487[4] , 
        \nScanOut1024[5] , \nOut19_24[2] , \nScanOut601[4] , \nOut23_20[2] , 
        \nScanOut735[7] , \nScanOut886[5] , \nScanOut135[3] , \nScanOut255[6] , 
        \nScanOut361[5] , \nScanOut455[2] , \nScanOut561[1] , \nOut7_17[4] , 
        \nScanOut907[7] , \nOut2_28[0] , \nScanOut780[6] , \nScanOut833[4] , 
        \nScanOut81[1] , \nScanOut180[2] , \nScanOut232[1] , \nScanOut306[2] , 
        \nScanOut666[3] , \nScanOut752[0] , \nOut13_22[6] , \nScanOut432[5] , 
        \nOut20_16[7] , \nScanOut506[6] , \nOut25_29[3] , \nScanOut82[2] , 
        \nScanOut152[4] , \nOut29_26[6] , \nScanOut231[2] , \nScanOut305[1] , 
        \nScanOut665[0] , \nScanOut751[3] , \nOut29_25[5] , \nScanOut50[4] , 
        \nScanOut151[7] , \nOut13_21[5] , \nScanOut431[6] , \nOut20_15[4] , 
        \nScanOut505[5] , \nScanOut183[1] , \nOut7_14[7] , \nScanOut783[5] , 
        \nScanOut904[4] , \nScanOut830[7] , \nOut13_3[0] , \nScanOut978[2] , 
        \nOut0_24[2] , \nOut0_27[1] , \nOut6_3[1] , \nOut14_12[3] , 
        \nOut27_26[2] , \nOut15_3[4] , \nOut22_19[6] , \nOut27_6[0] , 
        \nOut5_18[5] , \nOut9_17[0] , \nScanOut619[6] , \nScanOut379[7] , 
        \nOut9_14[3] , \nOut19_2[5] , \nScanOut579[3] , \nOut21_6[4] , 
        \nOut19_1[6] , \nOut21_5[7] , \nOut27_5[3] , \nOut0_4[6] , 
        \nScanOut10[6] , \nOut2_14[4] , \nScanOut48[6] , \nOut3_12[7] , 
        \nScanOut149[5] , \nOut6_0[2] , \nOut13_0[3] , \nOut14_11[0] , 
        \nOut15_0[7] , \nOut15_30[6] , \nScanOut229[0] , \nOut22_2[5] , 
        \nOut27_25[1] , \nOut12_18[1] , \nScanOut749[1] , \nOut24_13[4] , 
        \nOut9_6[1] , \nScanOut429[4] , \nOut17_27[5] , \nOut16_7[5] , 
        \nOut24_2[1] , \nOut28_3[0] , \nOut2_30[2] , \nOut3_7[4] , 
        \nOut5_7[0] , \nScanOut828[5] , \nOut3_11[4] , \nOut5_4[3] , 
        \nOut10_7[1] , \nOut28_0[3] , \nOut16_4[6] , \nScanOut798[4] , 
        \nOut3_4[7] , \nOut10_4[2] , \nScanOut99[3] , \nScanOut198[0] , 
        \nOut9_5[2] , \nOut17_24[6] , \nOut22_1[6] , \nOut24_1[2] , 
        \nOut24_10[7] , \nOut25_31[1] , \nOut2_17[7] , \nOut7_28[3] , 
        \nScanOut339[5] , \nOut16_21[6] , \nScanOut688[1] , \nOut25_15[7] , 
        \nOut16_22[5] , \nScanOut539[1] , \nOut20_29[0] , \nScanOut659[4] , 
        \nOut25_16[4] , \nOut29_19[1] , \nScanOut938[0] , \nOut1_21[2] , 
        \nOut1_22[1] , \nScanOut109[7] , \nOut8_11[3] , \nOut9_30[5] , 
        \nOut10_28[7] , \nOut15_14[0] , \nOut26_20[1] , \nOut15_17[3] , 
        \nOut19_18[6] , \nOut30_18[6] , \nOut26_23[2] , \nScanOut1018[1] , 
        \nScanOut868[7] , \nOut31_3[4] , \nOut8_12[0] , \nScanOut469[6] , 
        \nScanOut269[2] , \nScanOut709[3] , \nScanOut74[2] , \nOut6_11[7] , 
        \nScanOut175[1] , \nOut12_24[5] , \nScanOut415[0] , \nOut21_10[4] , 
        \nScanOut521[3] , \nOut20_31[2] , \nScanOut215[4] , \nScanOut321[7] , 
        \nScanOut641[6] , \nScanOut775[5] , \nOut28_20[5] , \nOut7_30[1] , 
        \nScanOut920[2] , \nScanOut77[1] , \nScanOut693[0] , \nScanOut814[1] , 
        \nOut6_12[4] , \nScanOut923[1] , \nScanOut176[2] , \nScanOut690[3] , 
        \nOut29_8[4] , \nScanOut817[2] , \nScanOut216[7] , \nScanOut322[4] , 
        \nOut12_27[6] , \nOut28_23[6] , \nScanOut416[3] , \nOut21_13[7] , 
        \nScanOut522[0] , \nOut17_18[2] , \nOut25_9[5] , \nOut23_9[1] , 
        \nOut10_30[5] , \nOut18_21[2] , \nScanOut642[5] , \nScanOut776[6] , 
        \nOut22_25[2] , \nScanOut597[1] , \nScanOut1000[3] , \nOut11_11[3] , 
        \nScanOut397[5] , \nOut31_22[1] , \nScanOut13[5] , \nOut0_18[6] , 
        \nScanOut111[5] , \nScanOut870[5] , \nScanOut944[6] , \nScanOut112[6] , 
        \nOut5_24[1] , \nScanOut345[3] , \nScanOut471[4] , \nScanOut545[7] , 
        \nScanOut271[0] , \nScanOut472[7] , \nScanOut625[2] , \nScanOut711[1] , 
        \nScanOut996[0] , \nScanOut546[4] , \nScanOut626[1] , \nScanOut712[2] , 
        \nScanOut995[3] , \nOut5_27[2] , \nScanOut346[0] , \nOut7_8[5] , 
        \nScanOut272[3] , \nOut9_28[7] , \nOut18_9[1] , \nScanOut594[2] , 
        \nScanOut1003[0] , \nOut11_12[0] , \nOut12_8[4] , \nOut14_8[0] , 
        \nOut18_22[1] , \nOut27_19[5] , \nOut22_26[1] , \nScanOut947[5] , 
        \nScanOut14[6] , \nScanOut17[5] , \nOut1_8[1] , \nScanOut394[6] , 
        \nScanOut873[6] , \nOut31_21[2] , \nOut2_8[0] , \nOut11_8[5] , 
        \nScanOut70[2] , \nScanOut73[1] , \nOut3_29[0] , \nOut4_8[4] , 
        \nOut6_16[4] , \nScanOut927[1] , \nScanOut694[3] , \nScanOut813[2] , 
        \nScanOut171[1] , \nScanOut172[2] , \nOut8_9[5] , \nScanOut412[3] , 
        \nOut17_8[1] , \nOut21_17[7] , \nScanOut526[0] , \nScanOut212[7] , 
        \nScanOut326[4] , \nOut12_23[6] , \nOut28_27[6] , \nScanOut646[5] , 
        \nOut24_28[3] , \nScanOut772[6] , \nOut12_20[5] , \nOut6_15[7] , 
        \nScanOut211[4] , \nScanOut325[7] , \nScanOut411[0] , \nOut28_24[5] , 
        \nScanOut525[3] , \nOut21_14[4] , \nScanOut645[6] , \nScanOut771[5] , 
        \nScanOut924[2] , \nScanOut116[6] , \nOut20_9[0] , \nScanOut697[0] , 
        \nScanOut810[1] , \nOut5_23[2] , \nScanOut476[7] , \nScanOut542[4] , 
        \nScanOut276[3] , \nScanOut342[0] , \nOut11_16[0] , \nOut14_29[4] , 
        \nOut18_26[1] , \nScanOut622[1] , \nScanOut716[2] , \nOut26_9[4] , 
        \nScanOut991[3] , \nOut22_22[1] , \nScanOut590[2] , \nScanOut1007[0] , 
        \nScanOut390[6] , \nOut31_25[2] , \nScanOut943[5] , \nOut11_15[3] , 
        \nScanOut593[1] , \nScanOut877[6] , \nScanOut1004[3] , \nOut18_25[2] , 
        \nOut22_21[2] , \nOut0_20[2] , \nOut2_10[4] , \nOut2_13[7] , 
        \nScanOut115[5] , \nScanOut393[5] , \nScanOut874[5] , \nScanOut940[6] , 
        \nScanOut475[4] , \nOut31_26[1] , \nScanOut541[7] , \nOut5_20[1] , 
        \nScanOut621[2] , \nScanOut715[1] , \nScanOut992[0] , \nScanOut169[3] , 
        \nScanOut275[0] , \nScanOut341[3] , \nScanOut209[6] , \nOut13_19[1] , 
        \nOut25_12[4] , \nScanOut409[2] , \nOut16_26[5] , \nScanOut769[7] , 
        \nScanOut68[0] , \nScanOut808[3] , \nOut1_25[2] , \nOut1_26[1] , 
        \nOut3_31[2] , \nOut15_13[3] , \nOut16_25[6] , \nOut24_30[1] , 
        \nOut25_11[7] , \nOut26_27[2] , \nScanOut559[5] , \nOut23_18[6] , 
        \nScanOut958[4] , \nScanOut639[0] , \nOut31_7[4] , \nOut4_19[5] , 
        \nScanOut359[1] , \nOut8_15[3] , \nOut8_16[0] , \nOut31_4[7] , 
        \nScanOut989[1] , \nScanOut388[4] , \nOut15_10[0] , \nOut14_31[6] , 
        \nScanOut588[0] , \nOut26_24[1] , \nScanOut899[4] , \nOut9_10[3] , 
        \nOut27_1[3] , \nOut8_31[5] , \nScanOut298[1] , \nOut13_4[3] , 
        \nOut19_5[6] , \nOut21_1[7] , \nOut31_19[6] , \nOut0_7[5] , 
        \nOut6_4[2] , \nScanOut498[5] , \nOut14_15[0] , \nOut15_4[7] , 
        \nOut27_21[1] , \nOut0_23[1] , \nScanOut28[2] , \nOut6_7[1] , 
        \nOut13_7[0] , \nOut14_16[3] , \nScanOut848[1] , \nOut15_7[4] , 
        \nOut18_19[6] , \nScanOut249[4] , \nOut9_13[0] , \nOut11_29[7] , 
        \nOut27_22[2] , \nOut19_6[5] , \nScanOut729[5] , \nOut27_2[0] , 
        \nScanOut30[0] , \nOut3_3[4] , \nOut3_15[4] , \nScanOut129[1] , 
        \nOut21_2[4] , \nScanOut449[0] , \nOut16_0[6] , \nOut3_16[7] , 
        \nOut3_0[7] , \nOut5_0[3] , \nOut28_4[3] , \nOut5_3[0] , \nOut6_29[3] , 
        \nOut9_1[2] , \nOut10_0[2] , \nOut17_20[6] , \nOut22_5[6] , 
        \nOut24_14[7] , \nOut24_5[2] , \nOut9_2[1] , \nScanOut319[3] , 
        \nScanOut679[2] , \nOut17_23[5] , \nOut22_6[5] , \nOut21_28[0] , 
        \nOut24_6[1] , \nScanOut519[7] , \nOut24_17[4] , \nOut28_18[1] , 
        \nScanOut918[6] , \nOut16_3[5] , \nOut28_7[0] , \nOut10_3[1] , 
        \nScanOut283[0] , \nOut30_23[1] , \nScanOut964[0] , \nScanOut33[3] , 
        \nOut1_19[6] , \nOut4_25[1] , \nOut10_10[3] , \nOut11_31[5] , 
        \nScanOut483[4] , \nOut19_20[2] , \nScanOut850[3] , \nOut23_24[2] , 
        \nScanOut1020[5] , \nScanOut131[3] , \nScanOut251[6] , 
        \nScanOut365[5] , \nScanOut605[4] , \nScanOut731[7] , \nScanOut882[5] , 
        \nScanOut451[2] , \nScanOut565[1] , \nScanOut732[4] , \nScanOut881[6] , 
        \nOut4_26[2] , \nOut8_29[7] , \nScanOut606[7] , \nScanOut132[0] , 
        \nScanOut252[5] , \nScanOut366[6] , \nScanOut452[1] , \nScanOut566[2] , 
        \nScanOut86[2] , \nScanOut280[3] , \nScanOut853[0] , \nScanOut967[3] , 
        \nOut30_20[2] , \nOut10_13[0] , \nScanOut480[7] , \nScanOut1023[6] , 
        \nOut19_23[1] , \nOut23_27[1] , \nOut26_18[5] , \nScanOut661[0] , 
        \nScanOut755[3] , \nScanOut1[6] , \nScanOut155[7] , \nScanOut235[2] , 
        \nScanOut301[1] , \nScanOut435[6] , \nOut20_11[4] , \nScanOut501[5] , 
        \nOut21_30[2] , \nOut29_21[5] , \nScanOut2[5] , \nScanOut54[4] , 
        \nOut13_25[5] , \nScanOut57[7] , \nScanOut187[1] , \nOut7_10[7] , 
        \nOut6_31[1] , \nScanOut787[5] , \nScanOut900[4] , \nScanOut834[7] , 
        \nOut7_13[4] , \nScanOut903[7] , \nScanOut85[1] , \nScanOut184[2] , 
        \nScanOut784[6] , \nScanOut837[4] , \nScanOut236[1] , \nScanOut302[2] , 
        \nScanOut156[4] , \nOut13_26[6] , \nScanOut662[3] , \nScanOut756[0] , 
        \nScanOut9[7] , \nOut0_9[3] , \nScanOut25[7] , \nScanOut41[3] , 
        \nScanOut93[5] , \nScanOut220[5] , \nScanOut314[6] , \nScanOut436[5] , 
        \nOut16_19[2] , \nOut20_12[7] , \nOut29_22[6] , \nScanOut502[6] , 
        \nScanOut140[0] , \nOut12_11[4] , \nOut13_30[2] , \nScanOut674[7] , 
        \nScanOut740[4] , \nOut28_15[4] , \nOut6_24[6] , \nScanOut420[1] , 
        \nScanOut514[2] , \nOut21_25[5] , \nScanOut915[3] , \nScanOut42[0] , 
        \nScanOut192[6] , \nScanOut792[2] , \nScanOut821[0] , \nOut28_9[6] , 
        \nOut3_18[1] , \nOut6_27[5] , \nScanOut791[1] , \nScanOut822[3] , 
        \nScanOut916[0] , \nScanOut90[6] , \nScanOut191[5] , \nScanOut143[3] , 
        \nScanOut223[6] , \nScanOut317[5] , \nScanOut677[4] , \nScanOut743[7] , 
        \nOut22_8[3] , \nScanOut423[2] , \nScanOut517[1] , \nOut21_26[6] , 
        \nOut24_8[7] , \nOut28_16[7] , \nOut12_12[7] , \nOut24_19[2] , 
        \nScanOut124[4] , \nOut4_30[6] , \nScanOut296[7] , \nScanOut845[4] , 
        \nScanOut971[7] , \nOut31_17[0] , \nOut11_24[2] , \nScanOut496[3] , 
        \nOut18_14[3] , \nOut22_10[3] , \nOut23_31[5] , \nScanOut610[3] , 
        \nScanOut724[0] , \nScanOut897[2] , \nOut5_11[0] , \nScanOut244[1] , 
        \nScanOut370[2] , \nScanOut444[5] , \nScanOut570[6] , \nScanOut127[7] , 
        \nOut5_12[3] , \nScanOut247[2] , \nScanOut373[1] , \nOut19_8[3] , 
        \nScanOut613[0] , \nScanOut727[3] , \nScanOut894[1] , \nScanOut295[4] , 
        \nScanOut447[6] , \nScanOut573[5] , \nOut31_14[3] , \nOut0_11[3] , 
        \nOut0_12[0] , \nScanOut19[3] , \nScanOut26[4] , \nScanOut972[4] , 
        \nOut1_2[7] , \nOut1_14[3] , \nOut2_21[5] , \nOut6_9[7] , 
        \nOut13_9[6] , \nScanOut846[7] , \nOut14_18[5] , \nOut15_9[2] , 
        \nOut18_17[0] , \nScanOut495[0] , \nOut22_13[0] , \nOut11_27[1] , 
        \nScanOut789[3] , \nOut2_22[6] , \nScanOut88[4] , \nScanOut189[7] , 
        \nScanOut158[2] , \nScanOut238[7] , \nOut16_14[7] , \nOut25_20[6] , 
        \nScanOut758[6] , \nOut13_28[0] , \nScanOut438[3] , \nOut16_17[4] , 
        \nOut25_23[5] , \nScanOut59[1] , \nOut8_24[2] , \nScanOut839[2] , 
        \nOut1_17[0] , \nOut15_21[1] , \nOut30_1[5] , \nOut15_22[2] , 
        \nOut23_29[7] , \nOut26_15[0] , \nOut26_16[3] , \nScanOut969[5] , 
        \nScanOut608[1] , \nOut4_28[4] , \nOut7_2[3] , \nOut8_27[1] , 
        \nScanOut368[0] , \nOut11_18[6] , \nOut14_2[6] , \nOut14_27[2] , 
        \nScanOut568[4] , \nOut30_2[6] , \nOut18_28[7] , \nScanOut1009[6] , 
        \nOut27_13[3] , \nOut12_2[2] , \nScanOut118[0] , \nScanOut879[0] , 
        \nScanOut278[5] , \nOut9_22[1] , \nScanOut478[1] , \nOut20_7[6] , 
        \nOut18_3[7] , \nScanOut718[4] , \nOut26_7[2] , \nOut20_4[5] , 
        \nOut26_4[1] , \nScanOut20[3] , \nScanOut23[0] , \nOut1_1[4] , 
        \nOut1_30[5] , \nOut7_1[0] , \nOut9_21[2] , \nOut18_0[4] , 
        \nOut27_10[0] , \nOut26_31[6] , \nOut12_1[1] , \nOut14_1[5] , 
        \nOut14_24[1] , \nOut31_28[7] , \nOut2_5[5] , \nOut2_6[6] , 
        \nOut8_7[3] , \nOut25_3[3] , \nOut11_6[3] , \nScanOut328[2] , 
        \nOut17_12[4] , \nOut21_19[1] , \nScanOut528[6] , \nScanOut648[3] , 
        \nOut24_26[5] , \nOut28_29[0] , \nOut23_3[7] , \nOut3_27[6] , 
        \nOut4_6[2] , \nOut6_18[2] , \nScanOut929[7] , \nOut29_2[2] , 
        \nOut17_6[7] , \nOut1_28[7] , \nOut3_24[5] , \nOut11_5[0] , 
        \nOut17_5[4] , \nOut4_5[1] , \nScanOut103[1] , \nOut8_4[0] , 
        \nOut16_30[1] , \nOut17_11[7] , \nScanOut699[6] , \nOut29_1[1] , 
        \nOut24_25[6] , \nOut25_0[0] , \nScanOut463[0] , \nOut23_0[4] , 
        \nScanOut557[3] , \nOut31_9[2] , \nScanOut703[5] , \nScanOut984[4] , 
        \nScanOut65[5] , \nScanOut66[6] , \nScanOut100[2] , \nOut4_17[3] , 
        \nOut8_18[6] , \nScanOut637[6] , \nScanOut357[7] , \nScanOut263[4] , 
        \nOut10_21[2] , \nOut10_22[1] , \nScanOut585[5] , \nOut26_29[4] , 
        \nScanOut1012[7] , \nScanOut385[1] , \nOut19_12[0] , \nOut23_16[0] , 
        \nScanOut862[1] , \nScanOut956[2] , \nOut18_30[5] , \nOut30_11[3] , 
        \nOut31_30[5] , \nOut19_11[3] , \nOut23_15[3] , \nScanOut1011[4] , 
        \nScanOut386[2] , \nScanOut586[6] , \nOut30_12[0] , \nScanOut861[2] , 
        \nScanOut955[1] , \nOut4_14[0] , \nScanOut354[4] , \nScanOut460[3] , 
        \nScanOut554[0] , \nOut7_22[5] , \nScanOut260[7] , \nScanOut634[5] , 
        \nScanOut700[6] , \nScanOut987[7] , \nScanOut932[6] , \nScanOut164[6] , 
        \nScanOut167[5] , \nOut13_17[7] , \nScanOut681[4] , \nScanOut806[5] , 
        \nScanOut207[0] , \nScanOut333[3] , \nScanOut407[4] , \nOut29_13[7] , 
        \nOut16_28[3] , \nScanOut533[7] , \nOut20_23[6] , \nScanOut404[7] , 
        \nScanOut653[2] , \nScanOut767[1] , \nScanOut530[4] , \nOut20_20[5] , 
        \nScanOut204[3] , \nScanOut330[0] , \nOut13_14[4] , \nOut29_10[4] , 
        \nOut28_31[2] , \nScanOut650[1] , \nScanOut764[2] , \nOut7_21[6] , 
        \nScanOut290[0] , \nOut11_22[5] , \nScanOut490[4] , \nOut18_12[4] , 
        \nScanOut682[7] , \nScanOut931[5] , \nOut22_16[4] , \nScanOut805[6] , 
        \nOut27_29[0] , \nOut30_30[1] , \nOut31_11[7] , \nOut0_28[3] , 
        \nScanOut122[3] , \nOut21_9[6] , \nScanOut843[3] , \nScanOut977[0] , 
        \nOut5_17[7] , \nOut9_18[2] , \nScanOut442[2] , \nScanOut576[1] , 
        \nScanOut242[6] , \nScanOut376[5] , \nScanOut722[7] , \nScanOut891[5] , 
        \nScanOut121[0] , \nScanOut441[1] , \nScanOut616[4] , \nOut27_9[2] , 
        \nScanOut575[2] , \nOut5_14[4] , \nScanOut615[7] , \nScanOut721[4] , 
        \nScanOut892[6] , \nScanOut241[5] , \nScanOut375[6] , \nOut11_21[6] , 
        \nScanOut493[7] , \nOut18_11[7] , \nOut19_30[1] , \nOut22_15[7] , 
        \nScanOut974[3] , \nOut0_30[1] , \nScanOut38[1] , \nOut1_12[4] , 
        \nScanOut44[7] , \nScanOut47[4] , \nOut3_8[6] , \nScanOut95[2] , 
        \nScanOut146[7] , \nOut9_9[3] , \nScanOut293[3] , \nScanOut840[0] , 
        \nOut31_12[4] , \nScanOut426[6] , \nOut17_28[7] , \nOut21_23[2] , 
        \nOut12_17[3] , \nScanOut512[5] , \nOut28_13[3] , \nScanOut226[2] , 
        \nScanOut312[1] , \nScanOut672[0] , \nScanOut746[3] , \nOut10_8[3] , 
        \nOut5_8[2] , \nOut6_22[1] , \nScanOut194[1] , \nScanOut913[4] , 
        \nScanOut197[2] , \nOut16_8[7] , \nScanOut794[5] , \nScanOut827[7] , 
        \nScanOut96[1] , \nScanOut145[4] , \nOut6_21[2] , \nScanOut797[6] , 
        \nScanOut824[4] , \nScanOut910[7] , \nOut28_10[0] , \nScanOut225[1] , 
        \nScanOut311[2] , \nOut12_14[0] , \nOut29_31[6] , \nScanOut425[5] , 
        \nScanOut511[6] , \nOut21_20[1] , \nScanOut139[2] , \nScanOut459[3] , 
        \nScanOut671[3] , \nScanOut745[0] , \nScanOut739[6] , \nOut30_7[2] , 
        \nOut8_22[5] , \nScanOut259[7] , \nOut10_18[2] , \nOut26_13[7] , 
        \nOut15_27[6] , \nOut19_28[3] , \nOut1_11[7] , \nOut8_21[6] , 
        \nScanOut288[2] , \nOut15_24[5] , \nScanOut858[2] , \nScanOut488[6] , 
        \nOut26_10[4] , \nOut27_31[2] , \nOut30_28[3] , \nOut30_4[1] , 
        \nScanOut889[7] , \nOut2_27[2] , \nOut7_18[6] , \nScanOut908[5] , 
        \nOut25_26[1] , \nOut29_29[4] , \nOut2_3[2] , \nOut2_24[1] , 
        \nScanOut309[0] , \nOut16_12[0] , \nScanOut509[4] , \nOut20_19[5] , 
        \nOut16_11[3] , \nScanOut669[1] , \nOut17_30[5] , \nOut25_25[2] , 
        \nOut2_0[1] , \nOut3_21[1] , \nOut8_1[4] , \nOut23_5[0] , 
        \nOut24_20[2] , \nOut25_5[4] , \nOut17_14[3] , \nOut4_0[5] , 
        \nOut17_0[0] , \nOut29_4[5] , \nScanOut78[3] , \nOut11_0[4] , 
        \nOut3_22[2] , \nOut4_3[6] , \nOut17_3[3] , \nScanOut818[0] , 
        \nOut29_7[6] , \nOut11_3[7] , \nScanOut179[0] , \nScanOut219[5] , 
        \nOut23_6[3] , \nScanOut779[4] , \nOut8_2[7] , \nScanOut419[1] , 
        \nOut17_17[0] , \nOut25_6[7] , \nOut12_4[5] , \nOut12_28[4] , 
        \nOut24_23[1] , \nScanOut11[2] , \nOut0_14[7] , \nOut1_4[0] , 
        \nScanOut398[7] , \nOut7_4[4] , \nScanOut598[3] , \nOut14_4[1] , 
        \nOut14_21[5] , \nOut27_15[4] , \nOut26_1[5] , \nScanOut999[2] , 
        \nOut0_17[4] , \nOut5_28[0] , \nOut9_24[6] , \nOut18_5[0] , 
        \nOut20_1[1] , \nOut9_27[5] , \nScanOut349[2] , \nOut18_6[3] , 
        \nScanOut629[3] , \nOut26_2[6] , \nOut1_7[3] , \nScanOut549[6] , 
        \nOut20_2[2] , \nOut2_18[5] , \nScanOut60[1] , \nOut7_7[7] , 
        \nOut12_7[6] , \nScanOut948[7] , \nOut14_7[2] , \nOut14_22[6] , 
        \nOut22_29[3] , \nOut27_16[7] , \nOut7_24[2] , \nScanOut934[1] , 
        \nScanOut161[2] , \nScanOut201[7] , \nScanOut335[4] , \nScanOut655[5] , 
        \nScanOut687[3] , \nScanOut800[2] , \nScanOut761[6] , \nOut12_30[6] , 
        \nScanOut401[3] , \nScanOut535[0] , \nOut20_25[1] , \nOut13_11[0] , 
        \nScanOut162[1] , \nScanOut202[4] , \nScanOut336[7] , \nOut29_15[0] , 
        \nScanOut656[6] , \nScanOut762[5] , \nOut13_12[3] , \nOut29_16[3] , 
        \nScanOut402[0] , \nOut25_19[6] , \nScanOut536[3] , \nOut20_26[2] , 
        \nScanOut63[2] , \nScanOut105[6] , \nOut4_11[4] , \nOut5_30[2] , 
        \nOut7_27[1] , \nScanOut684[0] , \nScanOut937[2] , \nScanOut803[1] , 
        \nScanOut351[0] , \nScanOut265[3] , \nScanOut631[1] , \nScanOut705[2] , 
        \nScanOut982[3] , \nScanOut106[5] , \nOut4_12[7] , \nOut10_24[6] , 
        \nScanOut383[6] , \nScanOut465[7] , \nScanOut551[4] , \nScanOut583[2] , 
        \nOut19_14[7] , \nOut23_10[7] , \nScanOut864[6] , \nOut30_17[4] , 
        \nScanOut950[5] , \nOut22_31[1] , \nScanOut1014[0] , \nOut10_27[5] , 
        \nScanOut380[5] , \nScanOut867[5] , \nScanOut953[6] , \nOut30_14[7] , 
        \nScanOut1017[3] , \nScanOut352[3] , \nOut15_18[1] , \nScanOut580[1] , 
        \nOut19_17[4] , \nOut23_13[4] , \nScanOut632[2] , \nScanOut706[1] , 
        \nScanOut981[0] , \nScanOut266[0] , \nScanOut466[4] , \nScanOut552[7] , 
        \nScanOut110[1] , \nOut5_25[5] , \nScanOut624[6] , \nScanOut710[5] , 
        \nScanOut997[4] , \nScanOut270[4] , \nScanOut344[7] , \nScanOut470[0] , 
        \nScanOut544[3] , \nScanOut945[2] , \nScanOut12[1] , \nOut1_9[5] , 
        \nOut11_10[7] , \nOut10_31[1] , \nScanOut396[1] , \nScanOut871[1] , 
        \nOut31_23[5] , \nScanOut1001[7] , \nScanOut596[5] , \nScanOut395[2] , 
        \nOut18_20[6] , \nOut22_24[6] , \nOut31_20[6] , \nOut0_19[2] , 
        \nOut5_26[6] , \nOut7_9[1] , \nOut11_13[4] , \nOut12_9[0] , 
        \nOut14_9[4] , \nOut18_23[5] , \nOut22_27[5] , \nScanOut872[2] , 
        \nScanOut946[1] , \nScanOut595[6] , \nScanOut1002[4] , \nOut27_18[1] , 
        \nOut9_29[3] , \nOut18_8[5] , \nScanOut273[7] , \nScanOut347[4] , 
        \nScanOut713[6] , \nScanOut994[7] , \nOut1_20[6] , \nScanOut75[6] , 
        \nScanOut113[2] , \nScanOut627[5] , \nScanOut473[3] , \nScanOut547[0] , 
        \nScanOut76[5] , \nOut6_10[3] , \nOut7_31[5] , \nOut6_13[0] , 
        \nScanOut174[5] , \nScanOut214[0] , \nScanOut320[3] , \nScanOut692[4] , 
        \nScanOut921[6] , \nScanOut815[5] , \nScanOut640[2] , \nScanOut774[1] , 
        \nScanOut177[6] , \nScanOut217[3] , \nScanOut323[0] , \nOut12_25[1] , 
        \nOut28_21[1] , \nScanOut414[4] , \nScanOut520[7] , \nOut20_30[6] , 
        \nOut21_11[0] , \nScanOut643[1] , \nScanOut777[2] , \nOut12_26[2] , 
        \nScanOut417[7] , \nOut17_19[6] , \nOut23_8[5] , \nOut25_8[1] , 
        \nScanOut523[4] , \nOut21_12[3] , \nOut28_22[2] , \nScanOut922[5] , 
        \nOut8_10[7] , \nOut15_15[4] , \nScanOut691[7] , \nScanOut816[6] , 
        \nOut29_9[0] , \nOut30_19[2] , \nOut26_21[5] , \nOut9_31[1] , 
        \nOut31_1[3] , \nOut1_23[5] , \nScanOut708[7] , \nScanOut108[3] , 
        \nOut8_13[4] , \nScanOut268[6] , \nScanOut468[2] , \nOut31_2[0] , 
        \nOut10_29[3] , \nScanOut869[3] , \nScanOut1019[5] , \nOut15_16[7] , 
        \nOut26_22[6] , \nOut19_19[2] , \nScanOut1[2] , \nOut0_1[2] , 
        \nOut0_2[1] , \nOut0_26[5] , \nOut2_15[0] , \nOut16_20[2] , 
        \nScanOut689[5] , \nOut25_14[3] , \nOut2_16[3] , \nScanOut49[2] , 
        \nOut3_6[0] , \nOut7_29[7] , \nOut10_6[5] , \nScanOut338[1] , 
        \nScanOut939[4] , \nOut16_23[1] , \nOut20_28[4] , \nScanOut658[0] , 
        \nOut25_17[0] , \nOut29_18[5] , \nScanOut538[5] , \nOut5_6[4] , 
        \nOut3_5[3] , \nOut3_13[3] , \nOut16_6[1] , \nScanOut829[1] , 
        \nOut28_2[4] , \nScanOut98[7] , \nScanOut148[1] , \nOut9_7[5] , 
        \nScanOut428[0] , \nOut17_26[1] , \nOut24_3[5] , \nScanOut228[4] , 
        \nOut12_19[5] , \nOut22_3[1] , \nScanOut748[5] , \nOut24_12[0] , 
        \nOut9_4[6] , \nOut17_25[2] , \nOut24_11[3] , \nOut25_30[5] , 
        \nOut24_0[6] , \nOut22_0[2] , \nOut3_10[0] , \nScanOut199[4] , 
        \nOut10_5[6] , \nOut16_5[2] , \nOut2_31[6] , \nOut5_5[7] , 
        \nOut5_19[1] , \nScanOut578[7] , \nOut21_7[0] , \nScanOut799[0] , 
        \nOut28_1[7] , \nOut9_16[4] , \nScanOut378[3] , \nOut19_3[1] , 
        \nScanOut618[2] , \nOut6_2[5] , \nOut14_13[7] , \nOut15_2[0] , 
        \nOut27_7[4] , \nOut22_18[2] , \nOut27_27[6] , \nOut6_1[6] , 
        \nOut13_2[4] , \nScanOut979[6] , \nOut13_1[7] , \nOut14_10[4] , 
        \nOut27_24[5] , \nOut15_1[3] , \nOut15_31[2] , \nScanOut2[1] , 
        \nScanOut4[2] , \nScanOut7[1] , \nOut0_25[6] , \nOut21_4[3] , 
        \nOut27_4[7] , \nScanOut153[0] , \nOut9_15[7] , \nOut19_0[2] , 
        \nOut29_27[2] , \nScanOut51[0] , \nScanOut52[3] , \nOut2_29[4] , 
        \nScanOut80[5] , \nScanOut233[5] , \nScanOut307[6] , \nOut13_23[2] , 
        \nOut25_28[7] , \nScanOut433[1] , \nOut20_17[3] , \nScanOut507[2] , 
        \nScanOut181[6] , \nScanOut667[7] , \nScanOut753[4] , \nScanOut182[5] , 
        \nOut7_16[0] , \nScanOut781[2] , \nScanOut906[3] , \nScanOut832[0] , 
        \nOut7_15[3] , \nScanOut905[0] , \nScanOut150[3] , \nOut13_20[1] , 
        \nScanOut430[2] , \nOut20_14[0] , \nScanOut782[1] , \nScanOut831[3] , 
        \nScanOut504[1] , \nOut0_9[7] , \nOut0_11[7] , \nOut1_1[0] , 
        \nScanOut35[4] , \nScanOut36[7] , \nScanOut83[6] , \nOut29_24[1] , 
        \nScanOut230[6] , \nScanOut304[5] , \nScanOut664[4] , \nScanOut750[7] , 
        \nOut10_16[4] , \nScanOut485[3] , \nOut15_29[0] , \nOut19_26[5] , 
        \nOut23_22[5] , \nScanOut962[7] , \nOut4_20[5] , \nOut4_23[6] , 
        \nScanOut137[4] , \nScanOut285[7] , \nScanOut856[4] , \nOut30_25[6] , 
        \nScanOut457[5] , \nScanOut563[6] , \nOut30_9[4] , \nScanOut603[3] , 
        \nScanOut737[0] , \nScanOut884[2] , \nScanOut134[7] , \nScanOut257[1] , 
        \nScanOut363[2] , \nScanOut454[6] , \nScanOut560[5] , \nScanOut254[2] , 
        \nScanOut360[1] , \nScanOut286[4] , \nOut10_15[7] , \nScanOut486[0] , 
        \nScanOut600[0] , \nScanOut734[3] , \nScanOut887[1] , \nOut19_25[6] , 
        \nOut23_21[6] , \nOut30_26[5] , \nOut1_28[3] , \nScanOut100[6] , 
        \nOut4_14[4] , \nScanOut354[0] , \nScanOut634[1] , \nScanOut700[2] , 
        \nScanOut855[7] , \nScanOut961[4] , \nScanOut987[3] , \nScanOut260[3] , 
        \nScanOut460[7] , \nScanOut554[4] , \nOut4_17[7] , \nOut8_18[2] , 
        \nOut10_21[6] , \nScanOut386[6] , \nScanOut861[6] , \nScanOut955[5] , 
        \nOut30_12[4] , \nScanOut586[2] , \nScanOut1011[0] , \nOut10_22[5] , 
        \nScanOut385[5] , \nOut18_30[1] , \nOut19_11[7] , \nOut23_15[7] , 
        \nOut19_12[4] , \nOut23_16[4] , \nScanOut862[5] , \nOut30_11[7] , 
        \nOut31_30[1] , \nScanOut956[6] , \nScanOut1012[3] , \nScanOut585[1] , 
        \nOut26_29[0] , \nScanOut357[3] , \nScanOut263[0] , \nScanOut703[1] , 
        \nScanOut984[0] , \nScanOut65[1] , \nScanOut103[5] , \nScanOut637[2] , 
        \nOut31_9[6] , \nScanOut463[4] , \nScanOut557[7] , \nScanOut66[2] , 
        \nScanOut164[2] , \nScanOut204[7] , \nOut7_21[2] , \nScanOut330[4] , 
        \nScanOut682[3] , \nScanOut931[1] , \nScanOut805[2] , \nScanOut650[5] , 
        \nScanOut764[6] , \nScanOut167[1] , \nScanOut207[4] , \nScanOut333[7] , 
        \nOut13_14[0] , \nOut29_10[0] , \nOut28_31[6] , \nScanOut404[3] , 
        \nScanOut530[0] , \nOut20_20[1] , \nScanOut653[6] , \nScanOut767[5] , 
        \nOut13_17[3] , \nScanOut407[0] , \nOut16_28[7] , \nOut20_23[2] , 
        \nScanOut533[3] , \nOut7_22[1] , \nOut29_13[3] , \nScanOut932[2] , 
        \nScanOut681[0] , \nScanOut806[1] , \nOut31_28[3] , \nOut7_1[4] , 
        \nOut12_1[5] , \nOut14_1[1] , \nOut14_24[5] , \nOut26_31[2] , 
        \nOut9_21[6] , \nOut18_0[0] , \nOut27_10[4] , \nOut26_4[5] , 
        \nOut0_12[4] , \nOut1_30[1] , \nOut20_4[1] , \nScanOut718[0] , 
        \nOut26_7[6] , \nScanOut19[7] , \nScanOut118[4] , \nScanOut278[1] , 
        \nOut9_22[5] , \nOut18_3[3] , \nScanOut478[5] , \nOut20_7[2] , 
        \nScanOut26[0] , \nOut1_2[3] , \nOut12_2[6] , \nScanOut879[4] , 
        \nOut2_5[1] , \nOut3_24[1] , \nOut4_5[5] , \nOut7_2[7] , 
        \nOut11_18[2] , \nOut27_13[7] , \nScanOut1009[2] , \nOut8_4[4] , 
        \nOut14_2[2] , \nOut14_27[6] , \nOut18_28[3] , \nOut16_30[5] , 
        \nOut17_11[3] , \nOut23_0[0] , \nOut25_0[4] , \nOut24_25[2] , 
        \nScanOut699[2] , \nOut29_1[5] , \nOut11_5[4] , \nOut17_5[0] , 
        \nOut2_6[2] , \nOut3_27[2] , \nOut17_6[3] , \nOut4_6[6] , 
        \nOut6_18[6] , \nScanOut929[3] , \nOut29_2[6] , \nScanOut41[7] , 
        \nScanOut42[4] , \nOut1_14[7] , \nOut1_17[4] , \nOut2_21[1] , 
        \nOut2_22[2] , \nScanOut59[5] , \nOut8_7[7] , \nOut11_6[7] , 
        \nScanOut328[6] , \nScanOut648[7] , \nOut23_3[3] , \nOut24_26[1] , 
        \nOut25_3[7] , \nOut28_29[4] , \nOut17_12[0] , \nScanOut528[2] , 
        \nOut21_19[5] , \nScanOut839[6] , \nScanOut88[0] , \nScanOut158[6] , 
        \nScanOut438[7] , \nOut16_17[0] , \nScanOut238[3] , \nOut13_28[4] , 
        \nOut25_23[1] , \nScanOut758[2] , \nOut16_14[3] , \nOut25_20[2] , 
        \nScanOut189[3] , \nOut4_28[0] , \nScanOut568[0] , \nScanOut789[7] , 
        \nOut30_2[2] , \nOut8_27[5] , \nScanOut368[4] , \nScanOut608[5] , 
        \nOut15_21[5] , \nOut15_22[6] , \nOut23_29[3] , \nOut26_15[4] , 
        \nOut26_16[7] , \nScanOut969[1] , \nOut30_1[1] , \nOut3_18[5] , 
        \nScanOut90[2] , \nScanOut143[7] , \nOut8_24[6] , \nOut28_16[3] , 
        \nScanOut223[2] , \nScanOut317[1] , \nOut12_12[3] , \nScanOut423[6] , 
        \nOut24_19[6] , \nScanOut517[5] , \nOut21_26[2] , \nOut22_8[7] , 
        \nOut24_8[3] , \nScanOut191[1] , \nScanOut677[0] , \nScanOut743[3] , 
        \nOut6_24[2] , \nOut6_27[1] , \nScanOut791[5] , \nOut28_9[2] , 
        \nScanOut192[2] , \nScanOut822[7] , \nScanOut916[4] , \nScanOut915[7] , 
        \nScanOut93[1] , \nScanOut140[4] , \nOut12_11[0] , \nOut13_30[6] , 
        \nScanOut420[5] , \nScanOut792[6] , \nScanOut821[4] , \nScanOut514[6] , 
        \nOut21_25[1] , \nOut28_15[0] , \nOut6_9[3] , \nScanOut220[1] , 
        \nScanOut314[2] , \nScanOut674[3] , \nScanOut740[0] , \nScanOut495[4] , 
        \nOut11_27[5] , \nOut14_18[1] , \nOut15_9[6] , \nOut18_17[4] , 
        \nOut22_13[4] , \nScanOut972[0] , \nScanOut295[0] , \nOut13_9[2] , 
        \nScanOut846[3] , \nOut31_14[7] , \nScanOut25[3] , \nScanOut124[0] , 
        \nScanOut127[3] , \nScanOut447[2] , \nScanOut573[1] , \nOut5_12[7] , 
        \nScanOut613[4] , \nScanOut727[7] , \nScanOut894[5] , \nScanOut247[6] , 
        \nScanOut373[5] , \nOut19_8[7] , \nOut4_30[2] , \nScanOut444[1] , 
        \nScanOut570[2] , \nOut5_11[4] , \nScanOut244[5] , \nScanOut370[6] , 
        \nScanOut296[3] , \nOut11_24[6] , \nScanOut496[7] , \nOut18_14[7] , 
        \nScanOut610[7] , \nScanOut724[4] , \nScanOut897[6] , \nOut22_10[7] , 
        \nOut23_31[1] , \nOut31_17[4] , \nScanOut30[4] , \nScanOut33[7] , 
        \nScanOut280[7] , \nOut10_13[4] , \nScanOut480[3] , \nOut19_23[5] , 
        \nOut23_27[5] , \nScanOut845[0] , \nScanOut971[3] , \nScanOut1023[2] , 
        \nOut26_18[1] , \nOut30_20[6] , \nOut1_19[2] , \nOut4_26[6] , 
        \nScanOut132[4] , \nScanOut853[4] , \nScanOut967[7] , \nOut8_29[3] , 
        \nScanOut452[5] , \nScanOut566[6] , \nScanOut252[1] , \nScanOut366[2] , 
        \nScanOut732[0] , \nScanOut881[2] , \nOut4_25[5] , \nScanOut131[7] , 
        \nScanOut451[6] , \nScanOut606[3] , \nScanOut565[5] , \nScanOut605[0] , 
        \nScanOut731[3] , \nScanOut882[1] , \nScanOut251[2] , \nScanOut365[1] , 
        \nOut10_10[7] , \nOut11_31[1] , \nScanOut483[0] , \nScanOut1020[1] , 
        \nOut19_20[6] , \nOut23_24[6] , \nScanOut964[4] , \nScanOut156[0] , 
        \nScanOut283[4] , \nScanOut850[7] , \nOut30_23[5] , \nOut13_26[2] , 
        \nScanOut436[1] , \nOut16_19[6] , \nOut20_12[3] , \nScanOut502[2] , 
        \nOut29_22[2] , \nScanOut54[0] , \nScanOut57[3] , \nScanOut85[5] , 
        \nScanOut184[6] , \nScanOut236[5] , \nScanOut302[6] , \nScanOut662[7] , 
        \nScanOut756[4] , \nOut7_13[0] , \nScanOut903[3] , \nScanOut187[5] , 
        \nScanOut784[2] , \nScanOut837[0] , \nScanOut155[3] , \nOut7_10[3] , 
        \nOut6_31[5] , \nScanOut787[1] , \nScanOut900[0] , \nScanOut834[3] , 
        \nOut13_25[1] , \nOut29_21[1] , \nScanOut435[2] , \nOut20_11[0] , 
        \nScanOut501[1] , \nOut21_30[6] , \nOut0_4[2] , \nOut0_7[1] , 
        \nOut0_23[5] , \nScanOut86[6] , \nScanOut235[6] , \nScanOut301[5] , 
        \nScanOut129[5] , \nScanOut449[4] , \nScanOut661[4] , \nScanOut755[7] , 
        \nOut21_2[0] , \nScanOut729[1] , \nScanOut28[6] , \nOut6_7[5] , 
        \nScanOut249[0] , \nOut9_13[4] , \nOut27_2[4] , \nOut19_6[1] , 
        \nOut11_29[3] , \nOut14_16[7] , \nOut27_22[6] , \nOut15_7[0] , 
        \nOut18_19[2] , \nOut13_7[4] , \nScanOut848[5] , \nOut6_4[6] , 
        \nOut14_15[4] , \nOut15_4[3] , \nScanOut498[1] , \nScanOut298[5] , 
        \nOut27_21[5] , \nOut31_19[2] , \nScanOut14[2] , \nOut0_20[6] , 
        \nOut9_10[7] , \nOut13_4[7] , \nOut21_1[3] , \nOut8_31[1] , 
        \nOut19_5[2] , \nOut27_1[7] , \nScanOut899[0] , \nOut2_8[4] , 
        \nOut2_10[0] , \nOut3_3[0] , \nOut3_15[0] , \nOut3_16[3] , 
        \nOut10_3[5] , \nOut16_3[1] , \nOut3_0[3] , \nOut5_3[4] , 
        \nOut6_29[7] , \nScanOut918[2] , \nOut9_1[6] , \nOut9_2[5] , 
        \nOut17_23[1] , \nOut21_28[4] , \nOut24_17[0] , \nOut28_7[4] , 
        \nOut28_18[5] , \nOut24_6[5] , \nScanOut319[7] , \nScanOut519[3] , 
        \nOut17_20[2] , \nOut22_6[1] , \nScanOut679[6] , \nOut24_5[6] , 
        \nOut10_0[6] , \nOut22_5[2] , \nOut24_14[3] , \nOut5_0[7] , 
        \nOut16_0[2] , \nOut28_4[7] , \nOut16_25[2] , \nOut24_30[5] , 
        \nOut25_11[3] , \nOut2_13[3] , \nScanOut68[4] , \nOut3_31[6] , 
        \nScanOut808[7] , \nOut1_25[6] , \nScanOut169[7] , \nScanOut209[2] , 
        \nScanOut769[3] , \nScanOut409[6] , \nOut16_26[1] , \nScanOut388[0] , 
        \nOut13_19[5] , \nOut25_12[0] , \nOut15_10[4] , \nScanOut588[4] , 
        \nOut26_24[5] , \nOut14_31[2] , \nScanOut989[5] , \nOut1_26[5] , 
        \nOut4_19[1] , \nOut8_15[7] , \nScanOut359[5] , \nOut31_4[3] , 
        \nOut8_16[4] , \nScanOut639[4] , \nScanOut70[6] , \nOut6_15[3] , 
        \nOut15_13[7] , \nScanOut559[1] , \nOut31_7[0] , \nOut23_18[2] , 
        \nScanOut958[0] , \nOut26_27[6] , \nScanOut924[6] , \nScanOut73[5] , 
        \nOut3_29[4] , \nScanOut171[5] , \nScanOut211[0] , \nScanOut325[3] , 
        \nScanOut645[2] , \nScanOut697[4] , \nScanOut810[5] , \nScanOut771[1] , 
        \nOut12_20[1] , \nScanOut411[4] , \nScanOut525[7] , \nOut21_14[0] , 
        \nScanOut172[6] , \nScanOut212[3] , \nScanOut326[0] , \nOut28_24[1] , 
        \nScanOut646[1] , \nScanOut772[2] , \nOut8_9[1] , \nOut12_23[2] , 
        \nOut24_28[7] , \nOut28_27[2] , \nScanOut412[7] , \nOut21_17[3] , 
        \nOut17_8[5] , \nScanOut526[4] , \nOut4_8[0] , \nOut6_16[0] , 
        \nScanOut927[5] , \nScanOut694[7] , \nScanOut813[6] , \nScanOut115[1] , 
        \nOut5_20[5] , \nOut11_8[1] , \nScanOut275[4] , \nScanOut341[7] , 
        \nScanOut621[6] , \nScanOut715[5] , \nScanOut992[4] , \nScanOut393[1] , 
        \nScanOut475[0] , \nScanOut541[3] , \nOut31_26[5] , \nScanOut17[1] , 
        \nOut11_15[7] , \nOut18_25[6] , \nOut22_21[6] , \nScanOut874[1] , 
        \nScanOut940[2] , \nScanOut593[5] , \nScanOut1004[7] , 
        \nScanOut943[1] , \nScanOut390[2] , \nScanOut877[2] , \nOut31_25[6] , 
        \nScanOut590[6] , \nScanOut1007[4] , \nOut11_16[4] , \nOut14_29[0] , 
        \nOut18_26[5] , \nOut22_22[5] , \nOut0_1[6] , \nScanOut4[6] , 
        \nScanOut83[2] , \nScanOut116[2] , \nOut5_23[6] , \nScanOut622[5] , 
        \nScanOut716[6] , \nOut26_9[0] , \nScanOut991[7] , \nScanOut276[7] , 
        \nScanOut342[4] , \nScanOut476[3] , \nScanOut542[0] , \nOut20_9[4] , 
        \nScanOut230[2] , \nScanOut304[1] , \nScanOut150[7] , \nOut13_20[5] , 
        \nScanOut664[0] , \nScanOut750[3] , \nOut29_24[5] , \nScanOut7[5] , 
        \nScanOut51[4] , \nOut7_15[7] , \nScanOut430[6] , \nOut20_14[4] , 
        \nScanOut504[5] , \nScanOut905[4] , \nScanOut52[7] , \nScanOut182[1] , 
        \nScanOut782[5] , \nScanOut831[7] , \nOut2_29[0] , \nOut7_16[4] , 
        \nScanOut781[6] , \nScanOut906[7] , \nScanOut832[4] , \nScanOut80[1] , 
        \nScanOut181[2] , \nScanOut153[4] , \nScanOut233[1] , \nScanOut307[2] , 
        \nScanOut667[3] , \nScanOut753[0] , \nScanOut433[5] , \nOut20_17[7] , 
        \nScanOut507[6] , \nOut0_25[2] , \nScanOut35[0] , \nOut13_23[6] , 
        \nOut29_27[6] , \nOut25_28[3] , \nScanOut36[3] , \nOut4_20[1] , 
        \nScanOut286[0] , \nScanOut855[3] , \nScanOut961[0] , \nOut30_26[1] , 
        \nOut10_15[3] , \nScanOut486[4] , \nScanOut600[4] , \nOut19_25[2] , 
        \nOut23_21[2] , \nScanOut734[7] , \nScanOut887[5] , \nOut4_23[2] , 
        \nScanOut134[3] , \nScanOut254[6] , \nScanOut360[5] , \nScanOut454[2] , 
        \nScanOut560[1] , \nScanOut137[0] , \nScanOut257[5] , \nScanOut363[6] , 
        \nScanOut603[7] , \nScanOut737[4] , \nScanOut884[6] , \nOut30_9[0] , 
        \nScanOut285[3] , \nScanOut457[1] , \nScanOut563[2] , \nOut30_25[2] , 
        \nScanOut962[3] , \nScanOut49[6] , \nOut3_5[7] , \nOut3_10[4] , 
        \nOut5_5[3] , \nOut10_16[0] , \nOut15_29[4] , \nOut19_26[1] , 
        \nScanOut856[0] , \nOut23_22[1] , \nScanOut485[7] , \nOut16_5[6] , 
        \nScanOut799[4] , \nOut28_1[3] , \nOut2_31[2] , \nOut10_5[2] , 
        \nOut3_13[7] , \nScanOut98[3] , \nScanOut199[0] , \nScanOut148[5] , 
        \nScanOut228[0] , \nOut9_4[2] , \nOut17_25[6] , \nOut22_0[6] , 
        \nOut24_0[2] , \nOut22_3[5] , \nOut24_11[7] , \nOut25_30[1] , 
        \nScanOut748[1] , \nOut9_7[1] , \nOut12_19[1] , \nOut24_12[4] , 
        \nScanOut428[4] , \nOut17_26[5] , \nOut24_3[1] , \nOut16_6[5] , 
        \nOut5_6[0] , \nOut28_2[0] , \nOut3_6[4] , \nScanOut829[5] , 
        \nOut9_15[3] , \nOut10_6[1] , \nOut19_0[6] , \nOut21_4[7] , 
        \nOut27_4[3] , \nOut0_2[5] , \nOut6_1[2] , \nOut13_1[3] , 
        \nOut14_10[0] , \nOut15_1[7] , \nOut15_31[6] , \nOut13_2[0] , 
        \nOut27_24[1] , \nScanOut979[2] , \nOut0_26[1] , \nOut6_2[1] , 
        \nOut14_13[3] , \nOut15_2[4] , \nOut27_27[2] , \nScanOut618[6] , 
        \nOut22_18[6] , \nOut27_7[0] , \nOut1_23[1] , \nScanOut108[7] , 
        \nOut5_19[5] , \nOut9_16[0] , \nScanOut378[7] , \nOut10_29[7] , 
        \nOut15_16[3] , \nScanOut578[3] , \nOut19_3[5] , \nOut21_7[4] , 
        \nOut19_19[6] , \nOut26_22[2] , \nScanOut1019[1] , \nScanOut869[7] , 
        \nOut31_2[4] , \nOut8_13[0] , \nScanOut468[6] , \nScanOut268[2] , 
        \nScanOut708[3] , \nOut31_1[7] , \nOut2_15[4] , \nOut2_16[7] , 
        \nOut1_20[2] , \nOut7_29[3] , \nOut8_10[3] , \nOut9_31[5] , 
        \nScanOut338[5] , \nOut15_15[0] , \nOut26_21[1] , \nOut16_23[5] , 
        \nOut30_19[6] , \nScanOut538[1] , \nOut20_28[0] , \nScanOut658[4] , 
        \nOut25_17[4] , \nOut29_18[1] , \nScanOut939[0] , \nOut16_20[6] , 
        \nScanOut689[1] , \nOut25_14[7] , \nScanOut11[6] , \nScanOut12[5] , 
        \nOut0_19[6] , \nScanOut113[6] , \nScanOut473[7] , \nScanOut547[4] , 
        \nScanOut713[2] , \nScanOut994[3] , \nOut5_26[2] , \nOut9_29[7] , 
        \nOut18_8[1] , \nScanOut627[1] , \nOut7_9[5] , \nScanOut273[3] , 
        \nScanOut347[0] , \nOut11_13[0] , \nScanOut595[2] , \nScanOut1002[0] , 
        \nOut12_9[4] , \nOut14_9[0] , \nOut18_23[1] , \nOut22_27[1] , 
        \nOut27_18[5] , \nOut1_9[1] , \nScanOut395[6] , \nScanOut872[6] , 
        \nScanOut946[5] , \nOut11_10[3] , \nOut10_31[5] , \nOut18_20[2] , 
        \nOut31_20[2] , \nScanOut596[1] , \nOut22_24[2] , \nScanOut1001[3] , 
        \nScanOut396[5] , \nOut31_23[1] , \nScanOut945[6] , \nOut0_14[3] , 
        \nOut0_17[0] , \nOut2_3[6] , \nOut2_18[1] , \nScanOut63[6] , 
        \nScanOut75[2] , \nScanOut76[1] , \nScanOut110[5] , \nScanOut871[5] , 
        \nOut5_25[1] , \nScanOut470[4] , \nScanOut544[7] , \nOut6_13[4] , 
        \nScanOut270[0] , \nScanOut344[3] , \nScanOut624[2] , \nScanOut710[1] , 
        \nScanOut997[0] , \nScanOut922[1] , \nScanOut174[1] , \nScanOut177[2] , 
        \nOut12_26[6] , \nScanOut691[3] , \nScanOut816[2] , \nOut29_9[4] , 
        \nScanOut217[7] , \nScanOut323[4] , \nScanOut417[3] , \nOut25_8[5] , 
        \nOut28_22[6] , \nScanOut523[0] , \nOut17_19[2] , \nOut21_12[7] , 
        \nScanOut414[0] , \nScanOut643[5] , \nOut23_8[1] , \nScanOut777[6] , 
        \nScanOut520[3] , \nOut20_30[2] , \nOut21_11[4] , \nScanOut214[4] , 
        \nScanOut320[7] , \nOut12_25[5] , \nOut28_21[5] , \nScanOut640[6] , 
        \nScanOut774[5] , \nOut6_10[7] , \nOut7_31[1] , \nScanOut692[0] , 
        \nScanOut921[2] , \nScanOut815[1] , \nOut7_27[5] , \nScanOut684[4] , 
        \nScanOut937[6] , \nScanOut803[5] , \nScanOut60[5] , \nScanOut161[6] , 
        \nScanOut162[5] , \nScanOut402[4] , \nScanOut536[7] , \nOut20_26[6] , 
        \nScanOut202[0] , \nScanOut336[3] , \nOut13_12[7] , \nOut25_19[2] , 
        \nOut29_16[7] , \nScanOut656[2] , \nScanOut762[1] , \nOut12_30[2] , 
        \nOut13_11[4] , \nScanOut201[3] , \nScanOut335[0] , \nScanOut401[7] , 
        \nOut29_15[4] , \nScanOut535[4] , \nOut20_25[5] , \nOut7_24[6] , 
        \nScanOut655[1] , \nScanOut761[2] , \nScanOut934[5] , \nScanOut105[2] , 
        \nScanOut106[1] , \nScanOut687[7] , \nScanOut800[6] , \nOut4_12[3] , 
        \nScanOut352[7] , \nScanOut466[0] , \nScanOut552[3] , \nScanOut266[4] , 
        \nOut10_24[2] , \nOut10_27[1] , \nOut15_18[5] , \nOut19_17[0] , 
        \nScanOut632[6] , \nScanOut706[5] , \nScanOut981[4] , \nScanOut580[5] , 
        \nOut23_13[0] , \nScanOut1017[7] , \nScanOut380[1] , \nOut30_14[3] , 
        \nScanOut867[1] , \nScanOut953[2] , \nScanOut1014[4] , 
        \nScanOut383[2] , \nScanOut583[6] , \nOut19_14[3] , \nOut23_10[3] , 
        \nOut22_31[5] , \nScanOut864[2] , \nScanOut950[1] , \nScanOut465[3] , 
        \nOut30_17[0] , \nScanOut551[0] , \nOut4_11[0] , \nOut5_30[6] , 
        \nScanOut631[5] , \nScanOut705[6] , \nScanOut982[7] , \nScanOut351[4] , 
        \nScanOut179[4] , \nScanOut265[7] , \nScanOut219[1] , \nOut8_2[3] , 
        \nOut12_28[0] , \nScanOut419[5] , \nOut24_23[5] , \nOut17_17[4] , 
        \nOut25_6[3] , \nOut23_6[7] , \nScanOut779[0] , \nOut1_7[7] , 
        \nOut2_0[5] , \nScanOut78[7] , \nOut3_22[6] , \nOut11_3[3] , 
        \nOut17_3[7] , \nOut4_3[2] , \nOut11_0[0] , \nScanOut818[4] , 
        \nOut29_7[2] , \nOut3_21[5] , \nOut4_0[1] , \nOut17_0[4] , 
        \nOut29_4[1] , \nOut7_7[3] , \nOut8_1[0] , \nOut25_5[0] , 
        \nOut17_14[7] , \nOut23_5[4] , \nOut24_20[6] , \nOut12_7[2] , 
        \nOut14_7[6] , \nOut14_22[2] , \nOut22_29[7] , \nOut27_16[3] , 
        \nScanOut948[3] , \nScanOut549[2] , \nOut20_2[6] , \nScanOut629[7] , 
        \nOut26_2[2] , \nOut5_28[4] , \nOut9_24[2] , \nOut9_27[1] , 
        \nScanOut349[6] , \nOut18_6[7] , \nOut18_5[4] , \nOut20_1[5] , 
        \nOut26_1[1] , \nScanOut999[6] , \nOut1_4[4] , \nOut7_4[0] , 
        \nOut14_4[5] , \nOut14_21[1] , \nScanOut598[7] , \nOut27_15[0] , 
        \nScanOut398[3] , \nOut12_4[1] , \nScanOut9[3] , \nOut0_30[5] , 
        \nOut1_11[3] , \nScanOut889[3] , \nScanOut38[5] , \nOut8_21[2] , 
        \nScanOut288[6] , \nOut30_4[5] , \nOut30_28[7] , \nOut15_24[1] , 
        \nScanOut488[2] , \nOut26_10[0] , \nOut27_31[6] , \nOut1_12[0] , 
        \nOut8_22[1] , \nOut10_18[6] , \nOut15_27[2] , \nScanOut858[6] , 
        \nOut19_28[7] , \nOut26_13[3] , \nScanOut259[3] , \nScanOut739[2] , 
        \nOut2_24[5] , \nScanOut139[6] , \nScanOut459[7] , \nOut30_7[6] , 
        \nScanOut309[4] , \nOut16_11[7] , \nOut25_25[6] , \nOut17_30[1] , 
        \nScanOut669[5] , \nOut16_12[4] , \nOut20_19[1] , \nScanOut509[0] , 
        \nOut25_26[5] , \nScanOut20[7] , \nOut2_27[6] , \nOut7_18[2] , 
        \nScanOut908[1] , \nOut29_29[0] , \nScanOut293[7] , \nOut31_12[0] , 
        \nScanOut974[7] , \nScanOut23[4] , \nOut0_28[7] , \nScanOut121[4] , 
        \nOut5_14[0] , \nOut11_21[2] , \nScanOut493[3] , \nOut18_11[3] , 
        \nOut19_30[5] , \nScanOut840[4] , \nOut22_15[3] , \nScanOut241[1] , 
        \nScanOut375[2] , \nScanOut615[3] , \nScanOut721[0] , \nScanOut892[2] , 
        \nScanOut441[5] , \nScanOut575[6] , \nScanOut722[3] , \nOut27_9[6] , 
        \nScanOut891[1] , \nScanOut122[7] , \nOut5_17[3] , \nOut9_18[6] , 
        \nScanOut616[0] , \nScanOut242[2] , \nScanOut376[1] , \nScanOut442[6] , 
        \nScanOut576[5] , \nOut21_9[2] , \nOut1_4[6] , \nOut2_3[4] , 
        \nScanOut44[3] , \nScanOut96[5] , \nScanOut290[4] , \nScanOut843[7] , 
        \nScanOut977[4] , \nOut30_30[5] , \nOut31_11[3] , \nOut11_22[1] , 
        \nScanOut490[0] , \nOut27_29[4] , \nOut18_12[0] , \nOut22_16[0] , 
        \nScanOut145[0] , \nScanOut225[5] , \nScanOut311[6] , \nScanOut671[7] , 
        \nScanOut745[4] , \nScanOut425[1] , \nScanOut511[2] , \nOut21_20[5] , 
        \nOut28_10[4] , \nOut12_14[4] , \nOut29_31[2] , \nScanOut47[0] , 
        \nOut5_8[6] , \nOut6_21[6] , \nScanOut797[2] , \nOut6_22[5] , 
        \nScanOut197[6] , \nScanOut824[0] , \nScanOut910[3] , \nOut16_8[3] , 
        \nScanOut913[0] , \nOut2_18[3] , \nScanOut60[7] , \nOut3_8[2] , 
        \nScanOut794[1] , \nScanOut827[3] , \nScanOut95[6] , \nScanOut194[5] , 
        \nScanOut226[6] , \nOut10_8[7] , \nScanOut312[5] , \nScanOut146[3] , 
        \nOut12_17[7] , \nScanOut672[4] , \nScanOut746[7] , \nOut28_13[7] , 
        \nOut7_24[4] , \nOut9_9[7] , \nScanOut426[2] , \nOut17_28[3] , 
        \nOut21_23[6] , \nScanOut512[1] , \nScanOut687[5] , \nScanOut800[4] , 
        \nScanOut934[7] , \nScanOut63[4] , \nScanOut161[4] , \nScanOut201[1] , 
        \nScanOut335[2] , \nOut12_30[0] , \nOut13_11[6] , \nScanOut655[3] , 
        \nScanOut761[0] , \nOut29_15[6] , \nScanOut162[7] , \nScanOut202[2] , 
        \nScanOut401[5] , \nScanOut535[6] , \nOut20_25[7] , \nScanOut656[0] , 
        \nScanOut762[3] , \nScanOut336[1] , \nScanOut402[6] , \nScanOut536[5] , 
        \nOut20_26[4] , \nOut29_16[5] , \nOut13_12[5] , \nScanOut684[6] , 
        \nOut25_19[0] , \nScanOut803[7] , \nOut7_27[7] , \nScanOut937[4] , 
        \nOut2_0[7] , \nOut3_21[7] , \nScanOut105[0] , \nOut4_11[2] , 
        \nScanOut265[5] , \nScanOut631[7] , \nScanOut705[4] , \nScanOut982[5] , 
        \nOut5_30[4] , \nScanOut351[6] , \nScanOut465[1] , \nScanOut551[2] , 
        \nScanOut106[3] , \nOut4_12[1] , \nScanOut266[6] , \nOut10_24[0] , 
        \nScanOut383[0] , \nScanOut864[0] , \nScanOut950[3] , \nScanOut583[4] , 
        \nOut30_17[2] , \nOut10_27[3] , \nScanOut380[3] , \nOut19_14[1] , 
        \nOut23_10[1] , \nOut22_31[7] , \nScanOut1014[6] , \nOut30_14[1] , 
        \nOut15_18[7] , \nOut19_17[2] , \nScanOut867[3] , \nScanOut953[0] , 
        \nOut23_13[2] , \nScanOut580[7] , \nScanOut1017[5] , \nScanOut352[5] , 
        \nScanOut632[4] , \nScanOut706[7] , \nScanOut981[6] , \nOut4_0[3] , 
        \nOut8_1[2] , \nScanOut466[2] , \nScanOut552[1] , \nOut23_5[6] , 
        \nOut17_14[5] , \nOut25_5[2] , \nOut24_20[4] , \nOut29_4[3] , 
        \nOut11_0[2] , \nOut17_0[6] , \nScanOut78[5] , \nOut3_22[4] , 
        \nOut17_3[5] , \nOut4_3[0] , \nOut29_7[0] , \nScanOut818[6] , 
        \nScanOut179[6] , \nScanOut219[3] , \nOut11_3[1] , \nOut23_6[5] , 
        \nScanOut779[2] , \nOut8_2[1] , \nOut12_28[2] , \nOut24_23[7] , 
        \nScanOut419[7] , \nOut17_17[6] , \nOut25_6[1] , \nScanOut398[1] , 
        \nOut0_1[4] , \nOut0_2[7] , \nScanOut4[4] , \nScanOut7[7] , 
        \nScanOut9[1] , \nOut0_14[1] , \nOut7_4[2] , \nOut12_4[3] , 
        \nOut14_4[7] , \nOut14_21[3] , \nOut9_24[0] , \nScanOut598[5] , 
        \nOut27_15[2] , \nOut18_5[6] , \nOut0_17[2] , \nOut20_1[7] , 
        \nOut26_1[3] , \nScanOut999[4] , \nScanOut629[5] , \nOut0_30[7] , 
        \nScanOut38[7] , \nOut1_7[5] , \nOut5_28[6] , \nScanOut349[4] , 
        \nOut26_2[0] , \nOut9_27[3] , \nOut12_7[0] , \nScanOut549[0] , 
        \nOut18_6[5] , \nOut20_2[4] , \nScanOut948[1] , \nOut1_12[2] , 
        \nScanOut139[4] , \nOut7_7[1] , \nOut27_16[1] , \nOut14_7[4] , 
        \nOut14_22[0] , \nOut22_29[5] , \nOut8_22[3] , \nScanOut259[1] , 
        \nScanOut459[5] , \nOut30_7[4] , \nOut10_18[4] , \nOut15_27[0] , 
        \nScanOut739[0] , \nOut19_28[5] , \nOut26_13[1] , \nScanOut858[4] , 
        \nScanOut288[4] , \nOut15_24[3] , \nScanOut488[0] , \nOut26_10[2] , 
        \nOut27_31[4] , \nOut30_4[7] , \nOut30_28[5] , \nOut1_11[1] , 
        \nOut2_27[4] , \nOut7_18[0] , \nOut8_21[0] , \nScanOut889[1] , 
        \nScanOut908[3] , \nOut16_12[6] , \nScanOut509[2] , \nOut20_19[3] , 
        \nOut25_26[7] , \nOut29_29[2] , \nScanOut20[5] , \nScanOut23[6] , 
        \nOut2_24[7] , \nScanOut309[6] , \nScanOut669[7] , \nOut16_11[5] , 
        \nOut17_30[3] , \nOut25_25[4] , \nOut11_22[3] , \nScanOut490[2] , 
        \nOut27_29[6] , \nOut18_12[2] , \nOut22_16[2] , \nScanOut843[5] , 
        \nOut0_28[5] , \nScanOut122[5] , \nScanOut290[6] , \nScanOut977[6] , 
        \nScanOut442[4] , \nScanOut576[7] , \nOut30_30[7] , \nOut31_11[1] , 
        \nOut21_9[0] , \nScanOut121[6] , \nOut5_17[1] , \nScanOut242[0] , 
        \nScanOut616[2] , \nOut27_9[4] , \nScanOut891[3] , \nScanOut722[1] , 
        \nOut9_18[4] , \nScanOut376[3] , \nOut5_14[2] , \nScanOut241[3] , 
        \nScanOut441[7] , \nScanOut575[4] , \nScanOut375[0] , \nScanOut293[5] , 
        \nOut11_21[0] , \nOut18_11[1] , \nScanOut615[1] , \nScanOut721[2] , 
        \nScanOut892[0] , \nOut19_30[7] , \nOut22_15[1] , \nScanOut493[1] , 
        \nScanOut840[6] , \nOut31_12[2] , \nScanOut974[5] , \nScanOut44[1] , 
        \nScanOut47[2] , \nOut3_8[0] , \nScanOut95[4] , \nScanOut146[1] , 
        \nOut12_17[5] , \nScanOut226[4] , \nOut9_9[5] , \nOut28_13[5] , 
        \nScanOut426[0] , \nScanOut512[3] , \nOut21_23[4] , \nOut17_28[1] , 
        \nScanOut312[7] , \nScanOut672[6] , \nScanOut746[5] , \nScanOut194[7] , 
        \nOut6_22[7] , \nOut10_8[5] , \nOut16_8[1] , \nScanOut827[1] , 
        \nScanOut913[2] , \nScanOut794[3] , \nOut5_8[4] , \nScanOut197[4] , 
        \nScanOut797[0] , \nScanOut824[2] , \nScanOut96[7] , \nScanOut145[2] , 
        \nOut6_21[4] , \nScanOut910[1] , \nScanOut425[3] , \nScanOut511[0] , 
        \nOut21_20[7] , \nOut29_31[0] , \nOut12_14[6] , \nOut28_10[6] , 
        \nScanOut671[5] , \nScanOut745[6] , \nScanOut225[7] , \nScanOut311[4] , 
        \nScanOut433[7] , \nScanOut507[4] , \nOut20_17[5] , \nOut29_27[4] , 
        \nScanOut51[6] , \nScanOut52[5] , \nScanOut80[3] , \nScanOut153[6] , 
        \nOut13_23[4] , \nOut25_28[1] , \nScanOut667[1] , \nScanOut753[2] , 
        \nScanOut181[0] , \nScanOut233[3] , \nScanOut307[0] , \nScanOut781[4] , 
        \nScanOut832[6] , \nOut2_29[2] , \nOut7_16[6] , \nScanOut906[5] , 
        \nScanOut182[3] , \nOut7_15[5] , \nScanOut831[5] , \nScanOut782[7] , 
        \nScanOut905[6] , \nOut13_20[7] , \nOut0_26[3] , \nScanOut35[2] , 
        \nScanOut36[1] , \nScanOut83[0] , \nScanOut150[5] , \nOut29_24[7] , 
        \nScanOut230[0] , \nScanOut430[4] , \nScanOut504[7] , \nOut20_14[6] , 
        \nScanOut304[3] , \nScanOut664[2] , \nScanOut750[1] , \nScanOut285[1] , 
        \nOut10_16[2] , \nOut15_29[6] , \nOut19_26[3] , \nOut23_22[3] , 
        \nScanOut485[5] , \nScanOut856[2] , \nOut30_25[0] , \nScanOut962[1] , 
        \nOut4_20[3] , \nOut4_23[0] , \nScanOut137[2] , \nOut30_9[2] , 
        \nScanOut257[7] , \nScanOut457[3] , \nScanOut563[0] , \nScanOut363[4] , 
        \nScanOut134[1] , \nScanOut454[0] , \nScanOut560[3] , \nScanOut603[5] , 
        \nScanOut737[6] , \nScanOut884[4] , \nScanOut254[4] , \nScanOut600[6] , 
        \nScanOut887[7] , \nScanOut734[5] , \nScanOut360[7] , \nOut10_15[1] , 
        \nScanOut486[6] , \nOut19_25[0] , \nOut23_21[0] , \nScanOut855[1] , 
        \nScanOut49[4] , \nOut3_6[6] , \nScanOut286[2] , \nScanOut961[2] , 
        \nOut30_26[3] , \nOut3_13[5] , \nOut10_6[3] , \nOut16_6[7] , 
        \nScanOut829[7] , \nOut3_5[5] , \nScanOut98[1] , \nOut5_6[2] , 
        \nOut28_2[2] , \nScanOut148[7] , \nScanOut228[2] , \nOut9_7[3] , 
        \nOut12_19[3] , \nOut24_12[6] , \nScanOut428[6] , \nOut24_3[3] , 
        \nOut17_26[7] , \nOut9_4[0] , \nOut22_3[7] , \nScanOut748[3] , 
        \nOut17_25[4] , \nOut24_0[0] , \nOut24_11[5] , \nOut25_30[3] , 
        \nScanOut199[2] , \nOut10_5[0] , \nOut22_0[4] , \nOut3_10[6] , 
        \nOut2_31[0] , \nOut5_5[1] , \nScanOut799[6] , \nOut28_1[1] , 
        \nOut16_5[4] , \nScanOut578[1] , \nScanOut618[4] , \nOut21_7[6] , 
        \nOut5_19[7] , \nScanOut378[5] , \nOut19_3[7] , \nOut27_7[2] , 
        \nOut6_2[3] , \nOut9_16[2] , \nOut27_27[0] , \nOut13_2[2] , 
        \nOut14_13[1] , \nOut15_2[6] , \nOut22_18[4] , \nScanOut979[0] , 
        \nOut6_1[0] , \nOut14_10[2] , \nOut15_31[4] , \nOut15_1[5] , 
        \nOut27_24[3] , \nOut0_25[0] , \nOut9_15[1] , \nOut13_1[1] , 
        \nOut19_0[4] , \nOut21_4[5] , \nOut27_4[1] , \nOut1_20[0] , 
        \nOut15_15[2] , \nOut26_21[3] , \nOut30_19[4] , \nOut8_10[1] , 
        \nOut9_31[7] , \nOut1_23[3] , \nOut8_13[2] , \nScanOut268[0] , 
        \nOut31_1[5] , \nScanOut108[5] , \nScanOut708[1] , \nOut10_29[5] , 
        \nOut15_16[1] , \nScanOut468[4] , \nOut31_2[6] , \nScanOut869[5] , 
        \nOut19_19[4] , \nOut26_22[0] , \nScanOut1019[3] , \nScanOut1[0] , 
        \nScanOut11[4] , \nOut2_15[6] , \nOut16_20[4] , \nOut25_14[5] , 
        \nOut2_16[5] , \nOut7_29[1] , \nScanOut689[3] , \nScanOut939[2] , 
        \nScanOut110[7] , \nOut5_25[3] , \nScanOut270[2] , \nScanOut338[7] , 
        \nScanOut658[6] , \nOut16_23[7] , \nScanOut538[3] , \nOut20_28[2] , 
        \nOut25_17[6] , \nOut29_18[3] , \nScanOut344[1] , \nScanOut624[0] , 
        \nScanOut710[3] , \nScanOut997[2] , \nScanOut396[7] , \nScanOut470[6] , 
        \nScanOut544[5] , \nOut31_23[3] , \nScanOut871[7] , \nScanOut945[4] , 
        \nScanOut12[7] , \nOut11_10[1] , \nOut18_20[0] , \nOut22_24[0] , 
        \nOut10_31[7] , \nScanOut596[3] , \nScanOut872[4] , \nScanOut1001[1] , 
        \nOut0_19[4] , \nOut1_9[3] , \nOut12_9[6] , \nScanOut946[7] , 
        \nOut7_9[7] , \nScanOut395[4] , \nOut27_18[7] , \nOut31_20[0] , 
        \nOut11_13[2] , \nOut14_9[2] , \nScanOut595[0] , \nScanOut1002[2] , 
        \nOut18_23[3] , \nOut22_27[3] , \nScanOut30[6] , \nScanOut75[0] , 
        \nScanOut113[4] , \nOut5_26[0] , \nScanOut273[1] , \nScanOut627[3] , 
        \nScanOut713[0] , \nScanOut994[1] , \nOut9_29[5] , \nScanOut347[2] , 
        \nOut18_8[3] , \nScanOut473[5] , \nScanOut547[6] , \nScanOut692[2] , 
        \nScanOut815[3] , \nScanOut76[3] , \nOut6_10[5] , \nScanOut921[0] , 
        \nOut6_13[6] , \nScanOut174[3] , \nScanOut214[6] , \nOut7_31[3] , 
        \nScanOut640[4] , \nScanOut774[7] , \nScanOut320[5] , \nScanOut414[2] , 
        \nScanOut520[1] , \nOut20_30[0] , \nOut21_11[6] , \nOut28_21[7] , 
        \nScanOut177[0] , \nScanOut217[5] , \nOut12_25[7] , \nScanOut323[6] , 
        \nOut23_8[3] , \nOut12_26[4] , \nScanOut643[7] , \nScanOut777[4] , 
        \nOut28_22[4] , \nScanOut417[1] , \nScanOut523[2] , \nOut17_19[0] , 
        \nOut25_8[7] , \nOut21_12[5] , \nScanOut691[1] , \nScanOut816[0] , 
        \nOut29_9[6] , \nScanOut922[3] , \nScanOut850[5] , \nScanOut964[6] , 
        \nScanOut33[5] , \nOut1_19[0] , \nOut4_25[7] , \nScanOut251[0] , 
        \nScanOut283[6] , \nOut10_10[5] , \nOut30_23[7] , \nOut11_31[3] , 
        \nScanOut483[2] , \nOut19_20[4] , \nScanOut1020[3] , \nScanOut605[2] , 
        \nOut23_24[4] , \nScanOut731[1] , \nScanOut882[3] , \nScanOut365[3] , 
        \nOut4_26[4] , \nScanOut131[5] , \nScanOut451[4] , \nScanOut565[7] , 
        \nScanOut252[3] , \nOut8_29[1] , \nScanOut366[0] , \nScanOut132[6] , 
        \nScanOut606[1] , \nScanOut881[0] , \nScanOut732[2] , \nScanOut280[5] , 
        \nScanOut452[7] , \nScanOut566[4] , \nScanOut853[6] , \nOut30_20[4] , 
        \nScanOut86[4] , \nScanOut235[4] , \nOut10_13[6] , \nOut19_23[7] , 
        \nOut23_27[7] , \nScanOut967[5] , \nScanOut480[1] , \nOut26_18[3] , 
        \nScanOut1023[0] , \nScanOut301[7] , \nScanOut661[6] , 
        \nScanOut755[5] , \nOut29_21[3] , \nScanOut2[3] , \nScanOut54[2] , 
        \nScanOut155[1] , \nOut13_25[3] , \nScanOut435[0] , \nScanOut501[3] , 
        \nOut21_30[4] , \nOut20_11[2] , \nScanOut787[3] , \nScanOut834[1] , 
        \nScanOut57[1] , \nScanOut187[7] , \nOut7_10[1] , \nOut6_31[7] , 
        \nScanOut900[2] , \nOut7_13[2] , \nScanOut837[2] , \nScanOut784[0] , 
        \nScanOut903[1] , \nScanOut85[7] , \nScanOut184[4] , \nScanOut662[5] , 
        \nScanOut756[6] , \nScanOut236[7] , \nScanOut302[4] , \nOut13_26[0] , 
        \nScanOut436[3] , \nScanOut502[0] , \nOut16_19[4] , \nOut20_12[1] , 
        \nOut0_4[0] , \nOut0_20[4] , \nScanOut156[2] , \nOut29_22[0] , 
        \nOut9_10[5] , \nOut8_31[3] , \nOut19_5[0] , \nOut21_1[1] , 
        \nOut27_1[5] , \nScanOut899[2] , \nOut0_7[3] , \nScanOut28[4] , 
        \nOut6_4[4] , \nScanOut298[7] , \nOut13_4[5] , \nOut31_19[0] , 
        \nOut14_15[6] , \nOut15_4[1] , \nOut27_21[7] , \nOut13_7[6] , 
        \nScanOut498[3] , \nScanOut848[7] , \nOut0_23[7] , \nOut6_7[7] , 
        \nOut11_29[1] , \nOut27_22[4] , \nOut14_16[5] , \nOut15_7[2] , 
        \nOut18_19[0] , \nOut27_2[6] , \nOut2_8[6] , \nOut2_10[2] , 
        \nOut2_13[1] , \nOut3_3[2] , \nOut3_15[2] , \nScanOut129[7] , 
        \nScanOut249[2] , \nOut19_6[3] , \nScanOut729[3] , \nOut9_13[6] , 
        \nScanOut449[6] , \nOut5_0[5] , \nOut21_2[2] , \nOut28_4[5] , 
        \nOut3_16[1] , \nOut3_0[1] , \nOut10_0[4] , \nOut16_0[0] , 
        \nOut9_1[4] , \nOut22_5[0] , \nOut9_2[7] , \nScanOut319[5] , 
        \nOut17_20[0] , \nOut24_5[4] , \nOut24_14[1] , \nOut22_6[3] , 
        \nScanOut679[4] , \nOut24_17[2] , \nOut28_18[7] , \nScanOut519[1] , 
        \nOut24_6[7] , \nOut17_23[3] , \nOut21_28[6] , \nOut5_3[6] , 
        \nOut6_29[5] , \nOut16_3[3] , \nScanOut918[0] , \nOut28_7[6] , 
        \nScanOut68[6] , \nScanOut169[5] , \nOut10_3[7] , \nScanOut409[4] , 
        \nOut16_26[3] , \nScanOut209[0] , \nOut13_19[7] , \nOut25_12[2] , 
        \nScanOut769[1] , \nScanOut808[5] , \nOut3_31[4] , \nOut1_25[4] , 
        \nOut1_26[7] , \nOut4_19[3] , \nOut15_13[5] , \nOut16_25[0] , 
        \nOut24_30[7] , \nOut25_11[1] , \nScanOut559[3] , \nOut23_18[0] , 
        \nOut26_27[4] , \nScanOut958[2] , \nOut31_7[2] , \nOut8_16[6] , 
        \nScanOut359[7] , \nScanOut639[6] , \nOut31_4[1] , \nOut8_15[5] , 
        \nScanOut989[7] , \nScanOut388[2] , \nOut15_10[6] , \nOut14_31[0] , 
        \nScanOut588[6] , \nOut26_24[7] , \nScanOut73[7] , \nOut3_29[6] , 
        \nOut11_8[3] , \nOut4_8[2] , \nOut17_8[7] , \nScanOut694[5] , 
        \nScanOut813[4] , \nScanOut14[0] , \nScanOut17[3] , \nScanOut70[4] , 
        \nScanOut171[7] , \nScanOut172[4] , \nOut6_16[2] , \nScanOut927[7] , 
        \nOut28_27[0] , \nScanOut212[1] , \nOut8_9[3] , \nOut12_23[0] , 
        \nScanOut412[5] , \nScanOut526[6] , \nOut24_28[5] , \nOut21_17[1] , 
        \nScanOut326[2] , \nOut12_20[3] , \nScanOut411[6] , \nScanOut525[5] , 
        \nScanOut646[3] , \nScanOut772[0] , \nOut21_14[2] , \nOut28_24[3] , 
        \nOut6_15[1] , \nScanOut211[2] , \nScanOut645[0] , \nScanOut771[3] , 
        \nScanOut325[1] , \nScanOut697[6] , \nScanOut810[7] , \nScanOut924[4] , 
        \nScanOut116[0] , \nScanOut476[1] , \nScanOut542[2] , \nOut20_9[6] , 
        \nOut5_23[4] , \nScanOut276[5] , \nScanOut622[7] , \nScanOut716[4] , 
        \nOut26_9[2] , \nScanOut991[5] , \nScanOut342[6] , \nOut11_16[6] , 
        \nOut14_29[2] , \nOut18_26[7] , \nScanOut590[4] , \nScanOut1007[6] , 
        \nOut22_22[7] , \nScanOut877[0] , \nScanOut943[3] , \nOut11_15[5] , 
        \nScanOut390[0] , \nOut31_25[4] , \nOut18_25[4] , \nOut22_21[4] , 
        \nScanOut393[3] , \nScanOut593[7] , \nScanOut1004[5] , 
        \nScanOut874[3] , \nOut31_26[7] , \nOut1_28[1] , \nScanOut103[7] , 
        \nScanOut115[3] , \nScanOut940[0] , \nOut5_20[7] , \nScanOut275[6] , 
        \nScanOut475[2] , \nScanOut541[1] , \nScanOut341[5] , \nScanOut621[4] , 
        \nScanOut715[7] , \nScanOut992[6] , \nOut4_17[5] , \nOut8_18[0] , 
        \nScanOut263[2] , \nScanOut463[6] , \nScanOut557[5] , \nOut31_9[4] , 
        \nScanOut357[1] , \nOut0_9[5] , \nOut0_11[5] , \nOut0_12[6] , 
        \nScanOut19[5] , \nScanOut65[3] , \nScanOut66[0] , \nScanOut100[4] , 
        \nOut10_21[4] , \nOut10_22[7] , \nScanOut585[3] , \nOut19_12[6] , 
        \nScanOut637[0] , \nScanOut703[3] , \nScanOut984[2] , \nOut23_16[6] , 
        \nOut26_29[2] , \nScanOut385[7] , \nScanOut1012[1] , \nScanOut862[7] , 
        \nOut30_11[5] , \nOut31_30[3] , \nScanOut956[4] , \nScanOut386[4] , 
        \nOut18_30[3] , \nScanOut586[0] , \nOut19_11[5] , \nScanOut1011[2] , 
        \nOut23_15[5] , \nScanOut861[4] , \nOut30_12[6] , \nScanOut955[7] , 
        \nScanOut460[5] , \nScanOut554[6] , \nOut4_14[6] , \nScanOut260[1] , 
        \nScanOut634[3] , \nScanOut700[0] , \nScanOut987[1] , \nOut7_22[3] , 
        \nScanOut354[2] , \nScanOut681[2] , \nScanOut806[3] , \nScanOut932[0] , 
        \nScanOut164[0] , \nScanOut167[3] , \nOut13_17[1] , \nScanOut407[2] , 
        \nOut16_28[5] , \nScanOut533[1] , \nOut20_23[0] , \nOut29_13[1] , 
        \nScanOut207[6] , \nScanOut653[4] , \nScanOut767[7] , \nScanOut333[5] , 
        \nOut29_10[2] , \nOut28_31[4] , \nScanOut204[5] , \nOut13_14[2] , 
        \nScanOut404[1] , \nScanOut530[2] , \nOut20_20[3] , \nScanOut330[6] , 
        \nScanOut650[7] , \nScanOut682[1] , \nScanOut764[4] , \nScanOut805[0] , 
        \nOut7_2[5] , \nOut7_21[0] , \nScanOut931[3] , \nOut11_18[0] , 
        \nOut12_2[4] , \nOut14_2[0] , \nOut27_13[5] , \nScanOut1009[0] , 
        \nOut14_27[4] , \nOut18_28[1] , \nScanOut879[6] , \nOut1_2[1] , 
        \nScanOut118[6] , \nScanOut478[7] , \nOut20_7[0] , \nOut1_30[3] , 
        \nOut9_21[4] , \nScanOut278[3] , \nScanOut718[2] , \nOut26_7[4] , 
        \nOut9_22[7] , \nOut18_3[1] , \nOut20_4[3] , \nOut18_0[2] , 
        \nScanOut25[1] , \nEnable[0] , \nOut1_1[2] , \nOut7_1[6] , 
        \nOut14_1[3] , \nOut26_4[7] , \nOut14_24[7] , \nOut27_10[6] , 
        \nOut26_31[0] , \nOut31_28[1] , \nOut2_5[3] , \nOut2_6[0] , 
        \nOut8_7[5] , \nOut12_1[7] , \nScanOut528[0] , \nOut24_26[3] , 
        \nOut28_29[6] , \nScanOut328[4] , \nOut17_12[2] , \nOut21_19[7] , 
        \nOut25_3[5] , \nOut23_3[1] , \nScanOut648[5] , \nOut3_27[0] , 
        \nOut11_6[5] , \nOut4_6[4] , \nOut17_6[1] , \nOut29_2[4] , 
        \nOut6_18[4] , \nScanOut929[1] , \nOut11_5[6] , \nOut2_21[3] , 
        \nOut3_24[3] , \nOut4_5[7] , \nScanOut699[0] , \nOut29_1[7] , 
        \nOut17_5[2] , \nOut8_4[6] , \nOut16_30[7] , \nOut17_11[1] , 
        \nOut23_0[2] , \nOut24_25[0] , \nOut25_0[6] , \nScanOut41[5] , 
        \nOut1_14[5] , \nOut2_22[0] , \nScanOut59[7] , \nScanOut88[2] , 
        \nScanOut189[1] , \nScanOut789[5] , \nScanOut158[4] , \nScanOut238[1] , 
        \nOut16_14[1] , \nOut25_20[0] , \nScanOut758[0] , \nScanOut438[5] , 
        \nOut16_17[2] , \nOut13_28[6] , \nOut25_23[3] , \nScanOut839[4] , 
        \nOut1_17[6] , \nOut4_28[2] , \nOut8_24[4] , \nScanOut368[6] , 
        \nOut15_21[7] , \nOut26_15[6] , \nOut30_1[3] , \nOut15_22[4] , 
        \nOut23_29[1] , \nScanOut969[3] , \nOut26_16[5] , \nOut8_27[7] , 
        \nScanOut608[7] , \nScanOut93[3] , \nScanOut568[2] , \nOut30_2[0] , 
        \nScanOut674[1] , \nScanOut740[2] , \nScanOut140[6] , \nScanOut220[3] , 
        \nScanOut314[0] , \nOut12_11[2] , \nScanOut420[7] , \nScanOut514[4] , 
        \nOut21_25[3] , \nOut13_30[4] , \nOut6_24[0] , \nScanOut821[6] , 
        \nOut28_15[2] , \nScanOut915[5] , \nScanOut792[4] , \nScanOut42[6] , 
        \nOut3_18[7] , \nScanOut192[0] , \nScanOut791[7] , \nScanOut822[5] , 
        \nOut28_9[0] , \nScanOut90[0] , \nOut6_27[3] , \nScanOut916[6] , 
        \nScanOut191[3] , \nScanOut223[0] , \nScanOut317[3] , \nOut22_8[5] , 
        \nScanOut677[2] , \nScanOut743[1] , \nScanOut143[5] , \nScanOut296[1] , 
        \nOut12_12[1] , \nOut24_19[4] , \nOut28_16[1] , \nScanOut423[4] , 
        \nScanOut517[7] , \nOut21_26[0] , \nOut24_8[1] , \nScanOut845[2] , 
        \nOut31_17[6] , \nScanOut26[2] , \nScanOut124[2] , \nOut4_30[0] , 
        \nOut5_11[6] , \nScanOut244[7] , \nOut11_24[4] , \nOut18_14[5] , 
        \nOut22_10[5] , \nOut23_31[3] , \nScanOut971[1] , \nScanOut496[5] , 
        \nScanOut370[4] , \nScanOut610[5] , \nScanOut897[4] , \nScanOut724[6] , 
        \nScanOut127[1] , \nOut5_12[5] , \nScanOut247[4] , \nScanOut444[3] , 
        \nScanOut570[0] , \nScanOut613[6] , \nScanOut727[5] , \nScanOut894[7] , 
        \nScanOut373[7] , \nOut19_8[5] , \nScanOut447[0] , \nScanOut573[3] , 
        \nOut13_9[0] , \nScanOut846[1] , \nScanOut972[2] , \nScanOut11[0] , 
        \nScanOut12[3] , \nOut0_19[0] , \nScanOut113[0] , \nOut6_9[1] , 
        \nScanOut295[2] , \nOut11_27[7] , \nOut31_14[5] , \nOut14_18[3] , 
        \nOut15_9[4] , \nScanOut495[6] , \nOut18_17[6] , \nOut22_13[6] , 
        \nOut5_26[4] , \nScanOut273[5] , \nScanOut473[1] , \nScanOut547[2] , 
        \nOut9_29[1] , \nScanOut347[6] , \nOut18_8[7] , \nOut1_9[7] , 
        \nOut7_9[3] , \nOut14_9[6] , \nScanOut627[7] , \nScanOut713[4] , 
        \nScanOut994[5] , \nOut18_23[7] , \nOut22_27[7] , \nOut11_13[6] , 
        \nScanOut595[4] , \nOut27_18[3] , \nScanOut1002[6] , \nOut12_9[2] , 
        \nScanOut395[0] , \nScanOut872[0] , \nOut31_20[4] , \nOut11_10[5] , 
        \nScanOut946[3] , \nOut10_31[3] , \nScanOut596[7] , \nOut18_20[4] , 
        \nScanOut1001[5] , \nOut22_24[4] , \nScanOut871[3] , \nScanOut945[0] , 
        \nOut1_23[7] , \nScanOut75[4] , \nScanOut76[7] , \nScanOut110[3] , 
        \nScanOut396[3] , \nOut31_23[7] , \nScanOut470[2] , \nScanOut544[1] , 
        \nOut5_25[7] , \nScanOut270[6] , \nScanOut624[4] , \nScanOut710[7] , 
        \nScanOut997[6] , \nScanOut344[5] , \nOut6_13[2] , \nScanOut691[5] , 
        \nScanOut816[4] , \nOut29_9[2] , \nScanOut922[7] , \nScanOut174[7] , 
        \nScanOut177[4] , \nOut12_26[0] , \nScanOut417[5] , \nScanOut523[6] , 
        \nOut21_12[1] , \nOut25_8[3] , \nOut17_19[4] , \nOut28_22[0] , 
        \nScanOut217[1] , \nScanOut643[3] , \nScanOut777[0] , \nScanOut323[2] , 
        \nOut23_8[7] , \nOut28_21[3] , \nScanOut214[2] , \nOut12_25[3] , 
        \nScanOut414[6] , \nScanOut520[5] , \nOut20_30[4] , \nOut21_11[2] , 
        \nScanOut320[1] , \nScanOut640[0] , \nScanOut692[6] , \nScanOut774[3] , 
        \nScanOut815[7] , \nScanOut108[1] , \nOut6_10[1] , \nScanOut921[4] , 
        \nOut7_31[7] , \nOut10_29[1] , \nOut26_22[4] , \nOut15_16[5] , 
        \nScanOut1019[7] , \nScanOut468[0] , \nOut19_19[0] , \nScanOut869[1] , 
        \nOut31_2[2] , \nOut8_13[6] , \nScanOut268[4] , \nScanOut708[5] , 
        \nOut2_15[2] , \nOut2_16[1] , \nOut1_20[4] , \nOut8_10[5] , 
        \nOut9_31[3] , \nOut31_1[1] , \nScanOut338[3] , \nOut15_15[6] , 
        \nOut16_23[3] , \nScanOut538[7] , \nOut25_17[2] , \nOut26_21[7] , 
        \nOut30_19[0] , \nOut29_18[7] , \nOut20_28[6] , \nScanOut658[2] , 
        \nOut7_29[5] , \nScanOut939[6] , \nScanOut689[7] , \nOut16_20[0] , 
        \nOut25_14[1] , \nOut0_1[0] , \nOut0_25[4] , \nScanOut49[0] , 
        \nOut3_5[1] , \nOut3_10[2] , \nOut2_31[4] , \nOut5_5[5] , 
        \nOut16_5[0] , \nScanOut799[2] , \nOut28_1[5] , \nScanOut199[6] , 
        \nScanOut98[5] , \nOut10_5[4] , \nOut22_0[0] , \nScanOut148[3] , 
        \nScanOut228[6] , \nOut9_4[4] , \nOut24_11[1] , \nOut25_30[7] , 
        \nOut17_25[0] , \nOut24_0[4] , \nScanOut748[7] , \nOut9_7[7] , 
        \nOut22_3[3] , \nScanOut428[2] , \nOut17_26[3] , \nOut24_3[7] , 
        \nOut12_19[7] , \nOut24_12[2] , \nScanOut829[3] , \nOut28_2[6] , 
        \nOut3_6[2] , \nOut3_13[1] , \nOut5_6[6] , \nOut10_6[7] , 
        \nOut16_6[3] , \nOut9_15[5] , \nOut19_0[0] , \nOut27_4[5] , 
        \nOut13_1[5] , \nOut21_4[1] , \nOut0_2[3] , \nOut6_1[4] , 
        \nOut27_24[7] , \nOut14_10[6] , \nOut15_31[0] , \nOut15_1[1] , 
        \nScanOut4[0] , \nOut0_26[7] , \nOut5_19[3] , \nOut6_2[7] , 
        \nOut13_2[6] , \nOut14_13[5] , \nOut15_2[2] , \nScanOut979[4] , 
        \nOut22_18[0] , \nOut27_27[4] , \nScanOut378[1] , \nOut19_3[3] , 
        \nOut9_16[6] , \nScanOut618[0] , \nOut27_7[6] , \nScanOut83[4] , 
        \nScanOut578[5] , \nOut21_7[2] , \nScanOut664[6] , \nScanOut750[5] , 
        \nScanOut230[4] , \nScanOut304[7] , \nOut13_20[3] , \nScanOut430[0] , 
        \nScanOut504[3] , \nOut20_14[2] , \nOut29_24[3] , \nScanOut7[3] , 
        \nScanOut51[2] , \nScanOut150[1] , \nOut7_15[1] , \nScanOut831[1] , 
        \nScanOut782[3] , \nScanOut905[2] , \nScanOut52[1] , \nOut2_29[6] , 
        \nScanOut182[7] , \nScanOut781[0] , \nScanOut832[2] , \nScanOut80[7] , 
        \nScanOut181[4] , \nOut7_16[2] , \nScanOut906[1] , \nScanOut233[7] , 
        \nScanOut307[4] , \nScanOut667[5] , \nScanOut753[6] , \nScanOut9[5] , 
        \nScanOut20[1] , \nScanOut35[6] , \nScanOut153[2] , \nOut29_27[0] , 
        \nScanOut286[6] , \nOut13_23[0] , \nScanOut433[3] , \nScanOut507[0] , 
        \nOut25_28[5] , \nOut20_17[1] , \nScanOut855[5] , \nOut30_26[7] , 
        \nScanOut36[5] , \nOut4_20[7] , \nScanOut254[0] , \nOut10_15[5] , 
        \nOut19_25[4] , \nOut23_21[4] , \nScanOut961[6] , \nScanOut486[2] , 
        \nScanOut360[3] , \nOut4_23[4] , \nScanOut134[5] , \nScanOut600[2] , 
        \nScanOut887[3] , \nScanOut734[1] , \nScanOut257[3] , \nScanOut454[4] , 
        \nScanOut560[7] , \nScanOut603[1] , \nScanOut737[2] , \nScanOut884[0] , 
        \nScanOut363[0] , \nScanOut137[6] , \nScanOut457[7] , \nScanOut563[4] , 
        \nOut30_9[6] , \nScanOut856[6] , \nScanOut962[5] , \nScanOut285[5] , 
        \nOut10_16[6] , \nOut30_25[4] , \nOut15_29[2] , \nScanOut485[1] , 
        \nOut19_26[7] , \nOut23_22[7] , \nScanOut840[2] , \nScanOut974[1] , 
        \nScanOut23[2] , \nOut0_28[1] , \nScanOut121[2] , \nOut5_14[6] , 
        \nScanOut241[7] , \nScanOut293[1] , \nOut11_21[4] , \nOut31_12[6] , 
        \nScanOut493[5] , \nOut18_11[5] , \nOut19_30[3] , \nScanOut615[5] , 
        \nOut22_15[5] , \nScanOut721[6] , \nScanOut892[4] , \nScanOut375[4] , 
        \nScanOut441[3] , \nScanOut575[0] , \nOut5_17[5] , \nScanOut242[4] , 
        \nOut9_18[0] , \nScanOut376[7] , \nOut27_9[0] , \nScanOut122[1] , 
        \nScanOut616[6] , \nScanOut891[7] , \nScanOut722[5] , \nScanOut290[2] , 
        \nScanOut442[0] , \nScanOut576[3] , \nOut21_9[4] , \nScanOut843[1] , 
        \nOut30_30[3] , \nOut31_11[5] , \nOut0_30[3] , \nScanOut44[5] , 
        \nScanOut96[3] , \nScanOut225[3] , \nOut11_22[7] , \nOut18_12[6] , 
        \nOut22_16[6] , \nScanOut977[2] , \nOut27_29[2] , \nScanOut490[6] , 
        \nScanOut311[0] , \nScanOut671[1] , \nScanOut745[2] , \nScanOut145[6] , 
        \nOut29_31[4] , \nOut12_14[2] , \nOut28_10[2] , \nScanOut425[7] , 
        \nScanOut511[4] , \nOut21_20[3] , \nScanOut797[4] , \nScanOut824[6] , 
        \nScanOut47[6] , \nOut6_21[0] , \nScanOut910[5] , \nOut6_22[3] , 
        \nScanOut197[0] , \nScanOut827[5] , \nScanOut913[6] , \nScanOut794[7] , 
        \nOut3_8[4] , \nOut5_8[0] , \nScanOut194[3] , \nOut10_8[1] , 
        \nOut16_8[5] , \nScanOut95[0] , \nScanOut672[2] , \nScanOut746[1] , 
        \nScanOut146[5] , \nScanOut226[0] , \nOut9_9[1] , \nScanOut312[3] , 
        \nOut12_17[1] , \nScanOut426[4] , \nScanOut512[7] , \nOut17_28[5] , 
        \nOut21_23[0] , \nOut8_21[4] , \nOut28_13[1] , \nScanOut38[3] , 
        \nOut1_11[5] , \nScanOut288[0] , \nScanOut889[5] , \nOut30_4[3] , 
        \nOut15_24[7] , \nOut30_28[1] , \nScanOut488[4] , \nOut26_10[6] , 
        \nOut27_31[0] , \nScanOut858[0] , \nOut1_12[6] , \nOut10_18[0] , 
        \nOut15_27[4] , \nOut26_13[5] , \nOut19_28[1] , \nOut2_24[3] , 
        \nScanOut139[0] , \nOut8_22[7] , \nScanOut259[5] , \nScanOut739[4] , 
        \nScanOut459[1] , \nOut30_7[0] , \nScanOut309[2] , \nOut16_11[1] , 
        \nOut17_30[7] , \nOut25_25[0] , \nScanOut669[3] , \nOut25_26[3] , 
        \nOut0_14[5] , \nOut0_17[6] , \nOut2_3[0] , \nOut2_27[0] , 
        \nOut16_12[2] , \nScanOut509[6] , \nOut29_29[6] , \nOut20_19[7] , 
        \nScanOut179[2] , \nOut7_18[4] , \nOut8_2[5] , \nScanOut419[3] , 
        \nScanOut908[7] , \nOut17_17[2] , \nOut25_6[5] , \nScanOut219[7] , 
        \nOut12_28[6] , \nOut23_6[1] , \nOut24_23[3] , \nScanOut779[6] , 
        \nOut11_3[5] , \nOut1_7[1] , \nOut2_0[3] , \nScanOut78[1] , 
        \nOut4_3[4] , \nOut29_7[4] , \nScanOut818[2] , \nOut3_22[0] , 
        \nOut17_3[1] , \nOut3_21[3] , \nOut11_0[6] , \nOut17_0[2] , 
        \nOut4_0[7] , \nOut29_4[7] , \nOut7_7[5] , \nOut8_1[6] , 
        \nOut24_20[0] , \nOut14_7[0] , \nOut17_14[1] , \nOut25_5[6] , 
        \nOut23_5[2] , \nOut14_22[4] , \nOut22_29[1] , \nOut27_16[5] , 
        \nOut5_28[2] , \nScanOut349[0] , \nOut12_7[4] , \nScanOut948[5] , 
        \nScanOut549[4] , \nOut20_2[0] , \nOut9_27[7] , \nOut18_6[1] , 
        \nScanOut629[1] , \nOut20_1[3] , \nOut26_2[4] , \nOut7_4[6] , 
        \nOut9_24[4] , \nOut26_1[7] , \nScanOut999[0] , \nOut18_5[2] , 
        \nOut27_15[6] , \nOut14_4[3] , \nScanOut598[1] , \nOut14_21[7] , 
        \nScanOut1[4] , \nScanOut2[7] , \nOut0_4[4] , \nOut0_7[7] , 
        \nOut0_9[1] , \nOut1_4[2] , \nOut12_4[7] , \nScanOut41[1] , 
        \nScanOut42[2] , \nOut2_18[7] , \nScanOut398[5] , \nScanOut60[3] , 
        \nScanOut63[0] , \nScanOut684[2] , \nScanOut803[3] , \nScanOut161[0] , 
        \nScanOut162[3] , \nOut7_27[3] , \nScanOut937[0] , \nOut29_16[1] , 
        \nScanOut202[6] , \nOut13_12[1] , \nOut25_19[4] , \nScanOut402[2] , 
        \nScanOut536[1] , \nOut20_26[0] , \nScanOut336[5] , \nOut12_30[4] , 
        \nOut13_11[2] , \nScanOut401[1] , \nScanOut535[2] , \nScanOut656[4] , 
        \nScanOut762[7] , \nOut20_25[3] , \nOut29_15[2] , \nScanOut201[5] , 
        \nScanOut655[7] , \nScanOut761[4] , \nOut7_24[0] , \nScanOut335[6] , 
        \nScanOut687[1] , \nScanOut800[0] , \nScanOut934[3] , \nScanOut90[4] , 
        \nScanOut105[4] , \nScanOut106[7] , \nScanOut466[6] , \nScanOut552[5] , 
        \nOut4_12[5] , \nScanOut266[2] , \nScanOut632[0] , \nScanOut706[3] , 
        \nScanOut981[2] , \nOut10_24[4] , \nOut10_27[7] , \nScanOut352[1] , 
        \nScanOut580[3] , \nScanOut380[7] , \nOut15_18[3] , \nOut19_17[6] , 
        \nScanOut1017[1] , \nOut23_13[6] , \nScanOut867[7] , \nOut30_14[5] , 
        \nScanOut953[4] , \nOut19_14[5] , \nOut23_10[5] , \nOut22_31[3] , 
        \nScanOut383[4] , \nScanOut583[0] , \nScanOut1014[2] , 
        \nScanOut864[4] , \nOut30_17[6] , \nScanOut950[7] , \nOut4_11[6] , 
        \nScanOut265[1] , \nScanOut465[5] , \nScanOut551[6] , \nScanOut143[1] , 
        \nOut5_30[0] , \nScanOut351[2] , \nScanOut423[0] , \nScanOut517[3] , 
        \nScanOut631[3] , \nScanOut705[0] , \nScanOut982[1] , \nOut21_26[4] , 
        \nOut24_8[5] , \nOut12_12[5] , \nOut28_16[5] , \nScanOut677[6] , 
        \nOut24_19[0] , \nScanOut743[5] , \nScanOut191[7] , \nScanOut223[4] , 
        \nScanOut317[7] , \nOut22_8[1] , \nScanOut791[3] , \nScanOut822[1] , 
        \nOut3_18[3] , \nOut6_27[7] , \nOut28_9[4] , \nScanOut916[2] , 
        \nOut6_24[4] , \nScanOut192[4] , \nScanOut821[2] , \nScanOut915[1] , 
        \nScanOut792[0] , \nScanOut93[7] , \nScanOut140[2] , \nOut12_11[6] , 
        \nOut13_30[0] , \nScanOut220[7] , \nScanOut420[3] , \nScanOut514[0] , 
        \nOut28_15[6] , \nOut21_25[7] , \nScanOut314[4] , \nScanOut674[5] , 
        \nScanOut740[6] , \nOut6_9[5] , \nOut11_27[3] , \nOut14_18[7] , 
        \nOut15_9[0] , \nOut18_17[2] , \nOut22_13[2] , \nScanOut495[2] , 
        \nOut0_11[1] , \nScanOut25[5] , \nScanOut26[6] , \nScanOut295[6] , 
        \nOut13_9[4] , \nScanOut846[5] , \nOut31_14[1] , \nScanOut972[6] , 
        \nScanOut124[6] , \nScanOut127[5] , \nOut5_12[1] , \nScanOut247[0] , 
        \nScanOut447[4] , \nScanOut573[7] , \nScanOut373[3] , \nOut19_8[1] , 
        \nScanOut444[7] , \nScanOut570[4] , \nScanOut613[2] , \nScanOut727[1] , 
        \nScanOut894[3] , \nOut4_30[4] , \nOut5_11[2] , \nScanOut244[3] , 
        \nScanOut610[1] , \nScanOut897[0] , \nScanOut724[2] , \nScanOut370[0] , 
        \nOut11_24[0] , \nScanOut496[1] , \nOut18_14[1] , \nOut22_10[1] , 
        \nOut23_31[7] , \nScanOut845[6] , \nOut1_1[6] , \nOut1_14[1] , 
        \nOut1_17[2] , \nOut2_21[7] , \nOut2_22[4] , \nScanOut296[5] , 
        \nScanOut971[5] , \nOut31_17[2] , \nScanOut59[3] , \nScanOut839[0] , 
        \nScanOut88[6] , \nScanOut158[0] , \nScanOut238[5] , \nOut13_28[2] , 
        \nOut25_23[7] , \nScanOut438[1] , \nOut16_17[6] , \nOut16_14[5] , 
        \nScanOut758[4] , \nOut25_20[4] , \nScanOut189[5] , \nScanOut789[1] , 
        \nScanOut568[6] , \nScanOut608[3] , \nOut30_2[4] , \nOut4_28[6] , 
        \nScanOut368[2] , \nOut8_24[0] , \nOut8_27[3] , \nOut15_21[3] , 
        \nOut15_22[0] , \nOut26_16[1] , \nOut23_29[5] , \nScanOut969[7] , 
        \nOut26_15[2] , \nOut30_1[7] , \nOut12_1[3] , \nOut31_28[5] , 
        \nOut1_30[7] , \nOut7_1[2] , \nOut14_1[7] , \nOut27_10[2] , 
        \nOut26_31[4] , \nOut14_24[3] , \nOut0_12[2] , \nOut9_21[0] , 
        \nOut26_4[3] , \nScanOut278[7] , \nOut18_0[6] , \nOut20_4[7] , 
        \nOut9_22[3] , \nOut18_3[5] , \nScanOut14[4] , \nScanOut19[1] , 
        \nOut1_2[5] , \nScanOut118[2] , \nScanOut718[6] , \nOut26_7[0] , 
        \nScanOut478[3] , \nOut20_7[4] , \nScanOut879[2] , \nOut2_5[7] , 
        \nOut3_24[7] , \nOut7_2[1] , \nOut12_2[0] , \nOut14_2[4] , 
        \nOut14_27[0] , \nOut18_28[5] , \nOut27_13[1] , \nOut8_4[2] , 
        \nOut11_18[4] , \nOut16_30[3] , \nOut23_0[6] , \nScanOut1009[4] , 
        \nOut24_25[4] , \nOut17_11[5] , \nOut25_0[2] , \nOut4_5[3] , 
        \nOut17_5[6] , \nScanOut699[4] , \nOut29_1[3] , \nOut2_6[4] , 
        \nOut3_27[4] , \nOut4_6[0] , \nOut11_5[2] , \nOut29_2[0] , 
        \nOut6_18[0] , \nScanOut929[5] , \nOut17_6[5] , \nOut11_6[1] , 
        \nOut2_8[2] , \nOut1_28[5] , \nScanOut100[0] , \nOut4_14[2] , 
        \nOut8_7[1] , \nScanOut328[0] , \nScanOut648[1] , \nOut23_3[5] , 
        \nScanOut528[4] , \nScanOut260[5] , \nOut17_12[6] , \nOut25_3[1] , 
        \nOut21_19[3] , \nOut24_26[7] , \nOut28_29[2] , \nScanOut354[6] , 
        \nScanOut634[7] , \nScanOut700[4] , \nScanOut987[5] , \nOut10_21[0] , 
        \nScanOut386[0] , \nScanOut460[1] , \nScanOut554[2] , \nOut30_12[2] , 
        \nOut18_30[7] , \nOut19_11[1] , \nScanOut861[0] , \nScanOut955[3] , 
        \nScanOut586[4] , \nOut23_15[1] , \nOut10_22[3] , \nScanOut385[3] , 
        \nScanOut862[3] , \nScanOut1011[6] , \nScanOut956[0] , \nOut30_11[1] , 
        \nOut31_30[7] , \nScanOut585[7] , \nOut19_12[2] , \nOut23_16[2] , 
        \nOut26_29[6] , \nScanOut1012[5] , \nScanOut65[7] , \nScanOut103[3] , 
        \nOut4_17[1] , \nOut8_18[4] , \nScanOut263[6] , \nScanOut637[4] , 
        \nScanOut703[7] , \nScanOut984[6] , \nScanOut357[5] , \nScanOut463[2] , 
        \nScanOut557[1] , \nScanOut682[5] , \nOut31_9[0] , \nScanOut805[4] , 
        \nScanOut66[4] , \nScanOut164[4] , \nScanOut204[1] , \nOut7_21[4] , 
        \nScanOut931[7] , \nScanOut650[3] , \nScanOut764[0] , \nScanOut330[2] , 
        \nScanOut404[5] , \nScanOut530[6] , \nOut20_20[7] , \nOut29_10[6] , 
        \nOut28_31[0] , \nScanOut167[7] , \nScanOut207[2] , \nOut13_14[6] , 
        \nScanOut333[1] , \nOut13_17[5] , \nScanOut653[0] , \nScanOut767[3] , 
        \nOut29_13[5] , \nOut7_22[7] , \nScanOut407[6] , \nOut16_28[1] , 
        \nScanOut533[5] , \nOut20_23[4] , \nScanOut681[6] , \nScanOut806[7] , 
        \nScanOut932[4] , \nScanOut70[0] , \nOut6_15[5] , \nScanOut697[2] , 
        \nScanOut810[3] , \nScanOut924[0] , \nScanOut73[3] , \nOut4_8[6] , 
        \nScanOut171[3] , \nScanOut211[6] , \nScanOut325[5] , \nOut12_20[7] , 
        \nScanOut645[4] , \nScanOut771[7] , \nOut28_24[7] , \nScanOut172[0] , 
        \nScanOut212[5] , \nScanOut411[2] , \nScanOut525[1] , \nOut21_14[6] , 
        \nScanOut646[7] , \nScanOut772[4] , \nOut8_9[7] , \nScanOut326[6] , 
        \nScanOut412[1] , \nScanOut526[2] , \nOut21_17[5] , \nOut28_27[4] , 
        \nOut12_23[4] , \nOut24_28[1] , \nScanOut694[1] , \nScanOut813[0] , 
        \nOut3_29[2] , \nOut6_16[6] , \nScanOut927[3] , \nOut17_8[3] , 
        \nOut11_8[7] , \nScanOut115[7] , \nOut5_20[3] , \nScanOut275[2] , 
        \nScanOut621[0] , \nScanOut715[3] , \nScanOut992[2] , \nScanOut341[1] , 
        \nScanOut475[6] , \nScanOut541[5] , \nScanOut874[7] , \nScanOut17[7] , 
        \nOut11_15[1] , \nScanOut393[7] , \nScanOut940[4] , \nOut31_26[3] , 
        \nScanOut390[4] , \nOut18_25[0] , \nScanOut593[3] , \nOut22_21[0] , 
        \nScanOut1004[1] , \nOut31_25[0] , \nScanOut877[4] , \nScanOut943[7] , 
        \nOut0_23[3] , \nOut2_10[6] , \nScanOut116[4] , \nOut5_23[0] , 
        \nScanOut276[1] , \nOut11_16[2] , \nOut14_29[6] , \nOut18_26[3] , 
        \nOut22_22[3] , \nScanOut590[0] , \nScanOut1007[2] , \nScanOut342[2] , 
        \nOut20_9[2] , \nScanOut622[3] , \nScanOut716[0] , \nOut26_9[6] , 
        \nScanOut991[1] , \nOut3_31[0] , \nScanOut476[5] , \nScanOut542[6] , 
        \nOut16_25[4] , \nOut24_30[3] , \nOut25_11[5] , \nOut2_13[5] , 
        \nOut1_25[0] , \nScanOut68[2] , \nScanOut808[1] , \nScanOut169[1] , 
        \nScanOut209[4] , \nScanOut769[5] , \nOut8_15[1] , \nScanOut388[6] , 
        \nOut13_19[3] , \nScanOut409[0] , \nOut16_26[7] , \nOut25_12[6] , 
        \nOut15_10[2] , \nOut14_31[4] , \nScanOut588[2] , \nOut26_24[3] , 
        \nOut1_26[3] , \nScanOut639[2] , \nOut31_4[5] , \nScanOut989[3] , 
        \nOut4_19[7] , \nScanOut129[3] , \nOut8_16[2] , \nScanOut359[3] , 
        \nOut15_13[1] , \nScanOut559[7] , \nOut23_18[4] , \nOut26_27[0] , 
        \nScanOut958[6] , \nOut31_7[6] , \nScanOut249[6] , \nScanOut449[2] , 
        \nOut21_2[6] , \nOut19_6[7] , \nOut9_13[2] , \nOut6_7[3] , 
        \nOut11_29[5] , \nOut14_16[1] , \nScanOut729[7] , \nOut27_2[2] , 
        \nOut15_7[6] , \nOut18_19[4] , \nOut27_22[0] , \nScanOut28[0] , 
        \nOut13_7[2] , \nScanOut848[3] , \nOut6_4[0] , \nOut27_21[3] , 
        \nOut13_4[1] , \nOut14_15[2] , \nOut15_4[5] , \nScanOut498[7] , 
        \nOut0_20[0] , \nScanOut298[3] , \nOut21_1[5] , \nOut31_19[4] , 
        \nOut27_1[1] , \nScanOut30[2] , \nScanOut33[1] , \nOut3_3[6] , 
        \nOut9_10[1] , \nOut8_31[7] , \nOut19_5[4] , \nScanOut899[6] , 
        \nOut10_3[3] , \nOut3_15[6] , \nOut3_16[5] , \nOut5_3[2] , 
        \nOut6_29[1] , \nScanOut918[4] , \nOut28_7[2] , \nOut3_0[5] , 
        \nOut9_1[0] , \nOut9_2[3] , \nOut16_3[7] , \nScanOut319[1] , 
        \nScanOut519[5] , \nOut24_6[3] , \nOut17_23[7] , \nOut21_28[2] , 
        \nScanOut679[0] , \nOut24_17[6] , \nOut28_18[3] , \nOut22_6[7] , 
        \nOut24_14[5] , \nOut17_20[4] , \nOut24_5[0] , \nOut22_5[4] , 
        \nOut10_0[0] , \nOut5_0[1] , \nOut16_0[4] , \nOut28_4[1] , 
        \nOut10_13[2] , \nOut26_18[7] , \nScanOut480[5] , \nScanOut1023[4] , 
        \nOut19_23[3] , \nOut23_27[3] , \nScanOut853[2] , \nOut1_19[4] , 
        \nScanOut132[2] , \nScanOut280[1] , \nScanOut967[1] , \nScanOut452[3] , 
        \nScanOut566[0] , \nOut30_20[0] , \nOut4_25[3] , \nOut4_26[0] , 
        \nScanOut252[7] , \nScanOut606[5] , \nScanOut881[4] , \nScanOut732[6] , 
        \nOut8_29[5] , \nScanOut366[4] , \nScanOut131[1] , \nScanOut251[4] , 
        \nScanOut451[0] , \nScanOut565[3] , \nScanOut365[7] , \nScanOut283[2] , 
        \nOut10_10[1] , \nOut19_20[0] , \nScanOut605[6] , \nScanOut731[5] , 
        \nScanOut882[7] , \nOut23_24[0] , \nOut11_31[7] , \nScanOut483[6] , 
        \nScanOut1020[7] , \nScanOut850[1] , \nOut30_23[3] , \nScanOut964[2] , 
        \nOut13_26[4] , \nOut29_22[4] , \nScanOut54[6] , \nScanOut57[5] , 
        \nScanOut85[3] , \nScanOut156[6] , \nScanOut236[3] , \nScanOut436[7] , 
        \nScanOut502[4] , \nOut16_19[0] , \nOut20_12[5] , \nScanOut302[0] , 
        \nScanOut662[1] , \nScanOut756[2] , \nScanOut184[0] , \nOut7_13[6] , 
        \nScanOut837[6] , \nScanOut784[4] , \nScanOut903[5] , \nScanOut187[3] , 
        \nScanOut787[7] , \nScanOut834[5] , \nOut7_10[5] , \nOut6_31[3] , 
        \nScanOut900[6] , \nScanOut435[4] , \nScanOut501[7] , \nOut21_30[0] , 
        \nOut20_11[6] , \nScanOut86[0] , \nScanOut155[5] , \nOut29_21[7] , 
        \nOut13_25[7] , \nScanOut661[2] , \nScanOut755[1] , \nScanOut235[0] , 
        \nScanOut301[3] ;
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_19 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut20[7] , \nScanOut20[6] , 
        \nScanOut20[5] , \nScanOut20[4] , \nScanOut20[3] , \nScanOut20[2] , 
        \nScanOut20[1] , \nScanOut20[0] }), .ScanOut({\nScanOut19[7] , 
        \nScanOut19[6] , \nScanOut19[5] , \nScanOut19[4] , \nScanOut19[3] , 
        \nScanOut19[2] , \nScanOut19[1] , \nScanOut19[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_19[7] , \nOut0_19[6] , 
        \nOut0_19[5] , \nOut0_19[4] , \nOut0_19[3] , \nOut0_19[2] , 
        \nOut0_19[1] , \nOut0_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_25 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut26[7] , \nScanOut26[6] , 
        \nScanOut26[5] , \nScanOut26[4] , \nScanOut26[3] , \nScanOut26[2] , 
        \nScanOut26[1] , \nScanOut26[0] }), .ScanOut({\nScanOut25[7] , 
        \nScanOut25[6] , \nScanOut25[5] , \nScanOut25[4] , \nScanOut25[3] , 
        \nScanOut25[2] , \nScanOut25[1] , \nScanOut25[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_25[7] , \nOut0_25[6] , 
        \nOut0_25[5] , \nOut0_25[4] , \nOut0_25[3] , \nOut0_25[2] , 
        \nOut0_25[1] , \nOut0_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_89 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut90[7] , \nScanOut90[6] , 
        \nScanOut90[5] , \nScanOut90[4] , \nScanOut90[3] , \nScanOut90[2] , 
        \nScanOut90[1] , \nScanOut90[0] }), .ScanOut({\nScanOut89[7] , 
        \nScanOut89[6] , \nScanOut89[5] , \nScanOut89[4] , \nScanOut89[3] , 
        \nScanOut89[2] , \nScanOut89[1] , \nScanOut89[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_24[7] , \nOut2_24[6] , \nOut2_24[5] , \nOut2_24[4] , 
        \nOut2_24[3] , \nOut2_24[2] , \nOut2_24[1] , \nOut2_24[0] }), 
        .SouthIn({\nOut2_26[7] , \nOut2_26[6] , \nOut2_26[5] , \nOut2_26[4] , 
        \nOut2_26[3] , \nOut2_26[2] , \nOut2_26[1] , \nOut2_26[0] }), .EastIn(
        {\nOut3_25[7] , \nOut3_25[6] , \nOut3_25[5] , \nOut3_25[4] , 
        \nOut3_25[3] , \nOut3_25[2] , \nOut3_25[1] , \nOut3_25[0] }), .WestIn(
        {\nOut1_25[7] , \nOut1_25[6] , \nOut1_25[5] , \nOut1_25[4] , 
        \nOut1_25[3] , \nOut1_25[2] , \nOut1_25[1] , \nOut1_25[0] }), .Out({
        \nOut2_25[7] , \nOut2_25[6] , \nOut2_25[5] , \nOut2_25[4] , 
        \nOut2_25[3] , \nOut2_25[2] , \nOut2_25[1] , \nOut2_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_869 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut870[7] , \nScanOut870[6] , 
        \nScanOut870[5] , \nScanOut870[4] , \nScanOut870[3] , \nScanOut870[2] , 
        \nScanOut870[1] , \nScanOut870[0] }), .ScanOut({\nScanOut869[7] , 
        \nScanOut869[6] , \nScanOut869[5] , \nScanOut869[4] , \nScanOut869[3] , 
        \nScanOut869[2] , \nScanOut869[1] , \nScanOut869[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_4[7] , \nOut27_4[6] , \nOut27_4[5] , \nOut27_4[4] , 
        \nOut27_4[3] , \nOut27_4[2] , \nOut27_4[1] , \nOut27_4[0] }), 
        .SouthIn({\nOut27_6[7] , \nOut27_6[6] , \nOut27_6[5] , \nOut27_6[4] , 
        \nOut27_6[3] , \nOut27_6[2] , \nOut27_6[1] , \nOut27_6[0] }), .EastIn(
        {\nOut28_5[7] , \nOut28_5[6] , \nOut28_5[5] , \nOut28_5[4] , 
        \nOut28_5[3] , \nOut28_5[2] , \nOut28_5[1] , \nOut28_5[0] }), .WestIn(
        {\nOut26_5[7] , \nOut26_5[6] , \nOut26_5[5] , \nOut26_5[4] , 
        \nOut26_5[3] , \nOut26_5[2] , \nOut26_5[1] , \nOut26_5[0] }), .Out({
        \nOut27_5[7] , \nOut27_5[6] , \nOut27_5[5] , \nOut27_5[4] , 
        \nOut27_5[3] , \nOut27_5[2] , \nOut27_5[1] , \nOut27_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_281 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut282[7] , \nScanOut282[6] , 
        \nScanOut282[5] , \nScanOut282[4] , \nScanOut282[3] , \nScanOut282[2] , 
        \nScanOut282[1] , \nScanOut282[0] }), .ScanOut({\nScanOut281[7] , 
        \nScanOut281[6] , \nScanOut281[5] , \nScanOut281[4] , \nScanOut281[3] , 
        \nScanOut281[2] , \nScanOut281[1] , \nScanOut281[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_24[7] , \nOut8_24[6] , \nOut8_24[5] , \nOut8_24[4] , 
        \nOut8_24[3] , \nOut8_24[2] , \nOut8_24[1] , \nOut8_24[0] }), 
        .SouthIn({\nOut8_26[7] , \nOut8_26[6] , \nOut8_26[5] , \nOut8_26[4] , 
        \nOut8_26[3] , \nOut8_26[2] , \nOut8_26[1] , \nOut8_26[0] }), .EastIn(
        {\nOut9_25[7] , \nOut9_25[6] , \nOut9_25[5] , \nOut9_25[4] , 
        \nOut9_25[3] , \nOut9_25[2] , \nOut9_25[1] , \nOut9_25[0] }), .WestIn(
        {\nOut7_25[7] , \nOut7_25[6] , \nOut7_25[5] , \nOut7_25[4] , 
        \nOut7_25[3] , \nOut7_25[2] , \nOut7_25[1] , \nOut7_25[0] }), .Out({
        \nOut8_25[7] , \nOut8_25[6] , \nOut8_25[5] , \nOut8_25[4] , 
        \nOut8_25[3] , \nOut8_25[2] , \nOut8_25[1] , \nOut8_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_500 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut501[7] , \nScanOut501[6] , 
        \nScanOut501[5] , \nScanOut501[4] , \nScanOut501[3] , \nScanOut501[2] , 
        \nScanOut501[1] , \nScanOut501[0] }), .ScanOut({\nScanOut500[7] , 
        \nScanOut500[6] , \nScanOut500[5] , \nScanOut500[4] , \nScanOut500[3] , 
        \nScanOut500[2] , \nScanOut500[1] , \nScanOut500[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_19[7] , \nOut15_19[6] , \nOut15_19[5] , \nOut15_19[4] , 
        \nOut15_19[3] , \nOut15_19[2] , \nOut15_19[1] , \nOut15_19[0] }), 
        .SouthIn({\nOut15_21[7] , \nOut15_21[6] , \nOut15_21[5] , 
        \nOut15_21[4] , \nOut15_21[3] , \nOut15_21[2] , \nOut15_21[1] , 
        \nOut15_21[0] }), .EastIn({\nOut16_20[7] , \nOut16_20[6] , 
        \nOut16_20[5] , \nOut16_20[4] , \nOut16_20[3] , \nOut16_20[2] , 
        \nOut16_20[1] , \nOut16_20[0] }), .WestIn({\nOut14_20[7] , 
        \nOut14_20[6] , \nOut14_20[5] , \nOut14_20[4] , \nOut14_20[3] , 
        \nOut14_20[2] , \nOut14_20[1] , \nOut14_20[0] }), .Out({\nOut15_20[7] , 
        \nOut15_20[6] , \nOut15_20[5] , \nOut15_20[4] , \nOut15_20[3] , 
        \nOut15_20[2] , \nOut15_20[1] , \nOut15_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_311 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut312[7] , \nScanOut312[6] , 
        \nScanOut312[5] , \nScanOut312[4] , \nScanOut312[3] , \nScanOut312[2] , 
        \nScanOut312[1] , \nScanOut312[0] }), .ScanOut({\nScanOut311[7] , 
        \nScanOut311[6] , \nScanOut311[5] , \nScanOut311[4] , \nScanOut311[3] , 
        \nScanOut311[2] , \nScanOut311[1] , \nScanOut311[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_22[7] , \nOut9_22[6] , \nOut9_22[5] , \nOut9_22[4] , 
        \nOut9_22[3] , \nOut9_22[2] , \nOut9_22[1] , \nOut9_22[0] }), 
        .SouthIn({\nOut9_24[7] , \nOut9_24[6] , \nOut9_24[5] , \nOut9_24[4] , 
        \nOut9_24[3] , \nOut9_24[2] , \nOut9_24[1] , \nOut9_24[0] }), .EastIn(
        {\nOut10_23[7] , \nOut10_23[6] , \nOut10_23[5] , \nOut10_23[4] , 
        \nOut10_23[3] , \nOut10_23[2] , \nOut10_23[1] , \nOut10_23[0] }), 
        .WestIn({\nOut8_23[7] , \nOut8_23[6] , \nOut8_23[5] , \nOut8_23[4] , 
        \nOut8_23[3] , \nOut8_23[2] , \nOut8_23[1] , \nOut8_23[0] }), .Out({
        \nOut9_23[7] , \nOut9_23[6] , \nOut9_23[5] , \nOut9_23[4] , 
        \nOut9_23[3] , \nOut9_23[2] , \nOut9_23[1] , \nOut9_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_490 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut491[7] , \nScanOut491[6] , 
        \nScanOut491[5] , \nScanOut491[4] , \nScanOut491[3] , \nScanOut491[2] , 
        \nScanOut491[1] , \nScanOut491[0] }), .ScanOut({\nScanOut490[7] , 
        \nScanOut490[6] , \nScanOut490[5] , \nScanOut490[4] , \nScanOut490[3] , 
        \nScanOut490[2] , \nScanOut490[1] , \nScanOut490[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_9[7] , \nOut15_9[6] , \nOut15_9[5] , \nOut15_9[4] , 
        \nOut15_9[3] , \nOut15_9[2] , \nOut15_9[1] , \nOut15_9[0] }), 
        .SouthIn({\nOut15_11[7] , \nOut15_11[6] , \nOut15_11[5] , 
        \nOut15_11[4] , \nOut15_11[3] , \nOut15_11[2] , \nOut15_11[1] , 
        \nOut15_11[0] }), .EastIn({\nOut16_10[7] , \nOut16_10[6] , 
        \nOut16_10[5] , \nOut16_10[4] , \nOut16_10[3] , \nOut16_10[2] , 
        \nOut16_10[1] , \nOut16_10[0] }), .WestIn({\nOut14_10[7] , 
        \nOut14_10[6] , \nOut14_10[5] , \nOut14_10[4] , \nOut14_10[3] , 
        \nOut14_10[2] , \nOut14_10[1] , \nOut14_10[0] }), .Out({\nOut15_10[7] , 
        \nOut15_10[6] , \nOut15_10[5] , \nOut15_10[4] , \nOut15_10[3] , 
        \nOut15_10[2] , \nOut15_10[1] , \nOut15_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_972 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut973[7] , \nScanOut973[6] , 
        \nScanOut973[5] , \nScanOut973[4] , \nScanOut973[3] , \nScanOut973[2] , 
        \nScanOut973[1] , \nScanOut973[0] }), .ScanOut({\nScanOut972[7] , 
        \nScanOut972[6] , \nScanOut972[5] , \nScanOut972[4] , \nScanOut972[3] , 
        \nScanOut972[2] , \nScanOut972[1] , \nScanOut972[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_11[7] , \nOut30_11[6] , \nOut30_11[5] , \nOut30_11[4] , 
        \nOut30_11[3] , \nOut30_11[2] , \nOut30_11[1] , \nOut30_11[0] }), 
        .SouthIn({\nOut30_13[7] , \nOut30_13[6] , \nOut30_13[5] , 
        \nOut30_13[4] , \nOut30_13[3] , \nOut30_13[2] , \nOut30_13[1] , 
        \nOut30_13[0] }), .EastIn({\nOut31_12[7] , \nOut31_12[6] , 
        \nOut31_12[5] , \nOut31_12[4] , \nOut31_12[3] , \nOut31_12[2] , 
        \nOut31_12[1] , \nOut31_12[0] }), .WestIn({\nOut29_12[7] , 
        \nOut29_12[6] , \nOut29_12[5] , \nOut29_12[4] , \nOut29_12[3] , 
        \nOut29_12[2] , \nOut29_12[1] , \nOut29_12[0] }), .Out({\nOut30_12[7] , 
        \nOut30_12[6] , \nOut30_12[5] , \nOut30_12[4] , \nOut30_12[3] , 
        \nOut30_12[2] , \nOut30_12[1] , \nOut30_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_50 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut51[7] , \nScanOut51[6] , 
        \nScanOut51[5] , \nScanOut51[4] , \nScanOut51[3] , \nScanOut51[2] , 
        \nScanOut51[1] , \nScanOut51[0] }), .ScanOut({\nScanOut50[7] , 
        \nScanOut50[6] , \nScanOut50[5] , \nScanOut50[4] , \nScanOut50[3] , 
        \nScanOut50[2] , \nScanOut50[1] , \nScanOut50[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_17[7] , \nOut1_17[6] , \nOut1_17[5] , \nOut1_17[4] , 
        \nOut1_17[3] , \nOut1_17[2] , \nOut1_17[1] , \nOut1_17[0] }), 
        .SouthIn({\nOut1_19[7] , \nOut1_19[6] , \nOut1_19[5] , \nOut1_19[4] , 
        \nOut1_19[3] , \nOut1_19[2] , \nOut1_19[1] , \nOut1_19[0] }), .EastIn(
        {\nOut2_18[7] , \nOut2_18[6] , \nOut2_18[5] , \nOut2_18[4] , 
        \nOut2_18[3] , \nOut2_18[2] , \nOut2_18[1] , \nOut2_18[0] }), .WestIn(
        {\nOut0_18[7] , \nOut0_18[6] , \nOut0_18[5] , \nOut0_18[4] , 
        \nOut0_18[3] , \nOut0_18[2] , \nOut0_18[1] , \nOut0_18[0] }), .Out({
        \nOut1_18[7] , \nOut1_18[6] , \nOut1_18[5] , \nOut1_18[4] , 
        \nOut1_18[3] , \nOut1_18[2] , \nOut1_18[1] , \nOut1_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_154 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut155[7] , \nScanOut155[6] , 
        \nScanOut155[5] , \nScanOut155[4] , \nScanOut155[3] , \nScanOut155[2] , 
        \nScanOut155[1] , \nScanOut155[0] }), .ScanOut({\nScanOut154[7] , 
        \nScanOut154[6] , \nScanOut154[5] , \nScanOut154[4] , \nScanOut154[3] , 
        \nScanOut154[2] , \nScanOut154[1] , \nScanOut154[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_25[7] , \nOut4_25[6] , \nOut4_25[5] , \nOut4_25[4] , 
        \nOut4_25[3] , \nOut4_25[2] , \nOut4_25[1] , \nOut4_25[0] }), 
        .SouthIn({\nOut4_27[7] , \nOut4_27[6] , \nOut4_27[5] , \nOut4_27[4] , 
        \nOut4_27[3] , \nOut4_27[2] , \nOut4_27[1] , \nOut4_27[0] }), .EastIn(
        {\nOut5_26[7] , \nOut5_26[6] , \nOut5_26[5] , \nOut5_26[4] , 
        \nOut5_26[3] , \nOut5_26[2] , \nOut5_26[1] , \nOut5_26[0] }), .WestIn(
        {\nOut3_26[7] , \nOut3_26[6] , \nOut3_26[5] , \nOut3_26[4] , 
        \nOut3_26[3] , \nOut3_26[2] , \nOut3_26[1] , \nOut3_26[0] }), .Out({
        \nOut4_26[7] , \nOut4_26[6] , \nOut4_26[5] , \nOut4_26[4] , 
        \nOut4_26[3] , \nOut4_26[2] , \nOut4_26[1] , \nOut4_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_173 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut174[7] , \nScanOut174[6] , 
        \nScanOut174[5] , \nScanOut174[4] , \nScanOut174[3] , \nScanOut174[2] , 
        \nScanOut174[1] , \nScanOut174[0] }), .ScanOut({\nScanOut173[7] , 
        \nScanOut173[6] , \nScanOut173[5] , \nScanOut173[4] , \nScanOut173[3] , 
        \nScanOut173[2] , \nScanOut173[1] , \nScanOut173[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }), 
        .SouthIn({\nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }), .EastIn(
        {\nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }), .WestIn(
        {\nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }), .Out({
        \nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_196 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut197[7] , \nScanOut197[6] , 
        \nScanOut197[5] , \nScanOut197[4] , \nScanOut197[3] , \nScanOut197[2] , 
        \nScanOut197[1] , \nScanOut197[0] }), .ScanOut({\nScanOut196[7] , 
        \nScanOut196[6] , \nScanOut196[5] , \nScanOut196[4] , \nScanOut196[3] , 
        \nScanOut196[2] , \nScanOut196[1] , \nScanOut196[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_3[7] , \nOut6_3[6] , \nOut6_3[5] , \nOut6_3[4] , \nOut6_3[3] , 
        \nOut6_3[2] , \nOut6_3[1] , \nOut6_3[0] }), .SouthIn({\nOut6_5[7] , 
        \nOut6_5[6] , \nOut6_5[5] , \nOut6_5[4] , \nOut6_5[3] , \nOut6_5[2] , 
        \nOut6_5[1] , \nOut6_5[0] }), .EastIn({\nOut7_4[7] , \nOut7_4[6] , 
        \nOut7_4[5] , \nOut7_4[4] , \nOut7_4[3] , \nOut7_4[2] , \nOut7_4[1] , 
        \nOut7_4[0] }), .WestIn({\nOut5_4[7] , \nOut5_4[6] , \nOut5_4[5] , 
        \nOut5_4[4] , \nOut5_4[3] , \nOut5_4[2] , \nOut5_4[1] , \nOut5_4[0] }), 
        .Out({\nOut6_4[7] , \nOut6_4[6] , \nOut6_4[5] , \nOut6_4[4] , 
        \nOut6_4[3] , \nOut6_4[2] , \nOut6_4[1] , \nOut6_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_630 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut631[7] , \nScanOut631[6] , 
        \nScanOut631[5] , \nScanOut631[4] , \nScanOut631[3] , \nScanOut631[2] , 
        \nScanOut631[1] , \nScanOut631[0] }), .ScanOut({\nScanOut630[7] , 
        \nScanOut630[6] , \nScanOut630[5] , \nScanOut630[4] , \nScanOut630[3] , 
        \nScanOut630[2] , \nScanOut630[1] , \nScanOut630[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_21[7] , \nOut19_21[6] , \nOut19_21[5] , \nOut19_21[4] , 
        \nOut19_21[3] , \nOut19_21[2] , \nOut19_21[1] , \nOut19_21[0] }), 
        .SouthIn({\nOut19_23[7] , \nOut19_23[6] , \nOut19_23[5] , 
        \nOut19_23[4] , \nOut19_23[3] , \nOut19_23[2] , \nOut19_23[1] , 
        \nOut19_23[0] }), .EastIn({\nOut20_22[7] , \nOut20_22[6] , 
        \nOut20_22[5] , \nOut20_22[4] , \nOut20_22[3] , \nOut20_22[2] , 
        \nOut20_22[1] , \nOut20_22[0] }), .WestIn({\nOut18_22[7] , 
        \nOut18_22[6] , \nOut18_22[5] , \nOut18_22[4] , \nOut18_22[3] , 
        \nOut18_22[2] , \nOut18_22[1] , \nOut18_22[0] }), .Out({\nOut19_22[7] , 
        \nOut19_22[6] , \nOut19_22[5] , \nOut19_22[4] , \nOut19_22[3] , 
        \nOut19_22[2] , \nOut19_22[1] , \nOut19_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_787 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut788[7] , \nScanOut788[6] , 
        \nScanOut788[5] , \nScanOut788[4] , \nScanOut788[3] , \nScanOut788[2] , 
        \nScanOut788[1] , \nScanOut788[0] }), .ScanOut({\nScanOut787[7] , 
        \nScanOut787[6] , \nScanOut787[5] , \nScanOut787[4] , \nScanOut787[3] , 
        \nScanOut787[2] , \nScanOut787[1] , \nScanOut787[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_18[7] , \nOut24_18[6] , \nOut24_18[5] , \nOut24_18[4] , 
        \nOut24_18[3] , \nOut24_18[2] , \nOut24_18[1] , \nOut24_18[0] }), 
        .SouthIn({\nOut24_20[7] , \nOut24_20[6] , \nOut24_20[5] , 
        \nOut24_20[4] , \nOut24_20[3] , \nOut24_20[2] , \nOut24_20[1] , 
        \nOut24_20[0] }), .EastIn({\nOut25_19[7] , \nOut25_19[6] , 
        \nOut25_19[5] , \nOut25_19[4] , \nOut25_19[3] , \nOut25_19[2] , 
        \nOut25_19[1] , \nOut25_19[0] }), .WestIn({\nOut23_19[7] , 
        \nOut23_19[6] , \nOut23_19[5] , \nOut23_19[4] , \nOut23_19[3] , 
        \nOut23_19[2] , \nOut23_19[1] , \nOut23_19[0] }), .Out({\nOut24_19[7] , 
        \nOut24_19[6] , \nOut24_19[5] , \nOut24_19[4] , \nOut24_19[3] , 
        \nOut24_19[2] , \nOut24_19[1] , \nOut24_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_336 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut337[7] , \nScanOut337[6] , 
        \nScanOut337[5] , \nScanOut337[4] , \nScanOut337[3] , \nScanOut337[2] , 
        \nScanOut337[1] , \nScanOut337[0] }), .ScanOut({\nScanOut336[7] , 
        \nScanOut336[6] , \nScanOut336[5] , \nScanOut336[4] , \nScanOut336[3] , 
        \nScanOut336[2] , \nScanOut336[1] , \nScanOut336[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_15[7] , \nOut10_15[6] , \nOut10_15[5] , \nOut10_15[4] , 
        \nOut10_15[3] , \nOut10_15[2] , \nOut10_15[1] , \nOut10_15[0] }), 
        .SouthIn({\nOut10_17[7] , \nOut10_17[6] , \nOut10_17[5] , 
        \nOut10_17[4] , \nOut10_17[3] , \nOut10_17[2] , \nOut10_17[1] , 
        \nOut10_17[0] }), .EastIn({\nOut11_16[7] , \nOut11_16[6] , 
        \nOut11_16[5] , \nOut11_16[4] , \nOut11_16[3] , \nOut11_16[2] , 
        \nOut11_16[1] , \nOut11_16[0] }), .WestIn({\nOut9_16[7] , 
        \nOut9_16[6] , \nOut9_16[5] , \nOut9_16[4] , \nOut9_16[3] , 
        \nOut9_16[2] , \nOut9_16[1] , \nOut9_16[0] }), .Out({\nOut10_16[7] , 
        \nOut10_16[6] , \nOut10_16[5] , \nOut10_16[4] , \nOut10_16[3] , 
        \nOut10_16[2] , \nOut10_16[1] , \nOut10_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_617 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut618[7] , \nScanOut618[6] , 
        \nScanOut618[5] , \nScanOut618[4] , \nScanOut618[3] , \nScanOut618[2] , 
        \nScanOut618[1] , \nScanOut618[0] }), .ScanOut({\nScanOut617[7] , 
        \nScanOut617[6] , \nScanOut617[5] , \nScanOut617[4] , \nScanOut617[3] , 
        \nScanOut617[2] , \nScanOut617[1] , \nScanOut617[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_8[7] , \nOut19_8[6] , \nOut19_8[5] , \nOut19_8[4] , 
        \nOut19_8[3] , \nOut19_8[2] , \nOut19_8[1] , \nOut19_8[0] }), 
        .SouthIn({\nOut19_10[7] , \nOut19_10[6] , \nOut19_10[5] , 
        \nOut19_10[4] , \nOut19_10[3] , \nOut19_10[2] , \nOut19_10[1] , 
        \nOut19_10[0] }), .EastIn({\nOut20_9[7] , \nOut20_9[6] , \nOut20_9[5] , 
        \nOut20_9[4] , \nOut20_9[3] , \nOut20_9[2] , \nOut20_9[1] , 
        \nOut20_9[0] }), .WestIn({\nOut18_9[7] , \nOut18_9[6] , \nOut18_9[5] , 
        \nOut18_9[4] , \nOut18_9[3] , \nOut18_9[2] , \nOut18_9[1] , 
        \nOut18_9[0] }), .Out({\nOut19_9[7] , \nOut19_9[6] , \nOut19_9[5] , 
        \nOut19_9[4] , \nOut19_9[3] , \nOut19_9[2] , \nOut19_9[1] , 
        \nOut19_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_358 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut359[7] , \nScanOut359[6] , 
        \nScanOut359[5] , \nScanOut359[4] , \nScanOut359[3] , \nScanOut359[2] , 
        \nScanOut359[1] , \nScanOut359[0] }), .ScanOut({\nScanOut358[7] , 
        \nScanOut358[6] , \nScanOut358[5] , \nScanOut358[4] , \nScanOut358[3] , 
        \nScanOut358[2] , \nScanOut358[1] , \nScanOut358[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }), 
        .SouthIn({\nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }), .EastIn(
        {\nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }), .WestIn(
        {\nOut10_6[7] , \nOut10_6[6] , \nOut10_6[5] , \nOut10_6[4] , 
        \nOut10_6[3] , \nOut10_6[2] , \nOut10_6[1] , \nOut10_6[0] }), .Out({
        \nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_527 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut528[7] , \nScanOut528[6] , 
        \nScanOut528[5] , \nScanOut528[4] , \nScanOut528[3] , \nScanOut528[2] , 
        \nScanOut528[1] , \nScanOut528[0] }), .ScanOut({\nScanOut527[7] , 
        \nScanOut527[6] , \nScanOut527[5] , \nScanOut527[4] , \nScanOut527[3] , 
        \nScanOut527[2] , \nScanOut527[1] , \nScanOut527[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_14[7] , \nOut16_14[6] , \nOut16_14[5] , \nOut16_14[4] , 
        \nOut16_14[3] , \nOut16_14[2] , \nOut16_14[1] , \nOut16_14[0] }), 
        .SouthIn({\nOut16_16[7] , \nOut16_16[6] , \nOut16_16[5] , 
        \nOut16_16[4] , \nOut16_16[3] , \nOut16_16[2] , \nOut16_16[1] , 
        \nOut16_16[0] }), .EastIn({\nOut17_15[7] , \nOut17_15[6] , 
        \nOut17_15[5] , \nOut17_15[4] , \nOut17_15[3] , \nOut17_15[2] , 
        \nOut17_15[1] , \nOut17_15[0] }), .WestIn({\nOut15_15[7] , 
        \nOut15_15[6] , \nOut15_15[5] , \nOut15_15[4] , \nOut15_15[3] , 
        \nOut15_15[2] , \nOut15_15[1] , \nOut15_15[0] }), .Out({\nOut16_15[7] , 
        \nOut16_15[6] , \nOut16_15[5] , \nOut16_15[4] , \nOut16_15[3] , 
        \nOut16_15[2] , \nOut16_15[1] , \nOut16_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_549 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut550[7] , \nScanOut550[6] , 
        \nScanOut550[5] , \nScanOut550[4] , \nScanOut550[3] , \nScanOut550[2] , 
        \nScanOut550[1] , \nScanOut550[0] }), .ScanOut({\nScanOut549[7] , 
        \nScanOut549[6] , \nScanOut549[5] , \nScanOut549[4] , \nScanOut549[3] , 
        \nScanOut549[2] , \nScanOut549[1] , \nScanOut549[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_4[7] , \nOut17_4[6] , \nOut17_4[5] , \nOut17_4[4] , 
        \nOut17_4[3] , \nOut17_4[2] , \nOut17_4[1] , \nOut17_4[0] }), 
        .SouthIn({\nOut17_6[7] , \nOut17_6[6] , \nOut17_6[5] , \nOut17_6[4] , 
        \nOut17_6[3] , \nOut17_6[2] , \nOut17_6[1] , \nOut17_6[0] }), .EastIn(
        {\nOut18_5[7] , \nOut18_5[6] , \nOut18_5[5] , \nOut18_5[4] , 
        \nOut18_5[3] , \nOut18_5[2] , \nOut18_5[1] , \nOut18_5[0] }), .WestIn(
        {\nOut16_5[7] , \nOut16_5[6] , \nOut16_5[5] , \nOut16_5[4] , 
        \nOut16_5[3] , \nOut16_5[2] , \nOut16_5[1] , \nOut16_5[0] }), .Out({
        \nOut17_5[7] , \nOut17_5[6] , \nOut17_5[5] , \nOut17_5[4] , 
        \nOut17_5[3] , \nOut17_5[2] , \nOut17_5[1] , \nOut17_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_679 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut680[7] , \nScanOut680[6] , 
        \nScanOut680[5] , \nScanOut680[4] , \nScanOut680[3] , \nScanOut680[2] , 
        \nScanOut680[1] , \nScanOut680[0] }), .ScanOut({\nScanOut679[7] , 
        \nScanOut679[6] , \nScanOut679[5] , \nScanOut679[4] , \nScanOut679[3] , 
        \nScanOut679[2] , \nScanOut679[1] , \nScanOut679[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_6[7] , \nOut21_6[6] , \nOut21_6[5] , \nOut21_6[4] , 
        \nOut21_6[3] , \nOut21_6[2] , \nOut21_6[1] , \nOut21_6[0] }), 
        .SouthIn({\nOut21_8[7] , \nOut21_8[6] , \nOut21_8[5] , \nOut21_8[4] , 
        \nOut21_8[3] , \nOut21_8[2] , \nOut21_8[1] , \nOut21_8[0] }), .EastIn(
        {\nOut22_7[7] , \nOut22_7[6] , \nOut22_7[5] , \nOut22_7[4] , 
        \nOut22_7[3] , \nOut22_7[2] , \nOut22_7[1] , \nOut22_7[0] }), .WestIn(
        {\nOut20_7[7] , \nOut20_7[6] , \nOut20_7[5] , \nOut20_7[4] , 
        \nOut20_7[3] , \nOut20_7[2] , \nOut20_7[1] , \nOut20_7[0] }), .Out({
        \nOut21_7[7] , \nOut21_7[6] , \nOut21_7[5] , \nOut21_7[4] , 
        \nOut21_7[3] , \nOut21_7[2] , \nOut21_7[1] , \nOut21_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_955 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut956[7] , \nScanOut956[6] , 
        \nScanOut956[5] , \nScanOut956[4] , \nScanOut956[3] , \nScanOut956[2] , 
        \nScanOut956[1] , \nScanOut956[0] }), .ScanOut({\nScanOut955[7] , 
        \nScanOut955[6] , \nScanOut955[5] , \nScanOut955[4] , \nScanOut955[3] , 
        \nScanOut955[2] , \nScanOut955[1] , \nScanOut955[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_26[7] , \nOut29_26[6] , \nOut29_26[5] , \nOut29_26[4] , 
        \nOut29_26[3] , \nOut29_26[2] , \nOut29_26[1] , \nOut29_26[0] }), 
        .SouthIn({\nOut29_28[7] , \nOut29_28[6] , \nOut29_28[5] , 
        \nOut29_28[4] , \nOut29_28[3] , \nOut29_28[2] , \nOut29_28[1] , 
        \nOut29_28[0] }), .EastIn({\nOut30_27[7] , \nOut30_27[6] , 
        \nOut30_27[5] , \nOut30_27[4] , \nOut30_27[3] , \nOut30_27[2] , 
        \nOut30_27[1] , \nOut30_27[0] }), .WestIn({\nOut28_27[7] , 
        \nOut28_27[6] , \nOut28_27[5] , \nOut28_27[4] , \nOut28_27[3] , 
        \nOut28_27[2] , \nOut28_27[1] , \nOut28_27[0] }), .Out({\nOut29_27[7] , 
        \nOut29_27[6] , \nOut29_27[5] , \nOut29_27[4] , \nOut29_27[3] , 
        \nOut29_27[2] , \nOut29_27[1] , \nOut29_27[0] }) );
    Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1 U_Jacobi_Control ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut0[7] , \nScanOut0[6] , 
        \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , \nScanOut0[2] , 
        \nScanOut0[1] , \nScanOut0[0] }), .ScanOut({\nScanOut1024[7] , 
        \nScanOut1024[6] , \nScanOut1024[5] , \nScanOut1024[4] , 
        \nScanOut1024[3] , \nScanOut1024[2] , \nScanOut1024[1] , 
        \nScanOut1024[0] }), .ScanEnable(\nScanEnable[0] ), .Id(1'b1), 
        .ScanId(1'b0), .Enable(\nEnable[0] ) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_243 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut244[7] , \nScanOut244[6] , 
        \nScanOut244[5] , \nScanOut244[4] , \nScanOut244[3] , \nScanOut244[2] , 
        \nScanOut244[1] , \nScanOut244[0] }), .ScanOut({\nScanOut243[7] , 
        \nScanOut243[6] , \nScanOut243[5] , \nScanOut243[4] , \nScanOut243[3] , 
        \nScanOut243[2] , \nScanOut243[1] , \nScanOut243[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_18[7] , \nOut7_18[6] , \nOut7_18[5] , \nOut7_18[4] , 
        \nOut7_18[3] , \nOut7_18[2] , \nOut7_18[1] , \nOut7_18[0] }), 
        .SouthIn({\nOut7_20[7] , \nOut7_20[6] , \nOut7_20[5] , \nOut7_20[4] , 
        \nOut7_20[3] , \nOut7_20[2] , \nOut7_20[1] , \nOut7_20[0] }), .EastIn(
        {\nOut8_19[7] , \nOut8_19[6] , \nOut8_19[5] , \nOut8_19[4] , 
        \nOut8_19[3] , \nOut8_19[2] , \nOut8_19[1] , \nOut8_19[0] }), .WestIn(
        {\nOut6_19[7] , \nOut6_19[6] , \nOut6_19[5] , \nOut6_19[4] , 
        \nOut6_19[3] , \nOut6_19[2] , \nOut6_19[1] , \nOut6_19[0] }), .Out({
        \nOut7_19[7] , \nOut7_19[6] , \nOut7_19[5] , \nOut7_19[4] , 
        \nOut7_19[3] , \nOut7_19[2] , \nOut7_19[1] , \nOut7_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_762 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut763[7] , \nScanOut763[6] , 
        \nScanOut763[5] , \nScanOut763[4] , \nScanOut763[3] , \nScanOut763[2] , 
        \nScanOut763[1] , \nScanOut763[0] }), .ScanOut({\nScanOut762[7] , 
        \nScanOut762[6] , \nScanOut762[5] , \nScanOut762[4] , \nScanOut762[3] , 
        \nScanOut762[2] , \nScanOut762[1] , \nScanOut762[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_25[7] , \nOut23_25[6] , \nOut23_25[5] , \nOut23_25[4] , 
        \nOut23_25[3] , \nOut23_25[2] , \nOut23_25[1] , \nOut23_25[0] }), 
        .SouthIn({\nOut23_27[7] , \nOut23_27[6] , \nOut23_27[5] , 
        \nOut23_27[4] , \nOut23_27[3] , \nOut23_27[2] , \nOut23_27[1] , 
        \nOut23_27[0] }), .EastIn({\nOut24_26[7] , \nOut24_26[6] , 
        \nOut24_26[5] , \nOut24_26[4] , \nOut24_26[3] , \nOut24_26[2] , 
        \nOut24_26[1] , \nOut24_26[0] }), .WestIn({\nOut22_26[7] , 
        \nOut22_26[6] , \nOut22_26[5] , \nOut22_26[4] , \nOut22_26[3] , 
        \nOut22_26[2] , \nOut22_26[1] , \nOut22_26[0] }), .Out({\nOut23_26[7] , 
        \nOut23_26[6] , \nOut23_26[5] , \nOut23_26[4] , \nOut23_26[3] , 
        \nOut23_26[2] , \nOut23_26[1] , \nOut23_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_264 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut265[7] , \nScanOut265[6] , 
        \nScanOut265[5] , \nScanOut265[4] , \nScanOut265[3] , \nScanOut265[2] , 
        \nScanOut265[1] , \nScanOut265[0] }), .ScanOut({\nScanOut264[7] , 
        \nScanOut264[6] , \nScanOut264[5] , \nScanOut264[4] , \nScanOut264[3] , 
        \nScanOut264[2] , \nScanOut264[1] , \nScanOut264[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_7[7] , \nOut8_7[6] , \nOut8_7[5] , \nOut8_7[4] , \nOut8_7[3] , 
        \nOut8_7[2] , \nOut8_7[1] , \nOut8_7[0] }), .SouthIn({\nOut8_9[7] , 
        \nOut8_9[6] , \nOut8_9[5] , \nOut8_9[4] , \nOut8_9[3] , \nOut8_9[2] , 
        \nOut8_9[1] , \nOut8_9[0] }), .EastIn({\nOut9_8[7] , \nOut9_8[6] , 
        \nOut9_8[5] , \nOut9_8[4] , \nOut9_8[3] , \nOut9_8[2] , \nOut9_8[1] , 
        \nOut9_8[0] }), .WestIn({\nOut7_8[7] , \nOut7_8[6] , \nOut7_8[5] , 
        \nOut7_8[4] , \nOut7_8[3] , \nOut7_8[2] , \nOut7_8[1] , \nOut7_8[0] }), 
        .Out({\nOut8_8[7] , \nOut8_8[6] , \nOut8_8[5] , \nOut8_8[4] , 
        \nOut8_8[3] , \nOut8_8[2] , \nOut8_8[1] , \nOut8_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_452 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut453[7] , \nScanOut453[6] , 
        \nScanOut453[5] , \nScanOut453[4] , \nScanOut453[3] , \nScanOut453[2] , 
        \nScanOut453[1] , \nScanOut453[0] }), .ScanOut({\nScanOut452[7] , 
        \nScanOut452[6] , \nScanOut452[5] , \nScanOut452[4] , \nScanOut452[3] , 
        \nScanOut452[2] , \nScanOut452[1] , \nScanOut452[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }), 
        .SouthIn({\nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }), .EastIn(
        {\nOut15_4[7] , \nOut15_4[6] , \nOut15_4[5] , \nOut15_4[4] , 
        \nOut15_4[3] , \nOut15_4[2] , \nOut15_4[1] , \nOut15_4[0] }), .WestIn(
        {\nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }), .Out({
        \nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_475 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut476[7] , \nScanOut476[6] , 
        \nScanOut476[5] , \nScanOut476[4] , \nScanOut476[3] , \nScanOut476[2] , 
        \nScanOut476[1] , \nScanOut476[0] }), .ScanOut({\nScanOut475[7] , 
        \nScanOut475[6] , \nScanOut475[5] , \nScanOut475[4] , \nScanOut475[3] , 
        \nScanOut475[2] , \nScanOut475[1] , \nScanOut475[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_26[7] , \nOut14_26[6] , \nOut14_26[5] , \nOut14_26[4] , 
        \nOut14_26[3] , \nOut14_26[2] , \nOut14_26[1] , \nOut14_26[0] }), 
        .SouthIn({\nOut14_28[7] , \nOut14_28[6] , \nOut14_28[5] , 
        \nOut14_28[4] , \nOut14_28[3] , \nOut14_28[2] , \nOut14_28[1] , 
        \nOut14_28[0] }), .EastIn({\nOut15_27[7] , \nOut15_27[6] , 
        \nOut15_27[5] , \nOut15_27[4] , \nOut15_27[3] , \nOut15_27[2] , 
        \nOut15_27[1] , \nOut15_27[0] }), .WestIn({\nOut13_27[7] , 
        \nOut13_27[6] , \nOut13_27[5] , \nOut13_27[4] , \nOut13_27[3] , 
        \nOut13_27[2] , \nOut13_27[1] , \nOut13_27[0] }), .Out({\nOut14_27[7] , 
        \nOut14_27[6] , \nOut14_27[5] , \nOut14_27[4] , \nOut14_27[3] , 
        \nOut14_27[2] , \nOut14_27[1] , \nOut14_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_820 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut821[7] , \nScanOut821[6] , 
        \nScanOut821[5] , \nScanOut821[4] , \nScanOut821[3] , \nScanOut821[2] , 
        \nScanOut821[1] , \nScanOut821[0] }), .ScanOut({\nScanOut820[7] , 
        \nScanOut820[6] , \nScanOut820[5] , \nScanOut820[4] , \nScanOut820[3] , 
        \nScanOut820[2] , \nScanOut820[1] , \nScanOut820[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_19[7] , \nOut25_19[6] , \nOut25_19[5] , \nOut25_19[4] , 
        \nOut25_19[3] , \nOut25_19[2] , \nOut25_19[1] , \nOut25_19[0] }), 
        .SouthIn({\nOut25_21[7] , \nOut25_21[6] , \nOut25_21[5] , 
        \nOut25_21[4] , \nOut25_21[3] , \nOut25_21[2] , \nOut25_21[1] , 
        \nOut25_21[0] }), .EastIn({\nOut26_20[7] , \nOut26_20[6] , 
        \nOut26_20[5] , \nOut26_20[4] , \nOut26_20[3] , \nOut26_20[2] , 
        \nOut26_20[1] , \nOut26_20[0] }), .WestIn({\nOut24_20[7] , 
        \nOut24_20[6] , \nOut24_20[5] , \nOut24_20[4] , \nOut24_20[3] , 
        \nOut24_20[2] , \nOut24_20[1] , \nOut24_20[0] }), .Out({\nOut25_20[7] , 
        \nOut25_20[6] , \nOut25_20[5] , \nOut25_20[4] , \nOut25_20[3] , 
        \nOut25_20[2] , \nOut25_20[1] , \nOut25_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_745 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut746[7] , \nScanOut746[6] , 
        \nScanOut746[5] , \nScanOut746[4] , \nScanOut746[3] , \nScanOut746[2] , 
        \nScanOut746[1] , \nScanOut746[0] }), .ScanOut({\nScanOut745[7] , 
        \nScanOut745[6] , \nScanOut745[5] , \nScanOut745[4] , \nScanOut745[3] , 
        \nScanOut745[2] , \nScanOut745[1] , \nScanOut745[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_8[7] , \nOut23_8[6] , \nOut23_8[5] , \nOut23_8[4] , 
        \nOut23_8[3] , \nOut23_8[2] , \nOut23_8[1] , \nOut23_8[0] }), 
        .SouthIn({\nOut23_10[7] , \nOut23_10[6] , \nOut23_10[5] , 
        \nOut23_10[4] , \nOut23_10[3] , \nOut23_10[2] , \nOut23_10[1] , 
        \nOut23_10[0] }), .EastIn({\nOut24_9[7] , \nOut24_9[6] , \nOut24_9[5] , 
        \nOut24_9[4] , \nOut24_9[3] , \nOut24_9[2] , \nOut24_9[1] , 
        \nOut24_9[0] }), .WestIn({\nOut22_9[7] , \nOut22_9[6] , \nOut22_9[5] , 
        \nOut22_9[4] , \nOut22_9[3] , \nOut22_9[2] , \nOut22_9[1] , 
        \nOut22_9[0] }), .Out({\nOut23_9[7] , \nOut23_9[6] , \nOut23_9[5] , 
        \nOut23_9[4] , \nOut23_9[3] , \nOut23_9[2] , \nOut23_9[1] , 
        \nOut23_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_807 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut808[7] , \nScanOut808[6] , 
        \nScanOut808[5] , \nScanOut808[4] , \nScanOut808[3] , \nScanOut808[2] , 
        \nScanOut808[1] , \nScanOut808[0] }), .ScanOut({\nScanOut807[7] , 
        \nScanOut807[6] , \nScanOut807[5] , \nScanOut807[4] , \nScanOut807[3] , 
        \nScanOut807[2] , \nScanOut807[1] , \nScanOut807[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_6[7] , \nOut25_6[6] , \nOut25_6[5] , \nOut25_6[4] , 
        \nOut25_6[3] , \nOut25_6[2] , \nOut25_6[1] , \nOut25_6[0] }), 
        .SouthIn({\nOut25_8[7] , \nOut25_8[6] , \nOut25_8[5] , \nOut25_8[4] , 
        \nOut25_8[3] , \nOut25_8[2] , \nOut25_8[1] , \nOut25_8[0] }), .EastIn(
        {\nOut26_7[7] , \nOut26_7[6] , \nOut26_7[5] , \nOut26_7[4] , 
        \nOut26_7[3] , \nOut26_7[2] , \nOut26_7[1] , \nOut26_7[0] }), .WestIn(
        {\nOut24_7[7] , \nOut24_7[6] , \nOut24_7[5] , \nOut24_7[4] , 
        \nOut24_7[3] , \nOut24_7[2] , \nOut24_7[1] , \nOut24_7[0] }), .Out({
        \nOut25_7[7] , \nOut25_7[6] , \nOut25_7[5] , \nOut25_7[4] , 
        \nOut25_7[3] , \nOut25_7[2] , \nOut25_7[1] , \nOut25_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_997 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut998[7] , \nScanOut998[6] , 
        \nScanOut998[5] , \nScanOut998[4] , \nScanOut998[3] , \nScanOut998[2] , 
        \nScanOut998[1] , \nScanOut998[0] }), .ScanOut({\nScanOut997[7] , 
        \nScanOut997[6] , \nScanOut997[5] , \nScanOut997[4] , \nScanOut997[3] , 
        \nScanOut997[2] , \nScanOut997[1] , \nScanOut997[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut31_5[7] , \nOut31_5[6] , 
        \nOut31_5[5] , \nOut31_5[4] , \nOut31_5[3] , \nOut31_5[2] , 
        \nOut31_5[1] , \nOut31_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_168 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut169[7] , \nScanOut169[6] , 
        \nScanOut169[5] , \nScanOut169[4] , \nScanOut169[3] , \nScanOut169[2] , 
        \nScanOut169[1] , \nScanOut169[0] }), .ScanOut({\nScanOut168[7] , 
        \nScanOut168[6] , \nScanOut168[5] , \nScanOut168[4] , \nScanOut168[3] , 
        \nScanOut168[2] , \nScanOut168[1] , \nScanOut168[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_7[7] , \nOut5_7[6] , \nOut5_7[5] , \nOut5_7[4] , \nOut5_7[3] , 
        \nOut5_7[2] , \nOut5_7[1] , \nOut5_7[0] }), .SouthIn({\nOut5_9[7] , 
        \nOut5_9[6] , \nOut5_9[5] , \nOut5_9[4] , \nOut5_9[3] , \nOut5_9[2] , 
        \nOut5_9[1] , \nOut5_9[0] }), .EastIn({\nOut6_8[7] , \nOut6_8[6] , 
        \nOut6_8[5] , \nOut6_8[4] , \nOut6_8[3] , \nOut6_8[2] , \nOut6_8[1] , 
        \nOut6_8[0] }), .WestIn({\nOut4_8[7] , \nOut4_8[6] , \nOut4_8[5] , 
        \nOut4_8[4] , \nOut4_8[3] , \nOut4_8[2] , \nOut4_8[1] , \nOut4_8[0] }), 
        .Out({\nOut5_8[7] , \nOut5_8[6] , \nOut5_8[5] , \nOut5_8[4] , 
        \nOut5_8[3] , \nOut5_8[2] , \nOut5_8[1] , \nOut5_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_258 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut259[7] , \nScanOut259[6] , 
        \nScanOut259[5] , \nScanOut259[4] , \nScanOut259[3] , \nScanOut259[2] , 
        \nScanOut259[1] , \nScanOut259[0] }), .ScanOut({\nScanOut258[7] , 
        \nScanOut258[6] , \nScanOut258[5] , \nScanOut258[4] , \nScanOut258[3] , 
        \nScanOut258[2] , \nScanOut258[1] , \nScanOut258[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_1[7] , \nOut8_1[6] , \nOut8_1[5] , \nOut8_1[4] , \nOut8_1[3] , 
        \nOut8_1[2] , \nOut8_1[1] , \nOut8_1[0] }), .SouthIn({\nOut8_3[7] , 
        \nOut8_3[6] , \nOut8_3[5] , \nOut8_3[4] , \nOut8_3[3] , \nOut8_3[2] , 
        \nOut8_3[1] , \nOut8_3[0] }), .EastIn({\nOut9_2[7] , \nOut9_2[6] , 
        \nOut9_2[5] , \nOut9_2[4] , \nOut9_2[3] , \nOut9_2[2] , \nOut9_2[1] , 
        \nOut9_2[0] }), .WestIn({\nOut7_2[7] , \nOut7_2[6] , \nOut7_2[5] , 
        \nOut7_2[4] , \nOut7_2[3] , \nOut7_2[2] , \nOut7_2[1] , \nOut7_2[0] }), 
        .Out({\nOut8_2[7] , \nOut8_2[6] , \nOut8_2[5] , \nOut8_2[4] , 
        \nOut8_2[3] , \nOut8_2[2] , \nOut8_2[1] , \nOut8_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_449 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut450[7] , \nScanOut450[6] , 
        \nScanOut450[5] , \nScanOut450[4] , \nScanOut450[3] , \nScanOut450[2] , 
        \nScanOut450[1] , \nScanOut450[0] }), .ScanOut({\nScanOut449[7] , 
        \nScanOut449[6] , \nScanOut449[5] , \nScanOut449[4] , \nScanOut449[3] , 
        \nScanOut449[2] , \nScanOut449[1] , \nScanOut449[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_0[7] , \nOut14_0[6] , \nOut14_0[5] , \nOut14_0[4] , 
        \nOut14_0[3] , \nOut14_0[2] , \nOut14_0[1] , \nOut14_0[0] }), 
        .SouthIn({\nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }), .EastIn(
        {\nOut15_1[7] , \nOut15_1[6] , \nOut15_1[5] , \nOut15_1[4] , 
        \nOut15_1[3] , \nOut15_1[2] , \nOut15_1[1] , \nOut15_1[0] }), .WestIn(
        {\nOut13_1[7] , \nOut13_1[6] , \nOut13_1[5] , \nOut13_1[4] , 
        \nOut13_1[3] , \nOut13_1[2] , \nOut13_1[1] , \nOut13_1[0] }), .Out({
        \nOut14_1[7] , \nOut14_1[6] , \nOut14_1[5] , \nOut14_1[4] , 
        \nOut14_1[3] , \nOut14_1[2] , \nOut14_1[1] , \nOut14_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_645 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut646[7] , \nScanOut646[6] , 
        \nScanOut646[5] , \nScanOut646[4] , \nScanOut646[3] , \nScanOut646[2] , 
        \nScanOut646[1] , \nScanOut646[0] }), .ScanOut({\nScanOut645[7] , 
        \nScanOut645[6] , \nScanOut645[5] , \nScanOut645[4] , \nScanOut645[3] , 
        \nScanOut645[2] , \nScanOut645[1] , \nScanOut645[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_4[7] , \nOut20_4[6] , \nOut20_4[5] , \nOut20_4[4] , 
        \nOut20_4[3] , \nOut20_4[2] , \nOut20_4[1] , \nOut20_4[0] }), 
        .SouthIn({\nOut20_6[7] , \nOut20_6[6] , \nOut20_6[5] , \nOut20_6[4] , 
        \nOut20_6[3] , \nOut20_6[2] , \nOut20_6[1] , \nOut20_6[0] }), .EastIn(
        {\nOut21_5[7] , \nOut21_5[6] , \nOut21_5[5] , \nOut21_5[4] , 
        \nOut21_5[3] , \nOut21_5[2] , \nOut21_5[1] , \nOut21_5[0] }), .WestIn(
        {\nOut19_5[7] , \nOut19_5[6] , \nOut19_5[5] , \nOut19_5[4] , 
        \nOut19_5[3] , \nOut19_5[2] , \nOut19_5[1] , \nOut19_5[0] }), .Out({
        \nOut20_5[7] , \nOut20_5[6] , \nOut20_5[5] , \nOut20_5[4] , 
        \nOut20_5[3] , \nOut20_5[2] , \nOut20_5[1] , \nOut20_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_779 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut780[7] , \nScanOut780[6] , 
        \nScanOut780[5] , \nScanOut780[4] , \nScanOut780[3] , \nScanOut780[2] , 
        \nScanOut780[1] , \nScanOut780[0] }), .ScanOut({\nScanOut779[7] , 
        \nScanOut779[6] , \nScanOut779[5] , \nScanOut779[4] , \nScanOut779[3] , 
        \nScanOut779[2] , \nScanOut779[1] , \nScanOut779[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_10[7] , \nOut24_10[6] , \nOut24_10[5] , \nOut24_10[4] , 
        \nOut24_10[3] , \nOut24_10[2] , \nOut24_10[1] , \nOut24_10[0] }), 
        .SouthIn({\nOut24_12[7] , \nOut24_12[6] , \nOut24_12[5] , 
        \nOut24_12[4] , \nOut24_12[3] , \nOut24_12[2] , \nOut24_12[1] , 
        \nOut24_12[0] }), .EastIn({\nOut25_11[7] , \nOut25_11[6] , 
        \nOut25_11[5] , \nOut25_11[4] , \nOut25_11[3] , \nOut25_11[2] , 
        \nOut25_11[1] , \nOut25_11[0] }), .WestIn({\nOut23_11[7] , 
        \nOut23_11[6] , \nOut23_11[5] , \nOut23_11[4] , \nOut23_11[3] , 
        \nOut23_11[2] , \nOut23_11[1] , \nOut23_11[0] }), .Out({\nOut24_11[7] , 
        \nOut24_11[6] , \nOut24_11[5] , \nOut24_11[4] , \nOut24_11[3] , 
        \nOut24_11[2] , \nOut24_11[1] , \nOut24_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_77 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut78[7] , \nScanOut78[6] , 
        \nScanOut78[5] , \nScanOut78[4] , \nScanOut78[3] , \nScanOut78[2] , 
        \nScanOut78[1] , \nScanOut78[0] }), .ScanOut({\nScanOut77[7] , 
        \nScanOut77[6] , \nScanOut77[5] , \nScanOut77[4] , \nScanOut77[3] , 
        \nScanOut77[2] , \nScanOut77[1] , \nScanOut77[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), 
        .SouthIn({\nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), .EastIn(
        {\nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }), .WestIn(
        {\nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), .Out({
        \nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_343 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut344[7] , \nScanOut344[6] , 
        \nScanOut344[5] , \nScanOut344[4] , \nScanOut344[3] , \nScanOut344[2] , 
        \nScanOut344[1] , \nScanOut344[0] }), .ScanOut({\nScanOut343[7] , 
        \nScanOut343[6] , \nScanOut343[5] , \nScanOut343[4] , \nScanOut343[3] , 
        \nScanOut343[2] , \nScanOut343[1] , \nScanOut343[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_22[7] , \nOut10_22[6] , \nOut10_22[5] , \nOut10_22[4] , 
        \nOut10_22[3] , \nOut10_22[2] , \nOut10_22[1] , \nOut10_22[0] }), 
        .SouthIn({\nOut10_24[7] , \nOut10_24[6] , \nOut10_24[5] , 
        \nOut10_24[4] , \nOut10_24[3] , \nOut10_24[2] , \nOut10_24[1] , 
        \nOut10_24[0] }), .EastIn({\nOut11_23[7] , \nOut11_23[6] , 
        \nOut11_23[5] , \nOut11_23[4] , \nOut11_23[3] , \nOut11_23[2] , 
        \nOut11_23[1] , \nOut11_23[0] }), .WestIn({\nOut9_23[7] , 
        \nOut9_23[6] , \nOut9_23[5] , \nOut9_23[4] , \nOut9_23[3] , 
        \nOut9_23[2] , \nOut9_23[1] , \nOut9_23[0] }), .Out({\nOut10_23[7] , 
        \nOut10_23[6] , \nOut10_23[5] , \nOut10_23[4] , \nOut10_23[3] , 
        \nOut10_23[2] , \nOut10_23[1] , \nOut10_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_364 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut365[7] , \nScanOut365[6] , 
        \nScanOut365[5] , \nScanOut365[4] , \nScanOut365[3] , \nScanOut365[2] , 
        \nScanOut365[1] , \nScanOut365[0] }), .ScanOut({\nScanOut364[7] , 
        \nScanOut364[6] , \nScanOut364[5] , \nScanOut364[4] , \nScanOut364[3] , 
        \nScanOut364[2] , \nScanOut364[1] , \nScanOut364[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_11[7] , \nOut11_11[6] , \nOut11_11[5] , \nOut11_11[4] , 
        \nOut11_11[3] , \nOut11_11[2] , \nOut11_11[1] , \nOut11_11[0] }), 
        .SouthIn({\nOut11_13[7] , \nOut11_13[6] , \nOut11_13[5] , 
        \nOut11_13[4] , \nOut11_13[3] , \nOut11_13[2] , \nOut11_13[1] , 
        \nOut11_13[0] }), .EastIn({\nOut12_12[7] , \nOut12_12[6] , 
        \nOut12_12[5] , \nOut12_12[4] , \nOut12_12[3] , \nOut12_12[2] , 
        \nOut12_12[1] , \nOut12_12[0] }), .WestIn({\nOut10_12[7] , 
        \nOut10_12[6] , \nOut10_12[5] , \nOut10_12[4] , \nOut10_12[3] , 
        \nOut10_12[2] , \nOut10_12[1] , \nOut10_12[0] }), .Out({\nOut11_12[7] , 
        \nOut11_12[6] , \nOut11_12[5] , \nOut11_12[4] , \nOut11_12[3] , 
        \nOut11_12[2] , \nOut11_12[1] , \nOut11_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_552 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut553[7] , \nScanOut553[6] , 
        \nScanOut553[5] , \nScanOut553[4] , \nScanOut553[3] , \nScanOut553[2] , 
        \nScanOut553[1] , \nScanOut553[0] }), .ScanOut({\nScanOut552[7] , 
        \nScanOut552[6] , \nScanOut552[5] , \nScanOut552[4] , \nScanOut552[3] , 
        \nScanOut552[2] , \nScanOut552[1] , \nScanOut552[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_7[7] , \nOut17_7[6] , \nOut17_7[5] , \nOut17_7[4] , 
        \nOut17_7[3] , \nOut17_7[2] , \nOut17_7[1] , \nOut17_7[0] }), 
        .SouthIn({\nOut17_9[7] , \nOut17_9[6] , \nOut17_9[5] , \nOut17_9[4] , 
        \nOut17_9[3] , \nOut17_9[2] , \nOut17_9[1] , \nOut17_9[0] }), .EastIn(
        {\nOut18_8[7] , \nOut18_8[6] , \nOut18_8[5] , \nOut18_8[4] , 
        \nOut18_8[3] , \nOut18_8[2] , \nOut18_8[1] , \nOut18_8[0] }), .WestIn(
        {\nOut16_8[7] , \nOut16_8[6] , \nOut16_8[5] , \nOut16_8[4] , 
        \nOut16_8[3] , \nOut16_8[2] , \nOut16_8[1] , \nOut16_8[0] }), .Out({
        \nOut17_8[7] , \nOut17_8[6] , \nOut17_8[5] , \nOut17_8[4] , 
        \nOut17_8[3] , \nOut17_8[2] , \nOut17_8[1] , \nOut17_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_575 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut576[7] , \nScanOut576[6] , 
        \nScanOut576[5] , \nScanOut576[4] , \nScanOut576[3] , \nScanOut576[2] , 
        \nScanOut576[1] , \nScanOut576[0] }), .ScanOut({\nScanOut575[7] , 
        \nScanOut575[6] , \nScanOut575[5] , \nScanOut575[4] , \nScanOut575[3] , 
        \nScanOut575[2] , \nScanOut575[1] , \nScanOut575[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut17_31[7] , \nOut17_31[6] , 
        \nOut17_31[5] , \nOut17_31[4] , \nOut17_31[3] , \nOut17_31[2] , 
        \nOut17_31[1] , \nOut17_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_897 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut898[7] , \nScanOut898[6] , 
        \nScanOut898[5] , \nScanOut898[4] , \nScanOut898[3] , \nScanOut898[2] , 
        \nScanOut898[1] , \nScanOut898[0] }), .ScanOut({\nScanOut897[7] , 
        \nScanOut897[6] , \nScanOut897[5] , \nScanOut897[4] , \nScanOut897[3] , 
        \nScanOut897[2] , \nScanOut897[1] , \nScanOut897[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_0[7] , \nOut28_0[6] , \nOut28_0[5] , \nOut28_0[4] , 
        \nOut28_0[3] , \nOut28_0[2] , \nOut28_0[1] , \nOut28_0[0] }), 
        .SouthIn({\nOut28_2[7] , \nOut28_2[6] , \nOut28_2[5] , \nOut28_2[4] , 
        \nOut28_2[3] , \nOut28_2[2] , \nOut28_2[1] , \nOut28_2[0] }), .EastIn(
        {\nOut29_1[7] , \nOut29_1[6] , \nOut29_1[5] , \nOut29_1[4] , 
        \nOut29_1[3] , \nOut29_1[2] , \nOut29_1[1] , \nOut29_1[0] }), .WestIn(
        {\nOut27_1[7] , \nOut27_1[6] , \nOut27_1[5] , \nOut27_1[4] , 
        \nOut27_1[3] , \nOut27_1[2] , \nOut27_1[1] , \nOut27_1[0] }), .Out({
        \nOut28_1[7] , \nOut28_1[6] , \nOut28_1[5] , \nOut28_1[4] , 
        \nOut28_1[3] , \nOut28_1[2] , \nOut28_1[1] , \nOut28_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_907 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut908[7] , \nScanOut908[6] , 
        \nScanOut908[5] , \nScanOut908[4] , \nScanOut908[3] , \nScanOut908[2] , 
        \nScanOut908[1] , \nScanOut908[0] }), .ScanOut({\nScanOut907[7] , 
        \nScanOut907[6] , \nScanOut907[5] , \nScanOut907[4] , \nScanOut907[3] , 
        \nScanOut907[2] , \nScanOut907[1] , \nScanOut907[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_10[7] , \nOut28_10[6] , \nOut28_10[5] , \nOut28_10[4] , 
        \nOut28_10[3] , \nOut28_10[2] , \nOut28_10[1] , \nOut28_10[0] }), 
        .SouthIn({\nOut28_12[7] , \nOut28_12[6] , \nOut28_12[5] , 
        \nOut28_12[4] , \nOut28_12[3] , \nOut28_12[2] , \nOut28_12[1] , 
        \nOut28_12[0] }), .EastIn({\nOut29_11[7] , \nOut29_11[6] , 
        \nOut29_11[5] , \nOut29_11[4] , \nOut29_11[3] , \nOut29_11[2] , 
        \nOut29_11[1] , \nOut29_11[0] }), .WestIn({\nOut27_11[7] , 
        \nOut27_11[6] , \nOut27_11[5] , \nOut27_11[4] , \nOut27_11[3] , 
        \nOut27_11[2] , \nOut27_11[1] , \nOut27_11[0] }), .Out({\nOut28_11[7] , 
        \nOut28_11[6] , \nOut28_11[5] , \nOut28_11[4] , \nOut28_11[3] , 
        \nOut28_11[2] , \nOut28_11[1] , \nOut28_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_662 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut663[7] , \nScanOut663[6] , 
        \nScanOut663[5] , \nScanOut663[4] , \nScanOut663[3] , \nScanOut663[2] , 
        \nScanOut663[1] , \nScanOut663[0] }), .ScanOut({\nScanOut662[7] , 
        \nScanOut662[6] , \nScanOut662[5] , \nScanOut662[4] , \nScanOut662[3] , 
        \nScanOut662[2] , \nScanOut662[1] , \nScanOut662[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_21[7] , \nOut20_21[6] , \nOut20_21[5] , \nOut20_21[4] , 
        \nOut20_21[3] , \nOut20_21[2] , \nOut20_21[1] , \nOut20_21[0] }), 
        .SouthIn({\nOut20_23[7] , \nOut20_23[6] , \nOut20_23[5] , 
        \nOut20_23[4] , \nOut20_23[3] , \nOut20_23[2] , \nOut20_23[1] , 
        \nOut20_23[0] }), .EastIn({\nOut21_22[7] , \nOut21_22[6] , 
        \nOut21_22[5] , \nOut21_22[4] , \nOut21_22[3] , \nOut21_22[2] , 
        \nOut21_22[1] , \nOut21_22[0] }), .WestIn({\nOut19_22[7] , 
        \nOut19_22[6] , \nOut19_22[5] , \nOut19_22[4] , \nOut19_22[3] , 
        \nOut19_22[2] , \nOut19_22[1] , \nOut19_22[0] }), .Out({\nOut20_22[7] , 
        \nOut20_22[6] , \nOut20_22[5] , \nOut20_22[4] , \nOut20_22[3] , 
        \nOut20_22[2] , \nOut20_22[1] , \nOut20_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_920 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut921[7] , \nScanOut921[6] , 
        \nScanOut921[5] , \nScanOut921[4] , \nScanOut921[3] , \nScanOut921[2] , 
        \nScanOut921[1] , \nScanOut921[0] }), .ScanOut({\nScanOut920[7] , 
        \nScanOut920[6] , \nScanOut920[5] , \nScanOut920[4] , \nScanOut920[3] , 
        \nScanOut920[2] , \nScanOut920[1] , \nScanOut920[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_23[7] , \nOut28_23[6] , \nOut28_23[5] , \nOut28_23[4] , 
        \nOut28_23[3] , \nOut28_23[2] , \nOut28_23[1] , \nOut28_23[0] }), 
        .SouthIn({\nOut28_25[7] , \nOut28_25[6] , \nOut28_25[5] , 
        \nOut28_25[4] , \nOut28_25[3] , \nOut28_25[2] , \nOut28_25[1] , 
        \nOut28_25[0] }), .EastIn({\nOut29_24[7] , \nOut29_24[6] , 
        \nOut29_24[5] , \nOut29_24[4] , \nOut29_24[3] , \nOut29_24[2] , 
        \nOut29_24[1] , \nOut29_24[0] }), .WestIn({\nOut27_24[7] , 
        \nOut27_24[6] , \nOut27_24[5] , \nOut27_24[4] , \nOut27_24[3] , 
        \nOut27_24[2] , \nOut27_24[1] , \nOut27_24[0] }), .Out({\nOut28_24[7] , 
        \nOut28_24[6] , \nOut28_24[5] , \nOut28_24[4] , \nOut28_24[3] , 
        \nOut28_24[2] , \nOut28_24[1] , \nOut28_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_80 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut81[7] , \nScanOut81[6] , 
        \nScanOut81[5] , \nScanOut81[4] , \nScanOut81[3] , \nScanOut81[2] , 
        \nScanOut81[1] , \nScanOut81[0] }), .ScanOut({\nScanOut80[7] , 
        \nScanOut80[6] , \nScanOut80[5] , \nScanOut80[4] , \nScanOut80[3] , 
        \nScanOut80[2] , \nScanOut80[1] , \nScanOut80[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_15[7] , \nOut2_15[6] , \nOut2_15[5] , \nOut2_15[4] , 
        \nOut2_15[3] , \nOut2_15[2] , \nOut2_15[1] , \nOut2_15[0] }), 
        .SouthIn({\nOut2_17[7] , \nOut2_17[6] , \nOut2_17[5] , \nOut2_17[4] , 
        \nOut2_17[3] , \nOut2_17[2] , \nOut2_17[1] , \nOut2_17[0] }), .EastIn(
        {\nOut3_16[7] , \nOut3_16[6] , \nOut3_16[5] , \nOut3_16[4] , 
        \nOut3_16[3] , \nOut3_16[2] , \nOut3_16[1] , \nOut3_16[0] }), .WestIn(
        {\nOut1_16[7] , \nOut1_16[6] , \nOut1_16[5] , \nOut1_16[4] , 
        \nOut1_16[3] , \nOut1_16[2] , \nOut1_16[1] , \nOut1_16[0] }), .Out({
        \nOut2_16[7] , \nOut2_16[6] , \nOut2_16[5] , \nOut2_16[4] , 
        \nOut2_16[3] , \nOut2_16[2] , \nOut2_16[1] , \nOut2_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_92 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut93[7] , \nScanOut93[6] , 
        \nScanOut93[5] , \nScanOut93[4] , \nScanOut93[3] , \nScanOut93[2] , 
        \nScanOut93[1] , \nScanOut93[0] }), .ScanOut({\nScanOut92[7] , 
        \nScanOut92[6] , \nScanOut92[5] , \nScanOut92[4] , \nScanOut92[3] , 
        \nScanOut92[2] , \nScanOut92[1] , \nScanOut92[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_27[7] , \nOut2_27[6] , \nOut2_27[5] , \nOut2_27[4] , 
        \nOut2_27[3] , \nOut2_27[2] , \nOut2_27[1] , \nOut2_27[0] }), 
        .SouthIn({\nOut2_29[7] , \nOut2_29[6] , \nOut2_29[5] , \nOut2_29[4] , 
        \nOut2_29[3] , \nOut2_29[2] , \nOut2_29[1] , \nOut2_29[0] }), .EastIn(
        {\nOut3_28[7] , \nOut3_28[6] , \nOut3_28[5] , \nOut3_28[4] , 
        \nOut3_28[3] , \nOut3_28[2] , \nOut3_28[1] , \nOut3_28[0] }), .WestIn(
        {\nOut1_28[7] , \nOut1_28[6] , \nOut1_28[5] , \nOut1_28[4] , 
        \nOut1_28[3] , \nOut1_28[2] , \nOut1_28[1] , \nOut1_28[0] }), .Out({
        \nOut2_28[7] , \nOut2_28[6] , \nOut2_28[5] , \nOut2_28[4] , 
        \nOut2_28[3] , \nOut2_28[2] , \nOut2_28[1] , \nOut2_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_236 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut237[7] , \nScanOut237[6] , 
        \nScanOut237[5] , \nScanOut237[4] , \nScanOut237[3] , \nScanOut237[2] , 
        \nScanOut237[1] , \nScanOut237[0] }), .ScanOut({\nScanOut236[7] , 
        \nScanOut236[6] , \nScanOut236[5] , \nScanOut236[4] , \nScanOut236[3] , 
        \nScanOut236[2] , \nScanOut236[1] , \nScanOut236[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_11[7] , \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , 
        \nOut7_11[3] , \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }), 
        .SouthIn({\nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }), .EastIn(
        {\nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }), .WestIn(
        {\nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }), .Out({
        \nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_427 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut428[7] , \nScanOut428[6] , 
        \nScanOut428[5] , \nScanOut428[4] , \nScanOut428[3] , \nScanOut428[2] , 
        \nScanOut428[1] , \nScanOut428[0] }), .ScanOut({\nScanOut427[7] , 
        \nScanOut427[6] , \nScanOut427[5] , \nScanOut427[4] , \nScanOut427[3] , 
        \nScanOut427[2] , \nScanOut427[1] , \nScanOut427[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_10[7] , \nOut13_10[6] , \nOut13_10[5] , \nOut13_10[4] , 
        \nOut13_10[3] , \nOut13_10[2] , \nOut13_10[1] , \nOut13_10[0] }), 
        .SouthIn({\nOut13_12[7] , \nOut13_12[6] , \nOut13_12[5] , 
        \nOut13_12[4] , \nOut13_12[3] , \nOut13_12[2] , \nOut13_12[1] , 
        \nOut13_12[0] }), .EastIn({\nOut14_11[7] , \nOut14_11[6] , 
        \nOut14_11[5] , \nOut14_11[4] , \nOut14_11[3] , \nOut14_11[2] , 
        \nOut14_11[1] , \nOut14_11[0] }), .WestIn({\nOut12_11[7] , 
        \nOut12_11[6] , \nOut12_11[5] , \nOut12_11[4] , \nOut12_11[3] , 
        \nOut12_11[2] , \nOut12_11[1] , \nOut12_11[0] }), .Out({\nOut13_11[7] , 
        \nOut13_11[6] , \nOut13_11[5] , \nOut13_11[4] , \nOut13_11[3] , 
        \nOut13_11[2] , \nOut13_11[1] , \nOut13_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_969 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut970[7] , \nScanOut970[6] , 
        \nScanOut970[5] , \nScanOut970[4] , \nScanOut970[3] , \nScanOut970[2] , 
        \nScanOut970[1] , \nScanOut970[0] }), .ScanOut({\nScanOut969[7] , 
        \nScanOut969[6] , \nScanOut969[5] , \nScanOut969[4] , \nScanOut969[3] , 
        \nScanOut969[2] , \nScanOut969[1] , \nScanOut969[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_8[7] , \nOut30_8[6] , \nOut30_8[5] , \nOut30_8[4] , 
        \nOut30_8[3] , \nOut30_8[2] , \nOut30_8[1] , \nOut30_8[0] }), 
        .SouthIn({\nOut30_10[7] , \nOut30_10[6] , \nOut30_10[5] , 
        \nOut30_10[4] , \nOut30_10[3] , \nOut30_10[2] , \nOut30_10[1] , 
        \nOut30_10[0] }), .EastIn({\nOut31_9[7] , \nOut31_9[6] , \nOut31_9[5] , 
        \nOut31_9[4] , \nOut31_9[3] , \nOut31_9[2] , \nOut31_9[1] , 
        \nOut31_9[0] }), .WestIn({\nOut29_9[7] , \nOut29_9[6] , \nOut29_9[5] , 
        \nOut29_9[4] , \nOut29_9[3] , \nOut29_9[2] , \nOut29_9[1] , 
        \nOut29_9[0] }), .Out({\nOut30_9[7] , \nOut30_9[6] , \nOut30_9[5] , 
        \nOut30_9[4] , \nOut30_9[3] , \nOut30_9[2] , \nOut30_9[1] , 
        \nOut30_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_855 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut856[7] , \nScanOut856[6] , 
        \nScanOut856[5] , \nScanOut856[4] , \nScanOut856[3] , \nScanOut856[2] , 
        \nScanOut856[1] , \nScanOut856[0] }), .ScanOut({\nScanOut855[7] , 
        \nScanOut855[6] , \nScanOut855[5] , \nScanOut855[4] , \nScanOut855[3] , 
        \nScanOut855[2] , \nScanOut855[1] , \nScanOut855[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_22[7] , \nOut26_22[6] , \nOut26_22[5] , \nOut26_22[4] , 
        \nOut26_22[3] , \nOut26_22[2] , \nOut26_22[1] , \nOut26_22[0] }), 
        .SouthIn({\nOut26_24[7] , \nOut26_24[6] , \nOut26_24[5] , 
        \nOut26_24[4] , \nOut26_24[3] , \nOut26_24[2] , \nOut26_24[1] , 
        \nOut26_24[0] }), .EastIn({\nOut27_23[7] , \nOut27_23[6] , 
        \nOut27_23[5] , \nOut27_23[4] , \nOut27_23[3] , \nOut27_23[2] , 
        \nOut27_23[1] , \nOut27_23[0] }), .WestIn({\nOut25_23[7] , 
        \nOut25_23[6] , \nOut25_23[5] , \nOut25_23[4] , \nOut25_23[3] , 
        \nOut25_23[2] , \nOut25_23[1] , \nOut25_23[0] }), .Out({\nOut26_23[7] , 
        \nOut26_23[6] , \nOut26_23[5] , \nOut26_23[4] , \nOut26_23[3] , 
        \nOut26_23[2] , \nOut26_23[1] , \nOut26_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_106 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut107[7] , \nScanOut107[6] , 
        \nScanOut107[5] , \nScanOut107[4] , \nScanOut107[3] , \nScanOut107[2] , 
        \nScanOut107[1] , \nScanOut107[0] }), .ScanOut({\nScanOut106[7] , 
        \nScanOut106[6] , \nScanOut106[5] , \nScanOut106[4] , \nScanOut106[3] , 
        \nScanOut106[2] , \nScanOut106[1] , \nScanOut106[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_9[7] , \nOut3_9[6] , \nOut3_9[5] , \nOut3_9[4] , \nOut3_9[3] , 
        \nOut3_9[2] , \nOut3_9[1] , \nOut3_9[0] }), .SouthIn({\nOut3_11[7] , 
        \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , \nOut3_11[3] , 
        \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }), .EastIn({\nOut4_10[7] , 
        \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , \nOut4_10[3] , 
        \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }), .WestIn({\nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), .Out({\nOut3_10[7] , 
        \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , \nOut3_10[3] , 
        \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_717 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut718[7] , \nScanOut718[6] , 
        \nScanOut718[5] , \nScanOut718[4] , \nScanOut718[3] , \nScanOut718[2] , 
        \nScanOut718[1] , \nScanOut718[0] }), .ScanOut({\nScanOut717[7] , 
        \nScanOut717[6] , \nScanOut717[5] , \nScanOut717[4] , \nScanOut717[3] , 
        \nScanOut717[2] , \nScanOut717[1] , \nScanOut717[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_12[7] , \nOut22_12[6] , \nOut22_12[5] , \nOut22_12[4] , 
        \nOut22_12[3] , \nOut22_12[2] , \nOut22_12[1] , \nOut22_12[0] }), 
        .SouthIn({\nOut22_14[7] , \nOut22_14[6] , \nOut22_14[5] , 
        \nOut22_14[4] , \nOut22_14[3] , \nOut22_14[2] , \nOut22_14[1] , 
        \nOut22_14[0] }), .EastIn({\nOut23_13[7] , \nOut23_13[6] , 
        \nOut23_13[5] , \nOut23_13[4] , \nOut23_13[3] , \nOut23_13[2] , 
        \nOut23_13[1] , \nOut23_13[0] }), .WestIn({\nOut21_13[7] , 
        \nOut21_13[6] , \nOut21_13[5] , \nOut21_13[4] , \nOut21_13[3] , 
        \nOut21_13[2] , \nOut21_13[1] , \nOut21_13[0] }), .Out({\nOut22_13[7] , 
        \nOut22_13[6] , \nOut22_13[5] , \nOut22_13[4] , \nOut22_13[3] , 
        \nOut22_13[2] , \nOut22_13[1] , \nOut22_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_121 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut122[7] , \nScanOut122[6] , 
        \nScanOut122[5] , \nScanOut122[4] , \nScanOut122[3] , \nScanOut122[2] , 
        \nScanOut122[1] , \nScanOut122[0] }), .ScanOut({\nScanOut121[7] , 
        \nScanOut121[6] , \nScanOut121[5] , \nScanOut121[4] , \nScanOut121[3] , 
        \nScanOut121[2] , \nScanOut121[1] , \nScanOut121[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_24[7] , \nOut3_24[6] , \nOut3_24[5] , \nOut3_24[4] , 
        \nOut3_24[3] , \nOut3_24[2] , \nOut3_24[1] , \nOut3_24[0] }), 
        .SouthIn({\nOut3_26[7] , \nOut3_26[6] , \nOut3_26[5] , \nOut3_26[4] , 
        \nOut3_26[3] , \nOut3_26[2] , \nOut3_26[1] , \nOut3_26[0] }), .EastIn(
        {\nOut4_25[7] , \nOut4_25[6] , \nOut4_25[5] , \nOut4_25[4] , 
        \nOut4_25[3] , \nOut4_25[2] , \nOut4_25[1] , \nOut4_25[0] }), .WestIn(
        {\nOut2_25[7] , \nOut2_25[6] , \nOut2_25[5] , \nOut2_25[4] , 
        \nOut2_25[3] , \nOut2_25[2] , \nOut2_25[1] , \nOut2_25[0] }), .Out({
        \nOut3_25[7] , \nOut3_25[6] , \nOut3_25[5] , \nOut3_25[4] , 
        \nOut3_25[3] , \nOut3_25[2] , \nOut3_25[1] , \nOut3_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_687 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut688[7] , \nScanOut688[6] , 
        \nScanOut688[5] , \nScanOut688[4] , \nScanOut688[3] , \nScanOut688[2] , 
        \nScanOut688[1] , \nScanOut688[0] }), .ScanOut({\nScanOut687[7] , 
        \nScanOut687[6] , \nScanOut687[5] , \nScanOut687[4] , \nScanOut687[3] , 
        \nScanOut687[2] , \nScanOut687[1] , \nScanOut687[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_14[7] , \nOut21_14[6] , \nOut21_14[5] , \nOut21_14[4] , 
        \nOut21_14[3] , \nOut21_14[2] , \nOut21_14[1] , \nOut21_14[0] }), 
        .SouthIn({\nOut21_16[7] , \nOut21_16[6] , \nOut21_16[5] , 
        \nOut21_16[4] , \nOut21_16[3] , \nOut21_16[2] , \nOut21_16[1] , 
        \nOut21_16[0] }), .EastIn({\nOut22_15[7] , \nOut22_15[6] , 
        \nOut22_15[5] , \nOut22_15[4] , \nOut22_15[3] , \nOut22_15[2] , 
        \nOut22_15[1] , \nOut22_15[0] }), .WestIn({\nOut20_15[7] , 
        \nOut20_15[6] , \nOut20_15[5] , \nOut20_15[4] , \nOut20_15[3] , 
        \nOut20_15[2] , \nOut20_15[1] , \nOut20_15[0] }), .Out({\nOut21_15[7] , 
        \nOut21_15[6] , \nOut21_15[5] , \nOut21_15[4] , \nOut21_15[3] , 
        \nOut21_15[2] , \nOut21_15[1] , \nOut21_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1011 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1012[7] , \nScanOut1012[6] , 
        \nScanOut1012[5] , \nScanOut1012[4] , \nScanOut1012[3] , 
        \nScanOut1012[2] , \nScanOut1012[1] , \nScanOut1012[0] }), .ScanOut({
        \nScanOut1011[7] , \nScanOut1011[6] , \nScanOut1011[5] , 
        \nScanOut1011[4] , \nScanOut1011[3] , \nScanOut1011[2] , 
        \nScanOut1011[1] , \nScanOut1011[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_19[7] , \nOut31_19[6] , \nOut31_19[5] , 
        \nOut31_19[4] , \nOut31_19[3] , \nOut31_19[2] , \nOut31_19[1] , 
        \nOut31_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_211 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut212[7] , \nScanOut212[6] , 
        \nScanOut212[5] , \nScanOut212[4] , \nScanOut212[3] , \nScanOut212[2] , 
        \nScanOut212[1] , \nScanOut212[0] }), .ScanOut({\nScanOut211[7] , 
        \nScanOut211[6] , \nScanOut211[5] , \nScanOut211[4] , \nScanOut211[3] , 
        \nScanOut211[2] , \nScanOut211[1] , \nScanOut211[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_18[7] , \nOut6_18[6] , \nOut6_18[5] , \nOut6_18[4] , 
        \nOut6_18[3] , \nOut6_18[2] , \nOut6_18[1] , \nOut6_18[0] }), 
        .SouthIn({\nOut6_20[7] , \nOut6_20[6] , \nOut6_20[5] , \nOut6_20[4] , 
        \nOut6_20[3] , \nOut6_20[2] , \nOut6_20[1] , \nOut6_20[0] }), .EastIn(
        {\nOut7_19[7] , \nOut7_19[6] , \nOut7_19[5] , \nOut7_19[4] , 
        \nOut7_19[3] , \nOut7_19[2] , \nOut7_19[1] , \nOut7_19[0] }), .WestIn(
        {\nOut5_19[7] , \nOut5_19[6] , \nOut5_19[5] , \nOut5_19[4] , 
        \nOut5_19[3] , \nOut5_19[2] , \nOut5_19[1] , \nOut5_19[0] }), .Out({
        \nOut6_19[7] , \nOut6_19[6] , \nOut6_19[5] , \nOut6_19[4] , 
        \nOut6_19[3] , \nOut6_19[2] , \nOut6_19[1] , \nOut6_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_590 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut591[7] , \nScanOut591[6] , 
        \nScanOut591[5] , \nScanOut591[4] , \nScanOut591[3] , \nScanOut591[2] , 
        \nScanOut591[1] , \nScanOut591[0] }), .ScanOut({\nScanOut590[7] , 
        \nScanOut590[6] , \nScanOut590[5] , \nScanOut590[4] , \nScanOut590[3] , 
        \nScanOut590[2] , \nScanOut590[1] , \nScanOut590[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_13[7] , \nOut18_13[6] , \nOut18_13[5] , \nOut18_13[4] , 
        \nOut18_13[3] , \nOut18_13[2] , \nOut18_13[1] , \nOut18_13[0] }), 
        .SouthIn({\nOut18_15[7] , \nOut18_15[6] , \nOut18_15[5] , 
        \nOut18_15[4] , \nOut18_15[3] , \nOut18_15[2] , \nOut18_15[1] , 
        \nOut18_15[0] }), .EastIn({\nOut19_14[7] , \nOut19_14[6] , 
        \nOut19_14[5] , \nOut19_14[4] , \nOut19_14[3] , \nOut19_14[2] , 
        \nOut19_14[1] , \nOut19_14[0] }), .WestIn({\nOut17_14[7] , 
        \nOut17_14[6] , \nOut17_14[5] , \nOut17_14[4] , \nOut17_14[3] , 
        \nOut17_14[2] , \nOut17_14[1] , \nOut17_14[0] }), .Out({\nOut18_14[7] , 
        \nOut18_14[6] , \nOut18_14[5] , \nOut18_14[4] , \nOut18_14[3] , 
        \nOut18_14[2] , \nOut18_14[1] , \nOut18_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_730 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut731[7] , \nScanOut731[6] , 
        \nScanOut731[5] , \nScanOut731[4] , \nScanOut731[3] , \nScanOut731[2] , 
        \nScanOut731[1] , \nScanOut731[0] }), .ScanOut({\nScanOut730[7] , 
        \nScanOut730[6] , \nScanOut730[5] , \nScanOut730[4] , \nScanOut730[3] , 
        \nScanOut730[2] , \nScanOut730[1] , \nScanOut730[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_25[7] , \nOut22_25[6] , \nOut22_25[5] , \nOut22_25[4] , 
        \nOut22_25[3] , \nOut22_25[2] , \nOut22_25[1] , \nOut22_25[0] }), 
        .SouthIn({\nOut22_27[7] , \nOut22_27[6] , \nOut22_27[5] , 
        \nOut22_27[4] , \nOut22_27[3] , \nOut22_27[2] , \nOut22_27[1] , 
        \nOut22_27[0] }), .EastIn({\nOut23_26[7] , \nOut23_26[6] , 
        \nOut23_26[5] , \nOut23_26[4] , \nOut23_26[3] , \nOut23_26[2] , 
        \nOut23_26[1] , \nOut23_26[0] }), .WestIn({\nOut21_26[7] , 
        \nOut21_26[6] , \nOut21_26[5] , \nOut21_26[4] , \nOut21_26[3] , 
        \nOut21_26[2] , \nOut21_26[1] , \nOut21_26[0] }), .Out({\nOut22_26[7] , 
        \nOut22_26[6] , \nOut22_26[5] , \nOut22_26[4] , \nOut22_26[3] , 
        \nOut22_26[2] , \nOut22_26[1] , \nOut22_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_224 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut225[7] , \nScanOut225[6] , 
        \nScanOut225[5] , \nScanOut225[4] , \nScanOut225[3] , \nScanOut225[2] , 
        \nScanOut225[1] , \nScanOut225[0] }), .ScanOut({\nScanOut224[7] , 
        \nScanOut224[6] , \nScanOut224[5] , \nScanOut224[4] , \nScanOut224[3] , 
        \nScanOut224[2] , \nScanOut224[1] , \nScanOut224[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut7_0[7] , \nOut7_0[6] , 
        \nOut7_0[5] , \nOut7_0[4] , \nOut7_0[3] , \nOut7_0[2] , \nOut7_0[1] , 
        \nOut7_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_381 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut382[7] , \nScanOut382[6] , 
        \nScanOut382[5] , \nScanOut382[4] , \nScanOut382[3] , \nScanOut382[2] , 
        \nScanOut382[1] , \nScanOut382[0] }), .ScanOut({\nScanOut381[7] , 
        \nScanOut381[6] , \nScanOut381[5] , \nScanOut381[4] , \nScanOut381[3] , 
        \nScanOut381[2] , \nScanOut381[1] , \nScanOut381[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_28[7] , \nOut11_28[6] , \nOut11_28[5] , \nOut11_28[4] , 
        \nOut11_28[3] , \nOut11_28[2] , \nOut11_28[1] , \nOut11_28[0] }), 
        .SouthIn({\nOut11_30[7] , \nOut11_30[6] , \nOut11_30[5] , 
        \nOut11_30[4] , \nOut11_30[3] , \nOut11_30[2] , \nOut11_30[1] , 
        \nOut11_30[0] }), .EastIn({\nOut12_29[7] , \nOut12_29[6] , 
        \nOut12_29[5] , \nOut12_29[4] , \nOut12_29[3] , \nOut12_29[2] , 
        \nOut12_29[1] , \nOut12_29[0] }), .WestIn({\nOut10_29[7] , 
        \nOut10_29[6] , \nOut10_29[5] , \nOut10_29[4] , \nOut10_29[3] , 
        \nOut10_29[2] , \nOut10_29[1] , \nOut10_29[0] }), .Out({\nOut11_29[7] , 
        \nOut11_29[6] , \nOut11_29[5] , \nOut11_29[4] , \nOut11_29[3] , 
        \nOut11_29[2] , \nOut11_29[1] , \nOut11_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_400 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut401[7] , \nScanOut401[6] , 
        \nScanOut401[5] , \nScanOut401[4] , \nScanOut401[3] , \nScanOut401[2] , 
        \nScanOut401[1] , \nScanOut401[0] }), .ScanOut({\nScanOut400[7] , 
        \nScanOut400[6] , \nScanOut400[5] , \nScanOut400[4] , \nScanOut400[3] , 
        \nScanOut400[2] , \nScanOut400[1] , \nScanOut400[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_15[7] , \nOut12_15[6] , \nOut12_15[5] , \nOut12_15[4] , 
        \nOut12_15[3] , \nOut12_15[2] , \nOut12_15[1] , \nOut12_15[0] }), 
        .SouthIn({\nOut12_17[7] , \nOut12_17[6] , \nOut12_17[5] , 
        \nOut12_17[4] , \nOut12_17[3] , \nOut12_17[2] , \nOut12_17[1] , 
        \nOut12_17[0] }), .EastIn({\nOut13_16[7] , \nOut13_16[6] , 
        \nOut13_16[5] , \nOut13_16[4] , \nOut13_16[3] , \nOut13_16[2] , 
        \nOut13_16[1] , \nOut13_16[0] }), .WestIn({\nOut11_16[7] , 
        \nOut11_16[6] , \nOut11_16[5] , \nOut11_16[4] , \nOut11_16[3] , 
        \nOut11_16[2] , \nOut11_16[1] , \nOut11_16[0] }), .Out({\nOut12_16[7] , 
        \nOut12_16[6] , \nOut12_16[5] , \nOut12_16[4] , \nOut12_16[3] , 
        \nOut12_16[2] , \nOut12_16[1] , \nOut12_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_847 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut848[7] , \nScanOut848[6] , 
        \nScanOut848[5] , \nScanOut848[4] , \nScanOut848[3] , \nScanOut848[2] , 
        \nScanOut848[1] , \nScanOut848[0] }), .ScanOut({\nScanOut847[7] , 
        \nScanOut847[6] , \nScanOut847[5] , \nScanOut847[4] , \nScanOut847[3] , 
        \nScanOut847[2] , \nScanOut847[1] , \nScanOut847[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_14[7] , \nOut26_14[6] , \nOut26_14[5] , \nOut26_14[4] , 
        \nOut26_14[3] , \nOut26_14[2] , \nOut26_14[1] , \nOut26_14[0] }), 
        .SouthIn({\nOut26_16[7] , \nOut26_16[6] , \nOut26_16[5] , 
        \nOut26_16[4] , \nOut26_16[3] , \nOut26_16[2] , \nOut26_16[1] , 
        \nOut26_16[0] }), .EastIn({\nOut27_15[7] , \nOut27_15[6] , 
        \nOut27_15[5] , \nOut27_15[4] , \nOut27_15[3] , \nOut27_15[2] , 
        \nOut27_15[1] , \nOut27_15[0] }), .WestIn({\nOut25_15[7] , 
        \nOut25_15[6] , \nOut25_15[5] , \nOut25_15[4] , \nOut25_15[3] , 
        \nOut25_15[2] , \nOut25_15[1] , \nOut25_15[0] }), .Out({\nOut26_15[7] , 
        \nOut26_15[6] , \nOut26_15[5] , \nOut26_15[4] , \nOut26_15[3] , 
        \nOut26_15[2] , \nOut26_15[1] , \nOut26_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_872 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut873[7] , \nScanOut873[6] , 
        \nScanOut873[5] , \nScanOut873[4] , \nScanOut873[3] , \nScanOut873[2] , 
        \nScanOut873[1] , \nScanOut873[0] }), .ScanOut({\nScanOut872[7] , 
        \nScanOut872[6] , \nScanOut872[5] , \nScanOut872[4] , \nScanOut872[3] , 
        \nScanOut872[2] , \nScanOut872[1] , \nScanOut872[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_7[7] , \nOut27_7[6] , \nOut27_7[5] , \nOut27_7[4] , 
        \nOut27_7[3] , \nOut27_7[2] , \nOut27_7[1] , \nOut27_7[0] }), 
        .SouthIn({\nOut27_9[7] , \nOut27_9[6] , \nOut27_9[5] , \nOut27_9[4] , 
        \nOut27_9[3] , \nOut27_9[2] , \nOut27_9[1] , \nOut27_9[0] }), .EastIn(
        {\nOut28_8[7] , \nOut28_8[6] , \nOut28_8[5] , \nOut28_8[4] , 
        \nOut28_8[3] , \nOut28_8[2] , \nOut28_8[1] , \nOut28_8[0] }), .WestIn(
        {\nOut26_8[7] , \nOut26_8[6] , \nOut26_8[5] , \nOut26_8[4] , 
        \nOut26_8[3] , \nOut26_8[2] , \nOut26_8[1] , \nOut26_8[0] }), .Out({
        \nOut27_8[7] , \nOut27_8[6] , \nOut27_8[5] , \nOut27_8[4] , 
        \nOut27_8[3] , \nOut27_8[2] , \nOut27_8[1] , \nOut27_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_435 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut436[7] , \nScanOut436[6] , 
        \nScanOut436[5] , \nScanOut436[4] , \nScanOut436[3] , \nScanOut436[2] , 
        \nScanOut436[1] , \nScanOut436[0] }), .ScanOut({\nScanOut435[7] , 
        \nScanOut435[6] , \nScanOut435[5] , \nScanOut435[4] , \nScanOut435[3] , 
        \nScanOut435[2] , \nScanOut435[1] , \nScanOut435[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_18[7] , \nOut13_18[6] , \nOut13_18[5] , \nOut13_18[4] , 
        \nOut13_18[3] , \nOut13_18[2] , \nOut13_18[1] , \nOut13_18[0] }), 
        .SouthIn({\nOut13_20[7] , \nOut13_20[6] , \nOut13_20[5] , 
        \nOut13_20[4] , \nOut13_20[3] , \nOut13_20[2] , \nOut13_20[1] , 
        \nOut13_20[0] }), .EastIn({\nOut14_19[7] , \nOut14_19[6] , 
        \nOut14_19[5] , \nOut14_19[4] , \nOut14_19[3] , \nOut14_19[2] , 
        \nOut14_19[1] , \nOut14_19[0] }), .WestIn({\nOut12_19[7] , 
        \nOut12_19[6] , \nOut12_19[5] , \nOut12_19[4] , \nOut12_19[3] , 
        \nOut12_19[2] , \nOut12_19[1] , \nOut12_19[0] }), .Out({\nOut13_19[7] , 
        \nOut13_19[6] , \nOut13_19[5] , \nOut13_19[4] , \nOut13_19[3] , 
        \nOut13_19[2] , \nOut13_19[1] , \nOut13_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_114 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut115[7] , \nScanOut115[6] , 
        \nScanOut115[5] , \nScanOut115[4] , \nScanOut115[3] , \nScanOut115[2] , 
        \nScanOut115[1] , \nScanOut115[0] }), .ScanOut({\nScanOut114[7] , 
        \nScanOut114[6] , \nScanOut114[5] , \nScanOut114[4] , \nScanOut114[3] , 
        \nScanOut114[2] , \nScanOut114[1] , \nScanOut114[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_17[7] , \nOut3_17[6] , \nOut3_17[5] , \nOut3_17[4] , 
        \nOut3_17[3] , \nOut3_17[2] , \nOut3_17[1] , \nOut3_17[0] }), 
        .SouthIn({\nOut3_19[7] , \nOut3_19[6] , \nOut3_19[5] , \nOut3_19[4] , 
        \nOut3_19[3] , \nOut3_19[2] , \nOut3_19[1] , \nOut3_19[0] }), .EastIn(
        {\nOut4_18[7] , \nOut4_18[6] , \nOut4_18[5] , \nOut4_18[4] , 
        \nOut4_18[3] , \nOut4_18[2] , \nOut4_18[1] , \nOut4_18[0] }), .WestIn(
        {\nOut2_18[7] , \nOut2_18[6] , \nOut2_18[5] , \nOut2_18[4] , 
        \nOut2_18[3] , \nOut2_18[2] , \nOut2_18[1] , \nOut2_18[0] }), .Out({
        \nOut3_18[7] , \nOut3_18[6] , \nOut3_18[5] , \nOut3_18[4] , 
        \nOut3_18[3] , \nOut3_18[2] , \nOut3_18[1] , \nOut3_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_695 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut696[7] , \nScanOut696[6] , 
        \nScanOut696[5] , \nScanOut696[4] , \nScanOut696[3] , \nScanOut696[2] , 
        \nScanOut696[1] , \nScanOut696[0] }), .ScanOut({\nScanOut695[7] , 
        \nScanOut695[6] , \nScanOut695[5] , \nScanOut695[4] , \nScanOut695[3] , 
        \nScanOut695[2] , \nScanOut695[1] , \nScanOut695[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_22[7] , \nOut21_22[6] , \nOut21_22[5] , \nOut21_22[4] , 
        \nOut21_22[3] , \nOut21_22[2] , \nOut21_22[1] , \nOut21_22[0] }), 
        .SouthIn({\nOut21_24[7] , \nOut21_24[6] , \nOut21_24[5] , 
        \nOut21_24[4] , \nOut21_24[3] , \nOut21_24[2] , \nOut21_24[1] , 
        \nOut21_24[0] }), .EastIn({\nOut22_23[7] , \nOut22_23[6] , 
        \nOut22_23[5] , \nOut22_23[4] , \nOut22_23[3] , \nOut22_23[2] , 
        \nOut22_23[1] , \nOut22_23[0] }), .WestIn({\nOut20_23[7] , 
        \nOut20_23[6] , \nOut20_23[5] , \nOut20_23[4] , \nOut20_23[3] , 
        \nOut20_23[2] , \nOut20_23[1] , \nOut20_23[0] }), .Out({\nOut21_23[7] , 
        \nOut21_23[6] , \nOut21_23[5] , \nOut21_23[4] , \nOut21_23[3] , 
        \nOut21_23[2] , \nOut21_23[1] , \nOut21_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1003 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1004[7] , \nScanOut1004[6] , 
        \nScanOut1004[5] , \nScanOut1004[4] , \nScanOut1004[3] , 
        \nScanOut1004[2] , \nScanOut1004[1] , \nScanOut1004[0] }), .ScanOut({
        \nScanOut1003[7] , \nScanOut1003[6] , \nScanOut1003[5] , 
        \nScanOut1003[4] , \nScanOut1003[3] , \nScanOut1003[2] , 
        \nScanOut1003[1] , \nScanOut1003[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_11[7] , \nOut31_11[6] , \nOut31_11[5] , 
        \nOut31_11[4] , \nOut31_11[3] , \nOut31_11[2] , \nOut31_11[1] , 
        \nOut31_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_705 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut706[7] , \nScanOut706[6] , 
        \nScanOut706[5] , \nScanOut706[4] , \nScanOut706[3] , \nScanOut706[2] , 
        \nScanOut706[1] , \nScanOut706[0] }), .ScanOut({\nScanOut705[7] , 
        \nScanOut705[6] , \nScanOut705[5] , \nScanOut705[4] , \nScanOut705[3] , 
        \nScanOut705[2] , \nScanOut705[1] , \nScanOut705[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_0[7] , \nOut22_0[6] , \nOut22_0[5] , \nOut22_0[4] , 
        \nOut22_0[3] , \nOut22_0[2] , \nOut22_0[1] , \nOut22_0[0] }), 
        .SouthIn({\nOut22_2[7] , \nOut22_2[6] , \nOut22_2[5] , \nOut22_2[4] , 
        \nOut22_2[3] , \nOut22_2[2] , \nOut22_2[1] , \nOut22_2[0] }), .EastIn(
        {\nOut23_1[7] , \nOut23_1[6] , \nOut23_1[5] , \nOut23_1[4] , 
        \nOut23_1[3] , \nOut23_1[2] , \nOut23_1[1] , \nOut23_1[0] }), .WestIn(
        {\nOut21_1[7] , \nOut21_1[6] , \nOut21_1[5] , \nOut21_1[4] , 
        \nOut21_1[3] , \nOut21_1[2] , \nOut21_1[1] , \nOut21_1[0] }), .Out({
        \nOut22_1[7] , \nOut22_1[6] , \nOut22_1[5] , \nOut22_1[4] , 
        \nOut22_1[3] , \nOut22_1[2] , \nOut22_1[1] , \nOut22_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1[7] , \nScanOut1[6] , 
        \nScanOut1[5] , \nScanOut1[4] , \nScanOut1[3] , \nScanOut1[2] , 
        \nScanOut1[1] , \nScanOut1[0] }), .ScanOut({\nScanOut0[7] , 
        \nScanOut0[6] , \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , 
        \nScanOut0[2] , \nScanOut0[1] , \nScanOut0[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_2 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut3[7] , \nScanOut3[6] , 
        \nScanOut3[5] , \nScanOut3[4] , \nScanOut3[3] , \nScanOut3[2] , 
        \nScanOut3[1] , \nScanOut3[0] }), .ScanOut({\nScanOut2[7] , 
        \nScanOut2[6] , \nScanOut2[5] , \nScanOut2[4] , \nScanOut2[3] , 
        \nScanOut2[2] , \nScanOut2[1] , \nScanOut2[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_2[7] , \nOut0_2[6] , 
        \nOut0_2[5] , \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , 
        \nOut0_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_3 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut4[7] , \nScanOut4[6] , 
        \nScanOut4[5] , \nScanOut4[4] , \nScanOut4[3] , \nScanOut4[2] , 
        \nScanOut4[1] , \nScanOut4[0] }), .ScanOut({\nScanOut3[7] , 
        \nScanOut3[6] , \nScanOut3[5] , \nScanOut3[4] , \nScanOut3[3] , 
        \nScanOut3[2] , \nScanOut3[1] , \nScanOut3[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_3[7] , \nOut0_3[6] , 
        \nOut0_3[5] , \nOut0_3[4] , \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , 
        \nOut0_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_4 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut5[7] , \nScanOut5[6] , 
        \nScanOut5[5] , \nScanOut5[4] , \nScanOut5[3] , \nScanOut5[2] , 
        \nScanOut5[1] , \nScanOut5[0] }), .ScanOut({\nScanOut4[7] , 
        \nScanOut4[6] , \nScanOut4[5] , \nScanOut4[4] , \nScanOut4[3] , 
        \nScanOut4[2] , \nScanOut4[1] , \nScanOut4[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_4[7] , \nOut0_4[6] , 
        \nOut0_4[5] , \nOut0_4[4] , \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , 
        \nOut0_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_133 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut134[7] , \nScanOut134[6] , 
        \nScanOut134[5] , \nScanOut134[4] , \nScanOut134[3] , \nScanOut134[2] , 
        \nScanOut134[1] , \nScanOut134[0] }), .ScanOut({\nScanOut133[7] , 
        \nScanOut133[6] , \nScanOut133[5] , \nScanOut133[4] , \nScanOut133[3] , 
        \nScanOut133[2] , \nScanOut133[1] , \nScanOut133[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_4[7] , \nOut4_4[6] , \nOut4_4[5] , \nOut4_4[4] , \nOut4_4[3] , 
        \nOut4_4[2] , \nOut4_4[1] , \nOut4_4[0] }), .SouthIn({\nOut4_6[7] , 
        \nOut4_6[6] , \nOut4_6[5] , \nOut4_6[4] , \nOut4_6[3] , \nOut4_6[2] , 
        \nOut4_6[1] , \nOut4_6[0] }), .EastIn({\nOut5_5[7] , \nOut5_5[6] , 
        \nOut5_5[5] , \nOut5_5[4] , \nOut5_5[3] , \nOut5_5[2] , \nOut5_5[1] , 
        \nOut5_5[0] }), .WestIn({\nOut3_5[7] , \nOut3_5[6] , \nOut3_5[5] , 
        \nOut3_5[4] , \nOut3_5[3] , \nOut3_5[2] , \nOut3_5[1] , \nOut3_5[0] }), 
        .Out({\nOut4_5[7] , \nOut4_5[6] , \nOut4_5[5] , \nOut4_5[4] , 
        \nOut4_5[3] , \nOut4_5[2] , \nOut4_5[1] , \nOut4_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_722 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut723[7] , \nScanOut723[6] , 
        \nScanOut723[5] , \nScanOut723[4] , \nScanOut723[3] , \nScanOut723[2] , 
        \nScanOut723[1] , \nScanOut723[0] }), .ScanOut({\nScanOut722[7] , 
        \nScanOut722[6] , \nScanOut722[5] , \nScanOut722[4] , \nScanOut722[3] , 
        \nScanOut722[2] , \nScanOut722[1] , \nScanOut722[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_17[7] , \nOut22_17[6] , \nOut22_17[5] , \nOut22_17[4] , 
        \nOut22_17[3] , \nOut22_17[2] , \nOut22_17[1] , \nOut22_17[0] }), 
        .SouthIn({\nOut22_19[7] , \nOut22_19[6] , \nOut22_19[5] , 
        \nOut22_19[4] , \nOut22_19[3] , \nOut22_19[2] , \nOut22_19[1] , 
        \nOut22_19[0] }), .EastIn({\nOut23_18[7] , \nOut23_18[6] , 
        \nOut23_18[5] , \nOut23_18[4] , \nOut23_18[3] , \nOut23_18[2] , 
        \nOut23_18[1] , \nOut23_18[0] }), .WestIn({\nOut21_18[7] , 
        \nOut21_18[6] , \nOut21_18[5] , \nOut21_18[4] , \nOut21_18[3] , 
        \nOut21_18[2] , \nOut21_18[1] , \nOut21_18[0] }), .Out({\nOut22_18[7] , 
        \nOut22_18[6] , \nOut22_18[5] , \nOut22_18[4] , \nOut22_18[3] , 
        \nOut22_18[2] , \nOut22_18[1] , \nOut22_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_203 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut204[7] , \nScanOut204[6] , 
        \nScanOut204[5] , \nScanOut204[4] , \nScanOut204[3] , \nScanOut204[2] , 
        \nScanOut204[1] , \nScanOut204[0] }), .ScanOut({\nScanOut203[7] , 
        \nScanOut203[6] , \nScanOut203[5] , \nScanOut203[4] , \nScanOut203[3] , 
        \nScanOut203[2] , \nScanOut203[1] , \nScanOut203[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_10[7] , \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , 
        \nOut6_10[3] , \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }), 
        .SouthIn({\nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }), .EastIn(
        {\nOut7_11[7] , \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , 
        \nOut7_11[3] , \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }), .WestIn(
        {\nOut5_11[7] , \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , 
        \nOut5_11[3] , \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }), .Out({
        \nOut6_11[7] , \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , 
        \nOut6_11[3] , \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_393 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut394[7] , \nScanOut394[6] , 
        \nScanOut394[5] , \nScanOut394[4] , \nScanOut394[3] , \nScanOut394[2] , 
        \nScanOut394[1] , \nScanOut394[0] }), .ScanOut({\nScanOut393[7] , 
        \nScanOut393[6] , \nScanOut393[5] , \nScanOut393[4] , \nScanOut393[3] , 
        \nScanOut393[2] , \nScanOut393[1] , \nScanOut393[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }), 
        .SouthIn({\nOut12_10[7] , \nOut12_10[6] , \nOut12_10[5] , 
        \nOut12_10[4] , \nOut12_10[3] , \nOut12_10[2] , \nOut12_10[1] , 
        \nOut12_10[0] }), .EastIn({\nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , 
        \nOut13_9[4] , \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , 
        \nOut13_9[0] }), .WestIn({\nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , 
        \nOut11_9[4] , \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , 
        \nOut11_9[0] }), .Out({\nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , 
        \nOut12_9[4] , \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , 
        \nOut12_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_412 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut413[7] , \nScanOut413[6] , 
        \nScanOut413[5] , \nScanOut413[4] , \nScanOut413[3] , \nScanOut413[2] , 
        \nScanOut413[1] , \nScanOut413[0] }), .ScanOut({\nScanOut412[7] , 
        \nScanOut412[6] , \nScanOut412[5] , \nScanOut412[4] , \nScanOut412[3] , 
        \nScanOut412[2] , \nScanOut412[1] , \nScanOut412[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_27[7] , \nOut12_27[6] , \nOut12_27[5] , \nOut12_27[4] , 
        \nOut12_27[3] , \nOut12_27[2] , \nOut12_27[1] , \nOut12_27[0] }), 
        .SouthIn({\nOut12_29[7] , \nOut12_29[6] , \nOut12_29[5] , 
        \nOut12_29[4] , \nOut12_29[3] , \nOut12_29[2] , \nOut12_29[1] , 
        \nOut12_29[0] }), .EastIn({\nOut13_28[7] , \nOut13_28[6] , 
        \nOut13_28[5] , \nOut13_28[4] , \nOut13_28[3] , \nOut13_28[2] , 
        \nOut13_28[1] , \nOut13_28[0] }), .WestIn({\nOut11_28[7] , 
        \nOut11_28[6] , \nOut11_28[5] , \nOut11_28[4] , \nOut11_28[3] , 
        \nOut11_28[2] , \nOut11_28[1] , \nOut11_28[0] }), .Out({\nOut12_28[7] , 
        \nOut12_28[6] , \nOut12_28[5] , \nOut12_28[4] , \nOut12_28[3] , 
        \nOut12_28[2] , \nOut12_28[1] , \nOut12_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_860 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut861[7] , \nScanOut861[6] , 
        \nScanOut861[5] , \nScanOut861[4] , \nScanOut861[3] , \nScanOut861[2] , 
        \nScanOut861[1] , \nScanOut861[0] }), .ScanOut({\nScanOut860[7] , 
        \nScanOut860[6] , \nScanOut860[5] , \nScanOut860[4] , \nScanOut860[3] , 
        \nScanOut860[2] , \nScanOut860[1] , \nScanOut860[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_27[7] , \nOut26_27[6] , \nOut26_27[5] , \nOut26_27[4] , 
        \nOut26_27[3] , \nOut26_27[2] , \nOut26_27[1] , \nOut26_27[0] }), 
        .SouthIn({\nOut26_29[7] , \nOut26_29[6] , \nOut26_29[5] , 
        \nOut26_29[4] , \nOut26_29[3] , \nOut26_29[2] , \nOut26_29[1] , 
        \nOut26_29[0] }), .EastIn({\nOut27_28[7] , \nOut27_28[6] , 
        \nOut27_28[5] , \nOut27_28[4] , \nOut27_28[3] , \nOut27_28[2] , 
        \nOut27_28[1] , \nOut27_28[0] }), .WestIn({\nOut25_28[7] , 
        \nOut25_28[6] , \nOut25_28[5] , \nOut25_28[4] , \nOut25_28[3] , 
        \nOut25_28[2] , \nOut25_28[1] , \nOut25_28[0] }), .Out({\nOut26_28[7] , 
        \nOut26_28[6] , \nOut26_28[5] , \nOut26_28[4] , \nOut26_28[3] , 
        \nOut26_28[2] , \nOut26_28[1] , \nOut26_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_582 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut583[7] , \nScanOut583[6] , 
        \nScanOut583[5] , \nScanOut583[4] , \nScanOut583[3] , \nScanOut583[2] , 
        \nScanOut583[1] , \nScanOut583[0] }), .ScanOut({\nScanOut582[7] , 
        \nScanOut582[6] , \nScanOut582[5] , \nScanOut582[4] , \nScanOut582[3] , 
        \nScanOut582[2] , \nScanOut582[1] , \nScanOut582[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_5[7] , \nOut18_5[6] , \nOut18_5[5] , \nOut18_5[4] , 
        \nOut18_5[3] , \nOut18_5[2] , \nOut18_5[1] , \nOut18_5[0] }), 
        .SouthIn({\nOut18_7[7] , \nOut18_7[6] , \nOut18_7[5] , \nOut18_7[4] , 
        \nOut18_7[3] , \nOut18_7[2] , \nOut18_7[1] , \nOut18_7[0] }), .EastIn(
        {\nOut19_6[7] , \nOut19_6[6] , \nOut19_6[5] , \nOut19_6[4] , 
        \nOut19_6[3] , \nOut19_6[2] , \nOut19_6[1] , \nOut19_6[0] }), .WestIn(
        {\nOut17_6[7] , \nOut17_6[6] , \nOut17_6[5] , \nOut17_6[4] , 
        \nOut17_6[3] , \nOut17_6[2] , \nOut17_6[1] , \nOut17_6[0] }), .Out({
        \nOut18_6[7] , \nOut18_6[6] , \nOut18_6[5] , \nOut18_6[4] , 
        \nOut18_6[3] , \nOut18_6[2] , \nOut18_6[1] , \nOut18_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_288 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut289[7] , \nScanOut289[6] , 
        \nScanOut289[5] , \nScanOut289[4] , \nScanOut289[3] , \nScanOut289[2] , 
        \nScanOut289[1] , \nScanOut289[0] }), .ScanOut({\nScanOut288[7] , 
        \nScanOut288[6] , \nScanOut288[5] , \nScanOut288[4] , \nScanOut288[3] , 
        \nScanOut288[2] , \nScanOut288[1] , \nScanOut288[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut9_0[7] , \nOut9_0[6] , 
        \nOut9_0[5] , \nOut9_0[4] , \nOut9_0[3] , \nOut9_0[2] , \nOut9_0[1] , 
        \nOut9_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_318 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut319[7] , \nScanOut319[6] , 
        \nScanOut319[5] , \nScanOut319[4] , \nScanOut319[3] , \nScanOut319[2] , 
        \nScanOut319[1] , \nScanOut319[0] }), .ScanOut({\nScanOut318[7] , 
        \nScanOut318[6] , \nScanOut318[5] , \nScanOut318[4] , \nScanOut318[3] , 
        \nScanOut318[2] , \nScanOut318[1] , \nScanOut318[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_29[7] , \nOut9_29[6] , \nOut9_29[5] , \nOut9_29[4] , 
        \nOut9_29[3] , \nOut9_29[2] , \nOut9_29[1] , \nOut9_29[0] }), 
        .SouthIn({\nOut9_31[7] , \nOut9_31[6] , \nOut9_31[5] , \nOut9_31[4] , 
        \nOut9_31[3] , \nOut9_31[2] , \nOut9_31[1] , \nOut9_31[0] }), .EastIn(
        {\nOut10_30[7] , \nOut10_30[6] , \nOut10_30[5] , \nOut10_30[4] , 
        \nOut10_30[3] , \nOut10_30[2] , \nOut10_30[1] , \nOut10_30[0] }), 
        .WestIn({\nOut8_30[7] , \nOut8_30[6] , \nOut8_30[5] , \nOut8_30[4] , 
        \nOut8_30[3] , \nOut8_30[2] , \nOut8_30[1] , \nOut8_30[0] }), .Out({
        \nOut9_30[7] , \nOut9_30[6] , \nOut9_30[5] , \nOut9_30[4] , 
        \nOut9_30[3] , \nOut9_30[2] , \nOut9_30[1] , \nOut9_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_499 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut500[7] , \nScanOut500[6] , 
        \nScanOut500[5] , \nScanOut500[4] , \nScanOut500[3] , \nScanOut500[2] , 
        \nScanOut500[1] , \nScanOut500[0] }), .ScanOut({\nScanOut499[7] , 
        \nScanOut499[6] , \nScanOut499[5] , \nScanOut499[4] , \nScanOut499[3] , 
        \nScanOut499[2] , \nScanOut499[1] , \nScanOut499[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_18[7] , \nOut15_18[6] , \nOut15_18[5] , \nOut15_18[4] , 
        \nOut15_18[3] , \nOut15_18[2] , \nOut15_18[1] , \nOut15_18[0] }), 
        .SouthIn({\nOut15_20[7] , \nOut15_20[6] , \nOut15_20[5] , 
        \nOut15_20[4] , \nOut15_20[3] , \nOut15_20[2] , \nOut15_20[1] , 
        \nOut15_20[0] }), .EastIn({\nOut16_19[7] , \nOut16_19[6] , 
        \nOut16_19[5] , \nOut16_19[4] , \nOut16_19[3] , \nOut16_19[2] , 
        \nOut16_19[1] , \nOut16_19[0] }), .WestIn({\nOut14_19[7] , 
        \nOut14_19[6] , \nOut14_19[5] , \nOut14_19[4] , \nOut14_19[3] , 
        \nOut14_19[2] , \nOut14_19[1] , \nOut14_19[0] }), .Out({\nOut15_19[7] , 
        \nOut15_19[6] , \nOut15_19[5] , \nOut15_19[4] , \nOut15_19[3] , 
        \nOut15_19[2] , \nOut15_19[1] , \nOut15_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_639 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut640[7] , \nScanOut640[6] , 
        \nScanOut640[5] , \nScanOut640[4] , \nScanOut640[3] , \nScanOut640[2] , 
        \nScanOut640[1] , \nScanOut640[0] }), .ScanOut({\nScanOut639[7] , 
        \nScanOut639[6] , \nScanOut639[5] , \nScanOut639[4] , \nScanOut639[3] , 
        \nScanOut639[2] , \nScanOut639[1] , \nScanOut639[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut19_31[7] , \nOut19_31[6] , 
        \nOut19_31[5] , \nOut19_31[4] , \nOut19_31[3] , \nOut19_31[2] , 
        \nOut19_31[1] , \nOut19_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_509 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut510[7] , \nScanOut510[6] , 
        \nScanOut510[5] , \nScanOut510[4] , \nScanOut510[3] , \nScanOut510[2] , 
        \nScanOut510[1] , \nScanOut510[0] }), .ScanOut({\nScanOut509[7] , 
        \nScanOut509[6] , \nScanOut509[5] , \nScanOut509[4] , \nScanOut509[3] , 
        \nScanOut509[2] , \nScanOut509[1] , \nScanOut509[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_28[7] , \nOut15_28[6] , \nOut15_28[5] , \nOut15_28[4] , 
        \nOut15_28[3] , \nOut15_28[2] , \nOut15_28[1] , \nOut15_28[0] }), 
        .SouthIn({\nOut15_30[7] , \nOut15_30[6] , \nOut15_30[5] , 
        \nOut15_30[4] , \nOut15_30[3] , \nOut15_30[2] , \nOut15_30[1] , 
        \nOut15_30[0] }), .EastIn({\nOut16_29[7] , \nOut16_29[6] , 
        \nOut16_29[5] , \nOut16_29[4] , \nOut16_29[3] , \nOut16_29[2] , 
        \nOut16_29[1] , \nOut16_29[0] }), .WestIn({\nOut14_29[7] , 
        \nOut14_29[6] , \nOut14_29[5] , \nOut14_29[4] , \nOut14_29[3] , 
        \nOut14_29[2] , \nOut14_29[1] , \nOut14_29[0] }), .Out({\nOut15_29[7] , 
        \nOut15_29[6] , \nOut15_29[5] , \nOut15_29[4] , \nOut15_29[3] , 
        \nOut15_29[2] , \nOut15_29[1] , \nOut15_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_10 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut11[7] , \nScanOut11[6] , 
        \nScanOut11[5] , \nScanOut11[4] , \nScanOut11[3] , \nScanOut11[2] , 
        \nScanOut11[1] , \nScanOut11[0] }), .ScanOut({\nScanOut10[7] , 
        \nScanOut10[6] , \nScanOut10[5] , \nScanOut10[4] , \nScanOut10[3] , 
        \nScanOut10[2] , \nScanOut10[1] , \nScanOut10[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_10[7] , \nOut0_10[6] , 
        \nOut0_10[5] , \nOut0_10[4] , \nOut0_10[3] , \nOut0_10[2] , 
        \nOut0_10[1] , \nOut0_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_37 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut38[7] , \nScanOut38[6] , 
        \nScanOut38[5] , \nScanOut38[4] , \nScanOut38[3] , \nScanOut38[2] , 
        \nScanOut38[1] , \nScanOut38[0] }), .ScanOut({\nScanOut37[7] , 
        \nScanOut37[6] , \nScanOut37[5] , \nScanOut37[4] , \nScanOut37[3] , 
        \nScanOut37[2] , \nScanOut37[1] , \nScanOut37[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , \nOut1_4[4] , \nOut1_4[3] , 
        \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }), .SouthIn({\nOut1_6[7] , 
        \nOut1_6[6] , \nOut1_6[5] , \nOut1_6[4] , \nOut1_6[3] , \nOut1_6[2] , 
        \nOut1_6[1] , \nOut1_6[0] }), .EastIn({\nOut2_5[7] , \nOut2_5[6] , 
        \nOut2_5[5] , \nOut2_5[4] , \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , 
        \nOut2_5[0] }), .WestIn({\nOut0_5[7] , \nOut0_5[6] , \nOut0_5[5] , 
        \nOut0_5[4] , \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , \nOut0_5[0] }), 
        .Out({\nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , \nOut1_5[4] , 
        \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_42 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut43[7] , \nScanOut43[6] , 
        \nScanOut43[5] , \nScanOut43[4] , \nScanOut43[3] , \nScanOut43[2] , 
        \nScanOut43[1] , \nScanOut43[0] }), .ScanOut({\nScanOut42[7] , 
        \nScanOut42[6] , \nScanOut42[5] , \nScanOut42[4] , \nScanOut42[3] , 
        \nScanOut42[2] , \nScanOut42[1] , \nScanOut42[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_9[7] , \nOut1_9[6] , \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , 
        \nOut1_9[2] , \nOut1_9[1] , \nOut1_9[0] }), .SouthIn({\nOut1_11[7] , 
        \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , \nOut1_11[3] , 
        \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), .EastIn({\nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), .WestIn({\nOut0_10[7] , 
        \nOut0_10[6] , \nOut0_10[5] , \nOut0_10[4] , \nOut0_10[3] , 
        \nOut0_10[2] , \nOut0_10[1] , \nOut0_10[0] }), .Out({\nOut1_10[7] , 
        \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , \nOut1_10[3] , 
        \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_657 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut658[7] , \nScanOut658[6] , 
        \nScanOut658[5] , \nScanOut658[4] , \nScanOut658[3] , \nScanOut658[2] , 
        \nScanOut658[1] , \nScanOut658[0] }), .ScanOut({\nScanOut657[7] , 
        \nScanOut657[6] , \nScanOut657[5] , \nScanOut657[4] , \nScanOut657[3] , 
        \nScanOut657[2] , \nScanOut657[1] , \nScanOut657[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_16[7] , \nOut20_16[6] , \nOut20_16[5] , \nOut20_16[4] , 
        \nOut20_16[3] , \nOut20_16[2] , \nOut20_16[1] , \nOut20_16[0] }), 
        .SouthIn({\nOut20_18[7] , \nOut20_18[6] , \nOut20_18[5] , 
        \nOut20_18[4] , \nOut20_18[3] , \nOut20_18[2] , \nOut20_18[1] , 
        \nOut20_18[0] }), .EastIn({\nOut21_17[7] , \nOut21_17[6] , 
        \nOut21_17[5] , \nOut21_17[4] , \nOut21_17[3] , \nOut21_17[2] , 
        \nOut21_17[1] , \nOut21_17[0] }), .WestIn({\nOut19_17[7] , 
        \nOut19_17[6] , \nOut19_17[5] , \nOut19_17[4] , \nOut19_17[3] , 
        \nOut19_17[2] , \nOut19_17[1] , \nOut19_17[0] }), .Out({\nOut20_17[7] , 
        \nOut20_17[6] , \nOut20_17[5] , \nOut20_17[4] , \nOut20_17[3] , 
        \nOut20_17[2] , \nOut20_17[1] , \nOut20_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_59 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut60[7] , \nScanOut60[6] , 
        \nScanOut60[5] , \nScanOut60[4] , \nScanOut60[3] , \nScanOut60[2] , 
        \nScanOut60[1] , \nScanOut60[0] }), .ScanOut({\nScanOut59[7] , 
        \nScanOut59[6] , \nScanOut59[5] , \nScanOut59[4] , \nScanOut59[3] , 
        \nScanOut59[2] , \nScanOut59[1] , \nScanOut59[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_26[7] , \nOut1_26[6] , \nOut1_26[5] , \nOut1_26[4] , 
        \nOut1_26[3] , \nOut1_26[2] , \nOut1_26[1] , \nOut1_26[0] }), 
        .SouthIn({\nOut1_28[7] , \nOut1_28[6] , \nOut1_28[5] , \nOut1_28[4] , 
        \nOut1_28[3] , \nOut1_28[2] , \nOut1_28[1] , \nOut1_28[0] }), .EastIn(
        {\nOut2_27[7] , \nOut2_27[6] , \nOut2_27[5] , \nOut2_27[4] , 
        \nOut2_27[3] , \nOut2_27[2] , \nOut2_27[1] , \nOut2_27[0] }), .WestIn(
        {\nOut0_27[7] , \nOut0_27[6] , \nOut0_27[5] , \nOut0_27[4] , 
        \nOut0_27[3] , \nOut0_27[2] , \nOut0_27[1] , \nOut0_27[0] }), .Out({
        \nOut1_27[7] , \nOut1_27[6] , \nOut1_27[5] , \nOut1_27[4] , 
        \nOut1_27[3] , \nOut1_27[2] , \nOut1_27[1] , \nOut1_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_65 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut66[7] , \nScanOut66[6] , 
        \nScanOut66[5] , \nScanOut66[4] , \nScanOut66[3] , \nScanOut66[2] , 
        \nScanOut66[1] , \nScanOut66[0] }), .ScanOut({\nScanOut65[7] , 
        \nScanOut65[6] , \nScanOut65[5] , \nScanOut65[4] , \nScanOut65[3] , 
        \nScanOut65[2] , \nScanOut65[1] , \nScanOut65[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_0[7] , \nOut2_0[6] , \nOut2_0[5] , \nOut2_0[4] , \nOut2_0[3] , 
        \nOut2_0[2] , \nOut2_0[1] , \nOut2_0[0] }), .SouthIn({\nOut2_2[7] , 
        \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , 
        \nOut2_2[1] , \nOut2_2[0] }), .EastIn({\nOut3_1[7] , \nOut3_1[6] , 
        \nOut3_1[5] , \nOut3_1[4] , \nOut3_1[3] , \nOut3_1[2] , \nOut3_1[1] , 
        \nOut3_1[0] }), .WestIn({\nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , 
        \nOut1_1[4] , \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), 
        .Out({\nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , \nOut2_1[4] , 
        \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_351 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut352[7] , \nScanOut352[6] , 
        \nScanOut352[5] , \nScanOut352[4] , \nScanOut352[3] , \nScanOut352[2] , 
        \nScanOut352[1] , \nScanOut352[0] }), .ScanOut({\nScanOut351[7] , 
        \nScanOut351[6] , \nScanOut351[5] , \nScanOut351[4] , \nScanOut351[3] , 
        \nScanOut351[2] , \nScanOut351[1] , \nScanOut351[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut10_31[7] , \nOut10_31[6] , 
        \nOut10_31[5] , \nOut10_31[4] , \nOut10_31[3] , \nOut10_31[2] , 
        \nOut10_31[1] , \nOut10_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_376 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut377[7] , \nScanOut377[6] , 
        \nScanOut377[5] , \nScanOut377[4] , \nScanOut377[3] , \nScanOut377[2] , 
        \nScanOut377[1] , \nScanOut377[0] }), .ScanOut({\nScanOut376[7] , 
        \nScanOut376[6] , \nScanOut376[5] , \nScanOut376[4] , \nScanOut376[3] , 
        \nScanOut376[2] , \nScanOut376[1] , \nScanOut376[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_23[7] , \nOut11_23[6] , \nOut11_23[5] , \nOut11_23[4] , 
        \nOut11_23[3] , \nOut11_23[2] , \nOut11_23[1] , \nOut11_23[0] }), 
        .SouthIn({\nOut11_25[7] , \nOut11_25[6] , \nOut11_25[5] , 
        \nOut11_25[4] , \nOut11_25[3] , \nOut11_25[2] , \nOut11_25[1] , 
        \nOut11_25[0] }), .EastIn({\nOut12_24[7] , \nOut12_24[6] , 
        \nOut12_24[5] , \nOut12_24[4] , \nOut12_24[3] , \nOut12_24[2] , 
        \nOut12_24[1] , \nOut12_24[0] }), .WestIn({\nOut10_24[7] , 
        \nOut10_24[6] , \nOut10_24[5] , \nOut10_24[4] , \nOut10_24[3] , 
        \nOut10_24[2] , \nOut10_24[1] , \nOut10_24[0] }), .Out({\nOut11_24[7] , 
        \nOut11_24[6] , \nOut11_24[5] , \nOut11_24[4] , \nOut11_24[3] , 
        \nOut11_24[2] , \nOut11_24[1] , \nOut11_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_567 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut568[7] , \nScanOut568[6] , 
        \nScanOut568[5] , \nScanOut568[4] , \nScanOut568[3] , \nScanOut568[2] , 
        \nScanOut568[1] , \nScanOut568[0] }), .ScanOut({\nScanOut567[7] , 
        \nScanOut567[6] , \nScanOut567[5] , \nScanOut567[4] , \nScanOut567[3] , 
        \nScanOut567[2] , \nScanOut567[1] , \nScanOut567[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_22[7] , \nOut17_22[6] , \nOut17_22[5] , \nOut17_22[4] , 
        \nOut17_22[3] , \nOut17_22[2] , \nOut17_22[1] , \nOut17_22[0] }), 
        .SouthIn({\nOut17_24[7] , \nOut17_24[6] , \nOut17_24[5] , 
        \nOut17_24[4] , \nOut17_24[3] , \nOut17_24[2] , \nOut17_24[1] , 
        \nOut17_24[0] }), .EastIn({\nOut18_23[7] , \nOut18_23[6] , 
        \nOut18_23[5] , \nOut18_23[4] , \nOut18_23[3] , \nOut18_23[2] , 
        \nOut18_23[1] , \nOut18_23[0] }), .WestIn({\nOut16_23[7] , 
        \nOut16_23[6] , \nOut16_23[5] , \nOut16_23[4] , \nOut16_23[3] , 
        \nOut16_23[2] , \nOut16_23[1] , \nOut16_23[0] }), .Out({\nOut17_23[7] , 
        \nOut17_23[6] , \nOut17_23[5] , \nOut17_23[4] , \nOut17_23[3] , 
        \nOut17_23[2] , \nOut17_23[1] , \nOut17_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_885 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut886[7] , \nScanOut886[6] , 
        \nScanOut886[5] , \nScanOut886[4] , \nScanOut886[3] , \nScanOut886[2] , 
        \nScanOut886[1] , \nScanOut886[0] }), .ScanOut({\nScanOut885[7] , 
        \nScanOut885[6] , \nScanOut885[5] , \nScanOut885[4] , \nScanOut885[3] , 
        \nScanOut885[2] , \nScanOut885[1] , \nScanOut885[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_20[7] , \nOut27_20[6] , \nOut27_20[5] , \nOut27_20[4] , 
        \nOut27_20[3] , \nOut27_20[2] , \nOut27_20[1] , \nOut27_20[0] }), 
        .SouthIn({\nOut27_22[7] , \nOut27_22[6] , \nOut27_22[5] , 
        \nOut27_22[4] , \nOut27_22[3] , \nOut27_22[2] , \nOut27_22[1] , 
        \nOut27_22[0] }), .EastIn({\nOut28_21[7] , \nOut28_21[6] , 
        \nOut28_21[5] , \nOut28_21[4] , \nOut28_21[3] , \nOut28_21[2] , 
        \nOut28_21[1] , \nOut28_21[0] }), .WestIn({\nOut26_21[7] , 
        \nOut26_21[6] , \nOut26_21[5] , \nOut26_21[4] , \nOut26_21[3] , 
        \nOut26_21[2] , \nOut26_21[1] , \nOut26_21[0] }), .Out({\nOut27_21[7] , 
        \nOut27_21[6] , \nOut27_21[5] , \nOut27_21[4] , \nOut27_21[3] , 
        \nOut27_21[2] , \nOut27_21[1] , \nOut27_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_915 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut916[7] , \nScanOut916[6] , 
        \nScanOut916[5] , \nScanOut916[4] , \nScanOut916[3] , \nScanOut916[2] , 
        \nScanOut916[1] , \nScanOut916[0] }), .ScanOut({\nScanOut915[7] , 
        \nScanOut915[6] , \nScanOut915[5] , \nScanOut915[4] , \nScanOut915[3] , 
        \nScanOut915[2] , \nScanOut915[1] , \nScanOut915[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_18[7] , \nOut28_18[6] , \nOut28_18[5] , \nOut28_18[4] , 
        \nOut28_18[3] , \nOut28_18[2] , \nOut28_18[1] , \nOut28_18[0] }), 
        .SouthIn({\nOut28_20[7] , \nOut28_20[6] , \nOut28_20[5] , 
        \nOut28_20[4] , \nOut28_20[3] , \nOut28_20[2] , \nOut28_20[1] , 
        \nOut28_20[0] }), .EastIn({\nOut29_19[7] , \nOut29_19[6] , 
        \nOut29_19[5] , \nOut29_19[4] , \nOut29_19[3] , \nOut29_19[2] , 
        \nOut29_19[1] , \nOut29_19[0] }), .WestIn({\nOut27_19[7] , 
        \nOut27_19[6] , \nOut27_19[5] , \nOut27_19[4] , \nOut27_19[3] , 
        \nOut27_19[2] , \nOut27_19[1] , \nOut27_19[0] }), .Out({\nOut28_19[7] , 
        \nOut28_19[6] , \nOut28_19[5] , \nOut28_19[4] , \nOut28_19[3] , 
        \nOut28_19[2] , \nOut28_19[1] , \nOut28_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_932 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut933[7] , \nScanOut933[6] , 
        \nScanOut933[5] , \nScanOut933[4] , \nScanOut933[3] , \nScanOut933[2] , 
        \nScanOut933[1] , \nScanOut933[0] }), .ScanOut({\nScanOut932[7] , 
        \nScanOut932[6] , \nScanOut932[5] , \nScanOut932[4] , \nScanOut932[3] , 
        \nScanOut932[2] , \nScanOut932[1] , \nScanOut932[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_3[7] , \nOut29_3[6] , \nOut29_3[5] , \nOut29_3[4] , 
        \nOut29_3[3] , \nOut29_3[2] , \nOut29_3[1] , \nOut29_3[0] }), 
        .SouthIn({\nOut29_5[7] , \nOut29_5[6] , \nOut29_5[5] , \nOut29_5[4] , 
        \nOut29_5[3] , \nOut29_5[2] , \nOut29_5[1] , \nOut29_5[0] }), .EastIn(
        {\nOut30_4[7] , \nOut30_4[6] , \nOut30_4[5] , \nOut30_4[4] , 
        \nOut30_4[3] , \nOut30_4[2] , \nOut30_4[1] , \nOut30_4[0] }), .WestIn(
        {\nOut28_4[7] , \nOut28_4[6] , \nOut28_4[5] , \nOut28_4[4] , 
        \nOut28_4[3] , \nOut28_4[2] , \nOut28_4[1] , \nOut28_4[0] }), .Out({
        \nOut29_4[7] , \nOut29_4[6] , \nOut29_4[5] , \nOut29_4[4] , 
        \nOut29_4[3] , \nOut29_4[2] , \nOut29_4[1] , \nOut29_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_540 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut541[7] , \nScanOut541[6] , 
        \nScanOut541[5] , \nScanOut541[4] , \nScanOut541[3] , \nScanOut541[2] , 
        \nScanOut541[1] , \nScanOut541[0] }), .ScanOut({\nScanOut540[7] , 
        \nScanOut540[6] , \nScanOut540[5] , \nScanOut540[4] , \nScanOut540[3] , 
        \nScanOut540[2] , \nScanOut540[1] , \nScanOut540[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_27[7] , \nOut16_27[6] , \nOut16_27[5] , \nOut16_27[4] , 
        \nOut16_27[3] , \nOut16_27[2] , \nOut16_27[1] , \nOut16_27[0] }), 
        .SouthIn({\nOut16_29[7] , \nOut16_29[6] , \nOut16_29[5] , 
        \nOut16_29[4] , \nOut16_29[3] , \nOut16_29[2] , \nOut16_29[1] , 
        \nOut16_29[0] }), .EastIn({\nOut17_28[7] , \nOut17_28[6] , 
        \nOut17_28[5] , \nOut17_28[4] , \nOut17_28[3] , \nOut17_28[2] , 
        \nOut17_28[1] , \nOut17_28[0] }), .WestIn({\nOut15_28[7] , 
        \nOut15_28[6] , \nOut15_28[5] , \nOut15_28[4] , \nOut15_28[3] , 
        \nOut15_28[2] , \nOut15_28[1] , \nOut15_28[0] }), .Out({\nOut16_28[7] , 
        \nOut16_28[6] , \nOut16_28[5] , \nOut16_28[4] , \nOut16_28[3] , 
        \nOut16_28[2] , \nOut16_28[1] , \nOut16_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_670 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut671[7] , \nScanOut671[6] , 
        \nScanOut671[5] , \nScanOut671[4] , \nScanOut671[3] , \nScanOut671[2] , 
        \nScanOut671[1] , \nScanOut671[0] }), .ScanOut({\nScanOut670[7] , 
        \nScanOut670[6] , \nScanOut670[5] , \nScanOut670[4] , \nScanOut670[3] , 
        \nScanOut670[2] , \nScanOut670[1] , \nScanOut670[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_29[7] , \nOut20_29[6] , \nOut20_29[5] , \nOut20_29[4] , 
        \nOut20_29[3] , \nOut20_29[2] , \nOut20_29[1] , \nOut20_29[0] }), 
        .SouthIn({\nOut20_31[7] , \nOut20_31[6] , \nOut20_31[5] , 
        \nOut20_31[4] , \nOut20_31[3] , \nOut20_31[2] , \nOut20_31[1] , 
        \nOut20_31[0] }), .EastIn({\nOut21_30[7] , \nOut21_30[6] , 
        \nOut21_30[5] , \nOut21_30[4] , \nOut21_30[3] , \nOut21_30[2] , 
        \nOut21_30[1] , \nOut21_30[0] }), .WestIn({\nOut19_30[7] , 
        \nOut19_30[6] , \nOut19_30[5] , \nOut19_30[4] , \nOut19_30[3] , 
        \nOut19_30[2] , \nOut19_30[1] , \nOut19_30[0] }), .Out({\nOut20_30[7] , 
        \nOut20_30[6] , \nOut20_30[5] , \nOut20_30[4] , \nOut20_30[3] , 
        \nOut20_30[2] , \nOut20_30[1] , \nOut20_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_146 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut147[7] , \nScanOut147[6] , 
        \nScanOut147[5] , \nScanOut147[4] , \nScanOut147[3] , \nScanOut147[2] , 
        \nScanOut147[1] , \nScanOut147[0] }), .ScanOut({\nScanOut146[7] , 
        \nScanOut146[6] , \nScanOut146[5] , \nScanOut146[4] , \nScanOut146[3] , 
        \nScanOut146[2] , \nScanOut146[1] , \nScanOut146[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_17[7] , \nOut4_17[6] , \nOut4_17[5] , \nOut4_17[4] , 
        \nOut4_17[3] , \nOut4_17[2] , \nOut4_17[1] , \nOut4_17[0] }), 
        .SouthIn({\nOut4_19[7] , \nOut4_19[6] , \nOut4_19[5] , \nOut4_19[4] , 
        \nOut4_19[3] , \nOut4_19[2] , \nOut4_19[1] , \nOut4_19[0] }), .EastIn(
        {\nOut5_18[7] , \nOut5_18[6] , \nOut5_18[5] , \nOut5_18[4] , 
        \nOut5_18[3] , \nOut5_18[2] , \nOut5_18[1] , \nOut5_18[0] }), .WestIn(
        {\nOut3_18[7] , \nOut3_18[6] , \nOut3_18[5] , \nOut3_18[4] , 
        \nOut3_18[3] , \nOut3_18[2] , \nOut3_18[1] , \nOut3_18[0] }), .Out({
        \nOut4_18[7] , \nOut4_18[6] , \nOut4_18[5] , \nOut4_18[4] , 
        \nOut4_18[3] , \nOut4_18[2] , \nOut4_18[1] , \nOut4_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_161 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut162[7] , \nScanOut162[6] , 
        \nScanOut162[5] , \nScanOut162[4] , \nScanOut162[3] , \nScanOut162[2] , 
        \nScanOut162[1] , \nScanOut162[0] }), .ScanOut({\nScanOut161[7] , 
        \nScanOut161[6] , \nScanOut161[5] , \nScanOut161[4] , \nScanOut161[3] , 
        \nScanOut161[2] , \nScanOut161[1] , \nScanOut161[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_0[7] , \nOut5_0[6] , \nOut5_0[5] , \nOut5_0[4] , \nOut5_0[3] , 
        \nOut5_0[2] , \nOut5_0[1] , \nOut5_0[0] }), .SouthIn({\nOut5_2[7] , 
        \nOut5_2[6] , \nOut5_2[5] , \nOut5_2[4] , \nOut5_2[3] , \nOut5_2[2] , 
        \nOut5_2[1] , \nOut5_2[0] }), .EastIn({\nOut6_1[7] , \nOut6_1[6] , 
        \nOut6_1[5] , \nOut6_1[4] , \nOut6_1[3] , \nOut6_1[2] , \nOut6_1[1] , 
        \nOut6_1[0] }), .WestIn({\nOut4_1[7] , \nOut4_1[6] , \nOut4_1[5] , 
        \nOut4_1[4] , \nOut4_1[3] , \nOut4_1[2] , \nOut4_1[1] , \nOut4_1[0] }), 
        .Out({\nOut5_1[7] , \nOut5_1[6] , \nOut5_1[5] , \nOut5_1[4] , 
        \nOut5_1[3] , \nOut5_1[2] , \nOut5_1[1] , \nOut5_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_770 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut771[7] , \nScanOut771[6] , 
        \nScanOut771[5] , \nScanOut771[4] , \nScanOut771[3] , \nScanOut771[2] , 
        \nScanOut771[1] , \nScanOut771[0] }), .ScanOut({\nScanOut770[7] , 
        \nScanOut770[6] , \nScanOut770[5] , \nScanOut770[4] , \nScanOut770[3] , 
        \nScanOut770[2] , \nScanOut770[1] , \nScanOut770[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_1[7] , \nOut24_1[6] , \nOut24_1[5] , \nOut24_1[4] , 
        \nOut24_1[3] , \nOut24_1[2] , \nOut24_1[1] , \nOut24_1[0] }), 
        .SouthIn({\nOut24_3[7] , \nOut24_3[6] , \nOut24_3[5] , \nOut24_3[4] , 
        \nOut24_3[3] , \nOut24_3[2] , \nOut24_3[1] , \nOut24_3[0] }), .EastIn(
        {\nOut25_2[7] , \nOut25_2[6] , \nOut25_2[5] , \nOut25_2[4] , 
        \nOut25_2[3] , \nOut25_2[2] , \nOut25_2[1] , \nOut25_2[0] }), .WestIn(
        {\nOut23_2[7] , \nOut23_2[6] , \nOut23_2[5] , \nOut23_2[4] , 
        \nOut23_2[3] , \nOut23_2[2] , \nOut23_2[1] , \nOut23_2[0] }), .Out({
        \nOut24_2[7] , \nOut24_2[6] , \nOut24_2[5] , \nOut24_2[4] , 
        \nOut24_2[3] , \nOut24_2[2] , \nOut24_2[1] , \nOut24_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_829 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut830[7] , \nScanOut830[6] , 
        \nScanOut830[5] , \nScanOut830[4] , \nScanOut830[3] , \nScanOut830[2] , 
        \nScanOut830[1] , \nScanOut830[0] }), .ScanOut({\nScanOut829[7] , 
        \nScanOut829[6] , \nScanOut829[5] , \nScanOut829[4] , \nScanOut829[3] , 
        \nScanOut829[2] , \nScanOut829[1] , \nScanOut829[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_28[7] , \nOut25_28[6] , \nOut25_28[5] , \nOut25_28[4] , 
        \nOut25_28[3] , \nOut25_28[2] , \nOut25_28[1] , \nOut25_28[0] }), 
        .SouthIn({\nOut25_30[7] , \nOut25_30[6] , \nOut25_30[5] , 
        \nOut25_30[4] , \nOut25_30[3] , \nOut25_30[2] , \nOut25_30[1] , 
        \nOut25_30[0] }), .EastIn({\nOut26_29[7] , \nOut26_29[6] , 
        \nOut26_29[5] , \nOut26_29[4] , \nOut26_29[3] , \nOut26_29[2] , 
        \nOut26_29[1] , \nOut26_29[0] }), .WestIn({\nOut24_29[7] , 
        \nOut24_29[6] , \nOut24_29[5] , \nOut24_29[4] , \nOut24_29[3] , 
        \nOut24_29[2] , \nOut24_29[1] , \nOut24_29[0] }), .Out({\nOut25_29[7] , 
        \nOut25_29[6] , \nOut25_29[5] , \nOut25_29[4] , \nOut25_29[3] , 
        \nOut25_29[2] , \nOut25_29[1] , \nOut25_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_251 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut252[7] , \nScanOut252[6] , 
        \nScanOut252[5] , \nScanOut252[4] , \nScanOut252[3] , \nScanOut252[2] , 
        \nScanOut252[1] , \nScanOut252[0] }), .ScanOut({\nScanOut251[7] , 
        \nScanOut251[6] , \nScanOut251[5] , \nScanOut251[4] , \nScanOut251[3] , 
        \nScanOut251[2] , \nScanOut251[1] , \nScanOut251[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_26[7] , \nOut7_26[6] , \nOut7_26[5] , \nOut7_26[4] , 
        \nOut7_26[3] , \nOut7_26[2] , \nOut7_26[1] , \nOut7_26[0] }), 
        .SouthIn({\nOut7_28[7] , \nOut7_28[6] , \nOut7_28[5] , \nOut7_28[4] , 
        \nOut7_28[3] , \nOut7_28[2] , \nOut7_28[1] , \nOut7_28[0] }), .EastIn(
        {\nOut8_27[7] , \nOut8_27[6] , \nOut8_27[5] , \nOut8_27[4] , 
        \nOut8_27[3] , \nOut8_27[2] , \nOut8_27[1] , \nOut8_27[0] }), .WestIn(
        {\nOut6_27[7] , \nOut6_27[6] , \nOut6_27[5] , \nOut6_27[4] , 
        \nOut6_27[3] , \nOut6_27[2] , \nOut6_27[1] , \nOut6_27[0] }), .Out({
        \nOut7_27[7] , \nOut7_27[6] , \nOut7_27[5] , \nOut7_27[4] , 
        \nOut7_27[3] , \nOut7_27[2] , \nOut7_27[1] , \nOut7_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_440 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut441[7] , \nScanOut441[6] , 
        \nScanOut441[5] , \nScanOut441[4] , \nScanOut441[3] , \nScanOut441[2] , 
        \nScanOut441[1] , \nScanOut441[0] }), .ScanOut({\nScanOut440[7] , 
        \nScanOut440[6] , \nScanOut440[5] , \nScanOut440[4] , \nScanOut440[3] , 
        \nScanOut440[2] , \nScanOut440[1] , \nScanOut440[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_23[7] , \nOut13_23[6] , \nOut13_23[5] , \nOut13_23[4] , 
        \nOut13_23[3] , \nOut13_23[2] , \nOut13_23[1] , \nOut13_23[0] }), 
        .SouthIn({\nOut13_25[7] , \nOut13_25[6] , \nOut13_25[5] , 
        \nOut13_25[4] , \nOut13_25[3] , \nOut13_25[2] , \nOut13_25[1] , 
        \nOut13_25[0] }), .EastIn({\nOut14_24[7] , \nOut14_24[6] , 
        \nOut14_24[5] , \nOut14_24[4] , \nOut14_24[3] , \nOut14_24[2] , 
        \nOut14_24[1] , \nOut14_24[0] }), .WestIn({\nOut12_24[7] , 
        \nOut12_24[6] , \nOut12_24[5] , \nOut12_24[4] , \nOut12_24[3] , 
        \nOut12_24[2] , \nOut12_24[1] , \nOut12_24[0] }), .Out({\nOut13_24[7] , 
        \nOut13_24[6] , \nOut13_24[5] , \nOut13_24[4] , \nOut13_24[3] , 
        \nOut13_24[2] , \nOut13_24[1] , \nOut13_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_832 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut833[7] , \nScanOut833[6] , 
        \nScanOut833[5] , \nScanOut833[4] , \nScanOut833[3] , \nScanOut833[2] , 
        \nScanOut833[1] , \nScanOut833[0] }), .ScanOut({\nScanOut832[7] , 
        \nScanOut832[6] , \nScanOut832[5] , \nScanOut832[4] , \nScanOut832[3] , 
        \nScanOut832[2] , \nScanOut832[1] , \nScanOut832[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut26_0[7] , \nOut26_0[6] , 
        \nOut26_0[5] , \nOut26_0[4] , \nOut26_0[3] , \nOut26_0[2] , 
        \nOut26_0[1] , \nOut26_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_276 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut277[7] , \nScanOut277[6] , 
        \nScanOut277[5] , \nScanOut277[4] , \nScanOut277[3] , \nScanOut277[2] , 
        \nScanOut277[1] , \nScanOut277[0] }), .ScanOut({\nScanOut276[7] , 
        \nScanOut276[6] , \nScanOut276[5] , \nScanOut276[4] , \nScanOut276[3] , 
        \nScanOut276[2] , \nScanOut276[1] , \nScanOut276[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_19[7] , \nOut8_19[6] , \nOut8_19[5] , \nOut8_19[4] , 
        \nOut8_19[3] , \nOut8_19[2] , \nOut8_19[1] , \nOut8_19[0] }), 
        .SouthIn({\nOut8_21[7] , \nOut8_21[6] , \nOut8_21[5] , \nOut8_21[4] , 
        \nOut8_21[3] , \nOut8_21[2] , \nOut8_21[1] , \nOut8_21[0] }), .EastIn(
        {\nOut9_20[7] , \nOut9_20[6] , \nOut9_20[5] , \nOut9_20[4] , 
        \nOut9_20[3] , \nOut9_20[2] , \nOut9_20[1] , \nOut9_20[0] }), .WestIn(
        {\nOut7_20[7] , \nOut7_20[6] , \nOut7_20[5] , \nOut7_20[4] , 
        \nOut7_20[3] , \nOut7_20[2] , \nOut7_20[1] , \nOut7_20[0] }), .Out({
        \nOut8_20[7] , \nOut8_20[6] , \nOut8_20[5] , \nOut8_20[4] , 
        \nOut8_20[3] , \nOut8_20[2] , \nOut8_20[1] , \nOut8_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_815 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut816[7] , \nScanOut816[6] , 
        \nScanOut816[5] , \nScanOut816[4] , \nScanOut816[3] , \nScanOut816[2] , 
        \nScanOut816[1] , \nScanOut816[0] }), .ScanOut({\nScanOut815[7] , 
        \nScanOut815[6] , \nScanOut815[5] , \nScanOut815[4] , \nScanOut815[3] , 
        \nScanOut815[2] , \nScanOut815[1] , \nScanOut815[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_14[7] , \nOut25_14[6] , \nOut25_14[5] , \nOut25_14[4] , 
        \nOut25_14[3] , \nOut25_14[2] , \nOut25_14[1] , \nOut25_14[0] }), 
        .SouthIn({\nOut25_16[7] , \nOut25_16[6] , \nOut25_16[5] , 
        \nOut25_16[4] , \nOut25_16[3] , \nOut25_16[2] , \nOut25_16[1] , 
        \nOut25_16[0] }), .EastIn({\nOut26_15[7] , \nOut26_15[6] , 
        \nOut26_15[5] , \nOut26_15[4] , \nOut26_15[3] , \nOut26_15[2] , 
        \nOut26_15[1] , \nOut26_15[0] }), .WestIn({\nOut24_15[7] , 
        \nOut24_15[6] , \nOut24_15[5] , \nOut24_15[4] , \nOut24_15[3] , 
        \nOut24_15[2] , \nOut24_15[1] , \nOut24_15[0] }), .Out({\nOut25_15[7] , 
        \nOut25_15[6] , \nOut25_15[5] , \nOut25_15[4] , \nOut25_15[3] , 
        \nOut25_15[2] , \nOut25_15[1] , \nOut25_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_985 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut986[7] , \nScanOut986[6] , 
        \nScanOut986[5] , \nScanOut986[4] , \nScanOut986[3] , \nScanOut986[2] , 
        \nScanOut986[1] , \nScanOut986[0] }), .ScanOut({\nScanOut985[7] , 
        \nScanOut985[6] , \nScanOut985[5] , \nScanOut985[4] , \nScanOut985[3] , 
        \nScanOut985[2] , \nScanOut985[1] , \nScanOut985[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_24[7] , \nOut30_24[6] , \nOut30_24[5] , \nOut30_24[4] , 
        \nOut30_24[3] , \nOut30_24[2] , \nOut30_24[1] , \nOut30_24[0] }), 
        .SouthIn({\nOut30_26[7] , \nOut30_26[6] , \nOut30_26[5] , 
        \nOut30_26[4] , \nOut30_26[3] , \nOut30_26[2] , \nOut30_26[1] , 
        \nOut30_26[0] }), .EastIn({\nOut31_25[7] , \nOut31_25[6] , 
        \nOut31_25[5] , \nOut31_25[4] , \nOut31_25[3] , \nOut31_25[2] , 
        \nOut31_25[1] , \nOut31_25[0] }), .WestIn({\nOut29_25[7] , 
        \nOut29_25[6] , \nOut29_25[5] , \nOut29_25[4] , \nOut29_25[3] , 
        \nOut29_25[2] , \nOut29_25[1] , \nOut29_25[0] }), .Out({\nOut30_25[7] , 
        \nOut30_25[6] , \nOut30_25[5] , \nOut30_25[4] , \nOut30_25[3] , 
        \nOut30_25[2] , \nOut30_25[1] , \nOut30_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_467 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut468[7] , \nScanOut468[6] , 
        \nScanOut468[5] , \nScanOut468[4] , \nScanOut468[3] , \nScanOut468[2] , 
        \nScanOut468[1] , \nScanOut468[0] }), .ScanOut({\nScanOut467[7] , 
        \nScanOut467[6] , \nScanOut467[5] , \nScanOut467[4] , \nScanOut467[3] , 
        \nScanOut467[2] , \nScanOut467[1] , \nScanOut467[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_18[7] , \nOut14_18[6] , \nOut14_18[5] , \nOut14_18[4] , 
        \nOut14_18[3] , \nOut14_18[2] , \nOut14_18[1] , \nOut14_18[0] }), 
        .SouthIn({\nOut14_20[7] , \nOut14_20[6] , \nOut14_20[5] , 
        \nOut14_20[4] , \nOut14_20[3] , \nOut14_20[2] , \nOut14_20[1] , 
        \nOut14_20[0] }), .EastIn({\nOut15_19[7] , \nOut15_19[6] , 
        \nOut15_19[5] , \nOut15_19[4] , \nOut15_19[3] , \nOut15_19[2] , 
        \nOut15_19[1] , \nOut15_19[0] }), .WestIn({\nOut13_19[7] , 
        \nOut13_19[6] , \nOut13_19[5] , \nOut13_19[4] , \nOut13_19[3] , 
        \nOut13_19[2] , \nOut13_19[1] , \nOut13_19[0] }), .Out({\nOut14_19[7] , 
        \nOut14_19[6] , \nOut14_19[5] , \nOut14_19[4] , \nOut14_19[3] , 
        \nOut14_19[2] , \nOut14_19[1] , \nOut14_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_757 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut758[7] , \nScanOut758[6] , 
        \nScanOut758[5] , \nScanOut758[4] , \nScanOut758[3] , \nScanOut758[2] , 
        \nScanOut758[1] , \nScanOut758[0] }), .ScanOut({\nScanOut757[7] , 
        \nScanOut757[6] , \nScanOut757[5] , \nScanOut757[4] , \nScanOut757[3] , 
        \nScanOut757[2] , \nScanOut757[1] , \nScanOut757[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_20[7] , \nOut23_20[6] , \nOut23_20[5] , \nOut23_20[4] , 
        \nOut23_20[3] , \nOut23_20[2] , \nOut23_20[1] , \nOut23_20[0] }), 
        .SouthIn({\nOut23_22[7] , \nOut23_22[6] , \nOut23_22[5] , 
        \nOut23_22[4] , \nOut23_22[3] , \nOut23_22[2] , \nOut23_22[1] , 
        \nOut23_22[0] }), .EastIn({\nOut24_21[7] , \nOut24_21[6] , 
        \nOut24_21[5] , \nOut24_21[4] , \nOut24_21[3] , \nOut24_21[2] , 
        \nOut24_21[1] , \nOut24_21[0] }), .WestIn({\nOut22_21[7] , 
        \nOut22_21[6] , \nOut22_21[5] , \nOut22_21[4] , \nOut22_21[3] , 
        \nOut22_21[2] , \nOut22_21[1] , \nOut22_21[0] }), .Out({\nOut23_21[7] , 
        \nOut23_21[6] , \nOut23_21[5] , \nOut23_21[4] , \nOut23_21[3] , 
        \nOut23_21[2] , \nOut23_21[1] , \nOut23_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_929 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut930[7] , \nScanOut930[6] , 
        \nScanOut930[5] , \nScanOut930[4] , \nScanOut930[3] , \nScanOut930[2] , 
        \nScanOut930[1] , \nScanOut930[0] }), .ScanOut({\nScanOut929[7] , 
        \nScanOut929[6] , \nScanOut929[5] , \nScanOut929[4] , \nScanOut929[3] , 
        \nScanOut929[2] , \nScanOut929[1] , \nScanOut929[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_0[7] , \nOut29_0[6] , \nOut29_0[5] , \nOut29_0[4] , 
        \nOut29_0[3] , \nOut29_0[2] , \nOut29_0[1] , \nOut29_0[0] }), 
        .SouthIn({\nOut29_2[7] , \nOut29_2[6] , \nOut29_2[5] , \nOut29_2[4] , 
        \nOut29_2[3] , \nOut29_2[2] , \nOut29_2[1] , \nOut29_2[0] }), .EastIn(
        {\nOut30_1[7] , \nOut30_1[6] , \nOut30_1[5] , \nOut30_1[4] , 
        \nOut30_1[3] , \nOut30_1[2] , \nOut30_1[1] , \nOut30_1[0] }), .WestIn(
        {\nOut28_1[7] , \nOut28_1[6] , \nOut28_1[5] , \nOut28_1[4] , 
        \nOut28_1[3] , \nOut28_1[2] , \nOut28_1[1] , \nOut28_1[0] }), .Out({
        \nOut29_1[7] , \nOut29_1[6] , \nOut29_1[5] , \nOut29_1[4] , 
        \nOut29_1[3] , \nOut29_1[2] , \nOut29_1[1] , \nOut29_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_293 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut294[7] , \nScanOut294[6] , 
        \nScanOut294[5] , \nScanOut294[4] , \nScanOut294[3] , \nScanOut294[2] , 
        \nScanOut294[1] , \nScanOut294[0] }), .ScanOut({\nScanOut293[7] , 
        \nScanOut293[6] , \nScanOut293[5] , \nScanOut293[4] , \nScanOut293[3] , 
        \nScanOut293[2] , \nScanOut293[1] , \nScanOut293[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_4[7] , \nOut9_4[6] , \nOut9_4[5] , \nOut9_4[4] , \nOut9_4[3] , 
        \nOut9_4[2] , \nOut9_4[1] , \nOut9_4[0] }), .SouthIn({\nOut9_6[7] , 
        \nOut9_6[6] , \nOut9_6[5] , \nOut9_6[4] , \nOut9_6[3] , \nOut9_6[2] , 
        \nOut9_6[1] , \nOut9_6[0] }), .EastIn({\nOut10_5[7] , \nOut10_5[6] , 
        \nOut10_5[5] , \nOut10_5[4] , \nOut10_5[3] , \nOut10_5[2] , 
        \nOut10_5[1] , \nOut10_5[0] }), .WestIn({\nOut8_5[7] , \nOut8_5[6] , 
        \nOut8_5[5] , \nOut8_5[4] , \nOut8_5[3] , \nOut8_5[2] , \nOut8_5[1] , 
        \nOut8_5[0] }), .Out({\nOut9_5[7] , \nOut9_5[6] , \nOut9_5[5] , 
        \nOut9_5[4] , \nOut9_5[3] , \nOut9_5[2] , \nOut9_5[1] , \nOut9_5[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_303 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut304[7] , \nScanOut304[6] , 
        \nScanOut304[5] , \nScanOut304[4] , \nScanOut304[3] , \nScanOut304[2] , 
        \nScanOut304[1] , \nScanOut304[0] }), .ScanOut({\nScanOut303[7] , 
        \nScanOut303[6] , \nScanOut303[5] , \nScanOut303[4] , \nScanOut303[3] , 
        \nScanOut303[2] , \nScanOut303[1] , \nScanOut303[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_14[7] , \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , 
        \nOut9_14[3] , \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }), 
        .SouthIn({\nOut9_16[7] , \nOut9_16[6] , \nOut9_16[5] , \nOut9_16[4] , 
        \nOut9_16[3] , \nOut9_16[2] , \nOut9_16[1] , \nOut9_16[0] }), .EastIn(
        {\nOut10_15[7] , \nOut10_15[6] , \nOut10_15[5] , \nOut10_15[4] , 
        \nOut10_15[3] , \nOut10_15[2] , \nOut10_15[1] , \nOut10_15[0] }), 
        .WestIn({\nOut8_15[7] , \nOut8_15[6] , \nOut8_15[5] , \nOut8_15[4] , 
        \nOut8_15[3] , \nOut8_15[2] , \nOut8_15[1] , \nOut8_15[0] }), .Out({
        \nOut9_15[7] , \nOut9_15[6] , \nOut9_15[5] , \nOut9_15[4] , 
        \nOut9_15[3] , \nOut9_15[2] , \nOut9_15[1] , \nOut9_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_482 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut483[7] , \nScanOut483[6] , 
        \nScanOut483[5] , \nScanOut483[4] , \nScanOut483[3] , \nScanOut483[2] , 
        \nScanOut483[1] , \nScanOut483[0] }), .ScanOut({\nScanOut482[7] , 
        \nScanOut482[6] , \nScanOut482[5] , \nScanOut482[4] , \nScanOut482[3] , 
        \nScanOut482[2] , \nScanOut482[1] , \nScanOut482[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_1[7] , \nOut15_1[6] , \nOut15_1[5] , \nOut15_1[4] , 
        \nOut15_1[3] , \nOut15_1[2] , \nOut15_1[1] , \nOut15_1[0] }), 
        .SouthIn({\nOut15_3[7] , \nOut15_3[6] , \nOut15_3[5] , \nOut15_3[4] , 
        \nOut15_3[3] , \nOut15_3[2] , \nOut15_3[1] , \nOut15_3[0] }), .EastIn(
        {\nOut16_2[7] , \nOut16_2[6] , \nOut16_2[5] , \nOut16_2[4] , 
        \nOut16_2[3] , \nOut16_2[2] , \nOut16_2[1] , \nOut16_2[0] }), .WestIn(
        {\nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }), .Out({
        \nOut15_2[7] , \nOut15_2[6] , \nOut15_2[5] , \nOut15_2[4] , 
        \nOut15_2[3] , \nOut15_2[2] , \nOut15_2[1] , \nOut15_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_960 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut961[7] , \nScanOut961[6] , 
        \nScanOut961[5] , \nScanOut961[4] , \nScanOut961[3] , \nScanOut961[2] , 
        \nScanOut961[1] , \nScanOut961[0] }), .ScanOut({\nScanOut960[7] , 
        \nScanOut960[6] , \nScanOut960[5] , \nScanOut960[4] , \nScanOut960[3] , 
        \nScanOut960[2] , \nScanOut960[1] , \nScanOut960[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut30_0[7] , \nOut30_0[6] , 
        \nOut30_0[5] , \nOut30_0[4] , \nOut30_0[3] , \nOut30_0[2] , 
        \nOut30_0[1] , \nOut30_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_512 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut513[7] , \nScanOut513[6] , 
        \nScanOut513[5] , \nScanOut513[4] , \nScanOut513[3] , \nScanOut513[2] , 
        \nScanOut513[1] , \nScanOut513[0] }), .ScanOut({\nScanOut512[7] , 
        \nScanOut512[6] , \nScanOut512[5] , \nScanOut512[4] , \nScanOut512[3] , 
        \nScanOut512[2] , \nScanOut512[1] , \nScanOut512[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut16_0[7] , \nOut16_0[6] , 
        \nOut16_0[5] , \nOut16_0[4] , \nOut16_0[3] , \nOut16_0[2] , 
        \nOut16_0[1] , \nOut16_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_622 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut623[7] , \nScanOut623[6] , 
        \nScanOut623[5] , \nScanOut623[4] , \nScanOut623[3] , \nScanOut623[2] , 
        \nScanOut623[1] , \nScanOut623[0] }), .ScanOut({\nScanOut622[7] , 
        \nScanOut622[6] , \nScanOut622[5] , \nScanOut622[4] , \nScanOut622[3] , 
        \nScanOut622[2] , \nScanOut622[1] , \nScanOut622[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_13[7] , \nOut19_13[6] , \nOut19_13[5] , \nOut19_13[4] , 
        \nOut19_13[3] , \nOut19_13[2] , \nOut19_13[1] , \nOut19_13[0] }), 
        .SouthIn({\nOut19_15[7] , \nOut19_15[6] , \nOut19_15[5] , 
        \nOut19_15[4] , \nOut19_15[3] , \nOut19_15[2] , \nOut19_15[1] , 
        \nOut19_15[0] }), .EastIn({\nOut20_14[7] , \nOut20_14[6] , 
        \nOut20_14[5] , \nOut20_14[4] , \nOut20_14[3] , \nOut20_14[2] , 
        \nOut20_14[1] , \nOut20_14[0] }), .WestIn({\nOut18_14[7] , 
        \nOut18_14[6] , \nOut18_14[5] , \nOut18_14[4] , \nOut18_14[3] , 
        \nOut18_14[2] , \nOut18_14[1] , \nOut18_14[0] }), .Out({\nOut19_14[7] , 
        \nOut19_14[6] , \nOut19_14[5] , \nOut19_14[4] , \nOut19_14[3] , 
        \nOut19_14[2] , \nOut19_14[1] , \nOut19_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_17 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut18[7] , \nScanOut18[6] , 
        \nScanOut18[5] , \nScanOut18[4] , \nScanOut18[3] , \nScanOut18[2] , 
        \nScanOut18[1] , \nScanOut18[0] }), .ScanOut({\nScanOut17[7] , 
        \nScanOut17[6] , \nScanOut17[5] , \nScanOut17[4] , \nScanOut17[3] , 
        \nScanOut17[2] , \nScanOut17[1] , \nScanOut17[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_17[7] , \nOut0_17[6] , 
        \nOut0_17[5] , \nOut0_17[4] , \nOut0_17[3] , \nOut0_17[2] , 
        \nOut0_17[1] , \nOut0_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_128 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut129[7] , \nScanOut129[6] , 
        \nScanOut129[5] , \nScanOut129[4] , \nScanOut129[3] , \nScanOut129[2] , 
        \nScanOut129[1] , \nScanOut129[0] }), .ScanOut({\nScanOut128[7] , 
        \nScanOut128[6] , \nScanOut128[5] , \nScanOut128[4] , \nScanOut128[3] , 
        \nScanOut128[2] , \nScanOut128[1] , \nScanOut128[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut4_0[7] , \nOut4_0[6] , 
        \nOut4_0[5] , \nOut4_0[4] , \nOut4_0[3] , \nOut4_0[2] , \nOut4_0[1] , 
        \nOut4_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_184 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut185[7] , \nScanOut185[6] , 
        \nScanOut185[5] , \nScanOut185[4] , \nScanOut185[3] , \nScanOut185[2] , 
        \nScanOut185[1] , \nScanOut185[0] }), .ScanOut({\nScanOut184[7] , 
        \nScanOut184[6] , \nScanOut184[5] , \nScanOut184[4] , \nScanOut184[3] , 
        \nScanOut184[2] , \nScanOut184[1] , \nScanOut184[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_23[7] , \nOut5_23[6] , \nOut5_23[5] , \nOut5_23[4] , 
        \nOut5_23[3] , \nOut5_23[2] , \nOut5_23[1] , \nOut5_23[0] }), 
        .SouthIn({\nOut5_25[7] , \nOut5_25[6] , \nOut5_25[5] , \nOut5_25[4] , 
        \nOut5_25[3] , \nOut5_25[2] , \nOut5_25[1] , \nOut5_25[0] }), .EastIn(
        {\nOut6_24[7] , \nOut6_24[6] , \nOut6_24[5] , \nOut6_24[4] , 
        \nOut6_24[3] , \nOut6_24[2] , \nOut6_24[1] , \nOut6_24[0] }), .WestIn(
        {\nOut4_24[7] , \nOut4_24[6] , \nOut4_24[5] , \nOut4_24[4] , 
        \nOut4_24[3] , \nOut4_24[2] , \nOut4_24[1] , \nOut4_24[0] }), .Out({
        \nOut5_24[7] , \nOut5_24[6] , \nOut5_24[5] , \nOut5_24[4] , 
        \nOut5_24[3] , \nOut5_24[2] , \nOut5_24[1] , \nOut5_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_218 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut219[7] , \nScanOut219[6] , 
        \nScanOut219[5] , \nScanOut219[4] , \nScanOut219[3] , \nScanOut219[2] , 
        \nScanOut219[1] , \nScanOut219[0] }), .ScanOut({\nScanOut218[7] , 
        \nScanOut218[6] , \nScanOut218[5] , \nScanOut218[4] , \nScanOut218[3] , 
        \nScanOut218[2] , \nScanOut218[1] , \nScanOut218[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_25[7] , \nOut6_25[6] , \nOut6_25[5] , \nOut6_25[4] , 
        \nOut6_25[3] , \nOut6_25[2] , \nOut6_25[1] , \nOut6_25[0] }), 
        .SouthIn({\nOut6_27[7] , \nOut6_27[6] , \nOut6_27[5] , \nOut6_27[4] , 
        \nOut6_27[3] , \nOut6_27[2] , \nOut6_27[1] , \nOut6_27[0] }), .EastIn(
        {\nOut7_26[7] , \nOut7_26[6] , \nOut7_26[5] , \nOut7_26[4] , 
        \nOut7_26[3] , \nOut7_26[2] , \nOut7_26[1] , \nOut7_26[0] }), .WestIn(
        {\nOut5_26[7] , \nOut5_26[6] , \nOut5_26[5] , \nOut5_26[4] , 
        \nOut5_26[3] , \nOut5_26[2] , \nOut5_26[1] , \nOut5_26[0] }), .Out({
        \nOut6_26[7] , \nOut6_26[6] , \nOut6_26[5] , \nOut6_26[4] , 
        \nOut6_26[3] , \nOut6_26[2] , \nOut6_26[1] , \nOut6_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_324 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut325[7] , \nScanOut325[6] , 
        \nScanOut325[5] , \nScanOut325[4] , \nScanOut325[3] , \nScanOut325[2] , 
        \nScanOut325[1] , \nScanOut325[0] }), .ScanOut({\nScanOut324[7] , 
        \nScanOut324[6] , \nScanOut324[5] , \nScanOut324[4] , \nScanOut324[3] , 
        \nScanOut324[2] , \nScanOut324[1] , \nScanOut324[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_3[7] , \nOut10_3[6] , \nOut10_3[5] , \nOut10_3[4] , 
        \nOut10_3[3] , \nOut10_3[2] , \nOut10_3[1] , \nOut10_3[0] }), 
        .SouthIn({\nOut10_5[7] , \nOut10_5[6] , \nOut10_5[5] , \nOut10_5[4] , 
        \nOut10_5[3] , \nOut10_5[2] , \nOut10_5[1] , \nOut10_5[0] }), .EastIn(
        {\nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }), .WestIn(
        {\nOut9_4[7] , \nOut9_4[6] , \nOut9_4[5] , \nOut9_4[4] , \nOut9_4[3] , 
        \nOut9_4[2] , \nOut9_4[1] , \nOut9_4[0] }), .Out({\nOut10_4[7] , 
        \nOut10_4[6] , \nOut10_4[5] , \nOut10_4[4] , \nOut10_4[3] , 
        \nOut10_4[2] , \nOut10_4[1] , \nOut10_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_535 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut536[7] , \nScanOut536[6] , 
        \nScanOut536[5] , \nScanOut536[4] , \nScanOut536[3] , \nScanOut536[2] , 
        \nScanOut536[1] , \nScanOut536[0] }), .ScanOut({\nScanOut535[7] , 
        \nScanOut535[6] , \nScanOut535[5] , \nScanOut535[4] , \nScanOut535[3] , 
        \nScanOut535[2] , \nScanOut535[1] , \nScanOut535[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_22[7] , \nOut16_22[6] , \nOut16_22[5] , \nOut16_22[4] , 
        \nOut16_22[3] , \nOut16_22[2] , \nOut16_22[1] , \nOut16_22[0] }), 
        .SouthIn({\nOut16_24[7] , \nOut16_24[6] , \nOut16_24[5] , 
        \nOut16_24[4] , \nOut16_24[3] , \nOut16_24[2] , \nOut16_24[1] , 
        \nOut16_24[0] }), .EastIn({\nOut17_23[7] , \nOut17_23[6] , 
        \nOut17_23[5] , \nOut17_23[4] , \nOut17_23[3] , \nOut17_23[2] , 
        \nOut17_23[1] , \nOut17_23[0] }), .WestIn({\nOut15_23[7] , 
        \nOut15_23[6] , \nOut15_23[5] , \nOut15_23[4] , \nOut15_23[3] , 
        \nOut15_23[2] , \nOut15_23[1] , \nOut15_23[0] }), .Out({\nOut16_23[7] , 
        \nOut16_23[6] , \nOut16_23[5] , \nOut16_23[4] , \nOut16_23[3] , 
        \nOut16_23[2] , \nOut16_23[1] , \nOut16_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_605 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut606[7] , \nScanOut606[6] , 
        \nScanOut606[5] , \nScanOut606[4] , \nScanOut606[3] , \nScanOut606[2] , 
        \nScanOut606[1] , \nScanOut606[0] }), .ScanOut({\nScanOut605[7] , 
        \nScanOut605[6] , \nScanOut605[5] , \nScanOut605[4] , \nScanOut605[3] , 
        \nScanOut605[2] , \nScanOut605[1] , \nScanOut605[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_28[7] , \nOut18_28[6] , \nOut18_28[5] , \nOut18_28[4] , 
        \nOut18_28[3] , \nOut18_28[2] , \nOut18_28[1] , \nOut18_28[0] }), 
        .SouthIn({\nOut18_30[7] , \nOut18_30[6] , \nOut18_30[5] , 
        \nOut18_30[4] , \nOut18_30[3] , \nOut18_30[2] , \nOut18_30[1] , 
        \nOut18_30[0] }), .EastIn({\nOut19_29[7] , \nOut19_29[6] , 
        \nOut19_29[5] , \nOut19_29[4] , \nOut19_29[3] , \nOut19_29[2] , 
        \nOut19_29[1] , \nOut19_29[0] }), .WestIn({\nOut17_29[7] , 
        \nOut17_29[6] , \nOut17_29[5] , \nOut17_29[4] , \nOut17_29[3] , 
        \nOut17_29[2] , \nOut17_29[1] , \nOut17_29[0] }), .Out({\nOut18_29[7] , 
        \nOut18_29[6] , \nOut18_29[5] , \nOut18_29[4] , \nOut18_29[3] , 
        \nOut18_29[2] , \nOut18_29[1] , \nOut18_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_795 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut796[7] , \nScanOut796[6] , 
        \nScanOut796[5] , \nScanOut796[4] , \nScanOut796[3] , \nScanOut796[2] , 
        \nScanOut796[1] , \nScanOut796[0] }), .ScanOut({\nScanOut795[7] , 
        \nScanOut795[6] , \nScanOut795[5] , \nScanOut795[4] , \nScanOut795[3] , 
        \nScanOut795[2] , \nScanOut795[1] , \nScanOut795[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_26[7] , \nOut24_26[6] , \nOut24_26[5] , \nOut24_26[4] , 
        \nOut24_26[3] , \nOut24_26[2] , \nOut24_26[1] , \nOut24_26[0] }), 
        .SouthIn({\nOut24_28[7] , \nOut24_28[6] , \nOut24_28[5] , 
        \nOut24_28[4] , \nOut24_28[3] , \nOut24_28[2] , \nOut24_28[1] , 
        \nOut24_28[0] }), .EastIn({\nOut25_27[7] , \nOut25_27[6] , 
        \nOut25_27[5] , \nOut25_27[4] , \nOut25_27[3] , \nOut25_27[2] , 
        \nOut25_27[1] , \nOut25_27[0] }), .WestIn({\nOut23_27[7] , 
        \nOut23_27[6] , \nOut23_27[5] , \nOut23_27[4] , \nOut23_27[3] , 
        \nOut23_27[2] , \nOut23_27[1] , \nOut23_27[0] }), .Out({\nOut24_27[7] , 
        \nOut24_27[6] , \nOut24_27[5] , \nOut24_27[4] , \nOut24_27[3] , 
        \nOut24_27[2] , \nOut24_27[1] , \nOut24_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_947 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut948[7] , \nScanOut948[6] , 
        \nScanOut948[5] , \nScanOut948[4] , \nScanOut948[3] , \nScanOut948[2] , 
        \nScanOut948[1] , \nScanOut948[0] }), .ScanOut({\nScanOut947[7] , 
        \nScanOut947[6] , \nScanOut947[5] , \nScanOut947[4] , \nScanOut947[3] , 
        \nScanOut947[2] , \nScanOut947[1] , \nScanOut947[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_18[7] , \nOut29_18[6] , \nOut29_18[5] , \nOut29_18[4] , 
        \nOut29_18[3] , \nOut29_18[2] , \nOut29_18[1] , \nOut29_18[0] }), 
        .SouthIn({\nOut29_20[7] , \nOut29_20[6] , \nOut29_20[5] , 
        \nOut29_20[4] , \nOut29_20[3] , \nOut29_20[2] , \nOut29_20[1] , 
        \nOut29_20[0] }), .EastIn({\nOut30_19[7] , \nOut30_19[6] , 
        \nOut30_19[5] , \nOut30_19[4] , \nOut30_19[3] , \nOut30_19[2] , 
        \nOut30_19[1] , \nOut30_19[0] }), .WestIn({\nOut28_19[7] , 
        \nOut28_19[6] , \nOut28_19[5] , \nOut28_19[4] , \nOut28_19[3] , 
        \nOut28_19[2] , \nOut28_19[1] , \nOut28_19[0] }), .Out({\nOut29_19[7] , 
        \nOut29_19[6] , \nOut29_19[5] , \nOut29_19[4] , \nOut29_19[3] , 
        \nOut29_19[2] , \nOut29_19[1] , \nOut29_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_388 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut389[7] , \nScanOut389[6] , 
        \nScanOut389[5] , \nScanOut389[4] , \nScanOut389[3] , \nScanOut389[2] , 
        \nScanOut389[1] , \nScanOut389[0] }), .ScanOut({\nScanOut388[7] , 
        \nScanOut388[6] , \nScanOut388[5] , \nScanOut388[4] , \nScanOut388[3] , 
        \nScanOut388[2] , \nScanOut388[1] , \nScanOut388[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }), 
        .SouthIn({\nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }), .EastIn(
        {\nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }), .WestIn(
        {\nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }), .Out({
        \nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_409 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut410[7] , \nScanOut410[6] , 
        \nScanOut410[5] , \nScanOut410[4] , \nScanOut410[3] , \nScanOut410[2] , 
        \nScanOut410[1] , \nScanOut410[0] }), .ScanOut({\nScanOut409[7] , 
        \nScanOut409[6] , \nScanOut409[5] , \nScanOut409[4] , \nScanOut409[3] , 
        \nScanOut409[2] , \nScanOut409[1] , \nScanOut409[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_24[7] , \nOut12_24[6] , \nOut12_24[5] , \nOut12_24[4] , 
        \nOut12_24[3] , \nOut12_24[2] , \nOut12_24[1] , \nOut12_24[0] }), 
        .SouthIn({\nOut12_26[7] , \nOut12_26[6] , \nOut12_26[5] , 
        \nOut12_26[4] , \nOut12_26[3] , \nOut12_26[2] , \nOut12_26[1] , 
        \nOut12_26[0] }), .EastIn({\nOut13_25[7] , \nOut13_25[6] , 
        \nOut13_25[5] , \nOut13_25[4] , \nOut13_25[3] , \nOut13_25[2] , 
        \nOut13_25[1] , \nOut13_25[0] }), .WestIn({\nOut11_25[7] , 
        \nOut11_25[6] , \nOut11_25[5] , \nOut11_25[4] , \nOut11_25[3] , 
        \nOut11_25[2] , \nOut11_25[1] , \nOut11_25[0] }), .Out({\nOut12_25[7] , 
        \nOut12_25[6] , \nOut12_25[5] , \nOut12_25[4] , \nOut12_25[3] , 
        \nOut12_25[2] , \nOut12_25[1] , \nOut12_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_599 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut600[7] , \nScanOut600[6] , 
        \nScanOut600[5] , \nScanOut600[4] , \nScanOut600[3] , \nScanOut600[2] , 
        \nScanOut600[1] , \nScanOut600[0] }), .ScanOut({\nScanOut599[7] , 
        \nScanOut599[6] , \nScanOut599[5] , \nScanOut599[4] , \nScanOut599[3] , 
        \nScanOut599[2] , \nScanOut599[1] , \nScanOut599[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_22[7] , \nOut18_22[6] , \nOut18_22[5] , \nOut18_22[4] , 
        \nOut18_22[3] , \nOut18_22[2] , \nOut18_22[1] , \nOut18_22[0] }), 
        .SouthIn({\nOut18_24[7] , \nOut18_24[6] , \nOut18_24[5] , 
        \nOut18_24[4] , \nOut18_24[3] , \nOut18_24[2] , \nOut18_24[1] , 
        \nOut18_24[0] }), .EastIn({\nOut19_23[7] , \nOut19_23[6] , 
        \nOut19_23[5] , \nOut19_23[4] , \nOut19_23[3] , \nOut19_23[2] , 
        \nOut19_23[1] , \nOut19_23[0] }), .WestIn({\nOut17_23[7] , 
        \nOut17_23[6] , \nOut17_23[5] , \nOut17_23[4] , \nOut17_23[3] , 
        \nOut17_23[2] , \nOut17_23[1] , \nOut17_23[0] }), .Out({\nOut18_23[7] , 
        \nOut18_23[6] , \nOut18_23[5] , \nOut18_23[4] , \nOut18_23[3] , 
        \nOut18_23[2] , \nOut18_23[1] , \nOut18_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_739 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut740[7] , \nScanOut740[6] , 
        \nScanOut740[5] , \nScanOut740[4] , \nScanOut740[3] , \nScanOut740[2] , 
        \nScanOut740[1] , \nScanOut740[0] }), .ScanOut({\nScanOut739[7] , 
        \nScanOut739[6] , \nScanOut739[5] , \nScanOut739[4] , \nScanOut739[3] , 
        \nScanOut739[2] , \nScanOut739[1] , \nScanOut739[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_2[7] , \nOut23_2[6] , \nOut23_2[5] , \nOut23_2[4] , 
        \nOut23_2[3] , \nOut23_2[2] , \nOut23_2[1] , \nOut23_2[0] }), 
        .SouthIn({\nOut23_4[7] , \nOut23_4[6] , \nOut23_4[5] , \nOut23_4[4] , 
        \nOut23_4[3] , \nOut23_4[2] , \nOut23_4[1] , \nOut23_4[0] }), .EastIn(
        {\nOut24_3[7] , \nOut24_3[6] , \nOut24_3[5] , \nOut24_3[4] , 
        \nOut24_3[3] , \nOut24_3[2] , \nOut24_3[1] , \nOut24_3[0] }), .WestIn(
        {\nOut22_3[7] , \nOut22_3[6] , \nOut22_3[5] , \nOut22_3[4] , 
        \nOut22_3[3] , \nOut22_3[2] , \nOut22_3[1] , \nOut22_3[0] }), .Out({
        \nOut23_3[7] , \nOut23_3[6] , \nOut23_3[5] , \nOut23_3[4] , 
        \nOut23_3[3] , \nOut23_3[2] , \nOut23_3[1] , \nOut23_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_183 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut184[7] , \nScanOut184[6] , 
        \nScanOut184[5] , \nScanOut184[4] , \nScanOut184[3] , \nScanOut184[2] , 
        \nScanOut184[1] , \nScanOut184[0] }), .ScanOut({\nScanOut183[7] , 
        \nScanOut183[6] , \nScanOut183[5] , \nScanOut183[4] , \nScanOut183[3] , 
        \nScanOut183[2] , \nScanOut183[1] , \nScanOut183[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_22[7] , \nOut5_22[6] , \nOut5_22[5] , \nOut5_22[4] , 
        \nOut5_22[3] , \nOut5_22[2] , \nOut5_22[1] , \nOut5_22[0] }), 
        .SouthIn({\nOut5_24[7] , \nOut5_24[6] , \nOut5_24[5] , \nOut5_24[4] , 
        \nOut5_24[3] , \nOut5_24[2] , \nOut5_24[1] , \nOut5_24[0] }), .EastIn(
        {\nOut6_23[7] , \nOut6_23[6] , \nOut6_23[5] , \nOut6_23[4] , 
        \nOut6_23[3] , \nOut6_23[2] , \nOut6_23[1] , \nOut6_23[0] }), .WestIn(
        {\nOut4_23[7] , \nOut4_23[6] , \nOut4_23[5] , \nOut4_23[4] , 
        \nOut4_23[3] , \nOut4_23[2] , \nOut4_23[1] , \nOut4_23[0] }), .Out({
        \nOut5_23[7] , \nOut5_23[6] , \nOut5_23[5] , \nOut5_23[4] , 
        \nOut5_23[3] , \nOut5_23[2] , \nOut5_23[1] , \nOut5_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_323 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut324[7] , \nScanOut324[6] , 
        \nScanOut324[5] , \nScanOut324[4] , \nScanOut324[3] , \nScanOut324[2] , 
        \nScanOut324[1] , \nScanOut324[0] }), .ScanOut({\nScanOut323[7] , 
        \nScanOut323[6] , \nScanOut323[5] , \nScanOut323[4] , \nScanOut323[3] , 
        \nScanOut323[2] , \nScanOut323[1] , \nScanOut323[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_2[7] , \nOut10_2[6] , \nOut10_2[5] , \nOut10_2[4] , 
        \nOut10_2[3] , \nOut10_2[2] , \nOut10_2[1] , \nOut10_2[0] }), 
        .SouthIn({\nOut10_4[7] , \nOut10_4[6] , \nOut10_4[5] , \nOut10_4[4] , 
        \nOut10_4[3] , \nOut10_4[2] , \nOut10_4[1] , \nOut10_4[0] }), .EastIn(
        {\nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }), .WestIn(
        {\nOut9_3[7] , \nOut9_3[6] , \nOut9_3[5] , \nOut9_3[4] , \nOut9_3[3] , 
        \nOut9_3[2] , \nOut9_3[1] , \nOut9_3[0] }), .Out({\nOut10_3[7] , 
        \nOut10_3[6] , \nOut10_3[5] , \nOut10_3[4] , \nOut10_3[3] , 
        \nOut10_3[2] , \nOut10_3[1] , \nOut10_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1018 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1019[7] , \nScanOut1019[6] , 
        \nScanOut1019[5] , \nScanOut1019[4] , \nScanOut1019[3] , 
        \nScanOut1019[2] , \nScanOut1019[1] , \nScanOut1019[0] }), .ScanOut({
        \nScanOut1018[7] , \nScanOut1018[6] , \nScanOut1018[5] , 
        \nScanOut1018[4] , \nScanOut1018[3] , \nScanOut1018[2] , 
        \nScanOut1018[1] , \nScanOut1018[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_26[7] , \nOut31_26[6] , \nOut31_26[5] , 
        \nOut31_26[4] , \nOut31_26[3] , \nOut31_26[2] , \nOut31_26[1] , 
        \nOut31_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_532 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut533[7] , \nScanOut533[6] , 
        \nScanOut533[5] , \nScanOut533[4] , \nScanOut533[3] , \nScanOut533[2] , 
        \nScanOut533[1] , \nScanOut533[0] }), .ScanOut({\nScanOut532[7] , 
        \nScanOut532[6] , \nScanOut532[5] , \nScanOut532[4] , \nScanOut532[3] , 
        \nScanOut532[2] , \nScanOut532[1] , \nScanOut532[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_19[7] , \nOut16_19[6] , \nOut16_19[5] , \nOut16_19[4] , 
        \nOut16_19[3] , \nOut16_19[2] , \nOut16_19[1] , \nOut16_19[0] }), 
        .SouthIn({\nOut16_21[7] , \nOut16_21[6] , \nOut16_21[5] , 
        \nOut16_21[4] , \nOut16_21[3] , \nOut16_21[2] , \nOut16_21[1] , 
        \nOut16_21[0] }), .EastIn({\nOut17_20[7] , \nOut17_20[6] , 
        \nOut17_20[5] , \nOut17_20[4] , \nOut17_20[3] , \nOut17_20[2] , 
        \nOut17_20[1] , \nOut17_20[0] }), .WestIn({\nOut15_20[7] , 
        \nOut15_20[6] , \nOut15_20[5] , \nOut15_20[4] , \nOut15_20[3] , 
        \nOut15_20[2] , \nOut15_20[1] , \nOut15_20[0] }), .Out({\nOut16_20[7] , 
        \nOut16_20[6] , \nOut16_20[5] , \nOut16_20[4] , \nOut16_20[3] , 
        \nOut16_20[2] , \nOut16_20[1] , \nOut16_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_602 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut603[7] , \nScanOut603[6] , 
        \nScanOut603[5] , \nScanOut603[4] , \nScanOut603[3] , \nScanOut603[2] , 
        \nScanOut603[1] , \nScanOut603[0] }), .ScanOut({\nScanOut602[7] , 
        \nScanOut602[6] , \nScanOut602[5] , \nScanOut602[4] , \nScanOut602[3] , 
        \nScanOut602[2] , \nScanOut602[1] , \nScanOut602[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_25[7] , \nOut18_25[6] , \nOut18_25[5] , \nOut18_25[4] , 
        \nOut18_25[3] , \nOut18_25[2] , \nOut18_25[1] , \nOut18_25[0] }), 
        .SouthIn({\nOut18_27[7] , \nOut18_27[6] , \nOut18_27[5] , 
        \nOut18_27[4] , \nOut18_27[3] , \nOut18_27[2] , \nOut18_27[1] , 
        \nOut18_27[0] }), .EastIn({\nOut19_26[7] , \nOut19_26[6] , 
        \nOut19_26[5] , \nOut19_26[4] , \nOut19_26[3] , \nOut19_26[2] , 
        \nOut19_26[1] , \nOut19_26[0] }), .WestIn({\nOut17_26[7] , 
        \nOut17_26[6] , \nOut17_26[5] , \nOut17_26[4] , \nOut17_26[3] , 
        \nOut17_26[2] , \nOut17_26[1] , \nOut17_26[0] }), .Out({\nOut18_26[7] , 
        \nOut18_26[6] , \nOut18_26[5] , \nOut18_26[4] , \nOut18_26[3] , 
        \nOut18_26[2] , \nOut18_26[1] , \nOut18_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_792 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut793[7] , \nScanOut793[6] , 
        \nScanOut793[5] , \nScanOut793[4] , \nScanOut793[3] , \nScanOut793[2] , 
        \nScanOut793[1] , \nScanOut793[0] }), .ScanOut({\nScanOut792[7] , 
        \nScanOut792[6] , \nScanOut792[5] , \nScanOut792[4] , \nScanOut792[3] , 
        \nScanOut792[2] , \nScanOut792[1] , \nScanOut792[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_23[7] , \nOut24_23[6] , \nOut24_23[5] , \nOut24_23[4] , 
        \nOut24_23[3] , \nOut24_23[2] , \nOut24_23[1] , \nOut24_23[0] }), 
        .SouthIn({\nOut24_25[7] , \nOut24_25[6] , \nOut24_25[5] , 
        \nOut24_25[4] , \nOut24_25[3] , \nOut24_25[2] , \nOut24_25[1] , 
        \nOut24_25[0] }), .EastIn({\nOut25_24[7] , \nOut25_24[6] , 
        \nOut25_24[5] , \nOut25_24[4] , \nOut25_24[3] , \nOut25_24[2] , 
        \nOut25_24[1] , \nOut25_24[0] }), .WestIn({\nOut23_24[7] , 
        \nOut23_24[6] , \nOut23_24[5] , \nOut23_24[4] , \nOut23_24[3] , 
        \nOut23_24[2] , \nOut23_24[1] , \nOut23_24[0] }), .Out({\nOut24_24[7] , 
        \nOut24_24[6] , \nOut24_24[5] , \nOut24_24[4] , \nOut24_24[3] , 
        \nOut24_24[2] , \nOut24_24[1] , \nOut24_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_940 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut941[7] , \nScanOut941[6] , 
        \nScanOut941[5] , \nScanOut941[4] , \nScanOut941[3] , \nScanOut941[2] , 
        \nScanOut941[1] , \nScanOut941[0] }), .ScanOut({\nScanOut940[7] , 
        \nScanOut940[6] , \nScanOut940[5] , \nScanOut940[4] , \nScanOut940[3] , 
        \nScanOut940[2] , \nScanOut940[1] , \nScanOut940[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_11[7] , \nOut29_11[6] , \nOut29_11[5] , \nOut29_11[4] , 
        \nOut29_11[3] , \nOut29_11[2] , \nOut29_11[1] , \nOut29_11[0] }), 
        .SouthIn({\nOut29_13[7] , \nOut29_13[6] , \nOut29_13[5] , 
        \nOut29_13[4] , \nOut29_13[3] , \nOut29_13[2] , \nOut29_13[1] , 
        \nOut29_13[0] }), .EastIn({\nOut30_12[7] , \nOut30_12[6] , 
        \nOut30_12[5] , \nOut30_12[4] , \nOut30_12[3] , \nOut30_12[2] , 
        \nOut30_12[1] , \nOut30_12[0] }), .WestIn({\nOut28_12[7] , 
        \nOut28_12[6] , \nOut28_12[5] , \nOut28_12[4] , \nOut28_12[3] , 
        \nOut28_12[2] , \nOut28_12[1] , \nOut28_12[0] }), .Out({\nOut29_12[7] , 
        \nOut29_12[6] , \nOut29_12[5] , \nOut29_12[4] , \nOut29_12[3] , 
        \nOut29_12[2] , \nOut29_12[1] , \nOut29_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_30 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut31[7] , \nScanOut31[6] , 
        \nScanOut31[5] , \nScanOut31[4] , \nScanOut31[3] , \nScanOut31[2] , 
        \nScanOut31[1] , \nScanOut31[0] }), .ScanOut({\nScanOut30[7] , 
        \nScanOut30[6] , \nScanOut30[5] , \nScanOut30[4] , \nScanOut30[3] , 
        \nScanOut30[2] , \nScanOut30[1] , \nScanOut30[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_30[7] , \nOut0_30[6] , 
        \nOut0_30[5] , \nOut0_30[4] , \nOut0_30[3] , \nOut0_30[2] , 
        \nOut0_30[1] , \nOut0_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_625 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut626[7] , \nScanOut626[6] , 
        \nScanOut626[5] , \nScanOut626[4] , \nScanOut626[3] , \nScanOut626[2] , 
        \nScanOut626[1] , \nScanOut626[0] }), .ScanOut({\nScanOut625[7] , 
        \nScanOut625[6] , \nScanOut625[5] , \nScanOut625[4] , \nScanOut625[3] , 
        \nScanOut625[2] , \nScanOut625[1] , \nScanOut625[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_16[7] , \nOut19_16[6] , \nOut19_16[5] , \nOut19_16[4] , 
        \nOut19_16[3] , \nOut19_16[2] , \nOut19_16[1] , \nOut19_16[0] }), 
        .SouthIn({\nOut19_18[7] , \nOut19_18[6] , \nOut19_18[5] , 
        \nOut19_18[4] , \nOut19_18[3] , \nOut19_18[2] , \nOut19_18[1] , 
        \nOut19_18[0] }), .EastIn({\nOut20_17[7] , \nOut20_17[6] , 
        \nOut20_17[5] , \nOut20_17[4] , \nOut20_17[3] , \nOut20_17[2] , 
        \nOut20_17[1] , \nOut20_17[0] }), .WestIn({\nOut18_17[7] , 
        \nOut18_17[6] , \nOut18_17[5] , \nOut18_17[4] , \nOut18_17[3] , 
        \nOut18_17[2] , \nOut18_17[1] , \nOut18_17[0] }), .Out({\nOut19_17[7] , 
        \nOut19_17[6] , \nOut19_17[5] , \nOut19_17[4] , \nOut19_17[3] , 
        \nOut19_17[2] , \nOut19_17[1] , \nOut19_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_45 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut46[7] , \nScanOut46[6] , 
        \nScanOut46[5] , \nScanOut46[4] , \nScanOut46[3] , \nScanOut46[2] , 
        \nScanOut46[1] , \nScanOut46[0] }), .ScanOut({\nScanOut45[7] , 
        \nScanOut45[6] , \nScanOut45[5] , \nScanOut45[4] , \nScanOut45[3] , 
        \nScanOut45[2] , \nScanOut45[1] , \nScanOut45[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), 
        .SouthIn({\nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), .EastIn(
        {\nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), .WestIn(
        {\nOut0_13[7] , \nOut0_13[6] , \nOut0_13[5] , \nOut0_13[4] , 
        \nOut0_13[3] , \nOut0_13[2] , \nOut0_13[1] , \nOut0_13[0] }), .Out({
        \nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_62 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut63[7] , \nScanOut63[6] , 
        \nScanOut63[5] , \nScanOut63[4] , \nScanOut63[3] , \nScanOut63[2] , 
        \nScanOut63[1] , \nScanOut63[0] }), .ScanOut({\nScanOut62[7] , 
        \nScanOut62[6] , \nScanOut62[5] , \nScanOut62[4] , \nScanOut62[3] , 
        \nScanOut62[2] , \nScanOut62[1] , \nScanOut62[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_29[7] , \nOut1_29[6] , \nOut1_29[5] , \nOut1_29[4] , 
        \nOut1_29[3] , \nOut1_29[2] , \nOut1_29[1] , \nOut1_29[0] }), 
        .SouthIn({\nOut1_31[7] , \nOut1_31[6] , \nOut1_31[5] , \nOut1_31[4] , 
        \nOut1_31[3] , \nOut1_31[2] , \nOut1_31[1] , \nOut1_31[0] }), .EastIn(
        {\nOut2_30[7] , \nOut2_30[6] , \nOut2_30[5] , \nOut2_30[4] , 
        \nOut2_30[3] , \nOut2_30[2] , \nOut2_30[1] , \nOut2_30[0] }), .WestIn(
        {\nOut0_30[7] , \nOut0_30[6] , \nOut0_30[5] , \nOut0_30[4] , 
        \nOut0_30[3] , \nOut0_30[2] , \nOut0_30[1] , \nOut0_30[0] }), .Out({
        \nOut1_30[7] , \nOut1_30[6] , \nOut1_30[5] , \nOut1_30[4] , 
        \nOut1_30[3] , \nOut1_30[2] , \nOut1_30[1] , \nOut1_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_79 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut80[7] , \nScanOut80[6] , 
        \nScanOut80[5] , \nScanOut80[4] , \nScanOut80[3] , \nScanOut80[2] , 
        \nScanOut80[1] , \nScanOut80[0] }), .ScanOut({\nScanOut79[7] , 
        \nScanOut79[6] , \nScanOut79[5] , \nScanOut79[4] , \nScanOut79[3] , 
        \nScanOut79[2] , \nScanOut79[1] , \nScanOut79[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), 
        .SouthIn({\nOut2_16[7] , \nOut2_16[6] , \nOut2_16[5] , \nOut2_16[4] , 
        \nOut2_16[3] , \nOut2_16[2] , \nOut2_16[1] , \nOut2_16[0] }), .EastIn(
        {\nOut3_15[7] , \nOut3_15[6] , \nOut3_15[5] , \nOut3_15[4] , 
        \nOut3_15[3] , \nOut3_15[2] , \nOut3_15[1] , \nOut3_15[0] }), .WestIn(
        {\nOut1_15[7] , \nOut1_15[6] , \nOut1_15[5] , \nOut1_15[4] , 
        \nOut1_15[3] , \nOut1_15[2] , \nOut1_15[1] , \nOut1_15[0] }), .Out({
        \nOut2_15[7] , \nOut2_15[6] , \nOut2_15[5] , \nOut2_15[4] , 
        \nOut2_15[3] , \nOut2_15[2] , \nOut2_15[1] , \nOut2_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_108 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut109[7] , \nScanOut109[6] , 
        \nScanOut109[5] , \nScanOut109[4] , \nScanOut109[3] , \nScanOut109[2] , 
        \nScanOut109[1] , \nScanOut109[0] }), .ScanOut({\nScanOut108[7] , 
        \nScanOut108[6] , \nScanOut108[5] , \nScanOut108[4] , \nScanOut108[3] , 
        \nScanOut108[2] , \nScanOut108[1] , \nScanOut108[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_11[7] , \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , 
        \nOut3_11[3] , \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }), 
        .SouthIn({\nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }), .EastIn(
        {\nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }), .WestIn(
        {\nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), .Out({
        \nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_238 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut239[7] , \nScanOut239[6] , 
        \nScanOut239[5] , \nScanOut239[4] , \nScanOut239[3] , \nScanOut239[2] , 
        \nScanOut239[1] , \nScanOut239[0] }), .ScanOut({\nScanOut238[7] , 
        \nScanOut238[6] , \nScanOut238[5] , \nScanOut238[4] , \nScanOut238[3] , 
        \nScanOut238[2] , \nScanOut238[1] , \nScanOut238[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }), 
        .SouthIn({\nOut7_15[7] , \nOut7_15[6] , \nOut7_15[5] , \nOut7_15[4] , 
        \nOut7_15[3] , \nOut7_15[2] , \nOut7_15[1] , \nOut7_15[0] }), .EastIn(
        {\nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }), .WestIn(
        {\nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }), .Out({
        \nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_294 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut295[7] , \nScanOut295[6] , 
        \nScanOut295[5] , \nScanOut295[4] , \nScanOut295[3] , \nScanOut295[2] , 
        \nScanOut295[1] , \nScanOut295[0] }), .ScanOut({\nScanOut294[7] , 
        \nScanOut294[6] , \nScanOut294[5] , \nScanOut294[4] , \nScanOut294[3] , 
        \nScanOut294[2] , \nScanOut294[1] , \nScanOut294[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_5[7] , \nOut9_5[6] , \nOut9_5[5] , \nOut9_5[4] , \nOut9_5[3] , 
        \nOut9_5[2] , \nOut9_5[1] , \nOut9_5[0] }), .SouthIn({\nOut9_7[7] , 
        \nOut9_7[6] , \nOut9_7[5] , \nOut9_7[4] , \nOut9_7[3] , \nOut9_7[2] , 
        \nOut9_7[1] , \nOut9_7[0] }), .EastIn({\nOut10_6[7] , \nOut10_6[6] , 
        \nOut10_6[5] , \nOut10_6[4] , \nOut10_6[3] , \nOut10_6[2] , 
        \nOut10_6[1] , \nOut10_6[0] }), .WestIn({\nOut8_6[7] , \nOut8_6[6] , 
        \nOut8_6[5] , \nOut8_6[4] , \nOut8_6[3] , \nOut8_6[2] , \nOut8_6[1] , 
        \nOut8_6[0] }), .Out({\nOut9_6[7] , \nOut9_6[6] , \nOut9_6[5] , 
        \nOut9_6[4] , \nOut9_6[3] , \nOut9_6[2] , \nOut9_6[1] , \nOut9_6[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_304 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut305[7] , \nScanOut305[6] , 
        \nScanOut305[5] , \nScanOut305[4] , \nScanOut305[3] , \nScanOut305[2] , 
        \nScanOut305[1] , \nScanOut305[0] }), .ScanOut({\nScanOut304[7] , 
        \nScanOut304[6] , \nScanOut304[5] , \nScanOut304[4] , \nScanOut304[3] , 
        \nScanOut304[2] , \nScanOut304[1] , \nScanOut304[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_15[7] , \nOut9_15[6] , \nOut9_15[5] , \nOut9_15[4] , 
        \nOut9_15[3] , \nOut9_15[2] , \nOut9_15[1] , \nOut9_15[0] }), 
        .SouthIn({\nOut9_17[7] , \nOut9_17[6] , \nOut9_17[5] , \nOut9_17[4] , 
        \nOut9_17[3] , \nOut9_17[2] , \nOut9_17[1] , \nOut9_17[0] }), .EastIn(
        {\nOut10_16[7] , \nOut10_16[6] , \nOut10_16[5] , \nOut10_16[4] , 
        \nOut10_16[3] , \nOut10_16[2] , \nOut10_16[1] , \nOut10_16[0] }), 
        .WestIn({\nOut8_16[7] , \nOut8_16[6] , \nOut8_16[5] , \nOut8_16[4] , 
        \nOut8_16[3] , \nOut8_16[2] , \nOut8_16[1] , \nOut8_16[0] }), .Out({
        \nOut9_16[7] , \nOut9_16[6] , \nOut9_16[5] , \nOut9_16[4] , 
        \nOut9_16[3] , \nOut9_16[2] , \nOut9_16[1] , \nOut9_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_515 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut516[7] , \nScanOut516[6] , 
        \nScanOut516[5] , \nScanOut516[4] , \nScanOut516[3] , \nScanOut516[2] , 
        \nScanOut516[1] , \nScanOut516[0] }), .ScanOut({\nScanOut515[7] , 
        \nScanOut515[6] , \nScanOut515[5] , \nScanOut515[4] , \nScanOut515[3] , 
        \nScanOut515[2] , \nScanOut515[1] , \nScanOut515[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_2[7] , \nOut16_2[6] , \nOut16_2[5] , \nOut16_2[4] , 
        \nOut16_2[3] , \nOut16_2[2] , \nOut16_2[1] , \nOut16_2[0] }), 
        .SouthIn({\nOut16_4[7] , \nOut16_4[6] , \nOut16_4[5] , \nOut16_4[4] , 
        \nOut16_4[3] , \nOut16_4[2] , \nOut16_4[1] , \nOut16_4[0] }), .EastIn(
        {\nOut17_3[7] , \nOut17_3[6] , \nOut17_3[5] , \nOut17_3[4] , 
        \nOut17_3[3] , \nOut17_3[2] , \nOut17_3[1] , \nOut17_3[0] }), .WestIn(
        {\nOut15_3[7] , \nOut15_3[6] , \nOut15_3[5] , \nOut15_3[4] , 
        \nOut15_3[3] , \nOut15_3[2] , \nOut15_3[1] , \nOut15_3[0] }), .Out({
        \nOut16_3[7] , \nOut16_3[6] , \nOut16_3[5] , \nOut16_3[4] , 
        \nOut16_3[3] , \nOut16_3[2] , \nOut16_3[1] , \nOut16_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_429 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut430[7] , \nScanOut430[6] , 
        \nScanOut430[5] , \nScanOut430[4] , \nScanOut430[3] , \nScanOut430[2] , 
        \nScanOut430[1] , \nScanOut430[0] }), .ScanOut({\nScanOut429[7] , 
        \nScanOut429[6] , \nScanOut429[5] , \nScanOut429[4] , \nScanOut429[3] , 
        \nScanOut429[2] , \nScanOut429[1] , \nScanOut429[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_12[7] , \nOut13_12[6] , \nOut13_12[5] , \nOut13_12[4] , 
        \nOut13_12[3] , \nOut13_12[2] , \nOut13_12[1] , \nOut13_12[0] }), 
        .SouthIn({\nOut13_14[7] , \nOut13_14[6] , \nOut13_14[5] , 
        \nOut13_14[4] , \nOut13_14[3] , \nOut13_14[2] , \nOut13_14[1] , 
        \nOut13_14[0] }), .EastIn({\nOut14_13[7] , \nOut14_13[6] , 
        \nOut14_13[5] , \nOut14_13[4] , \nOut14_13[3] , \nOut14_13[2] , 
        \nOut14_13[1] , \nOut14_13[0] }), .WestIn({\nOut12_13[7] , 
        \nOut12_13[6] , \nOut12_13[5] , \nOut12_13[4] , \nOut12_13[3] , 
        \nOut12_13[2] , \nOut12_13[1] , \nOut12_13[0] }), .Out({\nOut13_13[7] , 
        \nOut13_13[6] , \nOut13_13[5] , \nOut13_13[4] , \nOut13_13[3] , 
        \nOut13_13[2] , \nOut13_13[1] , \nOut13_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_485 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut486[7] , \nScanOut486[6] , 
        \nScanOut486[5] , \nScanOut486[4] , \nScanOut486[3] , \nScanOut486[2] , 
        \nScanOut486[1] , \nScanOut486[0] }), .ScanOut({\nScanOut485[7] , 
        \nScanOut485[6] , \nScanOut485[5] , \nScanOut485[4] , \nScanOut485[3] , 
        \nScanOut485[2] , \nScanOut485[1] , \nScanOut485[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_4[7] , \nOut15_4[6] , \nOut15_4[5] , \nOut15_4[4] , 
        \nOut15_4[3] , \nOut15_4[2] , \nOut15_4[1] , \nOut15_4[0] }), 
        .SouthIn({\nOut15_6[7] , \nOut15_6[6] , \nOut15_6[5] , \nOut15_6[4] , 
        \nOut15_6[3] , \nOut15_6[2] , \nOut15_6[1] , \nOut15_6[0] }), .EastIn(
        {\nOut16_5[7] , \nOut16_5[6] , \nOut16_5[5] , \nOut16_5[4] , 
        \nOut16_5[3] , \nOut16_5[2] , \nOut16_5[1] , \nOut16_5[0] }), .WestIn(
        {\nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }), .Out({
        \nOut15_5[7] , \nOut15_5[6] , \nOut15_5[5] , \nOut15_5[4] , 
        \nOut15_5[3] , \nOut15_5[2] , \nOut15_5[1] , \nOut15_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_967 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut968[7] , \nScanOut968[6] , 
        \nScanOut968[5] , \nScanOut968[4] , \nScanOut968[3] , \nScanOut968[2] , 
        \nScanOut968[1] , \nScanOut968[0] }), .ScanOut({\nScanOut967[7] , 
        \nScanOut967[6] , \nScanOut967[5] , \nScanOut967[4] , \nScanOut967[3] , 
        \nScanOut967[2] , \nScanOut967[1] , \nScanOut967[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_6[7] , \nOut30_6[6] , \nOut30_6[5] , \nOut30_6[4] , 
        \nOut30_6[3] , \nOut30_6[2] , \nOut30_6[1] , \nOut30_6[0] }), 
        .SouthIn({\nOut30_8[7] , \nOut30_8[6] , \nOut30_8[5] , \nOut30_8[4] , 
        \nOut30_8[3] , \nOut30_8[2] , \nOut30_8[1] , \nOut30_8[0] }), .EastIn(
        {\nOut31_7[7] , \nOut31_7[6] , \nOut31_7[5] , \nOut31_7[4] , 
        \nOut31_7[3] , \nOut31_7[2] , \nOut31_7[1] , \nOut31_7[0] }), .WestIn(
        {\nOut29_7[7] , \nOut29_7[6] , \nOut29_7[5] , \nOut29_7[4] , 
        \nOut29_7[3] , \nOut29_7[2] , \nOut29_7[1] , \nOut29_7[0] }), .Out({
        \nOut30_7[7] , \nOut30_7[6] , \nOut30_7[5] , \nOut30_7[4] , 
        \nOut30_7[3] , \nOut30_7[2] , \nOut30_7[1] , \nOut30_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_689 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut690[7] , \nScanOut690[6] , 
        \nScanOut690[5] , \nScanOut690[4] , \nScanOut690[3] , \nScanOut690[2] , 
        \nScanOut690[1] , \nScanOut690[0] }), .ScanOut({\nScanOut689[7] , 
        \nScanOut689[6] , \nScanOut689[5] , \nScanOut689[4] , \nScanOut689[3] , 
        \nScanOut689[2] , \nScanOut689[1] , \nScanOut689[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_16[7] , \nOut21_16[6] , \nOut21_16[5] , \nOut21_16[4] , 
        \nOut21_16[3] , \nOut21_16[2] , \nOut21_16[1] , \nOut21_16[0] }), 
        .SouthIn({\nOut21_18[7] , \nOut21_18[6] , \nOut21_18[5] , 
        \nOut21_18[4] , \nOut21_18[3] , \nOut21_18[2] , \nOut21_18[1] , 
        \nOut21_18[0] }), .EastIn({\nOut22_17[7] , \nOut22_17[6] , 
        \nOut22_17[5] , \nOut22_17[4] , \nOut22_17[3] , \nOut22_17[2] , 
        \nOut22_17[1] , \nOut22_17[0] }), .WestIn({\nOut20_17[7] , 
        \nOut20_17[6] , \nOut20_17[5] , \nOut20_17[4] , \nOut20_17[3] , 
        \nOut20_17[2] , \nOut20_17[1] , \nOut20_17[0] }), .Out({\nOut21_17[7] , 
        \nOut21_17[6] , \nOut21_17[5] , \nOut21_17[4] , \nOut21_17[3] , 
        \nOut21_17[2] , \nOut21_17[1] , \nOut21_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_719 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut720[7] , \nScanOut720[6] , 
        \nScanOut720[5] , \nScanOut720[4] , \nScanOut720[3] , \nScanOut720[2] , 
        \nScanOut720[1] , \nScanOut720[0] }), .ScanOut({\nScanOut719[7] , 
        \nScanOut719[6] , \nScanOut719[5] , \nScanOut719[4] , \nScanOut719[3] , 
        \nScanOut719[2] , \nScanOut719[1] , \nScanOut719[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_14[7] , \nOut22_14[6] , \nOut22_14[5] , \nOut22_14[4] , 
        \nOut22_14[3] , \nOut22_14[2] , \nOut22_14[1] , \nOut22_14[0] }), 
        .SouthIn({\nOut22_16[7] , \nOut22_16[6] , \nOut22_16[5] , 
        \nOut22_16[4] , \nOut22_16[3] , \nOut22_16[2] , \nOut22_16[1] , 
        \nOut22_16[0] }), .EastIn({\nOut23_15[7] , \nOut23_15[6] , 
        \nOut23_15[5] , \nOut23_15[4] , \nOut23_15[3] , \nOut23_15[2] , 
        \nOut23_15[1] , \nOut23_15[0] }), .WestIn({\nOut21_15[7] , 
        \nOut21_15[6] , \nOut21_15[5] , \nOut21_15[4] , \nOut21_15[3] , 
        \nOut21_15[2] , \nOut21_15[1] , \nOut21_15[0] }), .Out({\nOut22_15[7] , 
        \nOut22_15[6] , \nOut22_15[5] , \nOut22_15[4] , \nOut22_15[3] , 
        \nOut22_15[2] , \nOut22_15[1] , \nOut22_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_141 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut142[7] , \nScanOut142[6] , 
        \nScanOut142[5] , \nScanOut142[4] , \nScanOut142[3] , \nScanOut142[2] , 
        \nScanOut142[1] , \nScanOut142[0] }), .ScanOut({\nScanOut141[7] , 
        \nScanOut141[6] , \nScanOut141[5] , \nScanOut141[4] , \nScanOut141[3] , 
        \nScanOut141[2] , \nScanOut141[1] , \nScanOut141[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }), 
        .SouthIn({\nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }), .EastIn(
        {\nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }), .WestIn(
        {\nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }), .Out({
        \nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_750 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut751[7] , \nScanOut751[6] , 
        \nScanOut751[5] , \nScanOut751[4] , \nScanOut751[3] , \nScanOut751[2] , 
        \nScanOut751[1] , \nScanOut751[0] }), .ScanOut({\nScanOut750[7] , 
        \nScanOut750[6] , \nScanOut750[5] , \nScanOut750[4] , \nScanOut750[3] , 
        \nScanOut750[2] , \nScanOut750[1] , \nScanOut750[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_13[7] , \nOut23_13[6] , \nOut23_13[5] , \nOut23_13[4] , 
        \nOut23_13[3] , \nOut23_13[2] , \nOut23_13[1] , \nOut23_13[0] }), 
        .SouthIn({\nOut23_15[7] , \nOut23_15[6] , \nOut23_15[5] , 
        \nOut23_15[4] , \nOut23_15[3] , \nOut23_15[2] , \nOut23_15[1] , 
        \nOut23_15[0] }), .EastIn({\nOut24_14[7] , \nOut24_14[6] , 
        \nOut24_14[5] , \nOut24_14[4] , \nOut24_14[3] , \nOut24_14[2] , 
        \nOut24_14[1] , \nOut24_14[0] }), .WestIn({\nOut22_14[7] , 
        \nOut22_14[6] , \nOut22_14[5] , \nOut22_14[4] , \nOut22_14[3] , 
        \nOut22_14[2] , \nOut22_14[1] , \nOut22_14[0] }), .Out({\nOut23_14[7] , 
        \nOut23_14[6] , \nOut23_14[5] , \nOut23_14[4] , \nOut23_14[3] , 
        \nOut23_14[2] , \nOut23_14[1] , \nOut23_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_166 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut167[7] , \nScanOut167[6] , 
        \nScanOut167[5] , \nScanOut167[4] , \nScanOut167[3] , \nScanOut167[2] , 
        \nScanOut167[1] , \nScanOut167[0] }), .ScanOut({\nScanOut166[7] , 
        \nScanOut166[6] , \nScanOut166[5] , \nScanOut166[4] , \nScanOut166[3] , 
        \nScanOut166[2] , \nScanOut166[1] , \nScanOut166[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_5[7] , \nOut5_5[6] , \nOut5_5[5] , \nOut5_5[4] , \nOut5_5[3] , 
        \nOut5_5[2] , \nOut5_5[1] , \nOut5_5[0] }), .SouthIn({\nOut5_7[7] , 
        \nOut5_7[6] , \nOut5_7[5] , \nOut5_7[4] , \nOut5_7[3] , \nOut5_7[2] , 
        \nOut5_7[1] , \nOut5_7[0] }), .EastIn({\nOut6_6[7] , \nOut6_6[6] , 
        \nOut6_6[5] , \nOut6_6[4] , \nOut6_6[3] , \nOut6_6[2] , \nOut6_6[1] , 
        \nOut6_6[0] }), .WestIn({\nOut4_6[7] , \nOut4_6[6] , \nOut4_6[5] , 
        \nOut4_6[4] , \nOut4_6[3] , \nOut4_6[2] , \nOut4_6[1] , \nOut4_6[0] }), 
        .Out({\nOut5_6[7] , \nOut5_6[6] , \nOut5_6[5] , \nOut5_6[4] , 
        \nOut5_6[3] , \nOut5_6[2] , \nOut5_6[1] , \nOut5_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_256 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut257[7] , \nScanOut257[6] , 
        \nScanOut257[5] , \nScanOut257[4] , \nScanOut257[3] , \nScanOut257[2] , 
        \nScanOut257[1] , \nScanOut257[0] }), .ScanOut({\nScanOut256[7] , 
        \nScanOut256[6] , \nScanOut256[5] , \nScanOut256[4] , \nScanOut256[3] , 
        \nScanOut256[2] , \nScanOut256[1] , \nScanOut256[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut8_0[7] , \nOut8_0[6] , 
        \nOut8_0[5] , \nOut8_0[4] , \nOut8_0[3] , \nOut8_0[2] , \nOut8_0[1] , 
        \nOut8_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_271 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut272[7] , \nScanOut272[6] , 
        \nScanOut272[5] , \nScanOut272[4] , \nScanOut272[3] , \nScanOut272[2] , 
        \nScanOut272[1] , \nScanOut272[0] }), .ScanOut({\nScanOut271[7] , 
        \nScanOut271[6] , \nScanOut271[5] , \nScanOut271[4] , \nScanOut271[3] , 
        \nScanOut271[2] , \nScanOut271[1] , \nScanOut271[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }), 
        .SouthIn({\nOut8_16[7] , \nOut8_16[6] , \nOut8_16[5] , \nOut8_16[4] , 
        \nOut8_16[3] , \nOut8_16[2] , \nOut8_16[1] , \nOut8_16[0] }), .EastIn(
        {\nOut9_15[7] , \nOut9_15[6] , \nOut9_15[5] , \nOut9_15[4] , 
        \nOut9_15[3] , \nOut9_15[2] , \nOut9_15[1] , \nOut9_15[0] }), .WestIn(
        {\nOut7_15[7] , \nOut7_15[6] , \nOut7_15[5] , \nOut7_15[4] , 
        \nOut7_15[3] , \nOut7_15[2] , \nOut7_15[1] , \nOut7_15[0] }), .Out({
        \nOut8_15[7] , \nOut8_15[6] , \nOut8_15[5] , \nOut8_15[4] , 
        \nOut8_15[3] , \nOut8_15[2] , \nOut8_15[1] , \nOut8_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_460 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut461[7] , \nScanOut461[6] , 
        \nScanOut461[5] , \nScanOut461[4] , \nScanOut461[3] , \nScanOut461[2] , 
        \nScanOut461[1] , \nScanOut461[0] }), .ScanOut({\nScanOut460[7] , 
        \nScanOut460[6] , \nScanOut460[5] , \nScanOut460[4] , \nScanOut460[3] , 
        \nScanOut460[2] , \nScanOut460[1] , \nScanOut460[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_11[7] , \nOut14_11[6] , \nOut14_11[5] , \nOut14_11[4] , 
        \nOut14_11[3] , \nOut14_11[2] , \nOut14_11[1] , \nOut14_11[0] }), 
        .SouthIn({\nOut14_13[7] , \nOut14_13[6] , \nOut14_13[5] , 
        \nOut14_13[4] , \nOut14_13[3] , \nOut14_13[2] , \nOut14_13[1] , 
        \nOut14_13[0] }), .EastIn({\nOut15_12[7] , \nOut15_12[6] , 
        \nOut15_12[5] , \nOut15_12[4] , \nOut15_12[3] , \nOut15_12[2] , 
        \nOut15_12[1] , \nOut15_12[0] }), .WestIn({\nOut13_12[7] , 
        \nOut13_12[6] , \nOut13_12[5] , \nOut13_12[4] , \nOut13_12[3] , 
        \nOut13_12[2] , \nOut13_12[1] , \nOut13_12[0] }), .Out({\nOut14_12[7] , 
        \nOut14_12[6] , \nOut14_12[5] , \nOut14_12[4] , \nOut14_12[3] , 
        \nOut14_12[2] , \nOut14_12[1] , \nOut14_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_812 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut813[7] , \nScanOut813[6] , 
        \nScanOut813[5] , \nScanOut813[4] , \nScanOut813[3] , \nScanOut813[2] , 
        \nScanOut813[1] , \nScanOut813[0] }), .ScanOut({\nScanOut812[7] , 
        \nScanOut812[6] , \nScanOut812[5] , \nScanOut812[4] , \nScanOut812[3] , 
        \nScanOut812[2] , \nScanOut812[1] , \nScanOut812[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_11[7] , \nOut25_11[6] , \nOut25_11[5] , \nOut25_11[4] , 
        \nOut25_11[3] , \nOut25_11[2] , \nOut25_11[1] , \nOut25_11[0] }), 
        .SouthIn({\nOut25_13[7] , \nOut25_13[6] , \nOut25_13[5] , 
        \nOut25_13[4] , \nOut25_13[3] , \nOut25_13[2] , \nOut25_13[1] , 
        \nOut25_13[0] }), .EastIn({\nOut26_12[7] , \nOut26_12[6] , 
        \nOut26_12[5] , \nOut26_12[4] , \nOut26_12[3] , \nOut26_12[2] , 
        \nOut26_12[1] , \nOut26_12[0] }), .WestIn({\nOut24_12[7] , 
        \nOut24_12[6] , \nOut24_12[5] , \nOut24_12[4] , \nOut24_12[3] , 
        \nOut24_12[2] , \nOut24_12[1] , \nOut24_12[0] }), .Out({\nOut25_12[7] , 
        \nOut25_12[6] , \nOut25_12[5] , \nOut25_12[4] , \nOut25_12[3] , 
        \nOut25_12[2] , \nOut25_12[1] , \nOut25_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_982 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut983[7] , \nScanOut983[6] , 
        \nScanOut983[5] , \nScanOut983[4] , \nScanOut983[3] , \nScanOut983[2] , 
        \nScanOut983[1] , \nScanOut983[0] }), .ScanOut({\nScanOut982[7] , 
        \nScanOut982[6] , \nScanOut982[5] , \nScanOut982[4] , \nScanOut982[3] , 
        \nScanOut982[2] , \nScanOut982[1] , \nScanOut982[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_21[7] , \nOut30_21[6] , \nOut30_21[5] , \nOut30_21[4] , 
        \nOut30_21[3] , \nOut30_21[2] , \nOut30_21[1] , \nOut30_21[0] }), 
        .SouthIn({\nOut30_23[7] , \nOut30_23[6] , \nOut30_23[5] , 
        \nOut30_23[4] , \nOut30_23[3] , \nOut30_23[2] , \nOut30_23[1] , 
        \nOut30_23[0] }), .EastIn({\nOut31_22[7] , \nOut31_22[6] , 
        \nOut31_22[5] , \nOut31_22[4] , \nOut31_22[3] , \nOut31_22[2] , 
        \nOut31_22[1] , \nOut31_22[0] }), .WestIn({\nOut29_22[7] , 
        \nOut29_22[6] , \nOut29_22[5] , \nOut29_22[4] , \nOut29_22[3] , 
        \nOut29_22[2] , \nOut29_22[1] , \nOut29_22[0] }), .Out({\nOut30_22[7] , 
        \nOut30_22[6] , \nOut30_22[5] , \nOut30_22[4] , \nOut30_22[3] , 
        \nOut30_22[2] , \nOut30_22[1] , \nOut30_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_447 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut448[7] , \nScanOut448[6] , 
        \nScanOut448[5] , \nScanOut448[4] , \nScanOut448[3] , \nScanOut448[2] , 
        \nScanOut448[1] , \nScanOut448[0] }), .ScanOut({\nScanOut447[7] , 
        \nScanOut447[6] , \nScanOut447[5] , \nScanOut447[4] , \nScanOut447[3] , 
        \nScanOut447[2] , \nScanOut447[1] , \nScanOut447[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut13_31[7] , \nOut13_31[6] , 
        \nOut13_31[5] , \nOut13_31[4] , \nOut13_31[3] , \nOut13_31[2] , 
        \nOut13_31[1] , \nOut13_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_835 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut836[7] , \nScanOut836[6] , 
        \nScanOut836[5] , \nScanOut836[4] , \nScanOut836[3] , \nScanOut836[2] , 
        \nScanOut836[1] , \nScanOut836[0] }), .ScanOut({\nScanOut835[7] , 
        \nScanOut835[6] , \nScanOut835[5] , \nScanOut835[4] , \nScanOut835[3] , 
        \nScanOut835[2] , \nScanOut835[1] , \nScanOut835[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_2[7] , \nOut26_2[6] , \nOut26_2[5] , \nOut26_2[4] , 
        \nOut26_2[3] , \nOut26_2[2] , \nOut26_2[1] , \nOut26_2[0] }), 
        .SouthIn({\nOut26_4[7] , \nOut26_4[6] , \nOut26_4[5] , \nOut26_4[4] , 
        \nOut26_4[3] , \nOut26_4[2] , \nOut26_4[1] , \nOut26_4[0] }), .EastIn(
        {\nOut27_3[7] , \nOut27_3[6] , \nOut27_3[5] , \nOut27_3[4] , 
        \nOut27_3[3] , \nOut27_3[2] , \nOut27_3[1] , \nOut27_3[0] }), .WestIn(
        {\nOut25_3[7] , \nOut25_3[6] , \nOut25_3[5] , \nOut25_3[4] , 
        \nOut25_3[3] , \nOut25_3[2] , \nOut25_3[1] , \nOut25_3[0] }), .Out({
        \nOut26_3[7] , \nOut26_3[6] , \nOut26_3[5] , \nOut26_3[4] , 
        \nOut26_3[3] , \nOut26_3[2] , \nOut26_3[1] , \nOut26_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_777 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut778[7] , \nScanOut778[6] , 
        \nScanOut778[5] , \nScanOut778[4] , \nScanOut778[3] , \nScanOut778[2] , 
        \nScanOut778[1] , \nScanOut778[0] }), .ScanOut({\nScanOut777[7] , 
        \nScanOut777[6] , \nScanOut777[5] , \nScanOut777[4] , \nScanOut777[3] , 
        \nScanOut777[2] , \nScanOut777[1] , \nScanOut777[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_8[7] , \nOut24_8[6] , \nOut24_8[5] , \nOut24_8[4] , 
        \nOut24_8[3] , \nOut24_8[2] , \nOut24_8[1] , \nOut24_8[0] }), 
        .SouthIn({\nOut24_10[7] , \nOut24_10[6] , \nOut24_10[5] , 
        \nOut24_10[4] , \nOut24_10[3] , \nOut24_10[2] , \nOut24_10[1] , 
        \nOut24_10[0] }), .EastIn({\nOut25_9[7] , \nOut25_9[6] , \nOut25_9[5] , 
        \nOut25_9[4] , \nOut25_9[3] , \nOut25_9[2] , \nOut25_9[1] , 
        \nOut25_9[0] }), .WestIn({\nOut23_9[7] , \nOut23_9[6] , \nOut23_9[5] , 
        \nOut23_9[4] , \nOut23_9[3] , \nOut23_9[2] , \nOut23_9[1] , 
        \nOut23_9[0] }), .Out({\nOut24_9[7] , \nOut24_9[6] , \nOut24_9[5] , 
        \nOut24_9[4] , \nOut24_9[3] , \nOut24_9[2] , \nOut24_9[1] , 
        \nOut24_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_899 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut900[7] , \nScanOut900[6] , 
        \nScanOut900[5] , \nScanOut900[4] , \nScanOut900[3] , \nScanOut900[2] , 
        \nScanOut900[1] , \nScanOut900[0] }), .ScanOut({\nScanOut899[7] , 
        \nScanOut899[6] , \nScanOut899[5] , \nScanOut899[4] , \nScanOut899[3] , 
        \nScanOut899[2] , \nScanOut899[1] , \nScanOut899[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_2[7] , \nOut28_2[6] , \nOut28_2[5] , \nOut28_2[4] , 
        \nOut28_2[3] , \nOut28_2[2] , \nOut28_2[1] , \nOut28_2[0] }), 
        .SouthIn({\nOut28_4[7] , \nOut28_4[6] , \nOut28_4[5] , \nOut28_4[4] , 
        \nOut28_4[3] , \nOut28_4[2] , \nOut28_4[1] , \nOut28_4[0] }), .EastIn(
        {\nOut29_3[7] , \nOut29_3[6] , \nOut29_3[5] , \nOut29_3[4] , 
        \nOut29_3[3] , \nOut29_3[2] , \nOut29_3[1] , \nOut29_3[0] }), .WestIn(
        {\nOut27_3[7] , \nOut27_3[6] , \nOut27_3[5] , \nOut27_3[4] , 
        \nOut27_3[3] , \nOut27_3[2] , \nOut27_3[1] , \nOut27_3[0] }), .Out({
        \nOut28_3[7] , \nOut28_3[6] , \nOut28_3[5] , \nOut28_3[4] , 
        \nOut28_3[3] , \nOut28_3[2] , \nOut28_3[1] , \nOut28_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_909 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut910[7] , \nScanOut910[6] , 
        \nScanOut910[5] , \nScanOut910[4] , \nScanOut910[3] , \nScanOut910[2] , 
        \nScanOut910[1] , \nScanOut910[0] }), .ScanOut({\nScanOut909[7] , 
        \nScanOut909[6] , \nScanOut909[5] , \nScanOut909[4] , \nScanOut909[3] , 
        \nScanOut909[2] , \nScanOut909[1] , \nScanOut909[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_12[7] , \nOut28_12[6] , \nOut28_12[5] , \nOut28_12[4] , 
        \nOut28_12[3] , \nOut28_12[2] , \nOut28_12[1] , \nOut28_12[0] }), 
        .SouthIn({\nOut28_14[7] , \nOut28_14[6] , \nOut28_14[5] , 
        \nOut28_14[4] , \nOut28_14[3] , \nOut28_14[2] , \nOut28_14[1] , 
        \nOut28_14[0] }), .EastIn({\nOut29_13[7] , \nOut29_13[6] , 
        \nOut29_13[5] , \nOut29_13[4] , \nOut29_13[3] , \nOut29_13[2] , 
        \nOut29_13[1] , \nOut29_13[0] }), .WestIn({\nOut27_13[7] , 
        \nOut27_13[6] , \nOut27_13[5] , \nOut27_13[4] , \nOut27_13[3] , 
        \nOut27_13[2] , \nOut27_13[1] , \nOut27_13[0] }), .Out({\nOut28_13[7] , 
        \nOut28_13[6] , \nOut28_13[5] , \nOut28_13[4] , \nOut28_13[3] , 
        \nOut28_13[2] , \nOut28_13[1] , \nOut28_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_356 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut357[7] , \nScanOut357[6] , 
        \nScanOut357[5] , \nScanOut357[4] , \nScanOut357[3] , \nScanOut357[2] , 
        \nScanOut357[1] , \nScanOut357[0] }), .ScanOut({\nScanOut356[7] , 
        \nScanOut356[6] , \nScanOut356[5] , \nScanOut356[4] , \nScanOut356[3] , 
        \nScanOut356[2] , \nScanOut356[1] , \nScanOut356[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }), 
        .SouthIn({\nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }), .EastIn(
        {\nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }), .WestIn(
        {\nOut10_4[7] , \nOut10_4[6] , \nOut10_4[5] , \nOut10_4[4] , 
        \nOut10_4[3] , \nOut10_4[2] , \nOut10_4[1] , \nOut10_4[0] }), .Out({
        \nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_547 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut548[7] , \nScanOut548[6] , 
        \nScanOut548[5] , \nScanOut548[4] , \nScanOut548[3] , \nScanOut548[2] , 
        \nScanOut548[1] , \nScanOut548[0] }), .ScanOut({\nScanOut547[7] , 
        \nScanOut547[6] , \nScanOut547[5] , \nScanOut547[4] , \nScanOut547[3] , 
        \nScanOut547[2] , \nScanOut547[1] , \nScanOut547[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_2[7] , \nOut17_2[6] , \nOut17_2[5] , \nOut17_2[4] , 
        \nOut17_2[3] , \nOut17_2[2] , \nOut17_2[1] , \nOut17_2[0] }), 
        .SouthIn({\nOut17_4[7] , \nOut17_4[6] , \nOut17_4[5] , \nOut17_4[4] , 
        \nOut17_4[3] , \nOut17_4[2] , \nOut17_4[1] , \nOut17_4[0] }), .EastIn(
        {\nOut18_3[7] , \nOut18_3[6] , \nOut18_3[5] , \nOut18_3[4] , 
        \nOut18_3[3] , \nOut18_3[2] , \nOut18_3[1] , \nOut18_3[0] }), .WestIn(
        {\nOut16_3[7] , \nOut16_3[6] , \nOut16_3[5] , \nOut16_3[4] , 
        \nOut16_3[3] , \nOut16_3[2] , \nOut16_3[1] , \nOut16_3[0] }), .Out({
        \nOut17_3[7] , \nOut17_3[6] , \nOut17_3[5] , \nOut17_3[4] , 
        \nOut17_3[3] , \nOut17_3[2] , \nOut17_3[1] , \nOut17_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_677 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut678[7] , \nScanOut678[6] , 
        \nScanOut678[5] , \nScanOut678[4] , \nScanOut678[3] , \nScanOut678[2] , 
        \nScanOut678[1] , \nScanOut678[0] }), .ScanOut({\nScanOut677[7] , 
        \nScanOut677[6] , \nScanOut677[5] , \nScanOut677[4] , \nScanOut677[3] , 
        \nScanOut677[2] , \nScanOut677[1] , \nScanOut677[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_4[7] , \nOut21_4[6] , \nOut21_4[5] , \nOut21_4[4] , 
        \nOut21_4[3] , \nOut21_4[2] , \nOut21_4[1] , \nOut21_4[0] }), 
        .SouthIn({\nOut21_6[7] , \nOut21_6[6] , \nOut21_6[5] , \nOut21_6[4] , 
        \nOut21_6[3] , \nOut21_6[2] , \nOut21_6[1] , \nOut21_6[0] }), .EastIn(
        {\nOut22_5[7] , \nOut22_5[6] , \nOut22_5[5] , \nOut22_5[4] , 
        \nOut22_5[3] , \nOut22_5[2] , \nOut22_5[1] , \nOut22_5[0] }), .WestIn(
        {\nOut20_5[7] , \nOut20_5[6] , \nOut20_5[5] , \nOut20_5[4] , 
        \nOut20_5[3] , \nOut20_5[2] , \nOut20_5[1] , \nOut20_5[0] }), .Out({
        \nOut21_5[7] , \nOut21_5[6] , \nOut21_5[5] , \nOut21_5[4] , 
        \nOut21_5[3] , \nOut21_5[2] , \nOut21_5[1] , \nOut21_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_371 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut372[7] , \nScanOut372[6] , 
        \nScanOut372[5] , \nScanOut372[4] , \nScanOut372[3] , \nScanOut372[2] , 
        \nScanOut372[1] , \nScanOut372[0] }), .ScanOut({\nScanOut371[7] , 
        \nScanOut371[6] , \nScanOut371[5] , \nScanOut371[4] , \nScanOut371[3] , 
        \nScanOut371[2] , \nScanOut371[1] , \nScanOut371[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_18[7] , \nOut11_18[6] , \nOut11_18[5] , \nOut11_18[4] , 
        \nOut11_18[3] , \nOut11_18[2] , \nOut11_18[1] , \nOut11_18[0] }), 
        .SouthIn({\nOut11_20[7] , \nOut11_20[6] , \nOut11_20[5] , 
        \nOut11_20[4] , \nOut11_20[3] , \nOut11_20[2] , \nOut11_20[1] , 
        \nOut11_20[0] }), .EastIn({\nOut12_19[7] , \nOut12_19[6] , 
        \nOut12_19[5] , \nOut12_19[4] , \nOut12_19[3] , \nOut12_19[2] , 
        \nOut12_19[1] , \nOut12_19[0] }), .WestIn({\nOut10_19[7] , 
        \nOut10_19[6] , \nOut10_19[5] , \nOut10_19[4] , \nOut10_19[3] , 
        \nOut10_19[2] , \nOut10_19[1] , \nOut10_19[0] }), .Out({\nOut11_19[7] , 
        \nOut11_19[6] , \nOut11_19[5] , \nOut11_19[4] , \nOut11_19[3] , 
        \nOut11_19[2] , \nOut11_19[1] , \nOut11_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_935 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut936[7] , \nScanOut936[6] , 
        \nScanOut936[5] , \nScanOut936[4] , \nScanOut936[3] , \nScanOut936[2] , 
        \nScanOut936[1] , \nScanOut936[0] }), .ScanOut({\nScanOut935[7] , 
        \nScanOut935[6] , \nScanOut935[5] , \nScanOut935[4] , \nScanOut935[3] , 
        \nScanOut935[2] , \nScanOut935[1] , \nScanOut935[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_6[7] , \nOut29_6[6] , \nOut29_6[5] , \nOut29_6[4] , 
        \nOut29_6[3] , \nOut29_6[2] , \nOut29_6[1] , \nOut29_6[0] }), 
        .SouthIn({\nOut29_8[7] , \nOut29_8[6] , \nOut29_8[5] , \nOut29_8[4] , 
        \nOut29_8[3] , \nOut29_8[2] , \nOut29_8[1] , \nOut29_8[0] }), .EastIn(
        {\nOut30_7[7] , \nOut30_7[6] , \nOut30_7[5] , \nOut30_7[4] , 
        \nOut30_7[3] , \nOut30_7[2] , \nOut30_7[1] , \nOut30_7[0] }), .WestIn(
        {\nOut28_7[7] , \nOut28_7[6] , \nOut28_7[5] , \nOut28_7[4] , 
        \nOut28_7[3] , \nOut28_7[2] , \nOut28_7[1] , \nOut28_7[0] }), .Out({
        \nOut29_7[7] , \nOut29_7[6] , \nOut29_7[5] , \nOut29_7[4] , 
        \nOut29_7[3] , \nOut29_7[2] , \nOut29_7[1] , \nOut29_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_560 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut561[7] , \nScanOut561[6] , 
        \nScanOut561[5] , \nScanOut561[4] , \nScanOut561[3] , \nScanOut561[2] , 
        \nScanOut561[1] , \nScanOut561[0] }), .ScanOut({\nScanOut560[7] , 
        \nScanOut560[6] , \nScanOut560[5] , \nScanOut560[4] , \nScanOut560[3] , 
        \nScanOut560[2] , \nScanOut560[1] , \nScanOut560[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_15[7] , \nOut17_15[6] , \nOut17_15[5] , \nOut17_15[4] , 
        \nOut17_15[3] , \nOut17_15[2] , \nOut17_15[1] , \nOut17_15[0] }), 
        .SouthIn({\nOut17_17[7] , \nOut17_17[6] , \nOut17_17[5] , 
        \nOut17_17[4] , \nOut17_17[3] , \nOut17_17[2] , \nOut17_17[1] , 
        \nOut17_17[0] }), .EastIn({\nOut18_16[7] , \nOut18_16[6] , 
        \nOut18_16[5] , \nOut18_16[4] , \nOut18_16[3] , \nOut18_16[2] , 
        \nOut18_16[1] , \nOut18_16[0] }), .WestIn({\nOut16_16[7] , 
        \nOut16_16[6] , \nOut16_16[5] , \nOut16_16[4] , \nOut16_16[3] , 
        \nOut16_16[2] , \nOut16_16[1] , \nOut16_16[0] }), .Out({\nOut17_16[7] , 
        \nOut17_16[6] , \nOut17_16[5] , \nOut17_16[4] , \nOut17_16[3] , 
        \nOut17_16[2] , \nOut17_16[1] , \nOut17_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_882 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut883[7] , \nScanOut883[6] , 
        \nScanOut883[5] , \nScanOut883[4] , \nScanOut883[3] , \nScanOut883[2] , 
        \nScanOut883[1] , \nScanOut883[0] }), .ScanOut({\nScanOut882[7] , 
        \nScanOut882[6] , \nScanOut882[5] , \nScanOut882[4] , \nScanOut882[3] , 
        \nScanOut882[2] , \nScanOut882[1] , \nScanOut882[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_17[7] , \nOut27_17[6] , \nOut27_17[5] , \nOut27_17[4] , 
        \nOut27_17[3] , \nOut27_17[2] , \nOut27_17[1] , \nOut27_17[0] }), 
        .SouthIn({\nOut27_19[7] , \nOut27_19[6] , \nOut27_19[5] , 
        \nOut27_19[4] , \nOut27_19[3] , \nOut27_19[2] , \nOut27_19[1] , 
        \nOut27_19[0] }), .EastIn({\nOut28_18[7] , \nOut28_18[6] , 
        \nOut28_18[5] , \nOut28_18[4] , \nOut28_18[3] , \nOut28_18[2] , 
        \nOut28_18[1] , \nOut28_18[0] }), .WestIn({\nOut26_18[7] , 
        \nOut26_18[6] , \nOut26_18[5] , \nOut26_18[4] , \nOut26_18[3] , 
        \nOut26_18[2] , \nOut26_18[1] , \nOut26_18[0] }), .Out({\nOut27_18[7] , 
        \nOut27_18[6] , \nOut27_18[5] , \nOut27_18[4] , \nOut27_18[3] , 
        \nOut27_18[2] , \nOut27_18[1] , \nOut27_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_912 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut913[7] , \nScanOut913[6] , 
        \nScanOut913[5] , \nScanOut913[4] , \nScanOut913[3] , \nScanOut913[2] , 
        \nScanOut913[1] , \nScanOut913[0] }), .ScanOut({\nScanOut912[7] , 
        \nScanOut912[6] , \nScanOut912[5] , \nScanOut912[4] , \nScanOut912[3] , 
        \nScanOut912[2] , \nScanOut912[1] , \nScanOut912[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_15[7] , \nOut28_15[6] , \nOut28_15[5] , \nOut28_15[4] , 
        \nOut28_15[3] , \nOut28_15[2] , \nOut28_15[1] , \nOut28_15[0] }), 
        .SouthIn({\nOut28_17[7] , \nOut28_17[6] , \nOut28_17[5] , 
        \nOut28_17[4] , \nOut28_17[3] , \nOut28_17[2] , \nOut28_17[1] , 
        \nOut28_17[0] }), .EastIn({\nOut29_16[7] , \nOut29_16[6] , 
        \nOut29_16[5] , \nOut29_16[4] , \nOut29_16[3] , \nOut29_16[2] , 
        \nOut29_16[1] , \nOut29_16[0] }), .WestIn({\nOut27_16[7] , 
        \nOut27_16[6] , \nOut27_16[5] , \nOut27_16[4] , \nOut27_16[3] , 
        \nOut27_16[2] , \nOut27_16[1] , \nOut27_16[0] }), .Out({\nOut28_16[7] , 
        \nOut28_16[6] , \nOut28_16[5] , \nOut28_16[4] , \nOut28_16[3] , 
        \nOut28_16[2] , \nOut28_16[1] , \nOut28_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_650 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut651[7] , \nScanOut651[6] , 
        \nScanOut651[5] , \nScanOut651[4] , \nScanOut651[3] , \nScanOut651[2] , 
        \nScanOut651[1] , \nScanOut651[0] }), .ScanOut({\nScanOut650[7] , 
        \nScanOut650[6] , \nScanOut650[5] , \nScanOut650[4] , \nScanOut650[3] , 
        \nScanOut650[2] , \nScanOut650[1] , \nScanOut650[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_9[7] , \nOut20_9[6] , \nOut20_9[5] , \nOut20_9[4] , 
        \nOut20_9[3] , \nOut20_9[2] , \nOut20_9[1] , \nOut20_9[0] }), 
        .SouthIn({\nOut20_11[7] , \nOut20_11[6] , \nOut20_11[5] , 
        \nOut20_11[4] , \nOut20_11[3] , \nOut20_11[2] , \nOut20_11[1] , 
        \nOut20_11[0] }), .EastIn({\nOut21_10[7] , \nOut21_10[6] , 
        \nOut21_10[5] , \nOut21_10[4] , \nOut21_10[3] , \nOut21_10[2] , 
        \nOut21_10[1] , \nOut21_10[0] }), .WestIn({\nOut19_10[7] , 
        \nOut19_10[6] , \nOut19_10[5] , \nOut19_10[4] , \nOut19_10[3] , 
        \nOut19_10[2] , \nOut19_10[1] , \nOut19_10[0] }), .Out({\nOut20_10[7] , 
        \nOut20_10[6] , \nOut20_10[5] , \nOut20_10[4] , \nOut20_10[3] , 
        \nOut20_10[2] , \nOut20_10[1] , \nOut20_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_22 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut23[7] , \nScanOut23[6] , 
        \nScanOut23[5] , \nScanOut23[4] , \nScanOut23[3] , \nScanOut23[2] , 
        \nScanOut23[1] , \nScanOut23[0] }), .ScanOut({\nScanOut22[7] , 
        \nScanOut22[6] , \nScanOut22[5] , \nScanOut22[4] , \nScanOut22[3] , 
        \nScanOut22[2] , \nScanOut22[1] , \nScanOut22[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_22[7] , \nOut0_22[6] , 
        \nOut0_22[5] , \nOut0_22[4] , \nOut0_22[3] , \nOut0_22[2] , 
        \nOut0_22[1] , \nOut0_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_39 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut40[7] , \nScanOut40[6] , 
        \nScanOut40[5] , \nScanOut40[4] , \nScanOut40[3] , \nScanOut40[2] , 
        \nScanOut40[1] , \nScanOut40[0] }), .ScanOut({\nScanOut39[7] , 
        \nScanOut39[6] , \nScanOut39[5] , \nScanOut39[4] , \nScanOut39[3] , 
        \nScanOut39[2] , \nScanOut39[1] , \nScanOut39[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , \nOut1_6[4] , \nOut1_6[3] , 
        \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }), .SouthIn({\nOut1_8[7] , 
        \nOut1_8[6] , \nOut1_8[5] , \nOut1_8[4] , \nOut1_8[3] , \nOut1_8[2] , 
        \nOut1_8[1] , \nOut1_8[0] }), .EastIn({\nOut2_7[7] , \nOut2_7[6] , 
        \nOut2_7[5] , \nOut2_7[4] , \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , 
        \nOut2_7[0] }), .WestIn({\nOut0_7[7] , \nOut0_7[6] , \nOut0_7[5] , 
        \nOut0_7[4] , \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , \nOut0_7[0] }), 
        .Out({\nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , \nOut1_7[4] , 
        \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_87 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut88[7] , \nScanOut88[6] , 
        \nScanOut88[5] , \nScanOut88[4] , \nScanOut88[3] , \nScanOut88[2] , 
        \nScanOut88[1] , \nScanOut88[0] }), .ScanOut({\nScanOut87[7] , 
        \nScanOut87[6] , \nScanOut87[5] , \nScanOut87[4] , \nScanOut87[3] , 
        \nScanOut87[2] , \nScanOut87[1] , \nScanOut87[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_22[7] , \nOut2_22[6] , \nOut2_22[5] , \nOut2_22[4] , 
        \nOut2_22[3] , \nOut2_22[2] , \nOut2_22[1] , \nOut2_22[0] }), 
        .SouthIn({\nOut2_24[7] , \nOut2_24[6] , \nOut2_24[5] , \nOut2_24[4] , 
        \nOut2_24[3] , \nOut2_24[2] , \nOut2_24[1] , \nOut2_24[0] }), .EastIn(
        {\nOut3_23[7] , \nOut3_23[6] , \nOut3_23[5] , \nOut3_23[4] , 
        \nOut3_23[3] , \nOut3_23[2] , \nOut3_23[1] , \nOut3_23[0] }), .WestIn(
        {\nOut1_23[7] , \nOut1_23[6] , \nOut1_23[5] , \nOut1_23[4] , 
        \nOut1_23[3] , \nOut1_23[2] , \nOut1_23[1] , \nOut1_23[0] }), .Out({
        \nOut2_23[7] , \nOut2_23[6] , \nOut2_23[5] , \nOut2_23[4] , 
        \nOut2_23[3] , \nOut2_23[2] , \nOut2_23[1] , \nOut2_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_113 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut114[7] , \nScanOut114[6] , 
        \nScanOut114[5] , \nScanOut114[4] , \nScanOut114[3] , \nScanOut114[2] , 
        \nScanOut114[1] , \nScanOut114[0] }), .ScanOut({\nScanOut113[7] , 
        \nScanOut113[6] , \nScanOut113[5] , \nScanOut113[4] , \nScanOut113[3] , 
        \nScanOut113[2] , \nScanOut113[1] , \nScanOut113[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_16[7] , \nOut3_16[6] , \nOut3_16[5] , \nOut3_16[4] , 
        \nOut3_16[3] , \nOut3_16[2] , \nOut3_16[1] , \nOut3_16[0] }), 
        .SouthIn({\nOut3_18[7] , \nOut3_18[6] , \nOut3_18[5] , \nOut3_18[4] , 
        \nOut3_18[3] , \nOut3_18[2] , \nOut3_18[1] , \nOut3_18[0] }), .EastIn(
        {\nOut4_17[7] , \nOut4_17[6] , \nOut4_17[5] , \nOut4_17[4] , 
        \nOut4_17[3] , \nOut4_17[2] , \nOut4_17[1] , \nOut4_17[0] }), .WestIn(
        {\nOut2_17[7] , \nOut2_17[6] , \nOut2_17[5] , \nOut2_17[4] , 
        \nOut2_17[3] , \nOut2_17[2] , \nOut2_17[1] , \nOut2_17[0] }), .Out({
        \nOut3_17[7] , \nOut3_17[6] , \nOut3_17[5] , \nOut3_17[4] , 
        \nOut3_17[3] , \nOut3_17[2] , \nOut3_17[1] , \nOut3_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_134 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut135[7] , \nScanOut135[6] , 
        \nScanOut135[5] , \nScanOut135[4] , \nScanOut135[3] , \nScanOut135[2] , 
        \nScanOut135[1] , \nScanOut135[0] }), .ScanOut({\nScanOut134[7] , 
        \nScanOut134[6] , \nScanOut134[5] , \nScanOut134[4] , \nScanOut134[3] , 
        \nScanOut134[2] , \nScanOut134[1] , \nScanOut134[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_5[7] , \nOut4_5[6] , \nOut4_5[5] , \nOut4_5[4] , \nOut4_5[3] , 
        \nOut4_5[2] , \nOut4_5[1] , \nOut4_5[0] }), .SouthIn({\nOut4_7[7] , 
        \nOut4_7[6] , \nOut4_7[5] , \nOut4_7[4] , \nOut4_7[3] , \nOut4_7[2] , 
        \nOut4_7[1] , \nOut4_7[0] }), .EastIn({\nOut5_6[7] , \nOut5_6[6] , 
        \nOut5_6[5] , \nOut5_6[4] , \nOut5_6[3] , \nOut5_6[2] , \nOut5_6[1] , 
        \nOut5_6[0] }), .WestIn({\nOut3_6[7] , \nOut3_6[6] , \nOut3_6[5] , 
        \nOut3_6[4] , \nOut3_6[3] , \nOut3_6[2] , \nOut3_6[1] , \nOut3_6[0] }), 
        .Out({\nOut4_6[7] , \nOut4_6[6] , \nOut4_6[5] , \nOut4_6[4] , 
        \nOut4_6[3] , \nOut4_6[2] , \nOut4_6[1] , \nOut4_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_204 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut205[7] , \nScanOut205[6] , 
        \nScanOut205[5] , \nScanOut205[4] , \nScanOut205[3] , \nScanOut205[2] , 
        \nScanOut205[1] , \nScanOut205[0] }), .ScanOut({\nScanOut204[7] , 
        \nScanOut204[6] , \nScanOut204[5] , \nScanOut204[4] , \nScanOut204[3] , 
        \nScanOut204[2] , \nScanOut204[1] , \nScanOut204[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_11[7] , \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , 
        \nOut6_11[3] , \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }), 
        .SouthIn({\nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }), .EastIn(
        {\nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }), .WestIn(
        {\nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }), .Out({
        \nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_809 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut810[7] , \nScanOut810[6] , 
        \nScanOut810[5] , \nScanOut810[4] , \nScanOut810[3] , \nScanOut810[2] , 
        \nScanOut810[1] , \nScanOut810[0] }), .ScanOut({\nScanOut809[7] , 
        \nScanOut809[6] , \nScanOut809[5] , \nScanOut809[4] , \nScanOut809[3] , 
        \nScanOut809[2] , \nScanOut809[1] , \nScanOut809[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_8[7] , \nOut25_8[6] , \nOut25_8[5] , \nOut25_8[4] , 
        \nOut25_8[3] , \nOut25_8[2] , \nOut25_8[1] , \nOut25_8[0] }), 
        .SouthIn({\nOut25_10[7] , \nOut25_10[6] , \nOut25_10[5] , 
        \nOut25_10[4] , \nOut25_10[3] , \nOut25_10[2] , \nOut25_10[1] , 
        \nOut25_10[0] }), .EastIn({\nOut26_9[7] , \nOut26_9[6] , \nOut26_9[5] , 
        \nOut26_9[4] , \nOut26_9[3] , \nOut26_9[2] , \nOut26_9[1] , 
        \nOut26_9[0] }), .WestIn({\nOut24_9[7] , \nOut24_9[6] , \nOut24_9[5] , 
        \nOut24_9[4] , \nOut24_9[3] , \nOut24_9[2] , \nOut24_9[1] , 
        \nOut24_9[0] }), .Out({\nOut25_9[7] , \nOut25_9[6] , \nOut25_9[5] , 
        \nOut25_9[4] , \nOut25_9[3] , \nOut25_9[2] , \nOut25_9[1] , 
        \nOut25_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_999 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1000[7] , \nScanOut1000[6] , 
        \nScanOut1000[5] , \nScanOut1000[4] , \nScanOut1000[3] , 
        \nScanOut1000[2] , \nScanOut1000[1] , \nScanOut1000[0] }), .ScanOut({
        \nScanOut999[7] , \nScanOut999[6] , \nScanOut999[5] , \nScanOut999[4] , 
        \nScanOut999[3] , \nScanOut999[2] , \nScanOut999[1] , \nScanOut999[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Out({\nOut31_7[7] , 
        \nOut31_7[6] , \nOut31_7[5] , \nOut31_7[4] , \nOut31_7[3] , 
        \nOut31_7[2] , \nOut31_7[1] , \nOut31_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_394 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut395[7] , \nScanOut395[6] , 
        \nScanOut395[5] , \nScanOut395[4] , \nScanOut395[3] , \nScanOut395[2] , 
        \nScanOut395[1] , \nScanOut395[0] }), .ScanOut({\nScanOut394[7] , 
        \nScanOut394[6] , \nScanOut394[5] , \nScanOut394[4] , \nScanOut394[3] , 
        \nScanOut394[2] , \nScanOut394[1] , \nScanOut394[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , \nOut12_9[4] , 
        \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , \nOut12_9[0] }), 
        .SouthIn({\nOut12_11[7] , \nOut12_11[6] , \nOut12_11[5] , 
        \nOut12_11[4] , \nOut12_11[3] , \nOut12_11[2] , \nOut12_11[1] , 
        \nOut12_11[0] }), .EastIn({\nOut13_10[7] , \nOut13_10[6] , 
        \nOut13_10[5] , \nOut13_10[4] , \nOut13_10[3] , \nOut13_10[2] , 
        \nOut13_10[1] , \nOut13_10[0] }), .WestIn({\nOut11_10[7] , 
        \nOut11_10[6] , \nOut11_10[5] , \nOut11_10[4] , \nOut11_10[3] , 
        \nOut11_10[2] , \nOut11_10[1] , \nOut11_10[0] }), .Out({\nOut12_10[7] , 
        \nOut12_10[6] , \nOut12_10[5] , \nOut12_10[4] , \nOut12_10[3] , 
        \nOut12_10[2] , \nOut12_10[1] , \nOut12_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_585 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut586[7] , \nScanOut586[6] , 
        \nScanOut586[5] , \nScanOut586[4] , \nScanOut586[3] , \nScanOut586[2] , 
        \nScanOut586[1] , \nScanOut586[0] }), .ScanOut({\nScanOut585[7] , 
        \nScanOut585[6] , \nScanOut585[5] , \nScanOut585[4] , \nScanOut585[3] , 
        \nScanOut585[2] , \nScanOut585[1] , \nScanOut585[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_8[7] , \nOut18_8[6] , \nOut18_8[5] , \nOut18_8[4] , 
        \nOut18_8[3] , \nOut18_8[2] , \nOut18_8[1] , \nOut18_8[0] }), 
        .SouthIn({\nOut18_10[7] , \nOut18_10[6] , \nOut18_10[5] , 
        \nOut18_10[4] , \nOut18_10[3] , \nOut18_10[2] , \nOut18_10[1] , 
        \nOut18_10[0] }), .EastIn({\nOut19_9[7] , \nOut19_9[6] , \nOut19_9[5] , 
        \nOut19_9[4] , \nOut19_9[3] , \nOut19_9[2] , \nOut19_9[1] , 
        \nOut19_9[0] }), .WestIn({\nOut17_9[7] , \nOut17_9[6] , \nOut17_9[5] , 
        \nOut17_9[4] , \nOut17_9[3] , \nOut17_9[2] , \nOut17_9[1] , 
        \nOut17_9[0] }), .Out({\nOut18_9[7] , \nOut18_9[6] , \nOut18_9[5] , 
        \nOut18_9[4] , \nOut18_9[3] , \nOut18_9[2] , \nOut18_9[1] , 
        \nOut18_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_415 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut416[7] , \nScanOut416[6] , 
        \nScanOut416[5] , \nScanOut416[4] , \nScanOut416[3] , \nScanOut416[2] , 
        \nScanOut416[1] , \nScanOut416[0] }), .ScanOut({\nScanOut415[7] , 
        \nScanOut415[6] , \nScanOut415[5] , \nScanOut415[4] , \nScanOut415[3] , 
        \nScanOut415[2] , \nScanOut415[1] , \nScanOut415[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut12_31[7] , \nOut12_31[6] , 
        \nOut12_31[5] , \nOut12_31[4] , \nOut12_31[3] , \nOut12_31[2] , 
        \nOut12_31[1] , \nOut12_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_867 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut868[7] , \nScanOut868[6] , 
        \nScanOut868[5] , \nScanOut868[4] , \nScanOut868[3] , \nScanOut868[2] , 
        \nScanOut868[1] , \nScanOut868[0] }), .ScanOut({\nScanOut867[7] , 
        \nScanOut867[6] , \nScanOut867[5] , \nScanOut867[4] , \nScanOut867[3] , 
        \nScanOut867[2] , \nScanOut867[1] , \nScanOut867[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_2[7] , \nOut27_2[6] , \nOut27_2[5] , \nOut27_2[4] , 
        \nOut27_2[3] , \nOut27_2[2] , \nOut27_2[1] , \nOut27_2[0] }), 
        .SouthIn({\nOut27_4[7] , \nOut27_4[6] , \nOut27_4[5] , \nOut27_4[4] , 
        \nOut27_4[3] , \nOut27_4[2] , \nOut27_4[1] , \nOut27_4[0] }), .EastIn(
        {\nOut28_3[7] , \nOut28_3[6] , \nOut28_3[5] , \nOut28_3[4] , 
        \nOut28_3[3] , \nOut28_3[2] , \nOut28_3[1] , \nOut28_3[0] }), .WestIn(
        {\nOut26_3[7] , \nOut26_3[6] , \nOut26_3[5] , \nOut26_3[4] , 
        \nOut26_3[3] , \nOut26_3[2] , \nOut26_3[1] , \nOut26_3[0] }), .Out({
        \nOut27_3[7] , \nOut27_3[6] , \nOut27_3[5] , \nOut27_3[4] , 
        \nOut27_3[3] , \nOut27_3[2] , \nOut27_3[1] , \nOut27_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1023 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1024[7] , \nScanOut1024[6] , 
        \nScanOut1024[5] , \nScanOut1024[4] , \nScanOut1024[3] , 
        \nScanOut1024[2] , \nScanOut1024[1] , \nScanOut1024[0] }), .ScanOut({
        \nScanOut1023[7] , \nScanOut1023[6] , \nScanOut1023[5] , 
        \nScanOut1023[4] , \nScanOut1023[3] , \nScanOut1023[2] , 
        \nScanOut1023[1] , \nScanOut1023[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_692 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut693[7] , \nScanOut693[6] , 
        \nScanOut693[5] , \nScanOut693[4] , \nScanOut693[3] , \nScanOut693[2] , 
        \nScanOut693[1] , \nScanOut693[0] }), .ScanOut({\nScanOut692[7] , 
        \nScanOut692[6] , \nScanOut692[5] , \nScanOut692[4] , \nScanOut692[3] , 
        \nScanOut692[2] , \nScanOut692[1] , \nScanOut692[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_19[7] , \nOut21_19[6] , \nOut21_19[5] , \nOut21_19[4] , 
        \nOut21_19[3] , \nOut21_19[2] , \nOut21_19[1] , \nOut21_19[0] }), 
        .SouthIn({\nOut21_21[7] , \nOut21_21[6] , \nOut21_21[5] , 
        \nOut21_21[4] , \nOut21_21[3] , \nOut21_21[2] , \nOut21_21[1] , 
        \nOut21_21[0] }), .EastIn({\nOut22_20[7] , \nOut22_20[6] , 
        \nOut22_20[5] , \nOut22_20[4] , \nOut22_20[3] , \nOut22_20[2] , 
        \nOut22_20[1] , \nOut22_20[0] }), .WestIn({\nOut20_20[7] , 
        \nOut20_20[6] , \nOut20_20[5] , \nOut20_20[4] , \nOut20_20[3] , 
        \nOut20_20[2] , \nOut20_20[1] , \nOut20_20[0] }), .Out({\nOut21_20[7] , 
        \nOut21_20[6] , \nOut21_20[5] , \nOut21_20[4] , \nOut21_20[3] , 
        \nOut21_20[2] , \nOut21_20[1] , \nOut21_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_702 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut703[7] , \nScanOut703[6] , 
        \nScanOut703[5] , \nScanOut703[4] , \nScanOut703[3] , \nScanOut703[2] , 
        \nScanOut703[1] , \nScanOut703[0] }), .ScanOut({\nScanOut702[7] , 
        \nScanOut702[6] , \nScanOut702[5] , \nScanOut702[4] , \nScanOut702[3] , 
        \nScanOut702[2] , \nScanOut702[1] , \nScanOut702[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_29[7] , \nOut21_29[6] , \nOut21_29[5] , \nOut21_29[4] , 
        \nOut21_29[3] , \nOut21_29[2] , \nOut21_29[1] , \nOut21_29[0] }), 
        .SouthIn({\nOut21_31[7] , \nOut21_31[6] , \nOut21_31[5] , 
        \nOut21_31[4] , \nOut21_31[3] , \nOut21_31[2] , \nOut21_31[1] , 
        \nOut21_31[0] }), .EastIn({\nOut22_30[7] , \nOut22_30[6] , 
        \nOut22_30[5] , \nOut22_30[4] , \nOut22_30[3] , \nOut22_30[2] , 
        \nOut22_30[1] , \nOut22_30[0] }), .WestIn({\nOut20_30[7] , 
        \nOut20_30[6] , \nOut20_30[5] , \nOut20_30[4] , \nOut20_30[3] , 
        \nOut20_30[2] , \nOut20_30[1] , \nOut20_30[0] }), .Out({\nOut21_30[7] , 
        \nOut21_30[6] , \nOut21_30[5] , \nOut21_30[4] , \nOut21_30[3] , 
        \nOut21_30[2] , \nOut21_30[1] , \nOut21_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_725 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut726[7] , \nScanOut726[6] , 
        \nScanOut726[5] , \nScanOut726[4] , \nScanOut726[3] , \nScanOut726[2] , 
        \nScanOut726[1] , \nScanOut726[0] }), .ScanOut({\nScanOut725[7] , 
        \nScanOut725[6] , \nScanOut725[5] , \nScanOut725[4] , \nScanOut725[3] , 
        \nScanOut725[2] , \nScanOut725[1] , \nScanOut725[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_20[7] , \nOut22_20[6] , \nOut22_20[5] , \nOut22_20[4] , 
        \nOut22_20[3] , \nOut22_20[2] , \nOut22_20[1] , \nOut22_20[0] }), 
        .SouthIn({\nOut22_22[7] , \nOut22_22[6] , \nOut22_22[5] , 
        \nOut22_22[4] , \nOut22_22[3] , \nOut22_22[2] , \nOut22_22[1] , 
        \nOut22_22[0] }), .EastIn({\nOut23_21[7] , \nOut23_21[6] , 
        \nOut23_21[5] , \nOut23_21[4] , \nOut23_21[3] , \nOut23_21[2] , 
        \nOut23_21[1] , \nOut23_21[0] }), .WestIn({\nOut21_21[7] , 
        \nOut21_21[6] , \nOut21_21[5] , \nOut21_21[4] , \nOut21_21[3] , 
        \nOut21_21[2] , \nOut21_21[1] , \nOut21_21[0] }), .Out({\nOut22_21[7] , 
        \nOut22_21[6] , \nOut22_21[5] , \nOut22_21[4] , \nOut22_21[3] , 
        \nOut22_21[2] , \nOut22_21[1] , \nOut22_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1004 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1005[7] , \nScanOut1005[6] , 
        \nScanOut1005[5] , \nScanOut1005[4] , \nScanOut1005[3] , 
        \nScanOut1005[2] , \nScanOut1005[1] , \nScanOut1005[0] }), .ScanOut({
        \nScanOut1004[7] , \nScanOut1004[6] , \nScanOut1004[5] , 
        \nScanOut1004[4] , \nScanOut1004[3] , \nScanOut1004[2] , 
        \nScanOut1004[1] , \nScanOut1004[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_12[7] , \nOut31_12[6] , \nOut31_12[5] , 
        \nOut31_12[4] , \nOut31_12[3] , \nOut31_12[2] , \nOut31_12[1] , 
        \nOut31_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_198 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut199[7] , \nScanOut199[6] , 
        \nScanOut199[5] , \nScanOut199[4] , \nScanOut199[3] , \nScanOut199[2] , 
        \nScanOut199[1] , \nScanOut199[0] }), .ScanOut({\nScanOut198[7] , 
        \nScanOut198[6] , \nScanOut198[5] , \nScanOut198[4] , \nScanOut198[3] , 
        \nScanOut198[2] , \nScanOut198[1] , \nScanOut198[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_5[7] , \nOut6_5[6] , \nOut6_5[5] , \nOut6_5[4] , \nOut6_5[3] , 
        \nOut6_5[2] , \nOut6_5[1] , \nOut6_5[0] }), .SouthIn({\nOut6_7[7] , 
        \nOut6_7[6] , \nOut6_7[5] , \nOut6_7[4] , \nOut6_7[3] , \nOut6_7[2] , 
        \nOut6_7[1] , \nOut6_7[0] }), .EastIn({\nOut7_6[7] , \nOut7_6[6] , 
        \nOut7_6[5] , \nOut7_6[4] , \nOut7_6[3] , \nOut7_6[2] , \nOut7_6[1] , 
        \nOut7_6[0] }), .WestIn({\nOut5_6[7] , \nOut5_6[6] , \nOut5_6[5] , 
        \nOut5_6[4] , \nOut5_6[3] , \nOut5_6[2] , \nOut5_6[1] , \nOut5_6[0] }), 
        .Out({\nOut6_6[7] , \nOut6_6[6] , \nOut6_6[5] , \nOut6_6[4] , 
        \nOut6_6[3] , \nOut6_6[2] , \nOut6_6[1] , \nOut6_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_223 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut224[7] , \nScanOut224[6] , 
        \nScanOut224[5] , \nScanOut224[4] , \nScanOut224[3] , \nScanOut224[2] , 
        \nScanOut224[1] , \nScanOut224[0] }), .ScanOut({\nScanOut223[7] , 
        \nScanOut223[6] , \nScanOut223[5] , \nScanOut223[4] , \nScanOut223[3] , 
        \nScanOut223[2] , \nScanOut223[1] , \nScanOut223[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut6_31[7] , \nOut6_31[6] , 
        \nOut6_31[5] , \nOut6_31[4] , \nOut6_31[3] , \nOut6_31[2] , 
        \nOut6_31[1] , \nOut6_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_432 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut433[7] , \nScanOut433[6] , 
        \nScanOut433[5] , \nScanOut433[4] , \nScanOut433[3] , \nScanOut433[2] , 
        \nScanOut433[1] , \nScanOut433[0] }), .ScanOut({\nScanOut432[7] , 
        \nScanOut432[6] , \nScanOut432[5] , \nScanOut432[4] , \nScanOut432[3] , 
        \nScanOut432[2] , \nScanOut432[1] , \nScanOut432[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_15[7] , \nOut13_15[6] , \nOut13_15[5] , \nOut13_15[4] , 
        \nOut13_15[3] , \nOut13_15[2] , \nOut13_15[1] , \nOut13_15[0] }), 
        .SouthIn({\nOut13_17[7] , \nOut13_17[6] , \nOut13_17[5] , 
        \nOut13_17[4] , \nOut13_17[3] , \nOut13_17[2] , \nOut13_17[1] , 
        \nOut13_17[0] }), .EastIn({\nOut14_16[7] , \nOut14_16[6] , 
        \nOut14_16[5] , \nOut14_16[4] , \nOut14_16[3] , \nOut14_16[2] , 
        \nOut14_16[1] , \nOut14_16[0] }), .WestIn({\nOut12_16[7] , 
        \nOut12_16[6] , \nOut12_16[5] , \nOut12_16[4] , \nOut12_16[3] , 
        \nOut12_16[2] , \nOut12_16[1] , \nOut12_16[0] }), .Out({\nOut13_16[7] , 
        \nOut13_16[6] , \nOut13_16[5] , \nOut13_16[4] , \nOut13_16[3] , 
        \nOut13_16[2] , \nOut13_16[1] , \nOut13_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_619 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut620[7] , \nScanOut620[6] , 
        \nScanOut620[5] , \nScanOut620[4] , \nScanOut620[3] , \nScanOut620[2] , 
        \nScanOut620[1] , \nScanOut620[0] }), .ScanOut({\nScanOut619[7] , 
        \nScanOut619[6] , \nScanOut619[5] , \nScanOut619[4] , \nScanOut619[3] , 
        \nScanOut619[2] , \nScanOut619[1] , \nScanOut619[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_10[7] , \nOut19_10[6] , \nOut19_10[5] , \nOut19_10[4] , 
        \nOut19_10[3] , \nOut19_10[2] , \nOut19_10[1] , \nOut19_10[0] }), 
        .SouthIn({\nOut19_12[7] , \nOut19_12[6] , \nOut19_12[5] , 
        \nOut19_12[4] , \nOut19_12[3] , \nOut19_12[2] , \nOut19_12[1] , 
        \nOut19_12[0] }), .EastIn({\nOut20_11[7] , \nOut20_11[6] , 
        \nOut20_11[5] , \nOut20_11[4] , \nOut20_11[3] , \nOut20_11[2] , 
        \nOut20_11[1] , \nOut20_11[0] }), .WestIn({\nOut18_11[7] , 
        \nOut18_11[6] , \nOut18_11[5] , \nOut18_11[4] , \nOut18_11[3] , 
        \nOut18_11[2] , \nOut18_11[1] , \nOut18_11[0] }), .Out({\nOut19_11[7] , 
        \nOut19_11[6] , \nOut19_11[5] , \nOut19_11[4] , \nOut19_11[3] , 
        \nOut19_11[2] , \nOut19_11[1] , \nOut19_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_789 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut790[7] , \nScanOut790[6] , 
        \nScanOut790[5] , \nScanOut790[4] , \nScanOut790[3] , \nScanOut790[2] , 
        \nScanOut790[1] , \nScanOut790[0] }), .ScanOut({\nScanOut789[7] , 
        \nScanOut789[6] , \nScanOut789[5] , \nScanOut789[4] , \nScanOut789[3] , 
        \nScanOut789[2] , \nScanOut789[1] , \nScanOut789[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_20[7] , \nOut24_20[6] , \nOut24_20[5] , \nOut24_20[4] , 
        \nOut24_20[3] , \nOut24_20[2] , \nOut24_20[1] , \nOut24_20[0] }), 
        .SouthIn({\nOut24_22[7] , \nOut24_22[6] , \nOut24_22[5] , 
        \nOut24_22[4] , \nOut24_22[3] , \nOut24_22[2] , \nOut24_22[1] , 
        \nOut24_22[0] }), .EastIn({\nOut25_21[7] , \nOut25_21[6] , 
        \nOut25_21[5] , \nOut25_21[4] , \nOut25_21[3] , \nOut25_21[2] , 
        \nOut25_21[1] , \nOut25_21[0] }), .WestIn({\nOut23_21[7] , 
        \nOut23_21[6] , \nOut23_21[5] , \nOut23_21[4] , \nOut23_21[3] , 
        \nOut23_21[2] , \nOut23_21[1] , \nOut23_21[0] }), .Out({\nOut24_21[7] , 
        \nOut24_21[6] , \nOut24_21[5] , \nOut24_21[4] , \nOut24_21[3] , 
        \nOut24_21[2] , \nOut24_21[1] , \nOut24_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_840 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut841[7] , \nScanOut841[6] , 
        \nScanOut841[5] , \nScanOut841[4] , \nScanOut841[3] , \nScanOut841[2] , 
        \nScanOut841[1] , \nScanOut841[0] }), .ScanOut({\nScanOut840[7] , 
        \nScanOut840[6] , \nScanOut840[5] , \nScanOut840[4] , \nScanOut840[3] , 
        \nScanOut840[2] , \nScanOut840[1] , \nScanOut840[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_7[7] , \nOut26_7[6] , \nOut26_7[5] , \nOut26_7[4] , 
        \nOut26_7[3] , \nOut26_7[2] , \nOut26_7[1] , \nOut26_7[0] }), 
        .SouthIn({\nOut26_9[7] , \nOut26_9[6] , \nOut26_9[5] , \nOut26_9[4] , 
        \nOut26_9[3] , \nOut26_9[2] , \nOut26_9[1] , \nOut26_9[0] }), .EastIn(
        {\nOut27_8[7] , \nOut27_8[6] , \nOut27_8[5] , \nOut27_8[4] , 
        \nOut27_8[3] , \nOut27_8[2] , \nOut27_8[1] , \nOut27_8[0] }), .WestIn(
        {\nOut25_8[7] , \nOut25_8[6] , \nOut25_8[5] , \nOut25_8[4] , 
        \nOut25_8[3] , \nOut25_8[2] , \nOut25_8[1] , \nOut25_8[0] }), .Out({
        \nOut26_8[7] , \nOut26_8[6] , \nOut26_8[5] , \nOut26_8[4] , 
        \nOut26_8[3] , \nOut26_8[2] , \nOut26_8[1] , \nOut26_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_338 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut339[7] , \nScanOut339[6] , 
        \nScanOut339[5] , \nScanOut339[4] , \nScanOut339[3] , \nScanOut339[2] , 
        \nScanOut339[1] , \nScanOut339[0] }), .ScanOut({\nScanOut338[7] , 
        \nScanOut338[6] , \nScanOut338[5] , \nScanOut338[4] , \nScanOut338[3] , 
        \nScanOut338[2] , \nScanOut338[1] , \nScanOut338[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_17[7] , \nOut10_17[6] , \nOut10_17[5] , \nOut10_17[4] , 
        \nOut10_17[3] , \nOut10_17[2] , \nOut10_17[1] , \nOut10_17[0] }), 
        .SouthIn({\nOut10_19[7] , \nOut10_19[6] , \nOut10_19[5] , 
        \nOut10_19[4] , \nOut10_19[3] , \nOut10_19[2] , \nOut10_19[1] , 
        \nOut10_19[0] }), .EastIn({\nOut11_18[7] , \nOut11_18[6] , 
        \nOut11_18[5] , \nOut11_18[4] , \nOut11_18[3] , \nOut11_18[2] , 
        \nOut11_18[1] , \nOut11_18[0] }), .WestIn({\nOut9_18[7] , 
        \nOut9_18[6] , \nOut9_18[5] , \nOut9_18[4] , \nOut9_18[3] , 
        \nOut9_18[2] , \nOut9_18[1] , \nOut9_18[0] }), .Out({\nOut10_18[7] , 
        \nOut10_18[6] , \nOut10_18[5] , \nOut10_18[4] , \nOut10_18[3] , 
        \nOut10_18[2] , \nOut10_18[1] , \nOut10_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_529 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut530[7] , \nScanOut530[6] , 
        \nScanOut530[5] , \nScanOut530[4] , \nScanOut530[3] , \nScanOut530[2] , 
        \nScanOut530[1] , \nScanOut530[0] }), .ScanOut({\nScanOut529[7] , 
        \nScanOut529[6] , \nScanOut529[5] , \nScanOut529[4] , \nScanOut529[3] , 
        \nScanOut529[2] , \nScanOut529[1] , \nScanOut529[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_16[7] , \nOut16_16[6] , \nOut16_16[5] , \nOut16_16[4] , 
        \nOut16_16[3] , \nOut16_16[2] , \nOut16_16[1] , \nOut16_16[0] }), 
        .SouthIn({\nOut16_18[7] , \nOut16_18[6] , \nOut16_18[5] , 
        \nOut16_18[4] , \nOut16_18[3] , \nOut16_18[2] , \nOut16_18[1] , 
        \nOut16_18[0] }), .EastIn({\nOut17_17[7] , \nOut17_17[6] , 
        \nOut17_17[5] , \nOut17_17[4] , \nOut17_17[3] , \nOut17_17[2] , 
        \nOut17_17[1] , \nOut17_17[0] }), .WestIn({\nOut15_17[7] , 
        \nOut15_17[6] , \nOut15_17[5] , \nOut15_17[4] , \nOut15_17[3] , 
        \nOut15_17[2] , \nOut15_17[1] , \nOut15_17[0] }), .Out({\nOut16_17[7] , 
        \nOut16_17[6] , \nOut16_17[5] , \nOut16_17[4] , \nOut16_17[3] , 
        \nOut16_17[2] , \nOut16_17[1] , \nOut16_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_57 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut58[7] , \nScanOut58[6] , 
        \nScanOut58[5] , \nScanOut58[4] , \nScanOut58[3] , \nScanOut58[2] , 
        \nScanOut58[1] , \nScanOut58[0] }), .ScanOut({\nScanOut57[7] , 
        \nScanOut57[6] , \nScanOut57[5] , \nScanOut57[4] , \nScanOut57[3] , 
        \nScanOut57[2] , \nScanOut57[1] , \nScanOut57[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_24[7] , \nOut1_24[6] , \nOut1_24[5] , \nOut1_24[4] , 
        \nOut1_24[3] , \nOut1_24[2] , \nOut1_24[1] , \nOut1_24[0] }), 
        .SouthIn({\nOut1_26[7] , \nOut1_26[6] , \nOut1_26[5] , \nOut1_26[4] , 
        \nOut1_26[3] , \nOut1_26[2] , \nOut1_26[1] , \nOut1_26[0] }), .EastIn(
        {\nOut2_25[7] , \nOut2_25[6] , \nOut2_25[5] , \nOut2_25[4] , 
        \nOut2_25[3] , \nOut2_25[2] , \nOut2_25[1] , \nOut2_25[0] }), .WestIn(
        {\nOut0_25[7] , \nOut0_25[6] , \nOut0_25[5] , \nOut0_25[4] , 
        \nOut0_25[3] , \nOut0_25[2] , \nOut0_25[1] , \nOut0_25[0] }), .Out({
        \nOut1_25[7] , \nOut1_25[6] , \nOut1_25[5] , \nOut1_25[4] , 
        \nOut1_25[3] , \nOut1_25[2] , \nOut1_25[1] , \nOut1_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_70 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut71[7] , \nScanOut71[6] , 
        \nScanOut71[5] , \nScanOut71[4] , \nScanOut71[3] , \nScanOut71[2] , 
        \nScanOut71[1] , \nScanOut71[0] }), .ScanOut({\nScanOut70[7] , 
        \nScanOut70[6] , \nScanOut70[5] , \nScanOut70[4] , \nScanOut70[3] , 
        \nScanOut70[2] , \nScanOut70[1] , \nScanOut70[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_5[7] , \nOut2_5[6] , \nOut2_5[5] , \nOut2_5[4] , \nOut2_5[3] , 
        \nOut2_5[2] , \nOut2_5[1] , \nOut2_5[0] }), .SouthIn({\nOut2_7[7] , 
        \nOut2_7[6] , \nOut2_7[5] , \nOut2_7[4] , \nOut2_7[3] , \nOut2_7[2] , 
        \nOut2_7[1] , \nOut2_7[0] }), .EastIn({\nOut3_6[7] , \nOut3_6[6] , 
        \nOut3_6[5] , \nOut3_6[4] , \nOut3_6[3] , \nOut3_6[2] , \nOut3_6[1] , 
        \nOut3_6[0] }), .WestIn({\nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , 
        \nOut1_6[4] , \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }), 
        .Out({\nOut2_6[7] , \nOut2_6[6] , \nOut2_6[5] , \nOut2_6[4] , 
        \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , \nOut2_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_95 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut96[7] , \nScanOut96[6] , 
        \nScanOut96[5] , \nScanOut96[4] , \nScanOut96[3] , \nScanOut96[2] , 
        \nScanOut96[1] , \nScanOut96[0] }), .ScanOut({\nScanOut95[7] , 
        \nScanOut95[6] , \nScanOut95[5] , \nScanOut95[4] , \nScanOut95[3] , 
        \nScanOut95[2] , \nScanOut95[1] , \nScanOut95[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut2_31[7] , \nOut2_31[6] , 
        \nOut2_31[5] , \nOut2_31[4] , \nOut2_31[3] , \nOut2_31[2] , 
        \nOut2_31[1] , \nOut2_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_101 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut102[7] , \nScanOut102[6] , 
        \nScanOut102[5] , \nScanOut102[4] , \nScanOut102[3] , \nScanOut102[2] , 
        \nScanOut102[1] , \nScanOut102[0] }), .ScanOut({\nScanOut101[7] , 
        \nScanOut101[6] , \nScanOut101[5] , \nScanOut101[4] , \nScanOut101[3] , 
        \nScanOut101[2] , \nScanOut101[1] , \nScanOut101[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_4[7] , \nOut3_4[6] , \nOut3_4[5] , \nOut3_4[4] , \nOut3_4[3] , 
        \nOut3_4[2] , \nOut3_4[1] , \nOut3_4[0] }), .SouthIn({\nOut3_6[7] , 
        \nOut3_6[6] , \nOut3_6[5] , \nOut3_6[4] , \nOut3_6[3] , \nOut3_6[2] , 
        \nOut3_6[1] , \nOut3_6[0] }), .EastIn({\nOut4_5[7] , \nOut4_5[6] , 
        \nOut4_5[5] , \nOut4_5[4] , \nOut4_5[3] , \nOut4_5[2] , \nOut4_5[1] , 
        \nOut4_5[0] }), .WestIn({\nOut2_5[7] , \nOut2_5[6] , \nOut2_5[5] , 
        \nOut2_5[4] , \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , \nOut2_5[0] }), 
        .Out({\nOut3_5[7] , \nOut3_5[6] , \nOut3_5[5] , \nOut3_5[4] , 
        \nOut3_5[3] , \nOut3_5[2] , \nOut3_5[1] , \nOut3_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_126 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut127[7] , \nScanOut127[6] , 
        \nScanOut127[5] , \nScanOut127[4] , \nScanOut127[3] , \nScanOut127[2] , 
        \nScanOut127[1] , \nScanOut127[0] }), .ScanOut({\nScanOut126[7] , 
        \nScanOut126[6] , \nScanOut126[5] , \nScanOut126[4] , \nScanOut126[3] , 
        \nScanOut126[2] , \nScanOut126[1] , \nScanOut126[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_29[7] , \nOut3_29[6] , \nOut3_29[5] , \nOut3_29[4] , 
        \nOut3_29[3] , \nOut3_29[2] , \nOut3_29[1] , \nOut3_29[0] }), 
        .SouthIn({\nOut3_31[7] , \nOut3_31[6] , \nOut3_31[5] , \nOut3_31[4] , 
        \nOut3_31[3] , \nOut3_31[2] , \nOut3_31[1] , \nOut3_31[0] }), .EastIn(
        {\nOut4_30[7] , \nOut4_30[6] , \nOut4_30[5] , \nOut4_30[4] , 
        \nOut4_30[3] , \nOut4_30[2] , \nOut4_30[1] , \nOut4_30[0] }), .WestIn(
        {\nOut2_30[7] , \nOut2_30[6] , \nOut2_30[5] , \nOut2_30[4] , 
        \nOut2_30[3] , \nOut2_30[2] , \nOut2_30[1] , \nOut2_30[0] }), .Out({
        \nOut3_30[7] , \nOut3_30[6] , \nOut3_30[5] , \nOut3_30[4] , 
        \nOut3_30[3] , \nOut3_30[2] , \nOut3_30[1] , \nOut3_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_216 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut217[7] , \nScanOut217[6] , 
        \nScanOut217[5] , \nScanOut217[4] , \nScanOut217[3] , \nScanOut217[2] , 
        \nScanOut217[1] , \nScanOut217[0] }), .ScanOut({\nScanOut216[7] , 
        \nScanOut216[6] , \nScanOut216[5] , \nScanOut216[4] , \nScanOut216[3] , 
        \nScanOut216[2] , \nScanOut216[1] , \nScanOut216[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_23[7] , \nOut6_23[6] , \nOut6_23[5] , \nOut6_23[4] , 
        \nOut6_23[3] , \nOut6_23[2] , \nOut6_23[1] , \nOut6_23[0] }), 
        .SouthIn({\nOut6_25[7] , \nOut6_25[6] , \nOut6_25[5] , \nOut6_25[4] , 
        \nOut6_25[3] , \nOut6_25[2] , \nOut6_25[1] , \nOut6_25[0] }), .EastIn(
        {\nOut7_24[7] , \nOut7_24[6] , \nOut7_24[5] , \nOut7_24[4] , 
        \nOut7_24[3] , \nOut7_24[2] , \nOut7_24[1] , \nOut7_24[0] }), .WestIn(
        {\nOut5_24[7] , \nOut5_24[6] , \nOut5_24[5] , \nOut5_24[4] , 
        \nOut5_24[3] , \nOut5_24[2] , \nOut5_24[1] , \nOut5_24[0] }), .Out({
        \nOut6_24[7] , \nOut6_24[6] , \nOut6_24[5] , \nOut6_24[4] , 
        \nOut6_24[3] , \nOut6_24[2] , \nOut6_24[1] , \nOut6_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_386 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut387[7] , \nScanOut387[6] , 
        \nScanOut387[5] , \nScanOut387[4] , \nScanOut387[3] , \nScanOut387[2] , 
        \nScanOut387[1] , \nScanOut387[0] }), .ScanOut({\nScanOut386[7] , 
        \nScanOut386[6] , \nScanOut386[5] , \nScanOut386[4] , \nScanOut386[3] , 
        \nScanOut386[2] , \nScanOut386[1] , \nScanOut386[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_1[7] , \nOut12_1[6] , \nOut12_1[5] , \nOut12_1[4] , 
        \nOut12_1[3] , \nOut12_1[2] , \nOut12_1[1] , \nOut12_1[0] }), 
        .SouthIn({\nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }), .EastIn(
        {\nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }), .WestIn(
        {\nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }), .Out({
        \nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_875 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut876[7] , \nScanOut876[6] , 
        \nScanOut876[5] , \nScanOut876[4] , \nScanOut876[3] , \nScanOut876[2] , 
        \nScanOut876[1] , \nScanOut876[0] }), .ScanOut({\nScanOut875[7] , 
        \nScanOut875[6] , \nScanOut875[5] , \nScanOut875[4] , \nScanOut875[3] , 
        \nScanOut875[2] , \nScanOut875[1] , \nScanOut875[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_10[7] , \nOut27_10[6] , \nOut27_10[5] , \nOut27_10[4] , 
        \nOut27_10[3] , \nOut27_10[2] , \nOut27_10[1] , \nOut27_10[0] }), 
        .SouthIn({\nOut27_12[7] , \nOut27_12[6] , \nOut27_12[5] , 
        \nOut27_12[4] , \nOut27_12[3] , \nOut27_12[2] , \nOut27_12[1] , 
        \nOut27_12[0] }), .EastIn({\nOut28_11[7] , \nOut28_11[6] , 
        \nOut28_11[5] , \nOut28_11[4] , \nOut28_11[3] , \nOut28_11[2] , 
        \nOut28_11[1] , \nOut28_11[0] }), .WestIn({\nOut26_11[7] , 
        \nOut26_11[6] , \nOut26_11[5] , \nOut26_11[4] , \nOut26_11[3] , 
        \nOut26_11[2] , \nOut26_11[1] , \nOut26_11[0] }), .Out({\nOut27_11[7] , 
        \nOut27_11[6] , \nOut27_11[5] , \nOut27_11[4] , \nOut27_11[3] , 
        \nOut27_11[2] , \nOut27_11[1] , \nOut27_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_949 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut950[7] , \nScanOut950[6] , 
        \nScanOut950[5] , \nScanOut950[4] , \nScanOut950[3] , \nScanOut950[2] , 
        \nScanOut950[1] , \nScanOut950[0] }), .ScanOut({\nScanOut949[7] , 
        \nScanOut949[6] , \nScanOut949[5] , \nScanOut949[4] , \nScanOut949[3] , 
        \nScanOut949[2] , \nScanOut949[1] , \nScanOut949[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_20[7] , \nOut29_20[6] , \nOut29_20[5] , \nOut29_20[4] , 
        \nOut29_20[3] , \nOut29_20[2] , \nOut29_20[1] , \nOut29_20[0] }), 
        .SouthIn({\nOut29_22[7] , \nOut29_22[6] , \nOut29_22[5] , 
        \nOut29_22[4] , \nOut29_22[3] , \nOut29_22[2] , \nOut29_22[1] , 
        \nOut29_22[0] }), .EastIn({\nOut30_21[7] , \nOut30_21[6] , 
        \nOut30_21[5] , \nOut30_21[4] , \nOut30_21[3] , \nOut30_21[2] , 
        \nOut30_21[1] , \nOut30_21[0] }), .WestIn({\nOut28_21[7] , 
        \nOut28_21[6] , \nOut28_21[5] , \nOut28_21[4] , \nOut28_21[3] , 
        \nOut28_21[2] , \nOut28_21[1] , \nOut28_21[0] }), .Out({\nOut29_21[7] , 
        \nOut29_21[6] , \nOut29_21[5] , \nOut29_21[4] , \nOut29_21[3] , 
        \nOut29_21[2] , \nOut29_21[1] , \nOut29_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_407 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut408[7] , \nScanOut408[6] , 
        \nScanOut408[5] , \nScanOut408[4] , \nScanOut408[3] , \nScanOut408[2] , 
        \nScanOut408[1] , \nScanOut408[0] }), .ScanOut({\nScanOut407[7] , 
        \nScanOut407[6] , \nScanOut407[5] , \nScanOut407[4] , \nScanOut407[3] , 
        \nScanOut407[2] , \nScanOut407[1] , \nScanOut407[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_22[7] , \nOut12_22[6] , \nOut12_22[5] , \nOut12_22[4] , 
        \nOut12_22[3] , \nOut12_22[2] , \nOut12_22[1] , \nOut12_22[0] }), 
        .SouthIn({\nOut12_24[7] , \nOut12_24[6] , \nOut12_24[5] , 
        \nOut12_24[4] , \nOut12_24[3] , \nOut12_24[2] , \nOut12_24[1] , 
        \nOut12_24[0] }), .EastIn({\nOut13_23[7] , \nOut13_23[6] , 
        \nOut13_23[5] , \nOut13_23[4] , \nOut13_23[3] , \nOut13_23[2] , 
        \nOut13_23[1] , \nOut13_23[0] }), .WestIn({\nOut11_23[7] , 
        \nOut11_23[6] , \nOut11_23[5] , \nOut11_23[4] , \nOut11_23[3] , 
        \nOut11_23[2] , \nOut11_23[1] , \nOut11_23[0] }), .Out({\nOut12_23[7] , 
        \nOut12_23[6] , \nOut12_23[5] , \nOut12_23[4] , \nOut12_23[3] , 
        \nOut12_23[2] , \nOut12_23[1] , \nOut12_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_597 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut598[7] , \nScanOut598[6] , 
        \nScanOut598[5] , \nScanOut598[4] , \nScanOut598[3] , \nScanOut598[2] , 
        \nScanOut598[1] , \nScanOut598[0] }), .ScanOut({\nScanOut597[7] , 
        \nScanOut597[6] , \nScanOut597[5] , \nScanOut597[4] , \nScanOut597[3] , 
        \nScanOut597[2] , \nScanOut597[1] , \nScanOut597[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_20[7] , \nOut18_20[6] , \nOut18_20[5] , \nOut18_20[4] , 
        \nOut18_20[3] , \nOut18_20[2] , \nOut18_20[1] , \nOut18_20[0] }), 
        .SouthIn({\nOut18_22[7] , \nOut18_22[6] , \nOut18_22[5] , 
        \nOut18_22[4] , \nOut18_22[3] , \nOut18_22[2] , \nOut18_22[1] , 
        \nOut18_22[0] }), .EastIn({\nOut19_21[7] , \nOut19_21[6] , 
        \nOut19_21[5] , \nOut19_21[4] , \nOut19_21[3] , \nOut19_21[2] , 
        \nOut19_21[1] , \nOut19_21[0] }), .WestIn({\nOut17_21[7] , 
        \nOut17_21[6] , \nOut17_21[5] , \nOut17_21[4] , \nOut17_21[3] , 
        \nOut17_21[2] , \nOut17_21[1] , \nOut17_21[0] }), .Out({\nOut18_21[7] , 
        \nOut18_21[6] , \nOut18_21[5] , \nOut18_21[4] , \nOut18_21[3] , 
        \nOut18_21[2] , \nOut18_21[1] , \nOut18_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_737 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut738[7] , \nScanOut738[6] , 
        \nScanOut738[5] , \nScanOut738[4] , \nScanOut738[3] , \nScanOut738[2] , 
        \nScanOut738[1] , \nScanOut738[0] }), .ScanOut({\nScanOut737[7] , 
        \nScanOut737[6] , \nScanOut737[5] , \nScanOut737[4] , \nScanOut737[3] , 
        \nScanOut737[2] , \nScanOut737[1] , \nScanOut737[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_0[7] , \nOut23_0[6] , \nOut23_0[5] , \nOut23_0[4] , 
        \nOut23_0[3] , \nOut23_0[2] , \nOut23_0[1] , \nOut23_0[0] }), 
        .SouthIn({\nOut23_2[7] , \nOut23_2[6] , \nOut23_2[5] , \nOut23_2[4] , 
        \nOut23_2[3] , \nOut23_2[2] , \nOut23_2[1] , \nOut23_2[0] }), .EastIn(
        {\nOut24_1[7] , \nOut24_1[6] , \nOut24_1[5] , \nOut24_1[4] , 
        \nOut24_1[3] , \nOut24_1[2] , \nOut24_1[1] , \nOut24_1[0] }), .WestIn(
        {\nOut22_1[7] , \nOut22_1[6] , \nOut22_1[5] , \nOut22_1[4] , 
        \nOut22_1[3] , \nOut22_1[2] , \nOut22_1[1] , \nOut22_1[0] }), .Out({
        \nOut23_1[7] , \nOut23_1[6] , \nOut23_1[5] , \nOut23_1[4] , 
        \nOut23_1[3] , \nOut23_1[2] , \nOut23_1[1] , \nOut23_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_680 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut681[7] , \nScanOut681[6] , 
        \nScanOut681[5] , \nScanOut681[4] , \nScanOut681[3] , \nScanOut681[2] , 
        \nScanOut681[1] , \nScanOut681[0] }), .ScanOut({\nScanOut680[7] , 
        \nScanOut680[6] , \nScanOut680[5] , \nScanOut680[4] , \nScanOut680[3] , 
        \nScanOut680[2] , \nScanOut680[1] , \nScanOut680[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_7[7] , \nOut21_7[6] , \nOut21_7[5] , \nOut21_7[4] , 
        \nOut21_7[3] , \nOut21_7[2] , \nOut21_7[1] , \nOut21_7[0] }), 
        .SouthIn({\nOut21_9[7] , \nOut21_9[6] , \nOut21_9[5] , \nOut21_9[4] , 
        \nOut21_9[3] , \nOut21_9[2] , \nOut21_9[1] , \nOut21_9[0] }), .EastIn(
        {\nOut22_8[7] , \nOut22_8[6] , \nOut22_8[5] , \nOut22_8[4] , 
        \nOut22_8[3] , \nOut22_8[2] , \nOut22_8[1] , \nOut22_8[0] }), .WestIn(
        {\nOut20_8[7] , \nOut20_8[6] , \nOut20_8[5] , \nOut20_8[4] , 
        \nOut20_8[3] , \nOut20_8[2] , \nOut20_8[1] , \nOut20_8[0] }), .Out({
        \nOut21_8[7] , \nOut21_8[6] , \nOut21_8[5] , \nOut21_8[4] , 
        \nOut21_8[3] , \nOut21_8[2] , \nOut21_8[1] , \nOut21_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1016 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1017[7] , \nScanOut1017[6] , 
        \nScanOut1017[5] , \nScanOut1017[4] , \nScanOut1017[3] , 
        \nScanOut1017[2] , \nScanOut1017[1] , \nScanOut1017[0] }), .ScanOut({
        \nScanOut1016[7] , \nScanOut1016[6] , \nScanOut1016[5] , 
        \nScanOut1016[4] , \nScanOut1016[3] , \nScanOut1016[2] , 
        \nScanOut1016[1] , \nScanOut1016[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_24[7] , \nOut31_24[6] , \nOut31_24[5] , 
        \nOut31_24[4] , \nOut31_24[3] , \nOut31_24[2] , \nOut31_24[1] , 
        \nOut31_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_710 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut711[7] , \nScanOut711[6] , 
        \nScanOut711[5] , \nScanOut711[4] , \nScanOut711[3] , \nScanOut711[2] , 
        \nScanOut711[1] , \nScanOut711[0] }), .ScanOut({\nScanOut710[7] , 
        \nScanOut710[6] , \nScanOut710[5] , \nScanOut710[4] , \nScanOut710[3] , 
        \nScanOut710[2] , \nScanOut710[1] , \nScanOut710[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_5[7] , \nOut22_5[6] , \nOut22_5[5] , \nOut22_5[4] , 
        \nOut22_5[3] , \nOut22_5[2] , \nOut22_5[1] , \nOut22_5[0] }), 
        .SouthIn({\nOut22_7[7] , \nOut22_7[6] , \nOut22_7[5] , \nOut22_7[4] , 
        \nOut22_7[3] , \nOut22_7[2] , \nOut22_7[1] , \nOut22_7[0] }), .EastIn(
        {\nOut23_6[7] , \nOut23_6[6] , \nOut23_6[5] , \nOut23_6[4] , 
        \nOut23_6[3] , \nOut23_6[2] , \nOut23_6[1] , \nOut23_6[0] }), .WestIn(
        {\nOut21_6[7] , \nOut21_6[6] , \nOut21_6[5] , \nOut21_6[4] , 
        \nOut21_6[3] , \nOut21_6[2] , \nOut21_6[1] , \nOut21_6[0] }), .Out({
        \nOut22_6[7] , \nOut22_6[6] , \nOut22_6[5] , \nOut22_6[4] , 
        \nOut22_6[3] , \nOut22_6[2] , \nOut22_6[1] , \nOut22_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_148 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut149[7] , \nScanOut149[6] , 
        \nScanOut149[5] , \nScanOut149[4] , \nScanOut149[3] , \nScanOut149[2] , 
        \nScanOut149[1] , \nScanOut149[0] }), .ScanOut({\nScanOut148[7] , 
        \nScanOut148[6] , \nScanOut148[5] , \nScanOut148[4] , \nScanOut148[3] , 
        \nScanOut148[2] , \nScanOut148[1] , \nScanOut148[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_19[7] , \nOut4_19[6] , \nOut4_19[5] , \nOut4_19[4] , 
        \nOut4_19[3] , \nOut4_19[2] , \nOut4_19[1] , \nOut4_19[0] }), 
        .SouthIn({\nOut4_21[7] , \nOut4_21[6] , \nOut4_21[5] , \nOut4_21[4] , 
        \nOut4_21[3] , \nOut4_21[2] , \nOut4_21[1] , \nOut4_21[0] }), .EastIn(
        {\nOut5_20[7] , \nOut5_20[6] , \nOut5_20[5] , \nOut5_20[4] , 
        \nOut5_20[3] , \nOut5_20[2] , \nOut5_20[1] , \nOut5_20[0] }), .WestIn(
        {\nOut3_20[7] , \nOut3_20[6] , \nOut3_20[5] , \nOut3_20[4] , 
        \nOut3_20[3] , \nOut3_20[2] , \nOut3_20[1] , \nOut3_20[0] }), .Out({
        \nOut4_20[7] , \nOut4_20[6] , \nOut4_20[5] , \nOut4_20[4] , 
        \nOut4_20[3] , \nOut4_20[2] , \nOut4_20[1] , \nOut4_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_231 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut232[7] , \nScanOut232[6] , 
        \nScanOut232[5] , \nScanOut232[4] , \nScanOut232[3] , \nScanOut232[2] , 
        \nScanOut232[1] , \nScanOut232[0] }), .ScanOut({\nScanOut231[7] , 
        \nScanOut231[6] , \nScanOut231[5] , \nScanOut231[4] , \nScanOut231[3] , 
        \nScanOut231[2] , \nScanOut231[1] , \nScanOut231[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_6[7] , \nOut7_6[6] , \nOut7_6[5] , \nOut7_6[4] , \nOut7_6[3] , 
        \nOut7_6[2] , \nOut7_6[1] , \nOut7_6[0] }), .SouthIn({\nOut7_8[7] , 
        \nOut7_8[6] , \nOut7_8[5] , \nOut7_8[4] , \nOut7_8[3] , \nOut7_8[2] , 
        \nOut7_8[1] , \nOut7_8[0] }), .EastIn({\nOut8_7[7] , \nOut8_7[6] , 
        \nOut8_7[5] , \nOut8_7[4] , \nOut8_7[3] , \nOut8_7[2] , \nOut8_7[1] , 
        \nOut8_7[0] }), .WestIn({\nOut6_7[7] , \nOut6_7[6] , \nOut6_7[5] , 
        \nOut6_7[4] , \nOut6_7[3] , \nOut6_7[2] , \nOut6_7[1] , \nOut6_7[0] }), 
        .Out({\nOut7_7[7] , \nOut7_7[6] , \nOut7_7[5] , \nOut7_7[4] , 
        \nOut7_7[3] , \nOut7_7[2] , \nOut7_7[1] , \nOut7_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_852 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut853[7] , \nScanOut853[6] , 
        \nScanOut853[5] , \nScanOut853[4] , \nScanOut853[3] , \nScanOut853[2] , 
        \nScanOut853[1] , \nScanOut853[0] }), .ScanOut({\nScanOut852[7] , 
        \nScanOut852[6] , \nScanOut852[5] , \nScanOut852[4] , \nScanOut852[3] , 
        \nScanOut852[2] , \nScanOut852[1] , \nScanOut852[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_19[7] , \nOut26_19[6] , \nOut26_19[5] , \nOut26_19[4] , 
        \nOut26_19[3] , \nOut26_19[2] , \nOut26_19[1] , \nOut26_19[0] }), 
        .SouthIn({\nOut26_21[7] , \nOut26_21[6] , \nOut26_21[5] , 
        \nOut26_21[4] , \nOut26_21[3] , \nOut26_21[2] , \nOut26_21[1] , 
        \nOut26_21[0] }), .EastIn({\nOut27_20[7] , \nOut27_20[6] , 
        \nOut27_20[5] , \nOut27_20[4] , \nOut27_20[3] , \nOut27_20[2] , 
        \nOut27_20[1] , \nOut27_20[0] }), .WestIn({\nOut25_20[7] , 
        \nOut25_20[6] , \nOut25_20[5] , \nOut25_20[4] , \nOut25_20[3] , 
        \nOut25_20[2] , \nOut25_20[1] , \nOut25_20[0] }), .Out({\nOut26_20[7] , 
        \nOut26_20[6] , \nOut26_20[5] , \nOut26_20[4] , \nOut26_20[3] , 
        \nOut26_20[2] , \nOut26_20[1] , \nOut26_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_278 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut279[7] , \nScanOut279[6] , 
        \nScanOut279[5] , \nScanOut279[4] , \nScanOut279[3] , \nScanOut279[2] , 
        \nScanOut279[1] , \nScanOut279[0] }), .ScanOut({\nScanOut278[7] , 
        \nScanOut278[6] , \nScanOut278[5] , \nScanOut278[4] , \nScanOut278[3] , 
        \nScanOut278[2] , \nScanOut278[1] , \nScanOut278[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_21[7] , \nOut8_21[6] , \nOut8_21[5] , \nOut8_21[4] , 
        \nOut8_21[3] , \nOut8_21[2] , \nOut8_21[1] , \nOut8_21[0] }), 
        .SouthIn({\nOut8_23[7] , \nOut8_23[6] , \nOut8_23[5] , \nOut8_23[4] , 
        \nOut8_23[3] , \nOut8_23[2] , \nOut8_23[1] , \nOut8_23[0] }), .EastIn(
        {\nOut9_22[7] , \nOut9_22[6] , \nOut9_22[5] , \nOut9_22[4] , 
        \nOut9_22[3] , \nOut9_22[2] , \nOut9_22[1] , \nOut9_22[0] }), .WestIn(
        {\nOut7_22[7] , \nOut7_22[6] , \nOut7_22[5] , \nOut7_22[4] , 
        \nOut7_22[3] , \nOut7_22[2] , \nOut7_22[1] , \nOut7_22[0] }), .Out({
        \nOut8_22[7] , \nOut8_22[6] , \nOut8_22[5] , \nOut8_22[4] , 
        \nOut8_22[3] , \nOut8_22[2] , \nOut8_22[1] , \nOut8_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_420 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut421[7] , \nScanOut421[6] , 
        \nScanOut421[5] , \nScanOut421[4] , \nScanOut421[3] , \nScanOut421[2] , 
        \nScanOut421[1] , \nScanOut421[0] }), .ScanOut({\nScanOut420[7] , 
        \nScanOut420[6] , \nScanOut420[5] , \nScanOut420[4] , \nScanOut420[3] , 
        \nScanOut420[2] , \nScanOut420[1] , \nScanOut420[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }), 
        .SouthIn({\nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }), .EastIn(
        {\nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }), .WestIn(
        {\nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }), .Out({
        \nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_469 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut470[7] , \nScanOut470[6] , 
        \nScanOut470[5] , \nScanOut470[4] , \nScanOut470[3] , \nScanOut470[2] , 
        \nScanOut470[1] , \nScanOut470[0] }), .ScanOut({\nScanOut469[7] , 
        \nScanOut469[6] , \nScanOut469[5] , \nScanOut469[4] , \nScanOut469[3] , 
        \nScanOut469[2] , \nScanOut469[1] , \nScanOut469[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_20[7] , \nOut14_20[6] , \nOut14_20[5] , \nOut14_20[4] , 
        \nOut14_20[3] , \nOut14_20[2] , \nOut14_20[1] , \nOut14_20[0] }), 
        .SouthIn({\nOut14_22[7] , \nOut14_22[6] , \nOut14_22[5] , 
        \nOut14_22[4] , \nOut14_22[3] , \nOut14_22[2] , \nOut14_22[1] , 
        \nOut14_22[0] }), .EastIn({\nOut15_21[7] , \nOut15_21[6] , 
        \nOut15_21[5] , \nOut15_21[4] , \nOut15_21[3] , \nOut15_21[2] , 
        \nOut15_21[1] , \nOut15_21[0] }), .WestIn({\nOut13_21[7] , 
        \nOut13_21[6] , \nOut13_21[5] , \nOut13_21[4] , \nOut13_21[3] , 
        \nOut13_21[2] , \nOut13_21[1] , \nOut13_21[0] }), .Out({\nOut14_21[7] , 
        \nOut14_21[6] , \nOut14_21[5] , \nOut14_21[4] , \nOut14_21[3] , 
        \nOut14_21[2] , \nOut14_21[1] , \nOut14_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_759 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut760[7] , \nScanOut760[6] , 
        \nScanOut760[5] , \nScanOut760[4] , \nScanOut760[3] , \nScanOut760[2] , 
        \nScanOut760[1] , \nScanOut760[0] }), .ScanOut({\nScanOut759[7] , 
        \nScanOut759[6] , \nScanOut759[5] , \nScanOut759[4] , \nScanOut759[3] , 
        \nScanOut759[2] , \nScanOut759[1] , \nScanOut759[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_22[7] , \nOut23_22[6] , \nOut23_22[5] , \nOut23_22[4] , 
        \nOut23_22[3] , \nOut23_22[2] , \nOut23_22[1] , \nOut23_22[0] }), 
        .SouthIn({\nOut23_24[7] , \nOut23_24[6] , \nOut23_24[5] , 
        \nOut23_24[4] , \nOut23_24[3] , \nOut23_24[2] , \nOut23_24[1] , 
        \nOut23_24[0] }), .EastIn({\nOut24_23[7] , \nOut24_23[6] , 
        \nOut24_23[5] , \nOut24_23[4] , \nOut24_23[3] , \nOut24_23[2] , 
        \nOut24_23[1] , \nOut24_23[0] }), .WestIn({\nOut22_23[7] , 
        \nOut22_23[6] , \nOut22_23[5] , \nOut22_23[4] , \nOut22_23[3] , 
        \nOut22_23[2] , \nOut22_23[1] , \nOut22_23[0] }), .Out({\nOut23_23[7] , 
        \nOut23_23[6] , \nOut23_23[5] , \nOut23_23[4] , \nOut23_23[3] , 
        \nOut23_23[2] , \nOut23_23[1] , \nOut23_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_344 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut345[7] , \nScanOut345[6] , 
        \nScanOut345[5] , \nScanOut345[4] , \nScanOut345[3] , \nScanOut345[2] , 
        \nScanOut345[1] , \nScanOut345[0] }), .ScanOut({\nScanOut344[7] , 
        \nScanOut344[6] , \nScanOut344[5] , \nScanOut344[4] , \nScanOut344[3] , 
        \nScanOut344[2] , \nScanOut344[1] , \nScanOut344[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_23[7] , \nOut10_23[6] , \nOut10_23[5] , \nOut10_23[4] , 
        \nOut10_23[3] , \nOut10_23[2] , \nOut10_23[1] , \nOut10_23[0] }), 
        .SouthIn({\nOut10_25[7] , \nOut10_25[6] , \nOut10_25[5] , 
        \nOut10_25[4] , \nOut10_25[3] , \nOut10_25[2] , \nOut10_25[1] , 
        \nOut10_25[0] }), .EastIn({\nOut11_24[7] , \nOut11_24[6] , 
        \nOut11_24[5] , \nOut11_24[4] , \nOut11_24[3] , \nOut11_24[2] , 
        \nOut11_24[1] , \nOut11_24[0] }), .WestIn({\nOut9_24[7] , 
        \nOut9_24[6] , \nOut9_24[5] , \nOut9_24[4] , \nOut9_24[3] , 
        \nOut9_24[2] , \nOut9_24[1] , \nOut9_24[0] }), .Out({\nOut10_24[7] , 
        \nOut10_24[6] , \nOut10_24[5] , \nOut10_24[4] , \nOut10_24[3] , 
        \nOut10_24[2] , \nOut10_24[1] , \nOut10_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_665 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut666[7] , \nScanOut666[6] , 
        \nScanOut666[5] , \nScanOut666[4] , \nScanOut666[3] , \nScanOut666[2] , 
        \nScanOut666[1] , \nScanOut666[0] }), .ScanOut({\nScanOut665[7] , 
        \nScanOut665[6] , \nScanOut665[5] , \nScanOut665[4] , \nScanOut665[3] , 
        \nScanOut665[2] , \nScanOut665[1] , \nScanOut665[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_24[7] , \nOut20_24[6] , \nOut20_24[5] , \nOut20_24[4] , 
        \nOut20_24[3] , \nOut20_24[2] , \nOut20_24[1] , \nOut20_24[0] }), 
        .SouthIn({\nOut20_26[7] , \nOut20_26[6] , \nOut20_26[5] , 
        \nOut20_26[4] , \nOut20_26[3] , \nOut20_26[2] , \nOut20_26[1] , 
        \nOut20_26[0] }), .EastIn({\nOut21_25[7] , \nOut21_25[6] , 
        \nOut21_25[5] , \nOut21_25[4] , \nOut21_25[3] , \nOut21_25[2] , 
        \nOut21_25[1] , \nOut21_25[0] }), .WestIn({\nOut19_25[7] , 
        \nOut19_25[6] , \nOut19_25[5] , \nOut19_25[4] , \nOut19_25[3] , 
        \nOut19_25[2] , \nOut19_25[1] , \nOut19_25[0] }), .Out({\nOut20_25[7] , 
        \nOut20_25[6] , \nOut20_25[5] , \nOut20_25[4] , \nOut20_25[3] , 
        \nOut20_25[2] , \nOut20_25[1] , \nOut20_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_927 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut928[7] , \nScanOut928[6] , 
        \nScanOut928[5] , \nScanOut928[4] , \nScanOut928[3] , \nScanOut928[2] , 
        \nScanOut928[1] , \nScanOut928[0] }), .ScanOut({\nScanOut927[7] , 
        \nScanOut927[6] , \nScanOut927[5] , \nScanOut927[4] , \nScanOut927[3] , 
        \nScanOut927[2] , \nScanOut927[1] , \nScanOut927[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut28_31[7] , \nOut28_31[6] , 
        \nOut28_31[5] , \nOut28_31[4] , \nOut28_31[3] , \nOut28_31[2] , 
        \nOut28_31[1] , \nOut28_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_363 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut364[7] , \nScanOut364[6] , 
        \nScanOut364[5] , \nScanOut364[4] , \nScanOut364[3] , \nScanOut364[2] , 
        \nScanOut364[1] , \nScanOut364[0] }), .ScanOut({\nScanOut363[7] , 
        \nScanOut363[6] , \nScanOut363[5] , \nScanOut363[4] , \nScanOut363[3] , 
        \nScanOut363[2] , \nScanOut363[1] , \nScanOut363[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_10[7] , \nOut11_10[6] , \nOut11_10[5] , \nOut11_10[4] , 
        \nOut11_10[3] , \nOut11_10[2] , \nOut11_10[1] , \nOut11_10[0] }), 
        .SouthIn({\nOut11_12[7] , \nOut11_12[6] , \nOut11_12[5] , 
        \nOut11_12[4] , \nOut11_12[3] , \nOut11_12[2] , \nOut11_12[1] , 
        \nOut11_12[0] }), .EastIn({\nOut12_11[7] , \nOut12_11[6] , 
        \nOut12_11[5] , \nOut12_11[4] , \nOut12_11[3] , \nOut12_11[2] , 
        \nOut12_11[1] , \nOut12_11[0] }), .WestIn({\nOut10_11[7] , 
        \nOut10_11[6] , \nOut10_11[5] , \nOut10_11[4] , \nOut10_11[3] , 
        \nOut10_11[2] , \nOut10_11[1] , \nOut10_11[0] }), .Out({\nOut11_11[7] , 
        \nOut11_11[6] , \nOut11_11[5] , \nOut11_11[4] , \nOut11_11[3] , 
        \nOut11_11[2] , \nOut11_11[1] , \nOut11_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_555 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut556[7] , \nScanOut556[6] , 
        \nScanOut556[5] , \nScanOut556[4] , \nScanOut556[3] , \nScanOut556[2] , 
        \nScanOut556[1] , \nScanOut556[0] }), .ScanOut({\nScanOut555[7] , 
        \nScanOut555[6] , \nScanOut555[5] , \nScanOut555[4] , \nScanOut555[3] , 
        \nScanOut555[2] , \nScanOut555[1] , \nScanOut555[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_10[7] , \nOut17_10[6] , \nOut17_10[5] , \nOut17_10[4] , 
        \nOut17_10[3] , \nOut17_10[2] , \nOut17_10[1] , \nOut17_10[0] }), 
        .SouthIn({\nOut17_12[7] , \nOut17_12[6] , \nOut17_12[5] , 
        \nOut17_12[4] , \nOut17_12[3] , \nOut17_12[2] , \nOut17_12[1] , 
        \nOut17_12[0] }), .EastIn({\nOut18_11[7] , \nOut18_11[6] , 
        \nOut18_11[5] , \nOut18_11[4] , \nOut18_11[3] , \nOut18_11[2] , 
        \nOut18_11[1] , \nOut18_11[0] }), .WestIn({\nOut16_11[7] , 
        \nOut16_11[6] , \nOut16_11[5] , \nOut16_11[4] , \nOut16_11[3] , 
        \nOut16_11[2] , \nOut16_11[1] , \nOut16_11[0] }), .Out({\nOut17_11[7] , 
        \nOut17_11[6] , \nOut17_11[5] , \nOut17_11[4] , \nOut17_11[3] , 
        \nOut17_11[2] , \nOut17_11[1] , \nOut17_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_572 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut573[7] , \nScanOut573[6] , 
        \nScanOut573[5] , \nScanOut573[4] , \nScanOut573[3] , \nScanOut573[2] , 
        \nScanOut573[1] , \nScanOut573[0] }), .ScanOut({\nScanOut572[7] , 
        \nScanOut572[6] , \nScanOut572[5] , \nScanOut572[4] , \nScanOut572[3] , 
        \nScanOut572[2] , \nScanOut572[1] , \nScanOut572[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_27[7] , \nOut17_27[6] , \nOut17_27[5] , \nOut17_27[4] , 
        \nOut17_27[3] , \nOut17_27[2] , \nOut17_27[1] , \nOut17_27[0] }), 
        .SouthIn({\nOut17_29[7] , \nOut17_29[6] , \nOut17_29[5] , 
        \nOut17_29[4] , \nOut17_29[3] , \nOut17_29[2] , \nOut17_29[1] , 
        \nOut17_29[0] }), .EastIn({\nOut18_28[7] , \nOut18_28[6] , 
        \nOut18_28[5] , \nOut18_28[4] , \nOut18_28[3] , \nOut18_28[2] , 
        \nOut18_28[1] , \nOut18_28[0] }), .WestIn({\nOut16_28[7] , 
        \nOut16_28[6] , \nOut16_28[5] , \nOut16_28[4] , \nOut16_28[3] , 
        \nOut16_28[2] , \nOut16_28[1] , \nOut16_28[0] }), .Out({\nOut17_28[7] , 
        \nOut17_28[6] , \nOut17_28[5] , \nOut17_28[4] , \nOut17_28[3] , 
        \nOut17_28[2] , \nOut17_28[1] , \nOut17_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_890 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut891[7] , \nScanOut891[6] , 
        \nScanOut891[5] , \nScanOut891[4] , \nScanOut891[3] , \nScanOut891[2] , 
        \nScanOut891[1] , \nScanOut891[0] }), .ScanOut({\nScanOut890[7] , 
        \nScanOut890[6] , \nScanOut890[5] , \nScanOut890[4] , \nScanOut890[3] , 
        \nScanOut890[2] , \nScanOut890[1] , \nScanOut890[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_25[7] , \nOut27_25[6] , \nOut27_25[5] , \nOut27_25[4] , 
        \nOut27_25[3] , \nOut27_25[2] , \nOut27_25[1] , \nOut27_25[0] }), 
        .SouthIn({\nOut27_27[7] , \nOut27_27[6] , \nOut27_27[5] , 
        \nOut27_27[4] , \nOut27_27[3] , \nOut27_27[2] , \nOut27_27[1] , 
        \nOut27_27[0] }), .EastIn({\nOut28_26[7] , \nOut28_26[6] , 
        \nOut28_26[5] , \nOut28_26[4] , \nOut28_26[3] , \nOut28_26[2] , 
        \nOut28_26[1] , \nOut28_26[0] }), .WestIn({\nOut26_26[7] , 
        \nOut26_26[6] , \nOut26_26[5] , \nOut26_26[4] , \nOut26_26[3] , 
        \nOut26_26[2] , \nOut26_26[1] , \nOut26_26[0] }), .Out({\nOut27_26[7] , 
        \nOut27_26[6] , \nOut27_26[5] , \nOut27_26[4] , \nOut27_26[3] , 
        \nOut27_26[2] , \nOut27_26[1] , \nOut27_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_900 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut901[7] , \nScanOut901[6] , 
        \nScanOut901[5] , \nScanOut901[4] , \nScanOut901[3] , \nScanOut901[2] , 
        \nScanOut901[1] , \nScanOut901[0] }), .ScanOut({\nScanOut900[7] , 
        \nScanOut900[6] , \nScanOut900[5] , \nScanOut900[4] , \nScanOut900[3] , 
        \nScanOut900[2] , \nScanOut900[1] , \nScanOut900[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_3[7] , \nOut28_3[6] , \nOut28_3[5] , \nOut28_3[4] , 
        \nOut28_3[3] , \nOut28_3[2] , \nOut28_3[1] , \nOut28_3[0] }), 
        .SouthIn({\nOut28_5[7] , \nOut28_5[6] , \nOut28_5[5] , \nOut28_5[4] , 
        \nOut28_5[3] , \nOut28_5[2] , \nOut28_5[1] , \nOut28_5[0] }), .EastIn(
        {\nOut29_4[7] , \nOut29_4[6] , \nOut29_4[5] , \nOut29_4[4] , 
        \nOut29_4[3] , \nOut29_4[2] , \nOut29_4[1] , \nOut29_4[0] }), .WestIn(
        {\nOut27_4[7] , \nOut27_4[6] , \nOut27_4[5] , \nOut27_4[4] , 
        \nOut27_4[3] , \nOut27_4[2] , \nOut27_4[1] , \nOut27_4[0] }), .Out({
        \nOut28_4[7] , \nOut28_4[6] , \nOut28_4[5] , \nOut28_4[4] , 
        \nOut28_4[3] , \nOut28_4[2] , \nOut28_4[1] , \nOut28_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_153 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut154[7] , \nScanOut154[6] , 
        \nScanOut154[5] , \nScanOut154[4] , \nScanOut154[3] , \nScanOut154[2] , 
        \nScanOut154[1] , \nScanOut154[0] }), .ScanOut({\nScanOut153[7] , 
        \nScanOut153[6] , \nScanOut153[5] , \nScanOut153[4] , \nScanOut153[3] , 
        \nScanOut153[2] , \nScanOut153[1] , \nScanOut153[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_24[7] , \nOut4_24[6] , \nOut4_24[5] , \nOut4_24[4] , 
        \nOut4_24[3] , \nOut4_24[2] , \nOut4_24[1] , \nOut4_24[0] }), 
        .SouthIn({\nOut4_26[7] , \nOut4_26[6] , \nOut4_26[5] , \nOut4_26[4] , 
        \nOut4_26[3] , \nOut4_26[2] , \nOut4_26[1] , \nOut4_26[0] }), .EastIn(
        {\nOut5_25[7] , \nOut5_25[6] , \nOut5_25[5] , \nOut5_25[4] , 
        \nOut5_25[3] , \nOut5_25[2] , \nOut5_25[1] , \nOut5_25[0] }), .WestIn(
        {\nOut3_25[7] , \nOut3_25[6] , \nOut3_25[5] , \nOut3_25[4] , 
        \nOut3_25[3] , \nOut3_25[2] , \nOut3_25[1] , \nOut3_25[0] }), .Out({
        \nOut4_25[7] , \nOut4_25[6] , \nOut4_25[5] , \nOut4_25[4] , 
        \nOut4_25[3] , \nOut4_25[2] , \nOut4_25[1] , \nOut4_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_378 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut379[7] , \nScanOut379[6] , 
        \nScanOut379[5] , \nScanOut379[4] , \nScanOut379[3] , \nScanOut379[2] , 
        \nScanOut379[1] , \nScanOut379[0] }), .ScanOut({\nScanOut378[7] , 
        \nScanOut378[6] , \nScanOut378[5] , \nScanOut378[4] , \nScanOut378[3] , 
        \nScanOut378[2] , \nScanOut378[1] , \nScanOut378[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_25[7] , \nOut11_25[6] , \nOut11_25[5] , \nOut11_25[4] , 
        \nOut11_25[3] , \nOut11_25[2] , \nOut11_25[1] , \nOut11_25[0] }), 
        .SouthIn({\nOut11_27[7] , \nOut11_27[6] , \nOut11_27[5] , 
        \nOut11_27[4] , \nOut11_27[3] , \nOut11_27[2] , \nOut11_27[1] , 
        \nOut11_27[0] }), .EastIn({\nOut12_26[7] , \nOut12_26[6] , 
        \nOut12_26[5] , \nOut12_26[4] , \nOut12_26[3] , \nOut12_26[2] , 
        \nOut12_26[1] , \nOut12_26[0] }), .WestIn({\nOut10_26[7] , 
        \nOut10_26[6] , \nOut10_26[5] , \nOut10_26[4] , \nOut10_26[3] , 
        \nOut10_26[2] , \nOut10_26[1] , \nOut10_26[0] }), .Out({\nOut11_26[7] , 
        \nOut11_26[6] , \nOut11_26[5] , \nOut11_26[4] , \nOut11_26[3] , 
        \nOut11_26[2] , \nOut11_26[1] , \nOut11_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_569 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut570[7] , \nScanOut570[6] , 
        \nScanOut570[5] , \nScanOut570[4] , \nScanOut570[3] , \nScanOut570[2] , 
        \nScanOut570[1] , \nScanOut570[0] }), .ScanOut({\nScanOut569[7] , 
        \nScanOut569[6] , \nScanOut569[5] , \nScanOut569[4] , \nScanOut569[3] , 
        \nScanOut569[2] , \nScanOut569[1] , \nScanOut569[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_24[7] , \nOut17_24[6] , \nOut17_24[5] , \nOut17_24[4] , 
        \nOut17_24[3] , \nOut17_24[2] , \nOut17_24[1] , \nOut17_24[0] }), 
        .SouthIn({\nOut17_26[7] , \nOut17_26[6] , \nOut17_26[5] , 
        \nOut17_26[4] , \nOut17_26[3] , \nOut17_26[2] , \nOut17_26[1] , 
        \nOut17_26[0] }), .EastIn({\nOut18_25[7] , \nOut18_25[6] , 
        \nOut18_25[5] , \nOut18_25[4] , \nOut18_25[3] , \nOut18_25[2] , 
        \nOut18_25[1] , \nOut18_25[0] }), .WestIn({\nOut16_25[7] , 
        \nOut16_25[6] , \nOut16_25[5] , \nOut16_25[4] , \nOut16_25[3] , 
        \nOut16_25[2] , \nOut16_25[1] , \nOut16_25[0] }), .Out({\nOut17_25[7] , 
        \nOut17_25[6] , \nOut17_25[5] , \nOut17_25[4] , \nOut17_25[3] , 
        \nOut17_25[2] , \nOut17_25[1] , \nOut17_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_642 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut643[7] , \nScanOut643[6] , 
        \nScanOut643[5] , \nScanOut643[4] , \nScanOut643[3] , \nScanOut643[2] , 
        \nScanOut643[1] , \nScanOut643[0] }), .ScanOut({\nScanOut642[7] , 
        \nScanOut642[6] , \nScanOut642[5] , \nScanOut642[4] , \nScanOut642[3] , 
        \nScanOut642[2] , \nScanOut642[1] , \nScanOut642[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_1[7] , \nOut20_1[6] , \nOut20_1[5] , \nOut20_1[4] , 
        \nOut20_1[3] , \nOut20_1[2] , \nOut20_1[1] , \nOut20_1[0] }), 
        .SouthIn({\nOut20_3[7] , \nOut20_3[6] , \nOut20_3[5] , \nOut20_3[4] , 
        \nOut20_3[3] , \nOut20_3[2] , \nOut20_3[1] , \nOut20_3[0] }), .EastIn(
        {\nOut21_2[7] , \nOut21_2[6] , \nOut21_2[5] , \nOut21_2[4] , 
        \nOut21_2[3] , \nOut21_2[2] , \nOut21_2[1] , \nOut21_2[0] }), .WestIn(
        {\nOut19_2[7] , \nOut19_2[6] , \nOut19_2[5] , \nOut19_2[4] , 
        \nOut19_2[3] , \nOut19_2[2] , \nOut19_2[1] , \nOut19_2[0] }), .Out({
        \nOut20_2[7] , \nOut20_2[6] , \nOut20_2[5] , \nOut20_2[4] , 
        \nOut20_2[3] , \nOut20_2[2] , \nOut20_2[1] , \nOut20_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_659 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut660[7] , \nScanOut660[6] , 
        \nScanOut660[5] , \nScanOut660[4] , \nScanOut660[3] , \nScanOut660[2] , 
        \nScanOut660[1] , \nScanOut660[0] }), .ScanOut({\nScanOut659[7] , 
        \nScanOut659[6] , \nScanOut659[5] , \nScanOut659[4] , \nScanOut659[3] , 
        \nScanOut659[2] , \nScanOut659[1] , \nScanOut659[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_18[7] , \nOut20_18[6] , \nOut20_18[5] , \nOut20_18[4] , 
        \nOut20_18[3] , \nOut20_18[2] , \nOut20_18[1] , \nOut20_18[0] }), 
        .SouthIn({\nOut20_20[7] , \nOut20_20[6] , \nOut20_20[5] , 
        \nOut20_20[4] , \nOut20_20[3] , \nOut20_20[2] , \nOut20_20[1] , 
        \nOut20_20[0] }), .EastIn({\nOut21_19[7] , \nOut21_19[6] , 
        \nOut21_19[5] , \nOut21_19[4] , \nOut21_19[3] , \nOut21_19[2] , 
        \nOut21_19[1] , \nOut21_19[0] }), .WestIn({\nOut19_19[7] , 
        \nOut19_19[6] , \nOut19_19[5] , \nOut19_19[4] , \nOut19_19[3] , 
        \nOut19_19[2] , \nOut19_19[1] , \nOut19_19[0] }), .Out({\nOut20_19[7] , 
        \nOut20_19[6] , \nOut20_19[5] , \nOut20_19[4] , \nOut20_19[3] , 
        \nOut20_19[2] , \nOut20_19[1] , \nOut20_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_174 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut175[7] , \nScanOut175[6] , 
        \nScanOut175[5] , \nScanOut175[4] , \nScanOut175[3] , \nScanOut175[2] , 
        \nScanOut175[1] , \nScanOut175[0] }), .ScanOut({\nScanOut174[7] , 
        \nScanOut174[6] , \nScanOut174[5] , \nScanOut174[4] , \nScanOut174[3] , 
        \nScanOut174[2] , \nScanOut174[1] , \nScanOut174[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }), 
        .SouthIn({\nOut5_15[7] , \nOut5_15[6] , \nOut5_15[5] , \nOut5_15[4] , 
        \nOut5_15[3] , \nOut5_15[2] , \nOut5_15[1] , \nOut5_15[0] }), .EastIn(
        {\nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }), .WestIn(
        {\nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }), .Out({
        \nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_244 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut245[7] , \nScanOut245[6] , 
        \nScanOut245[5] , \nScanOut245[4] , \nScanOut245[3] , \nScanOut245[2] , 
        \nScanOut245[1] , \nScanOut245[0] }), .ScanOut({\nScanOut244[7] , 
        \nScanOut244[6] , \nScanOut244[5] , \nScanOut244[4] , \nScanOut244[3] , 
        \nScanOut244[2] , \nScanOut244[1] , \nScanOut244[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_19[7] , \nOut7_19[6] , \nOut7_19[5] , \nOut7_19[4] , 
        \nOut7_19[3] , \nOut7_19[2] , \nOut7_19[1] , \nOut7_19[0] }), 
        .SouthIn({\nOut7_21[7] , \nOut7_21[6] , \nOut7_21[5] , \nOut7_21[4] , 
        \nOut7_21[3] , \nOut7_21[2] , \nOut7_21[1] , \nOut7_21[0] }), .EastIn(
        {\nOut8_20[7] , \nOut8_20[6] , \nOut8_20[5] , \nOut8_20[4] , 
        \nOut8_20[3] , \nOut8_20[2] , \nOut8_20[1] , \nOut8_20[0] }), .WestIn(
        {\nOut6_20[7] , \nOut6_20[6] , \nOut6_20[5] , \nOut6_20[4] , 
        \nOut6_20[3] , \nOut6_20[2] , \nOut6_20[1] , \nOut6_20[0] }), .Out({
        \nOut7_20[7] , \nOut7_20[6] , \nOut7_20[5] , \nOut7_20[4] , 
        \nOut7_20[3] , \nOut7_20[2] , \nOut7_20[1] , \nOut7_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_263 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut264[7] , \nScanOut264[6] , 
        \nScanOut264[5] , \nScanOut264[4] , \nScanOut264[3] , \nScanOut264[2] , 
        \nScanOut264[1] , \nScanOut264[0] }), .ScanOut({\nScanOut263[7] , 
        \nScanOut263[6] , \nScanOut263[5] , \nScanOut263[4] , \nScanOut263[3] , 
        \nScanOut263[2] , \nScanOut263[1] , \nScanOut263[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_6[7] , \nOut8_6[6] , \nOut8_6[5] , \nOut8_6[4] , \nOut8_6[3] , 
        \nOut8_6[2] , \nOut8_6[1] , \nOut8_6[0] }), .SouthIn({\nOut8_8[7] , 
        \nOut8_8[6] , \nOut8_8[5] , \nOut8_8[4] , \nOut8_8[3] , \nOut8_8[2] , 
        \nOut8_8[1] , \nOut8_8[0] }), .EastIn({\nOut9_7[7] , \nOut9_7[6] , 
        \nOut9_7[5] , \nOut9_7[4] , \nOut9_7[3] , \nOut9_7[2] , \nOut9_7[1] , 
        \nOut9_7[0] }), .WestIn({\nOut7_7[7] , \nOut7_7[6] , \nOut7_7[5] , 
        \nOut7_7[4] , \nOut7_7[3] , \nOut7_7[2] , \nOut7_7[1] , \nOut7_7[0] }), 
        .Out({\nOut8_7[7] , \nOut8_7[6] , \nOut8_7[5] , \nOut8_7[4] , 
        \nOut8_7[3] , \nOut8_7[2] , \nOut8_7[1] , \nOut8_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_742 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut743[7] , \nScanOut743[6] , 
        \nScanOut743[5] , \nScanOut743[4] , \nScanOut743[3] , \nScanOut743[2] , 
        \nScanOut743[1] , \nScanOut743[0] }), .ScanOut({\nScanOut742[7] , 
        \nScanOut742[6] , \nScanOut742[5] , \nScanOut742[4] , \nScanOut742[3] , 
        \nScanOut742[2] , \nScanOut742[1] , \nScanOut742[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_5[7] , \nOut23_5[6] , \nOut23_5[5] , \nOut23_5[4] , 
        \nOut23_5[3] , \nOut23_5[2] , \nOut23_5[1] , \nOut23_5[0] }), 
        .SouthIn({\nOut23_7[7] , \nOut23_7[6] , \nOut23_7[5] , \nOut23_7[4] , 
        \nOut23_7[3] , \nOut23_7[2] , \nOut23_7[1] , \nOut23_7[0] }), .EastIn(
        {\nOut24_6[7] , \nOut24_6[6] , \nOut24_6[5] , \nOut24_6[4] , 
        \nOut24_6[3] , \nOut24_6[2] , \nOut24_6[1] , \nOut24_6[0] }), .WestIn(
        {\nOut22_6[7] , \nOut22_6[6] , \nOut22_6[5] , \nOut22_6[4] , 
        \nOut22_6[3] , \nOut22_6[2] , \nOut22_6[1] , \nOut22_6[0] }), .Out({
        \nOut23_6[7] , \nOut23_6[6] , \nOut23_6[5] , \nOut23_6[4] , 
        \nOut23_6[3] , \nOut23_6[2] , \nOut23_6[1] , \nOut23_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_800 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut801[7] , \nScanOut801[6] , 
        \nScanOut801[5] , \nScanOut801[4] , \nScanOut801[3] , \nScanOut801[2] , 
        \nScanOut801[1] , \nScanOut801[0] }), .ScanOut({\nScanOut800[7] , 
        \nScanOut800[6] , \nScanOut800[5] , \nScanOut800[4] , \nScanOut800[3] , 
        \nScanOut800[2] , \nScanOut800[1] , \nScanOut800[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut25_0[7] , \nOut25_0[6] , 
        \nOut25_0[5] , \nOut25_0[4] , \nOut25_0[3] , \nOut25_0[2] , 
        \nOut25_0[1] , \nOut25_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_990 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut991[7] , \nScanOut991[6] , 
        \nScanOut991[5] , \nScanOut991[4] , \nScanOut991[3] , \nScanOut991[2] , 
        \nScanOut991[1] , \nScanOut991[0] }), .ScanOut({\nScanOut990[7] , 
        \nScanOut990[6] , \nScanOut990[5] , \nScanOut990[4] , \nScanOut990[3] , 
        \nScanOut990[2] , \nScanOut990[1] , \nScanOut990[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_29[7] , \nOut30_29[6] , \nOut30_29[5] , \nOut30_29[4] , 
        \nOut30_29[3] , \nOut30_29[2] , \nOut30_29[1] , \nOut30_29[0] }), 
        .SouthIn({\nOut30_31[7] , \nOut30_31[6] , \nOut30_31[5] , 
        \nOut30_31[4] , \nOut30_31[3] , \nOut30_31[2] , \nOut30_31[1] , 
        \nOut30_31[0] }), .EastIn({\nOut31_30[7] , \nOut31_30[6] , 
        \nOut31_30[5] , \nOut31_30[4] , \nOut31_30[3] , \nOut31_30[2] , 
        \nOut31_30[1] , \nOut31_30[0] }), .WestIn({\nOut29_30[7] , 
        \nOut29_30[6] , \nOut29_30[5] , \nOut29_30[4] , \nOut29_30[3] , 
        \nOut29_30[2] , \nOut29_30[1] , \nOut29_30[0] }), .Out({\nOut30_30[7] , 
        \nOut30_30[6] , \nOut30_30[5] , \nOut30_30[4] , \nOut30_30[3] , 
        \nOut30_30[2] , \nOut30_30[1] , \nOut30_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_455 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut456[7] , \nScanOut456[6] , 
        \nScanOut456[5] , \nScanOut456[4] , \nScanOut456[3] , \nScanOut456[2] , 
        \nScanOut456[1] , \nScanOut456[0] }), .ScanOut({\nScanOut455[7] , 
        \nScanOut455[6] , \nScanOut455[5] , \nScanOut455[4] , \nScanOut455[3] , 
        \nScanOut455[2] , \nScanOut455[1] , \nScanOut455[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }), 
        .SouthIn({\nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }), .EastIn(
        {\nOut15_7[7] , \nOut15_7[6] , \nOut15_7[5] , \nOut15_7[4] , 
        \nOut15_7[3] , \nOut15_7[2] , \nOut15_7[1] , \nOut15_7[0] }), .WestIn(
        {\nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }), .Out({
        \nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_472 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut473[7] , \nScanOut473[6] , 
        \nScanOut473[5] , \nScanOut473[4] , \nScanOut473[3] , \nScanOut473[2] , 
        \nScanOut473[1] , \nScanOut473[0] }), .ScanOut({\nScanOut472[7] , 
        \nScanOut472[6] , \nScanOut472[5] , \nScanOut472[4] , \nScanOut472[3] , 
        \nScanOut472[2] , \nScanOut472[1] , \nScanOut472[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_23[7] , \nOut14_23[6] , \nOut14_23[5] , \nOut14_23[4] , 
        \nOut14_23[3] , \nOut14_23[2] , \nOut14_23[1] , \nOut14_23[0] }), 
        .SouthIn({\nOut14_25[7] , \nOut14_25[6] , \nOut14_25[5] , 
        \nOut14_25[4] , \nOut14_25[3] , \nOut14_25[2] , \nOut14_25[1] , 
        \nOut14_25[0] }), .EastIn({\nOut15_24[7] , \nOut15_24[6] , 
        \nOut15_24[5] , \nOut15_24[4] , \nOut15_24[3] , \nOut15_24[2] , 
        \nOut15_24[1] , \nOut15_24[0] }), .WestIn({\nOut13_24[7] , 
        \nOut13_24[6] , \nOut13_24[5] , \nOut13_24[4] , \nOut13_24[3] , 
        \nOut13_24[2] , \nOut13_24[1] , \nOut13_24[0] }), .Out({\nOut14_24[7] , 
        \nOut14_24[6] , \nOut14_24[5] , \nOut14_24[4] , \nOut14_24[3] , 
        \nOut14_24[2] , \nOut14_24[1] , \nOut14_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_827 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut828[7] , \nScanOut828[6] , 
        \nScanOut828[5] , \nScanOut828[4] , \nScanOut828[3] , \nScanOut828[2] , 
        \nScanOut828[1] , \nScanOut828[0] }), .ScanOut({\nScanOut827[7] , 
        \nScanOut827[6] , \nScanOut827[5] , \nScanOut827[4] , \nScanOut827[3] , 
        \nScanOut827[2] , \nScanOut827[1] , \nScanOut827[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_26[7] , \nOut25_26[6] , \nOut25_26[5] , \nOut25_26[4] , 
        \nOut25_26[3] , \nOut25_26[2] , \nOut25_26[1] , \nOut25_26[0] }), 
        .SouthIn({\nOut25_28[7] , \nOut25_28[6] , \nOut25_28[5] , 
        \nOut25_28[4] , \nOut25_28[3] , \nOut25_28[2] , \nOut25_28[1] , 
        \nOut25_28[0] }), .EastIn({\nOut26_27[7] , \nOut26_27[6] , 
        \nOut26_27[5] , \nOut26_27[4] , \nOut26_27[3] , \nOut26_27[2] , 
        \nOut26_27[1] , \nOut26_27[0] }), .WestIn({\nOut24_27[7] , 
        \nOut24_27[6] , \nOut24_27[5] , \nOut24_27[4] , \nOut24_27[3] , 
        \nOut24_27[2] , \nOut24_27[1] , \nOut24_27[0] }), .Out({\nOut25_27[7] , 
        \nOut25_27[6] , \nOut25_27[5] , \nOut25_27[4] , \nOut25_27[3] , 
        \nOut25_27[2] , \nOut25_27[1] , \nOut25_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_765 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut766[7] , \nScanOut766[6] , 
        \nScanOut766[5] , \nScanOut766[4] , \nScanOut766[3] , \nScanOut766[2] , 
        \nScanOut766[1] , \nScanOut766[0] }), .ScanOut({\nScanOut765[7] , 
        \nScanOut765[6] , \nScanOut765[5] , \nScanOut765[4] , \nScanOut765[3] , 
        \nScanOut765[2] , \nScanOut765[1] , \nScanOut765[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_28[7] , \nOut23_28[6] , \nOut23_28[5] , \nOut23_28[4] , 
        \nOut23_28[3] , \nOut23_28[2] , \nOut23_28[1] , \nOut23_28[0] }), 
        .SouthIn({\nOut23_30[7] , \nOut23_30[6] , \nOut23_30[5] , 
        \nOut23_30[4] , \nOut23_30[3] , \nOut23_30[2] , \nOut23_30[1] , 
        \nOut23_30[0] }), .EastIn({\nOut24_29[7] , \nOut24_29[6] , 
        \nOut24_29[5] , \nOut24_29[4] , \nOut24_29[3] , \nOut24_29[2] , 
        \nOut24_29[1] , \nOut24_29[0] }), .WestIn({\nOut22_29[7] , 
        \nOut22_29[6] , \nOut22_29[5] , \nOut22_29[4] , \nOut22_29[3] , 
        \nOut22_29[2] , \nOut22_29[1] , \nOut22_29[0] }), .Out({\nOut23_29[7] , 
        \nOut23_29[6] , \nOut23_29[5] , \nOut23_29[4] , \nOut23_29[3] , 
        \nOut23_29[2] , \nOut23_29[1] , \nOut23_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_191 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut192[7] , \nScanOut192[6] , 
        \nScanOut192[5] , \nScanOut192[4] , \nScanOut192[3] , \nScanOut192[2] , 
        \nScanOut192[1] , \nScanOut192[0] }), .ScanOut({\nScanOut191[7] , 
        \nScanOut191[6] , \nScanOut191[5] , \nScanOut191[4] , \nScanOut191[3] , 
        \nScanOut191[2] , \nScanOut191[1] , \nScanOut191[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut5_31[7] , \nOut5_31[6] , 
        \nOut5_31[5] , \nOut5_31[4] , \nOut5_31[3] , \nOut5_31[2] , 
        \nOut5_31[1] , \nOut5_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_331 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut332[7] , \nScanOut332[6] , 
        \nScanOut332[5] , \nScanOut332[4] , \nScanOut332[3] , \nScanOut332[2] , 
        \nScanOut332[1] , \nScanOut332[0] }), .ScanOut({\nScanOut331[7] , 
        \nScanOut331[6] , \nScanOut331[5] , \nScanOut331[4] , \nScanOut331[3] , 
        \nScanOut331[2] , \nScanOut331[1] , \nScanOut331[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_10[7] , \nOut10_10[6] , \nOut10_10[5] , \nOut10_10[4] , 
        \nOut10_10[3] , \nOut10_10[2] , \nOut10_10[1] , \nOut10_10[0] }), 
        .SouthIn({\nOut10_12[7] , \nOut10_12[6] , \nOut10_12[5] , 
        \nOut10_12[4] , \nOut10_12[3] , \nOut10_12[2] , \nOut10_12[1] , 
        \nOut10_12[0] }), .EastIn({\nOut11_11[7] , \nOut11_11[6] , 
        \nOut11_11[5] , \nOut11_11[4] , \nOut11_11[3] , \nOut11_11[2] , 
        \nOut11_11[1] , \nOut11_11[0] }), .WestIn({\nOut9_11[7] , 
        \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , \nOut9_11[3] , 
        \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }), .Out({\nOut10_11[7] , 
        \nOut10_11[6] , \nOut10_11[5] , \nOut10_11[4] , \nOut10_11[3] , 
        \nOut10_11[2] , \nOut10_11[1] , \nOut10_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_520 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut521[7] , \nScanOut521[6] , 
        \nScanOut521[5] , \nScanOut521[4] , \nScanOut521[3] , \nScanOut521[2] , 
        \nScanOut521[1] , \nScanOut521[0] }), .ScanOut({\nScanOut520[7] , 
        \nScanOut520[6] , \nScanOut520[5] , \nScanOut520[4] , \nScanOut520[3] , 
        \nScanOut520[2] , \nScanOut520[1] , \nScanOut520[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_7[7] , \nOut16_7[6] , \nOut16_7[5] , \nOut16_7[4] , 
        \nOut16_7[3] , \nOut16_7[2] , \nOut16_7[1] , \nOut16_7[0] }), 
        .SouthIn({\nOut16_9[7] , \nOut16_9[6] , \nOut16_9[5] , \nOut16_9[4] , 
        \nOut16_9[3] , \nOut16_9[2] , \nOut16_9[1] , \nOut16_9[0] }), .EastIn(
        {\nOut17_8[7] , \nOut17_8[6] , \nOut17_8[5] , \nOut17_8[4] , 
        \nOut17_8[3] , \nOut17_8[2] , \nOut17_8[1] , \nOut17_8[0] }), .WestIn(
        {\nOut15_8[7] , \nOut15_8[6] , \nOut15_8[5] , \nOut15_8[4] , 
        \nOut15_8[3] , \nOut15_8[2] , \nOut15_8[1] , \nOut15_8[0] }), .Out({
        \nOut16_8[7] , \nOut16_8[6] , \nOut16_8[5] , \nOut16_8[4] , 
        \nOut16_8[3] , \nOut16_8[2] , \nOut16_8[1] , \nOut16_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_849 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut850[7] , \nScanOut850[6] , 
        \nScanOut850[5] , \nScanOut850[4] , \nScanOut850[3] , \nScanOut850[2] , 
        \nScanOut850[1] , \nScanOut850[0] }), .ScanOut({\nScanOut849[7] , 
        \nScanOut849[6] , \nScanOut849[5] , \nScanOut849[4] , \nScanOut849[3] , 
        \nScanOut849[2] , \nScanOut849[1] , \nScanOut849[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_16[7] , \nOut26_16[6] , \nOut26_16[5] , \nOut26_16[4] , 
        \nOut26_16[3] , \nOut26_16[2] , \nOut26_16[1] , \nOut26_16[0] }), 
        .SouthIn({\nOut26_18[7] , \nOut26_18[6] , \nOut26_18[5] , 
        \nOut26_18[4] , \nOut26_18[3] , \nOut26_18[2] , \nOut26_18[1] , 
        \nOut26_18[0] }), .EastIn({\nOut27_17[7] , \nOut27_17[6] , 
        \nOut27_17[5] , \nOut27_17[4] , \nOut27_17[3] , \nOut27_17[2] , 
        \nOut27_17[1] , \nOut27_17[0] }), .WestIn({\nOut25_17[7] , 
        \nOut25_17[6] , \nOut25_17[5] , \nOut25_17[4] , \nOut25_17[3] , 
        \nOut25_17[2] , \nOut25_17[1] , \nOut25_17[0] }), .Out({\nOut26_17[7] , 
        \nOut26_17[6] , \nOut26_17[5] , \nOut26_17[4] , \nOut26_17[3] , 
        \nOut26_17[2] , \nOut26_17[1] , \nOut26_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_952 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut953[7] , \nScanOut953[6] , 
        \nScanOut953[5] , \nScanOut953[4] , \nScanOut953[3] , \nScanOut953[2] , 
        \nScanOut953[1] , \nScanOut953[0] }), .ScanOut({\nScanOut952[7] , 
        \nScanOut952[6] , \nScanOut952[5] , \nScanOut952[4] , \nScanOut952[3] , 
        \nScanOut952[2] , \nScanOut952[1] , \nScanOut952[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_23[7] , \nOut29_23[6] , \nOut29_23[5] , \nOut29_23[4] , 
        \nOut29_23[3] , \nOut29_23[2] , \nOut29_23[1] , \nOut29_23[0] }), 
        .SouthIn({\nOut29_25[7] , \nOut29_25[6] , \nOut29_25[5] , 
        \nOut29_25[4] , \nOut29_25[3] , \nOut29_25[2] , \nOut29_25[1] , 
        \nOut29_25[0] }), .EastIn({\nOut30_24[7] , \nOut30_24[6] , 
        \nOut30_24[5] , \nOut30_24[4] , \nOut30_24[3] , \nOut30_24[2] , 
        \nOut30_24[1] , \nOut30_24[0] }), .WestIn({\nOut28_24[7] , 
        \nOut28_24[6] , \nOut28_24[5] , \nOut28_24[4] , \nOut28_24[3] , 
        \nOut28_24[2] , \nOut28_24[1] , \nOut28_24[0] }), .Out({\nOut29_24[7] , 
        \nOut29_24[6] , \nOut29_24[5] , \nOut29_24[4] , \nOut29_24[3] , 
        \nOut29_24[2] , \nOut29_24[1] , \nOut29_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_610 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut611[7] , \nScanOut611[6] , 
        \nScanOut611[5] , \nScanOut611[4] , \nScanOut611[3] , \nScanOut611[2] , 
        \nScanOut611[1] , \nScanOut611[0] }), .ScanOut({\nScanOut610[7] , 
        \nScanOut610[6] , \nScanOut610[5] , \nScanOut610[4] , \nScanOut610[3] , 
        \nScanOut610[2] , \nScanOut610[1] , \nScanOut610[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_1[7] , \nOut19_1[6] , \nOut19_1[5] , \nOut19_1[4] , 
        \nOut19_1[3] , \nOut19_1[2] , \nOut19_1[1] , \nOut19_1[0] }), 
        .SouthIn({\nOut19_3[7] , \nOut19_3[6] , \nOut19_3[5] , \nOut19_3[4] , 
        \nOut19_3[3] , \nOut19_3[2] , \nOut19_3[1] , \nOut19_3[0] }), .EastIn(
        {\nOut20_2[7] , \nOut20_2[6] , \nOut20_2[5] , \nOut20_2[4] , 
        \nOut20_2[3] , \nOut20_2[2] , \nOut20_2[1] , \nOut20_2[0] }), .WestIn(
        {\nOut18_2[7] , \nOut18_2[6] , \nOut18_2[5] , \nOut18_2[4] , 
        \nOut18_2[3] , \nOut18_2[2] , \nOut18_2[1] , \nOut18_2[0] }), .Out({
        \nOut19_2[7] , \nOut19_2[6] , \nOut19_2[5] , \nOut19_2[4] , 
        \nOut19_2[3] , \nOut19_2[2] , \nOut19_2[1] , \nOut19_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_637 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut638[7] , \nScanOut638[6] , 
        \nScanOut638[5] , \nScanOut638[4] , \nScanOut638[3] , \nScanOut638[2] , 
        \nScanOut638[1] , \nScanOut638[0] }), .ScanOut({\nScanOut637[7] , 
        \nScanOut637[6] , \nScanOut637[5] , \nScanOut637[4] , \nScanOut637[3] , 
        \nScanOut637[2] , \nScanOut637[1] , \nScanOut637[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_28[7] , \nOut19_28[6] , \nOut19_28[5] , \nOut19_28[4] , 
        \nOut19_28[3] , \nOut19_28[2] , \nOut19_28[1] , \nOut19_28[0] }), 
        .SouthIn({\nOut19_30[7] , \nOut19_30[6] , \nOut19_30[5] , 
        \nOut19_30[4] , \nOut19_30[3] , \nOut19_30[2] , \nOut19_30[1] , 
        \nOut19_30[0] }), .EastIn({\nOut20_29[7] , \nOut20_29[6] , 
        \nOut20_29[5] , \nOut20_29[4] , \nOut20_29[3] , \nOut20_29[2] , 
        \nOut20_29[1] , \nOut20_29[0] }), .WestIn({\nOut18_29[7] , 
        \nOut18_29[6] , \nOut18_29[5] , \nOut18_29[4] , \nOut18_29[3] , 
        \nOut18_29[2] , \nOut18_29[1] , \nOut18_29[0] }), .Out({\nOut19_29[7] , 
        \nOut19_29[6] , \nOut19_29[5] , \nOut19_29[4] , \nOut19_29[3] , 
        \nOut19_29[2] , \nOut19_29[1] , \nOut19_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_780 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut781[7] , \nScanOut781[6] , 
        \nScanOut781[5] , \nScanOut781[4] , \nScanOut781[3] , \nScanOut781[2] , 
        \nScanOut781[1] , \nScanOut781[0] }), .ScanOut({\nScanOut780[7] , 
        \nScanOut780[6] , \nScanOut780[5] , \nScanOut780[4] , \nScanOut780[3] , 
        \nScanOut780[2] , \nScanOut780[1] , \nScanOut780[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_11[7] , \nOut24_11[6] , \nOut24_11[5] , \nOut24_11[4] , 
        \nOut24_11[3] , \nOut24_11[2] , \nOut24_11[1] , \nOut24_11[0] }), 
        .SouthIn({\nOut24_13[7] , \nOut24_13[6] , \nOut24_13[5] , 
        \nOut24_13[4] , \nOut24_13[3] , \nOut24_13[2] , \nOut24_13[1] , 
        \nOut24_13[0] }), .EastIn({\nOut25_12[7] , \nOut25_12[6] , 
        \nOut25_12[5] , \nOut25_12[4] , \nOut25_12[3] , \nOut25_12[2] , 
        \nOut25_12[1] , \nOut25_12[0] }), .WestIn({\nOut23_12[7] , 
        \nOut23_12[6] , \nOut23_12[5] , \nOut23_12[4] , \nOut23_12[3] , 
        \nOut23_12[2] , \nOut23_12[1] , \nOut23_12[0] }), .Out({\nOut24_12[7] , 
        \nOut24_12[6] , \nOut24_12[5] , \nOut24_12[4] , \nOut24_12[3] , 
        \nOut24_12[2] , \nOut24_12[1] , \nOut24_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_63 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut64[7] , \nScanOut64[6] , 
        \nScanOut64[5] , \nScanOut64[4] , \nScanOut64[3] , \nScanOut64[2] , 
        \nScanOut64[1] , \nScanOut64[0] }), .ScanOut({\nScanOut63[7] , 
        \nScanOut63[6] , \nScanOut63[5] , \nScanOut63[4] , \nScanOut63[3] , 
        \nScanOut63[2] , \nScanOut63[1] , \nScanOut63[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut1_31[7] , \nOut1_31[6] , 
        \nOut1_31[5] , \nOut1_31[4] , \nOut1_31[3] , \nOut1_31[2] , 
        \nOut1_31[1] , \nOut1_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_86 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut87[7] , \nScanOut87[6] , 
        \nScanOut87[5] , \nScanOut87[4] , \nScanOut87[3] , \nScanOut87[2] , 
        \nScanOut87[1] , \nScanOut87[0] }), .ScanOut({\nScanOut86[7] , 
        \nScanOut86[6] , \nScanOut86[5] , \nScanOut86[4] , \nScanOut86[3] , 
        \nScanOut86[2] , \nScanOut86[1] , \nScanOut86[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_21[7] , \nOut2_21[6] , \nOut2_21[5] , \nOut2_21[4] , 
        \nOut2_21[3] , \nOut2_21[2] , \nOut2_21[1] , \nOut2_21[0] }), 
        .SouthIn({\nOut2_23[7] , \nOut2_23[6] , \nOut2_23[5] , \nOut2_23[4] , 
        \nOut2_23[3] , \nOut2_23[2] , \nOut2_23[1] , \nOut2_23[0] }), .EastIn(
        {\nOut3_22[7] , \nOut3_22[6] , \nOut3_22[5] , \nOut3_22[4] , 
        \nOut3_22[3] , \nOut3_22[2] , \nOut3_22[1] , \nOut3_22[0] }), .WestIn(
        {\nOut1_22[7] , \nOut1_22[6] , \nOut1_22[5] , \nOut1_22[4] , 
        \nOut1_22[3] , \nOut1_22[2] , \nOut1_22[1] , \nOut1_22[0] }), .Out({
        \nOut2_22[7] , \nOut2_22[6] , \nOut2_22[5] , \nOut2_22[4] , 
        \nOut2_22[3] , \nOut2_22[2] , \nOut2_22[1] , \nOut2_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_135 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut136[7] , \nScanOut136[6] , 
        \nScanOut136[5] , \nScanOut136[4] , \nScanOut136[3] , \nScanOut136[2] , 
        \nScanOut136[1] , \nScanOut136[0] }), .ScanOut({\nScanOut135[7] , 
        \nScanOut135[6] , \nScanOut135[5] , \nScanOut135[4] , \nScanOut135[3] , 
        \nScanOut135[2] , \nScanOut135[1] , \nScanOut135[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_6[7] , \nOut4_6[6] , \nOut4_6[5] , \nOut4_6[4] , \nOut4_6[3] , 
        \nOut4_6[2] , \nOut4_6[1] , \nOut4_6[0] }), .SouthIn({\nOut4_8[7] , 
        \nOut4_8[6] , \nOut4_8[5] , \nOut4_8[4] , \nOut4_8[3] , \nOut4_8[2] , 
        \nOut4_8[1] , \nOut4_8[0] }), .EastIn({\nOut5_7[7] , \nOut5_7[6] , 
        \nOut5_7[5] , \nOut5_7[4] , \nOut5_7[3] , \nOut5_7[2] , \nOut5_7[1] , 
        \nOut5_7[0] }), .WestIn({\nOut3_7[7] , \nOut3_7[6] , \nOut3_7[5] , 
        \nOut3_7[4] , \nOut3_7[3] , \nOut3_7[2] , \nOut3_7[1] , \nOut3_7[0] }), 
        .Out({\nOut4_7[7] , \nOut4_7[6] , \nOut4_7[5] , \nOut4_7[4] , 
        \nOut4_7[3] , \nOut4_7[2] , \nOut4_7[1] , \nOut4_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_205 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut206[7] , \nScanOut206[6] , 
        \nScanOut206[5] , \nScanOut206[4] , \nScanOut206[3] , \nScanOut206[2] , 
        \nScanOut206[1] , \nScanOut206[0] }), .ScanOut({\nScanOut205[7] , 
        \nScanOut205[6] , \nScanOut205[5] , \nScanOut205[4] , \nScanOut205[3] , 
        \nScanOut205[2] , \nScanOut205[1] , \nScanOut205[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }), 
        .SouthIn({\nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }), .EastIn(
        {\nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }), .WestIn(
        {\nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }), .Out({
        \nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_286 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut287[7] , \nScanOut287[6] , 
        \nScanOut287[5] , \nScanOut287[4] , \nScanOut287[3] , \nScanOut287[2] , 
        \nScanOut287[1] , \nScanOut287[0] }), .ScanOut({\nScanOut286[7] , 
        \nScanOut286[6] , \nScanOut286[5] , \nScanOut286[4] , \nScanOut286[3] , 
        \nScanOut286[2] , \nScanOut286[1] , \nScanOut286[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_29[7] , \nOut8_29[6] , \nOut8_29[5] , \nOut8_29[4] , 
        \nOut8_29[3] , \nOut8_29[2] , \nOut8_29[1] , \nOut8_29[0] }), 
        .SouthIn({\nOut8_31[7] , \nOut8_31[6] , \nOut8_31[5] , \nOut8_31[4] , 
        \nOut8_31[3] , \nOut8_31[2] , \nOut8_31[1] , \nOut8_31[0] }), .EastIn(
        {\nOut9_30[7] , \nOut9_30[6] , \nOut9_30[5] , \nOut9_30[4] , 
        \nOut9_30[3] , \nOut9_30[2] , \nOut9_30[1] , \nOut9_30[0] }), .WestIn(
        {\nOut7_30[7] , \nOut7_30[6] , \nOut7_30[5] , \nOut7_30[4] , 
        \nOut7_30[3] , \nOut7_30[2] , \nOut7_30[1] , \nOut7_30[0] }), .Out({
        \nOut8_30[7] , \nOut8_30[6] , \nOut8_30[5] , \nOut8_30[4] , 
        \nOut8_30[3] , \nOut8_30[2] , \nOut8_30[1] , \nOut8_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_316 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut317[7] , \nScanOut317[6] , 
        \nScanOut317[5] , \nScanOut317[4] , \nScanOut317[3] , \nScanOut317[2] , 
        \nScanOut317[1] , \nScanOut317[0] }), .ScanOut({\nScanOut316[7] , 
        \nScanOut316[6] , \nScanOut316[5] , \nScanOut316[4] , \nScanOut316[3] , 
        \nScanOut316[2] , \nScanOut316[1] , \nScanOut316[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_27[7] , \nOut9_27[6] , \nOut9_27[5] , \nOut9_27[4] , 
        \nOut9_27[3] , \nOut9_27[2] , \nOut9_27[1] , \nOut9_27[0] }), 
        .SouthIn({\nOut9_29[7] , \nOut9_29[6] , \nOut9_29[5] , \nOut9_29[4] , 
        \nOut9_29[3] , \nOut9_29[2] , \nOut9_29[1] , \nOut9_29[0] }), .EastIn(
        {\nOut10_28[7] , \nOut10_28[6] , \nOut10_28[5] , \nOut10_28[4] , 
        \nOut10_28[3] , \nOut10_28[2] , \nOut10_28[1] , \nOut10_28[0] }), 
        .WestIn({\nOut8_28[7] , \nOut8_28[6] , \nOut8_28[5] , \nOut8_28[4] , 
        \nOut8_28[3] , \nOut8_28[2] , \nOut8_28[1] , \nOut8_28[0] }), .Out({
        \nOut9_28[7] , \nOut9_28[6] , \nOut9_28[5] , \nOut9_28[4] , 
        \nOut9_28[3] , \nOut9_28[2] , \nOut9_28[1] , \nOut9_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_975 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut976[7] , \nScanOut976[6] , 
        \nScanOut976[5] , \nScanOut976[4] , \nScanOut976[3] , \nScanOut976[2] , 
        \nScanOut976[1] , \nScanOut976[0] }), .ScanOut({\nScanOut975[7] , 
        \nScanOut975[6] , \nScanOut975[5] , \nScanOut975[4] , \nScanOut975[3] , 
        \nScanOut975[2] , \nScanOut975[1] , \nScanOut975[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_14[7] , \nOut30_14[6] , \nOut30_14[5] , \nOut30_14[4] , 
        \nOut30_14[3] , \nOut30_14[2] , \nOut30_14[1] , \nOut30_14[0] }), 
        .SouthIn({\nOut30_16[7] , \nOut30_16[6] , \nOut30_16[5] , 
        \nOut30_16[4] , \nOut30_16[3] , \nOut30_16[2] , \nOut30_16[1] , 
        \nOut30_16[0] }), .EastIn({\nOut31_15[7] , \nOut31_15[6] , 
        \nOut31_15[5] , \nOut31_15[4] , \nOut31_15[3] , \nOut31_15[2] , 
        \nOut31_15[1] , \nOut31_15[0] }), .WestIn({\nOut29_15[7] , 
        \nOut29_15[6] , \nOut29_15[5] , \nOut29_15[4] , \nOut29_15[3] , 
        \nOut29_15[2] , \nOut29_15[1] , \nOut29_15[0] }), .Out({\nOut30_15[7] , 
        \nOut30_15[6] , \nOut30_15[5] , \nOut30_15[4] , \nOut30_15[3] , 
        \nOut30_15[2] , \nOut30_15[1] , \nOut30_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_497 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut498[7] , \nScanOut498[6] , 
        \nScanOut498[5] , \nScanOut498[4] , \nScanOut498[3] , \nScanOut498[2] , 
        \nScanOut498[1] , \nScanOut498[0] }), .ScanOut({\nScanOut497[7] , 
        \nScanOut497[6] , \nScanOut497[5] , \nScanOut497[4] , \nScanOut497[3] , 
        \nScanOut497[2] , \nScanOut497[1] , \nScanOut497[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_16[7] , \nOut15_16[6] , \nOut15_16[5] , \nOut15_16[4] , 
        \nOut15_16[3] , \nOut15_16[2] , \nOut15_16[1] , \nOut15_16[0] }), 
        .SouthIn({\nOut15_18[7] , \nOut15_18[6] , \nOut15_18[5] , 
        \nOut15_18[4] , \nOut15_18[3] , \nOut15_18[2] , \nOut15_18[1] , 
        \nOut15_18[0] }), .EastIn({\nOut16_17[7] , \nOut16_17[6] , 
        \nOut16_17[5] , \nOut16_17[4] , \nOut16_17[3] , \nOut16_17[2] , 
        \nOut16_17[1] , \nOut16_17[0] }), .WestIn({\nOut14_17[7] , 
        \nOut14_17[6] , \nOut14_17[5] , \nOut14_17[4] , \nOut14_17[3] , 
        \nOut14_17[2] , \nOut14_17[1] , \nOut14_17[0] }), .Out({\nOut15_17[7] , 
        \nOut15_17[6] , \nOut15_17[5] , \nOut15_17[4] , \nOut15_17[3] , 
        \nOut15_17[2] , \nOut15_17[1] , \nOut15_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_395 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut396[7] , \nScanOut396[6] , 
        \nScanOut396[5] , \nScanOut396[4] , \nScanOut396[3] , \nScanOut396[2] , 
        \nScanOut396[1] , \nScanOut396[0] }), .ScanOut({\nScanOut395[7] , 
        \nScanOut395[6] , \nScanOut395[5] , \nScanOut395[4] , \nScanOut395[3] , 
        \nScanOut395[2] , \nScanOut395[1] , \nScanOut395[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_10[7] , \nOut12_10[6] , \nOut12_10[5] , \nOut12_10[4] , 
        \nOut12_10[3] , \nOut12_10[2] , \nOut12_10[1] , \nOut12_10[0] }), 
        .SouthIn({\nOut12_12[7] , \nOut12_12[6] , \nOut12_12[5] , 
        \nOut12_12[4] , \nOut12_12[3] , \nOut12_12[2] , \nOut12_12[1] , 
        \nOut12_12[0] }), .EastIn({\nOut13_11[7] , \nOut13_11[6] , 
        \nOut13_11[5] , \nOut13_11[4] , \nOut13_11[3] , \nOut13_11[2] , 
        \nOut13_11[1] , \nOut13_11[0] }), .WestIn({\nOut11_11[7] , 
        \nOut11_11[6] , \nOut11_11[5] , \nOut11_11[4] , \nOut11_11[3] , 
        \nOut11_11[2] , \nOut11_11[1] , \nOut11_11[0] }), .Out({\nOut12_11[7] , 
        \nOut12_11[6] , \nOut12_11[5] , \nOut12_11[4] , \nOut12_11[3] , 
        \nOut12_11[2] , \nOut12_11[1] , \nOut12_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_414 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut415[7] , \nScanOut415[6] , 
        \nScanOut415[5] , \nScanOut415[4] , \nScanOut415[3] , \nScanOut415[2] , 
        \nScanOut415[1] , \nScanOut415[0] }), .ScanOut({\nScanOut414[7] , 
        \nScanOut414[6] , \nScanOut414[5] , \nScanOut414[4] , \nScanOut414[3] , 
        \nScanOut414[2] , \nScanOut414[1] , \nScanOut414[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_29[7] , \nOut12_29[6] , \nOut12_29[5] , \nOut12_29[4] , 
        \nOut12_29[3] , \nOut12_29[2] , \nOut12_29[1] , \nOut12_29[0] }), 
        .SouthIn({\nOut12_31[7] , \nOut12_31[6] , \nOut12_31[5] , 
        \nOut12_31[4] , \nOut12_31[3] , \nOut12_31[2] , \nOut12_31[1] , 
        \nOut12_31[0] }), .EastIn({\nOut13_30[7] , \nOut13_30[6] , 
        \nOut13_30[5] , \nOut13_30[4] , \nOut13_30[3] , \nOut13_30[2] , 
        \nOut13_30[1] , \nOut13_30[0] }), .WestIn({\nOut11_30[7] , 
        \nOut11_30[6] , \nOut11_30[5] , \nOut11_30[4] , \nOut11_30[3] , 
        \nOut11_30[2] , \nOut11_30[1] , \nOut11_30[0] }), .Out({\nOut12_30[7] , 
        \nOut12_30[6] , \nOut12_30[5] , \nOut12_30[4] , \nOut12_30[3] , 
        \nOut12_30[2] , \nOut12_30[1] , \nOut12_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_507 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut508[7] , \nScanOut508[6] , 
        \nScanOut508[5] , \nScanOut508[4] , \nScanOut508[3] , \nScanOut508[2] , 
        \nScanOut508[1] , \nScanOut508[0] }), .ScanOut({\nScanOut507[7] , 
        \nScanOut507[6] , \nScanOut507[5] , \nScanOut507[4] , \nScanOut507[3] , 
        \nScanOut507[2] , \nScanOut507[1] , \nScanOut507[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_26[7] , \nOut15_26[6] , \nOut15_26[5] , \nOut15_26[4] , 
        \nOut15_26[3] , \nOut15_26[2] , \nOut15_26[1] , \nOut15_26[0] }), 
        .SouthIn({\nOut15_28[7] , \nOut15_28[6] , \nOut15_28[5] , 
        \nOut15_28[4] , \nOut15_28[3] , \nOut15_28[2] , \nOut15_28[1] , 
        \nOut15_28[0] }), .EastIn({\nOut16_27[7] , \nOut16_27[6] , 
        \nOut16_27[5] , \nOut16_27[4] , \nOut16_27[3] , \nOut16_27[2] , 
        \nOut16_27[1] , \nOut16_27[0] }), .WestIn({\nOut14_27[7] , 
        \nOut14_27[6] , \nOut14_27[5] , \nOut14_27[4] , \nOut14_27[3] , 
        \nOut14_27[2] , \nOut14_27[1] , \nOut14_27[0] }), .Out({\nOut15_27[7] , 
        \nOut15_27[6] , \nOut15_27[5] , \nOut15_27[4] , \nOut15_27[3] , 
        \nOut15_27[2] , \nOut15_27[1] , \nOut15_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_584 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut585[7] , \nScanOut585[6] , 
        \nScanOut585[5] , \nScanOut585[4] , \nScanOut585[3] , \nScanOut585[2] , 
        \nScanOut585[1] , \nScanOut585[0] }), .ScanOut({\nScanOut584[7] , 
        \nScanOut584[6] , \nScanOut584[5] , \nScanOut584[4] , \nScanOut584[3] , 
        \nScanOut584[2] , \nScanOut584[1] , \nScanOut584[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_7[7] , \nOut18_7[6] , \nOut18_7[5] , \nOut18_7[4] , 
        \nOut18_7[3] , \nOut18_7[2] , \nOut18_7[1] , \nOut18_7[0] }), 
        .SouthIn({\nOut18_9[7] , \nOut18_9[6] , \nOut18_9[5] , \nOut18_9[4] , 
        \nOut18_9[3] , \nOut18_9[2] , \nOut18_9[1] , \nOut18_9[0] }), .EastIn(
        {\nOut19_8[7] , \nOut19_8[6] , \nOut19_8[5] , \nOut19_8[4] , 
        \nOut19_8[3] , \nOut19_8[2] , \nOut19_8[1] , \nOut19_8[0] }), .WestIn(
        {\nOut17_8[7] , \nOut17_8[6] , \nOut17_8[5] , \nOut17_8[4] , 
        \nOut17_8[3] , \nOut17_8[2] , \nOut17_8[1] , \nOut17_8[0] }), .Out({
        \nOut18_8[7] , \nOut18_8[6] , \nOut18_8[5] , \nOut18_8[4] , 
        \nOut18_8[3] , \nOut18_8[2] , \nOut18_8[1] , \nOut18_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_724 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut725[7] , \nScanOut725[6] , 
        \nScanOut725[5] , \nScanOut725[4] , \nScanOut725[3] , \nScanOut725[2] , 
        \nScanOut725[1] , \nScanOut725[0] }), .ScanOut({\nScanOut724[7] , 
        \nScanOut724[6] , \nScanOut724[5] , \nScanOut724[4] , \nScanOut724[3] , 
        \nScanOut724[2] , \nScanOut724[1] , \nScanOut724[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_19[7] , \nOut22_19[6] , \nOut22_19[5] , \nOut22_19[4] , 
        \nOut22_19[3] , \nOut22_19[2] , \nOut22_19[1] , \nOut22_19[0] }), 
        .SouthIn({\nOut22_21[7] , \nOut22_21[6] , \nOut22_21[5] , 
        \nOut22_21[4] , \nOut22_21[3] , \nOut22_21[2] , \nOut22_21[1] , 
        \nOut22_21[0] }), .EastIn({\nOut23_20[7] , \nOut23_20[6] , 
        \nOut23_20[5] , \nOut23_20[4] , \nOut23_20[3] , \nOut23_20[2] , 
        \nOut23_20[1] , \nOut23_20[0] }), .WestIn({\nOut21_20[7] , 
        \nOut21_20[6] , \nOut21_20[5] , \nOut21_20[4] , \nOut21_20[3] , 
        \nOut21_20[2] , \nOut21_20[1] , \nOut21_20[0] }), .Out({\nOut22_20[7] , 
        \nOut22_20[6] , \nOut22_20[5] , \nOut22_20[4] , \nOut22_20[3] , 
        \nOut22_20[2] , \nOut22_20[1] , \nOut22_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_866 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut867[7] , \nScanOut867[6] , 
        \nScanOut867[5] , \nScanOut867[4] , \nScanOut867[3] , \nScanOut867[2] , 
        \nScanOut867[1] , \nScanOut867[0] }), .ScanOut({\nScanOut866[7] , 
        \nScanOut866[6] , \nScanOut866[5] , \nScanOut866[4] , \nScanOut866[3] , 
        \nScanOut866[2] , \nScanOut866[1] , \nScanOut866[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_1[7] , \nOut27_1[6] , \nOut27_1[5] , \nOut27_1[4] , 
        \nOut27_1[3] , \nOut27_1[2] , \nOut27_1[1] , \nOut27_1[0] }), 
        .SouthIn({\nOut27_3[7] , \nOut27_3[6] , \nOut27_3[5] , \nOut27_3[4] , 
        \nOut27_3[3] , \nOut27_3[2] , \nOut27_3[1] , \nOut27_3[0] }), .EastIn(
        {\nOut28_2[7] , \nOut28_2[6] , \nOut28_2[5] , \nOut28_2[4] , 
        \nOut28_2[3] , \nOut28_2[2] , \nOut28_2[1] , \nOut28_2[0] }), .WestIn(
        {\nOut26_2[7] , \nOut26_2[6] , \nOut26_2[5] , \nOut26_2[4] , 
        \nOut26_2[3] , \nOut26_2[2] , \nOut26_2[1] , \nOut26_2[0] }), .Out({
        \nOut27_2[7] , \nOut27_2[6] , \nOut27_2[5] , \nOut27_2[4] , 
        \nOut27_2[3] , \nOut27_2[2] , \nOut27_2[1] , \nOut27_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1022 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1023[7] , \nScanOut1023[6] , 
        \nScanOut1023[5] , \nScanOut1023[4] , \nScanOut1023[3] , 
        \nScanOut1023[2] , \nScanOut1023[1] , \nScanOut1023[0] }), .ScanOut({
        \nScanOut1022[7] , \nScanOut1022[6] , \nScanOut1022[5] , 
        \nScanOut1022[4] , \nScanOut1022[3] , \nScanOut1022[2] , 
        \nScanOut1022[1] , \nScanOut1022[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_30[7] , \nOut31_30[6] , \nOut31_30[5] , 
        \nOut31_30[4] , \nOut31_30[3] , \nOut31_30[2] , \nOut31_30[1] , 
        \nOut31_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_112 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut113[7] , \nScanOut113[6] , 
        \nScanOut113[5] , \nScanOut113[4] , \nScanOut113[3] , \nScanOut113[2] , 
        \nScanOut113[1] , \nScanOut113[0] }), .ScanOut({\nScanOut112[7] , 
        \nScanOut112[6] , \nScanOut112[5] , \nScanOut112[4] , \nScanOut112[3] , 
        \nScanOut112[2] , \nScanOut112[1] , \nScanOut112[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_15[7] , \nOut3_15[6] , \nOut3_15[5] , \nOut3_15[4] , 
        \nOut3_15[3] , \nOut3_15[2] , \nOut3_15[1] , \nOut3_15[0] }), 
        .SouthIn({\nOut3_17[7] , \nOut3_17[6] , \nOut3_17[5] , \nOut3_17[4] , 
        \nOut3_17[3] , \nOut3_17[2] , \nOut3_17[1] , \nOut3_17[0] }), .EastIn(
        {\nOut4_16[7] , \nOut4_16[6] , \nOut4_16[5] , \nOut4_16[4] , 
        \nOut4_16[3] , \nOut4_16[2] , \nOut4_16[1] , \nOut4_16[0] }), .WestIn(
        {\nOut2_16[7] , \nOut2_16[6] , \nOut2_16[5] , \nOut2_16[4] , 
        \nOut2_16[3] , \nOut2_16[2] , \nOut2_16[1] , \nOut2_16[0] }), .Out({
        \nOut3_16[7] , \nOut3_16[6] , \nOut3_16[5] , \nOut3_16[4] , 
        \nOut3_16[3] , \nOut3_16[2] , \nOut3_16[1] , \nOut3_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_199 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut200[7] , \nScanOut200[6] , 
        \nScanOut200[5] , \nScanOut200[4] , \nScanOut200[3] , \nScanOut200[2] , 
        \nScanOut200[1] , \nScanOut200[0] }), .ScanOut({\nScanOut199[7] , 
        \nScanOut199[6] , \nScanOut199[5] , \nScanOut199[4] , \nScanOut199[3] , 
        \nScanOut199[2] , \nScanOut199[1] , \nScanOut199[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_6[7] , \nOut6_6[6] , \nOut6_6[5] , \nOut6_6[4] , \nOut6_6[3] , 
        \nOut6_6[2] , \nOut6_6[1] , \nOut6_6[0] }), .SouthIn({\nOut6_8[7] , 
        \nOut6_8[6] , \nOut6_8[5] , \nOut6_8[4] , \nOut6_8[3] , \nOut6_8[2] , 
        \nOut6_8[1] , \nOut6_8[0] }), .EastIn({\nOut7_7[7] , \nOut7_7[6] , 
        \nOut7_7[5] , \nOut7_7[4] , \nOut7_7[3] , \nOut7_7[2] , \nOut7_7[1] , 
        \nOut7_7[0] }), .WestIn({\nOut5_7[7] , \nOut5_7[6] , \nOut5_7[5] , 
        \nOut5_7[4] , \nOut5_7[3] , \nOut5_7[2] , \nOut5_7[1] , \nOut5_7[0] }), 
        .Out({\nOut6_7[7] , \nOut6_7[6] , \nOut6_7[5] , \nOut6_7[4] , 
        \nOut6_7[3] , \nOut6_7[2] , \nOut6_7[1] , \nOut6_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_222 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut223[7] , \nScanOut223[6] , 
        \nScanOut223[5] , \nScanOut223[4] , \nScanOut223[3] , \nScanOut223[2] , 
        \nScanOut223[1] , \nScanOut223[0] }), .ScanOut({\nScanOut222[7] , 
        \nScanOut222[6] , \nScanOut222[5] , \nScanOut222[4] , \nScanOut222[3] , 
        \nScanOut222[2] , \nScanOut222[1] , \nScanOut222[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_29[7] , \nOut6_29[6] , \nOut6_29[5] , \nOut6_29[4] , 
        \nOut6_29[3] , \nOut6_29[2] , \nOut6_29[1] , \nOut6_29[0] }), 
        .SouthIn({\nOut6_31[7] , \nOut6_31[6] , \nOut6_31[5] , \nOut6_31[4] , 
        \nOut6_31[3] , \nOut6_31[2] , \nOut6_31[1] , \nOut6_31[0] }), .EastIn(
        {\nOut7_30[7] , \nOut7_30[6] , \nOut7_30[5] , \nOut7_30[4] , 
        \nOut7_30[3] , \nOut7_30[2] , \nOut7_30[1] , \nOut7_30[0] }), .WestIn(
        {\nOut5_30[7] , \nOut5_30[6] , \nOut5_30[5] , \nOut5_30[4] , 
        \nOut5_30[3] , \nOut5_30[2] , \nOut5_30[1] , \nOut5_30[0] }), .Out({
        \nOut6_30[7] , \nOut6_30[6] , \nOut6_30[5] , \nOut6_30[4] , 
        \nOut6_30[3] , \nOut6_30[2] , \nOut6_30[1] , \nOut6_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_693 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut694[7] , \nScanOut694[6] , 
        \nScanOut694[5] , \nScanOut694[4] , \nScanOut694[3] , \nScanOut694[2] , 
        \nScanOut694[1] , \nScanOut694[0] }), .ScanOut({\nScanOut693[7] , 
        \nScanOut693[6] , \nScanOut693[5] , \nScanOut693[4] , \nScanOut693[3] , 
        \nScanOut693[2] , \nScanOut693[1] , \nScanOut693[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_20[7] , \nOut21_20[6] , \nOut21_20[5] , \nOut21_20[4] , 
        \nOut21_20[3] , \nOut21_20[2] , \nOut21_20[1] , \nOut21_20[0] }), 
        .SouthIn({\nOut21_22[7] , \nOut21_22[6] , \nOut21_22[5] , 
        \nOut21_22[4] , \nOut21_22[3] , \nOut21_22[2] , \nOut21_22[1] , 
        \nOut21_22[0] }), .EastIn({\nOut22_21[7] , \nOut22_21[6] , 
        \nOut22_21[5] , \nOut22_21[4] , \nOut22_21[3] , \nOut22_21[2] , 
        \nOut22_21[1] , \nOut22_21[0] }), .WestIn({\nOut20_21[7] , 
        \nOut20_21[6] , \nOut20_21[5] , \nOut20_21[4] , \nOut20_21[3] , 
        \nOut20_21[2] , \nOut20_21[1] , \nOut20_21[0] }), .Out({\nOut21_21[7] , 
        \nOut21_21[6] , \nOut21_21[5] , \nOut21_21[4] , \nOut21_21[3] , 
        \nOut21_21[2] , \nOut21_21[1] , \nOut21_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1005 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1006[7] , \nScanOut1006[6] , 
        \nScanOut1006[5] , \nScanOut1006[4] , \nScanOut1006[3] , 
        \nScanOut1006[2] , \nScanOut1006[1] , \nScanOut1006[0] }), .ScanOut({
        \nScanOut1005[7] , \nScanOut1005[6] , \nScanOut1005[5] , 
        \nScanOut1005[4] , \nScanOut1005[3] , \nScanOut1005[2] , 
        \nScanOut1005[1] , \nScanOut1005[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_13[7] , \nOut31_13[6] , \nOut31_13[5] , 
        \nOut31_13[4] , \nOut31_13[3] , \nOut31_13[2] , \nOut31_13[1] , 
        \nOut31_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_703 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut704[7] , \nScanOut704[6] , 
        \nScanOut704[5] , \nScanOut704[4] , \nScanOut704[3] , \nScanOut704[2] , 
        \nScanOut704[1] , \nScanOut704[0] }), .ScanOut({\nScanOut703[7] , 
        \nScanOut703[6] , \nScanOut703[5] , \nScanOut703[4] , \nScanOut703[3] , 
        \nScanOut703[2] , \nScanOut703[1] , \nScanOut703[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut21_31[7] , \nOut21_31[6] , 
        \nOut21_31[5] , \nOut21_31[4] , \nOut21_31[3] , \nOut21_31[2] , 
        \nOut21_31[1] , \nOut21_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_433 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut434[7] , \nScanOut434[6] , 
        \nScanOut434[5] , \nScanOut434[4] , \nScanOut434[3] , \nScanOut434[2] , 
        \nScanOut434[1] , \nScanOut434[0] }), .ScanOut({\nScanOut433[7] , 
        \nScanOut433[6] , \nScanOut433[5] , \nScanOut433[4] , \nScanOut433[3] , 
        \nScanOut433[2] , \nScanOut433[1] , \nScanOut433[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_16[7] , \nOut13_16[6] , \nOut13_16[5] , \nOut13_16[4] , 
        \nOut13_16[3] , \nOut13_16[2] , \nOut13_16[1] , \nOut13_16[0] }), 
        .SouthIn({\nOut13_18[7] , \nOut13_18[6] , \nOut13_18[5] , 
        \nOut13_18[4] , \nOut13_18[3] , \nOut13_18[2] , \nOut13_18[1] , 
        \nOut13_18[0] }), .EastIn({\nOut14_17[7] , \nOut14_17[6] , 
        \nOut14_17[5] , \nOut14_17[4] , \nOut14_17[3] , \nOut14_17[2] , 
        \nOut14_17[1] , \nOut14_17[0] }), .WestIn({\nOut12_17[7] , 
        \nOut12_17[6] , \nOut12_17[5] , \nOut12_17[4] , \nOut12_17[3] , 
        \nOut12_17[2] , \nOut12_17[1] , \nOut12_17[0] }), .Out({\nOut13_17[7] , 
        \nOut13_17[6] , \nOut13_17[5] , \nOut13_17[4] , \nOut13_17[3] , 
        \nOut13_17[2] , \nOut13_17[1] , \nOut13_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_841 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut842[7] , \nScanOut842[6] , 
        \nScanOut842[5] , \nScanOut842[4] , \nScanOut842[3] , \nScanOut842[2] , 
        \nScanOut842[1] , \nScanOut842[0] }), .ScanOut({\nScanOut841[7] , 
        \nScanOut841[6] , \nScanOut841[5] , \nScanOut841[4] , \nScanOut841[3] , 
        \nScanOut841[2] , \nScanOut841[1] , \nScanOut841[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_8[7] , \nOut26_8[6] , \nOut26_8[5] , \nOut26_8[4] , 
        \nOut26_8[3] , \nOut26_8[2] , \nOut26_8[1] , \nOut26_8[0] }), 
        .SouthIn({\nOut26_10[7] , \nOut26_10[6] , \nOut26_10[5] , 
        \nOut26_10[4] , \nOut26_10[3] , \nOut26_10[2] , \nOut26_10[1] , 
        \nOut26_10[0] }), .EastIn({\nOut27_9[7] , \nOut27_9[6] , \nOut27_9[5] , 
        \nOut27_9[4] , \nOut27_9[3] , \nOut27_9[2] , \nOut27_9[1] , 
        \nOut27_9[0] }), .WestIn({\nOut25_9[7] , \nOut25_9[6] , \nOut25_9[5] , 
        \nOut25_9[4] , \nOut25_9[3] , \nOut25_9[2] , \nOut25_9[1] , 
        \nOut25_9[0] }), .Out({\nOut26_9[7] , \nOut26_9[6] , \nOut26_9[5] , 
        \nOut26_9[4] , \nOut26_9[3] , \nOut26_9[2] , \nOut26_9[1] , 
        \nOut26_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_339 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut340[7] , \nScanOut340[6] , 
        \nScanOut340[5] , \nScanOut340[4] , \nScanOut340[3] , \nScanOut340[2] , 
        \nScanOut340[1] , \nScanOut340[0] }), .ScanOut({\nScanOut339[7] , 
        \nScanOut339[6] , \nScanOut339[5] , \nScanOut339[4] , \nScanOut339[3] , 
        \nScanOut339[2] , \nScanOut339[1] , \nScanOut339[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_18[7] , \nOut10_18[6] , \nOut10_18[5] , \nOut10_18[4] , 
        \nOut10_18[3] , \nOut10_18[2] , \nOut10_18[1] , \nOut10_18[0] }), 
        .SouthIn({\nOut10_20[7] , \nOut10_20[6] , \nOut10_20[5] , 
        \nOut10_20[4] , \nOut10_20[3] , \nOut10_20[2] , \nOut10_20[1] , 
        \nOut10_20[0] }), .EastIn({\nOut11_19[7] , \nOut11_19[6] , 
        \nOut11_19[5] , \nOut11_19[4] , \nOut11_19[3] , \nOut11_19[2] , 
        \nOut11_19[1] , \nOut11_19[0] }), .WestIn({\nOut9_19[7] , 
        \nOut9_19[6] , \nOut9_19[5] , \nOut9_19[4] , \nOut9_19[3] , 
        \nOut9_19[2] , \nOut9_19[1] , \nOut9_19[0] }), .Out({\nOut10_19[7] , 
        \nOut10_19[6] , \nOut10_19[5] , \nOut10_19[4] , \nOut10_19[3] , 
        \nOut10_19[2] , \nOut10_19[1] , \nOut10_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_528 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut529[7] , \nScanOut529[6] , 
        \nScanOut529[5] , \nScanOut529[4] , \nScanOut529[3] , \nScanOut529[2] , 
        \nScanOut529[1] , \nScanOut529[0] }), .ScanOut({\nScanOut528[7] , 
        \nScanOut528[6] , \nScanOut528[5] , \nScanOut528[4] , \nScanOut528[3] , 
        \nScanOut528[2] , \nScanOut528[1] , \nScanOut528[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_15[7] , \nOut16_15[6] , \nOut16_15[5] , \nOut16_15[4] , 
        \nOut16_15[3] , \nOut16_15[2] , \nOut16_15[1] , \nOut16_15[0] }), 
        .SouthIn({\nOut16_17[7] , \nOut16_17[6] , \nOut16_17[5] , 
        \nOut16_17[4] , \nOut16_17[3] , \nOut16_17[2] , \nOut16_17[1] , 
        \nOut16_17[0] }), .EastIn({\nOut17_16[7] , \nOut17_16[6] , 
        \nOut17_16[5] , \nOut17_16[4] , \nOut17_16[3] , \nOut17_16[2] , 
        \nOut17_16[1] , \nOut17_16[0] }), .WestIn({\nOut15_16[7] , 
        \nOut15_16[6] , \nOut15_16[5] , \nOut15_16[4] , \nOut15_16[3] , 
        \nOut15_16[2] , \nOut15_16[1] , \nOut15_16[0] }), .Out({\nOut16_16[7] , 
        \nOut16_16[6] , \nOut16_16[5] , \nOut16_16[4] , \nOut16_16[3] , 
        \nOut16_16[2] , \nOut16_16[1] , \nOut16_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_618 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut619[7] , \nScanOut619[6] , 
        \nScanOut619[5] , \nScanOut619[4] , \nScanOut619[3] , \nScanOut619[2] , 
        \nScanOut619[1] , \nScanOut619[0] }), .ScanOut({\nScanOut618[7] , 
        \nScanOut618[6] , \nScanOut618[5] , \nScanOut618[4] , \nScanOut618[3] , 
        \nScanOut618[2] , \nScanOut618[1] , \nScanOut618[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_9[7] , \nOut19_9[6] , \nOut19_9[5] , \nOut19_9[4] , 
        \nOut19_9[3] , \nOut19_9[2] , \nOut19_9[1] , \nOut19_9[0] }), 
        .SouthIn({\nOut19_11[7] , \nOut19_11[6] , \nOut19_11[5] , 
        \nOut19_11[4] , \nOut19_11[3] , \nOut19_11[2] , \nOut19_11[1] , 
        \nOut19_11[0] }), .EastIn({\nOut20_10[7] , \nOut20_10[6] , 
        \nOut20_10[5] , \nOut20_10[4] , \nOut20_10[3] , \nOut20_10[2] , 
        \nOut20_10[1] , \nOut20_10[0] }), .WestIn({\nOut18_10[7] , 
        \nOut18_10[6] , \nOut18_10[5] , \nOut18_10[4] , \nOut18_10[3] , 
        \nOut18_10[2] , \nOut18_10[1] , \nOut18_10[0] }), .Out({\nOut19_10[7] , 
        \nOut19_10[6] , \nOut19_10[5] , \nOut19_10[4] , \nOut19_10[3] , 
        \nOut19_10[2] , \nOut19_10[1] , \nOut19_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_788 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut789[7] , \nScanOut789[6] , 
        \nScanOut789[5] , \nScanOut789[4] , \nScanOut789[3] , \nScanOut789[2] , 
        \nScanOut789[1] , \nScanOut789[0] }), .ScanOut({\nScanOut788[7] , 
        \nScanOut788[6] , \nScanOut788[5] , \nScanOut788[4] , \nScanOut788[3] , 
        \nScanOut788[2] , \nScanOut788[1] , \nScanOut788[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_19[7] , \nOut24_19[6] , \nOut24_19[5] , \nOut24_19[4] , 
        \nOut24_19[3] , \nOut24_19[2] , \nOut24_19[1] , \nOut24_19[0] }), 
        .SouthIn({\nOut24_21[7] , \nOut24_21[6] , \nOut24_21[5] , 
        \nOut24_21[4] , \nOut24_21[3] , \nOut24_21[2] , \nOut24_21[1] , 
        \nOut24_21[0] }), .EastIn({\nOut25_20[7] , \nOut25_20[6] , 
        \nOut25_20[5] , \nOut25_20[4] , \nOut25_20[3] , \nOut25_20[2] , 
        \nOut25_20[1] , \nOut25_20[0] }), .WestIn({\nOut23_20[7] , 
        \nOut23_20[6] , \nOut23_20[5] , \nOut23_20[4] , \nOut23_20[3] , 
        \nOut23_20[2] , \nOut23_20[1] , \nOut23_20[0] }), .Out({\nOut24_20[7] , 
        \nOut24_20[6] , \nOut24_20[5] , \nOut24_20[4] , \nOut24_20[3] , 
        \nOut24_20[2] , \nOut24_20[1] , \nOut24_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_676 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut677[7] , \nScanOut677[6] , 
        \nScanOut677[5] , \nScanOut677[4] , \nScanOut677[3] , \nScanOut677[2] , 
        \nScanOut677[1] , \nScanOut677[0] }), .ScanOut({\nScanOut676[7] , 
        \nScanOut676[6] , \nScanOut676[5] , \nScanOut676[4] , \nScanOut676[3] , 
        \nScanOut676[2] , \nScanOut676[1] , \nScanOut676[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_3[7] , \nOut21_3[6] , \nOut21_3[5] , \nOut21_3[4] , 
        \nOut21_3[3] , \nOut21_3[2] , \nOut21_3[1] , \nOut21_3[0] }), 
        .SouthIn({\nOut21_5[7] , \nOut21_5[6] , \nOut21_5[5] , \nOut21_5[4] , 
        \nOut21_5[3] , \nOut21_5[2] , \nOut21_5[1] , \nOut21_5[0] }), .EastIn(
        {\nOut22_4[7] , \nOut22_4[6] , \nOut22_4[5] , \nOut22_4[4] , 
        \nOut22_4[3] , \nOut22_4[2] , \nOut22_4[1] , \nOut22_4[0] }), .WestIn(
        {\nOut20_4[7] , \nOut20_4[6] , \nOut20_4[5] , \nOut20_4[4] , 
        \nOut20_4[3] , \nOut20_4[2] , \nOut20_4[1] , \nOut20_4[0] }), .Out({
        \nOut21_4[7] , \nOut21_4[6] , \nOut21_4[5] , \nOut21_4[4] , 
        \nOut21_4[3] , \nOut21_4[2] , \nOut21_4[1] , \nOut21_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_357 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut358[7] , \nScanOut358[6] , 
        \nScanOut358[5] , \nScanOut358[4] , \nScanOut358[3] , \nScanOut358[2] , 
        \nScanOut358[1] , \nScanOut358[0] }), .ScanOut({\nScanOut357[7] , 
        \nScanOut357[6] , \nScanOut357[5] , \nScanOut357[4] , \nScanOut357[3] , 
        \nScanOut357[2] , \nScanOut357[1] , \nScanOut357[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }), 
        .SouthIn({\nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }), .EastIn(
        {\nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }), .WestIn(
        {\nOut10_5[7] , \nOut10_5[6] , \nOut10_5[5] , \nOut10_5[4] , 
        \nOut10_5[3] , \nOut10_5[2] , \nOut10_5[1] , \nOut10_5[0] }), .Out({
        \nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_370 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut371[7] , \nScanOut371[6] , 
        \nScanOut371[5] , \nScanOut371[4] , \nScanOut371[3] , \nScanOut371[2] , 
        \nScanOut371[1] , \nScanOut371[0] }), .ScanOut({\nScanOut370[7] , 
        \nScanOut370[6] , \nScanOut370[5] , \nScanOut370[4] , \nScanOut370[3] , 
        \nScanOut370[2] , \nScanOut370[1] , \nScanOut370[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_17[7] , \nOut11_17[6] , \nOut11_17[5] , \nOut11_17[4] , 
        \nOut11_17[3] , \nOut11_17[2] , \nOut11_17[1] , \nOut11_17[0] }), 
        .SouthIn({\nOut11_19[7] , \nOut11_19[6] , \nOut11_19[5] , 
        \nOut11_19[4] , \nOut11_19[3] , \nOut11_19[2] , \nOut11_19[1] , 
        \nOut11_19[0] }), .EastIn({\nOut12_18[7] , \nOut12_18[6] , 
        \nOut12_18[5] , \nOut12_18[4] , \nOut12_18[3] , \nOut12_18[2] , 
        \nOut12_18[1] , \nOut12_18[0] }), .WestIn({\nOut10_18[7] , 
        \nOut10_18[6] , \nOut10_18[5] , \nOut10_18[4] , \nOut10_18[3] , 
        \nOut10_18[2] , \nOut10_18[1] , \nOut10_18[0] }), .Out({\nOut11_18[7] , 
        \nOut11_18[6] , \nOut11_18[5] , \nOut11_18[4] , \nOut11_18[3] , 
        \nOut11_18[2] , \nOut11_18[1] , \nOut11_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_546 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut547[7] , \nScanOut547[6] , 
        \nScanOut547[5] , \nScanOut547[4] , \nScanOut547[3] , \nScanOut547[2] , 
        \nScanOut547[1] , \nScanOut547[0] }), .ScanOut({\nScanOut546[7] , 
        \nScanOut546[6] , \nScanOut546[5] , \nScanOut546[4] , \nScanOut546[3] , 
        \nScanOut546[2] , \nScanOut546[1] , \nScanOut546[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_1[7] , \nOut17_1[6] , \nOut17_1[5] , \nOut17_1[4] , 
        \nOut17_1[3] , \nOut17_1[2] , \nOut17_1[1] , \nOut17_1[0] }), 
        .SouthIn({\nOut17_3[7] , \nOut17_3[6] , \nOut17_3[5] , \nOut17_3[4] , 
        \nOut17_3[3] , \nOut17_3[2] , \nOut17_3[1] , \nOut17_3[0] }), .EastIn(
        {\nOut18_2[7] , \nOut18_2[6] , \nOut18_2[5] , \nOut18_2[4] , 
        \nOut18_2[3] , \nOut18_2[2] , \nOut18_2[1] , \nOut18_2[0] }), .WestIn(
        {\nOut16_2[7] , \nOut16_2[6] , \nOut16_2[5] , \nOut16_2[4] , 
        \nOut16_2[3] , \nOut16_2[2] , \nOut16_2[1] , \nOut16_2[0] }), .Out({
        \nOut17_2[7] , \nOut17_2[6] , \nOut17_2[5] , \nOut17_2[4] , 
        \nOut17_2[3] , \nOut17_2[2] , \nOut17_2[1] , \nOut17_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_561 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut562[7] , \nScanOut562[6] , 
        \nScanOut562[5] , \nScanOut562[4] , \nScanOut562[3] , \nScanOut562[2] , 
        \nScanOut562[1] , \nScanOut562[0] }), .ScanOut({\nScanOut561[7] , 
        \nScanOut561[6] , \nScanOut561[5] , \nScanOut561[4] , \nScanOut561[3] , 
        \nScanOut561[2] , \nScanOut561[1] , \nScanOut561[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_16[7] , \nOut17_16[6] , \nOut17_16[5] , \nOut17_16[4] , 
        \nOut17_16[3] , \nOut17_16[2] , \nOut17_16[1] , \nOut17_16[0] }), 
        .SouthIn({\nOut17_18[7] , \nOut17_18[6] , \nOut17_18[5] , 
        \nOut17_18[4] , \nOut17_18[3] , \nOut17_18[2] , \nOut17_18[1] , 
        \nOut17_18[0] }), .EastIn({\nOut18_17[7] , \nOut18_17[6] , 
        \nOut18_17[5] , \nOut18_17[4] , \nOut18_17[3] , \nOut18_17[2] , 
        \nOut18_17[1] , \nOut18_17[0] }), .WestIn({\nOut16_17[7] , 
        \nOut16_17[6] , \nOut16_17[5] , \nOut16_17[4] , \nOut16_17[3] , 
        \nOut16_17[2] , \nOut16_17[1] , \nOut16_17[0] }), .Out({\nOut17_17[7] , 
        \nOut17_17[6] , \nOut17_17[5] , \nOut17_17[4] , \nOut17_17[3] , 
        \nOut17_17[2] , \nOut17_17[1] , \nOut17_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_934 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut935[7] , \nScanOut935[6] , 
        \nScanOut935[5] , \nScanOut935[4] , \nScanOut935[3] , \nScanOut935[2] , 
        \nScanOut935[1] , \nScanOut935[0] }), .ScanOut({\nScanOut934[7] , 
        \nScanOut934[6] , \nScanOut934[5] , \nScanOut934[4] , \nScanOut934[3] , 
        \nScanOut934[2] , \nScanOut934[1] , \nScanOut934[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_5[7] , \nOut29_5[6] , \nOut29_5[5] , \nOut29_5[4] , 
        \nOut29_5[3] , \nOut29_5[2] , \nOut29_5[1] , \nOut29_5[0] }), 
        .SouthIn({\nOut29_7[7] , \nOut29_7[6] , \nOut29_7[5] , \nOut29_7[4] , 
        \nOut29_7[3] , \nOut29_7[2] , \nOut29_7[1] , \nOut29_7[0] }), .EastIn(
        {\nOut30_6[7] , \nOut30_6[6] , \nOut30_6[5] , \nOut30_6[4] , 
        \nOut30_6[3] , \nOut30_6[2] , \nOut30_6[1] , \nOut30_6[0] }), .WestIn(
        {\nOut28_6[7] , \nOut28_6[6] , \nOut28_6[5] , \nOut28_6[4] , 
        \nOut28_6[3] , \nOut28_6[2] , \nOut28_6[1] , \nOut28_6[0] }), .Out({
        \nOut29_6[7] , \nOut29_6[6] , \nOut29_6[5] , \nOut29_6[4] , 
        \nOut29_6[3] , \nOut29_6[2] , \nOut29_6[1] , \nOut29_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_883 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut884[7] , \nScanOut884[6] , 
        \nScanOut884[5] , \nScanOut884[4] , \nScanOut884[3] , \nScanOut884[2] , 
        \nScanOut884[1] , \nScanOut884[0] }), .ScanOut({\nScanOut883[7] , 
        \nScanOut883[6] , \nScanOut883[5] , \nScanOut883[4] , \nScanOut883[3] , 
        \nScanOut883[2] , \nScanOut883[1] , \nScanOut883[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_18[7] , \nOut27_18[6] , \nOut27_18[5] , \nOut27_18[4] , 
        \nOut27_18[3] , \nOut27_18[2] , \nOut27_18[1] , \nOut27_18[0] }), 
        .SouthIn({\nOut27_20[7] , \nOut27_20[6] , \nOut27_20[5] , 
        \nOut27_20[4] , \nOut27_20[3] , \nOut27_20[2] , \nOut27_20[1] , 
        \nOut27_20[0] }), .EastIn({\nOut28_19[7] , \nOut28_19[6] , 
        \nOut28_19[5] , \nOut28_19[4] , \nOut28_19[3] , \nOut28_19[2] , 
        \nOut28_19[1] , \nOut28_19[0] }), .WestIn({\nOut26_19[7] , 
        \nOut26_19[6] , \nOut26_19[5] , \nOut26_19[4] , \nOut26_19[3] , 
        \nOut26_19[2] , \nOut26_19[1] , \nOut26_19[0] }), .Out({\nOut27_19[7] , 
        \nOut27_19[6] , \nOut27_19[5] , \nOut27_19[4] , \nOut27_19[3] , 
        \nOut27_19[2] , \nOut27_19[1] , \nOut27_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_913 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut914[7] , \nScanOut914[6] , 
        \nScanOut914[5] , \nScanOut914[4] , \nScanOut914[3] , \nScanOut914[2] , 
        \nScanOut914[1] , \nScanOut914[0] }), .ScanOut({\nScanOut913[7] , 
        \nScanOut913[6] , \nScanOut913[5] , \nScanOut913[4] , \nScanOut913[3] , 
        \nScanOut913[2] , \nScanOut913[1] , \nScanOut913[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_16[7] , \nOut28_16[6] , \nOut28_16[5] , \nOut28_16[4] , 
        \nOut28_16[3] , \nOut28_16[2] , \nOut28_16[1] , \nOut28_16[0] }), 
        .SouthIn({\nOut28_18[7] , \nOut28_18[6] , \nOut28_18[5] , 
        \nOut28_18[4] , \nOut28_18[3] , \nOut28_18[2] , \nOut28_18[1] , 
        \nOut28_18[0] }), .EastIn({\nOut29_17[7] , \nOut29_17[6] , 
        \nOut29_17[5] , \nOut29_17[4] , \nOut29_17[3] , \nOut29_17[2] , 
        \nOut29_17[1] , \nOut29_17[0] }), .WestIn({\nOut27_17[7] , 
        \nOut27_17[6] , \nOut27_17[5] , \nOut27_17[4] , \nOut27_17[3] , 
        \nOut27_17[2] , \nOut27_17[1] , \nOut27_17[0] }), .Out({\nOut28_17[7] , 
        \nOut28_17[6] , \nOut28_17[5] , \nOut28_17[4] , \nOut28_17[3] , 
        \nOut28_17[2] , \nOut28_17[1] , \nOut28_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_5 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut6[7] , \nScanOut6[6] , 
        \nScanOut6[5] , \nScanOut6[4] , \nScanOut6[3] , \nScanOut6[2] , 
        \nScanOut6[1] , \nScanOut6[0] }), .ScanOut({\nScanOut5[7] , 
        \nScanOut5[6] , \nScanOut5[5] , \nScanOut5[4] , \nScanOut5[3] , 
        \nScanOut5[2] , \nScanOut5[1] , \nScanOut5[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_5[7] , \nOut0_5[6] , 
        \nOut0_5[5] , \nOut0_5[4] , \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , 
        \nOut0_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_11 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut12[7] , \nScanOut12[6] , 
        \nScanOut12[5] , \nScanOut12[4] , \nScanOut12[3] , \nScanOut12[2] , 
        \nScanOut12[1] , \nScanOut12[0] }), .ScanOut({\nScanOut11[7] , 
        \nScanOut11[6] , \nScanOut11[5] , \nScanOut11[4] , \nScanOut11[3] , 
        \nScanOut11[2] , \nScanOut11[1] , \nScanOut11[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_11[7] , \nOut0_11[6] , 
        \nOut0_11[5] , \nOut0_11[4] , \nOut0_11[3] , \nOut0_11[2] , 
        \nOut0_11[1] , \nOut0_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_16 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut17[7] , \nScanOut17[6] , 
        \nScanOut17[5] , \nScanOut17[4] , \nScanOut17[3] , \nScanOut17[2] , 
        \nScanOut17[1] , \nScanOut17[0] }), .ScanOut({\nScanOut16[7] , 
        \nScanOut16[6] , \nScanOut16[5] , \nScanOut16[4] , \nScanOut16[3] , 
        \nScanOut16[2] , \nScanOut16[1] , \nScanOut16[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_16[7] , \nOut0_16[6] , 
        \nOut0_16[5] , \nOut0_16[4] , \nOut0_16[3] , \nOut0_16[2] , 
        \nOut0_16[1] , \nOut0_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_44 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut45[7] , \nScanOut45[6] , 
        \nScanOut45[5] , \nScanOut45[4] , \nScanOut45[3] , \nScanOut45[2] , 
        \nScanOut45[1] , \nScanOut45[0] }), .ScanOut({\nScanOut44[7] , 
        \nScanOut44[6] , \nScanOut44[5] , \nScanOut44[4] , \nScanOut44[3] , 
        \nScanOut44[2] , \nScanOut44[1] , \nScanOut44[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_11[7] , \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , 
        \nOut1_11[3] , \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), 
        .SouthIn({\nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), .EastIn(
        {\nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), .WestIn(
        {\nOut0_12[7] , \nOut0_12[6] , \nOut0_12[5] , \nOut0_12[4] , 
        \nOut0_12[3] , \nOut0_12[2] , \nOut0_12[1] , \nOut0_12[0] }), .Out({
        \nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_651 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut652[7] , \nScanOut652[6] , 
        \nScanOut652[5] , \nScanOut652[4] , \nScanOut652[3] , \nScanOut652[2] , 
        \nScanOut652[1] , \nScanOut652[0] }), .ScanOut({\nScanOut651[7] , 
        \nScanOut651[6] , \nScanOut651[5] , \nScanOut651[4] , \nScanOut651[3] , 
        \nScanOut651[2] , \nScanOut651[1] , \nScanOut651[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_10[7] , \nOut20_10[6] , \nOut20_10[5] , \nOut20_10[4] , 
        \nOut20_10[3] , \nOut20_10[2] , \nOut20_10[1] , \nOut20_10[0] }), 
        .SouthIn({\nOut20_12[7] , \nOut20_12[6] , \nOut20_12[5] , 
        \nOut20_12[4] , \nOut20_12[3] , \nOut20_12[2] , \nOut20_12[1] , 
        \nOut20_12[0] }), .EastIn({\nOut21_11[7] , \nOut21_11[6] , 
        \nOut21_11[5] , \nOut21_11[4] , \nOut21_11[3] , \nOut21_11[2] , 
        \nOut21_11[1] , \nOut21_11[0] }), .WestIn({\nOut19_11[7] , 
        \nOut19_11[6] , \nOut19_11[5] , \nOut19_11[4] , \nOut19_11[3] , 
        \nOut19_11[2] , \nOut19_11[1] , \nOut19_11[0] }), .Out({\nOut20_11[7] , 
        \nOut20_11[6] , \nOut20_11[5] , \nOut20_11[4] , \nOut20_11[3] , 
        \nOut20_11[2] , \nOut20_11[1] , \nOut20_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_78 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut79[7] , \nScanOut79[6] , 
        \nScanOut79[5] , \nScanOut79[4] , \nScanOut79[3] , \nScanOut79[2] , 
        \nScanOut79[1] , \nScanOut79[0] }), .ScanOut({\nScanOut78[7] , 
        \nScanOut78[6] , \nScanOut78[5] , \nScanOut78[4] , \nScanOut78[3] , 
        \nScanOut78[2] , \nScanOut78[1] , \nScanOut78[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), 
        .SouthIn({\nOut2_15[7] , \nOut2_15[6] , \nOut2_15[5] , \nOut2_15[4] , 
        \nOut2_15[3] , \nOut2_15[2] , \nOut2_15[1] , \nOut2_15[0] }), .EastIn(
        {\nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }), .WestIn(
        {\nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), .Out({
        \nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_140 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut141[7] , \nScanOut141[6] , 
        \nScanOut141[5] , \nScanOut141[4] , \nScanOut141[3] , \nScanOut141[2] , 
        \nScanOut141[1] , \nScanOut141[0] }), .ScanOut({\nScanOut140[7] , 
        \nScanOut140[6] , \nScanOut140[5] , \nScanOut140[4] , \nScanOut140[3] , 
        \nScanOut140[2] , \nScanOut140[1] , \nScanOut140[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_11[7] , \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , 
        \nOut4_11[3] , \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }), 
        .SouthIn({\nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }), .EastIn(
        {\nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }), .WestIn(
        {\nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }), .Out({
        \nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_808 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut809[7] , \nScanOut809[6] , 
        \nScanOut809[5] , \nScanOut809[4] , \nScanOut809[3] , \nScanOut809[2] , 
        \nScanOut809[1] , \nScanOut809[0] }), .ScanOut({\nScanOut808[7] , 
        \nScanOut808[6] , \nScanOut808[5] , \nScanOut808[4] , \nScanOut808[3] , 
        \nScanOut808[2] , \nScanOut808[1] , \nScanOut808[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_7[7] , \nOut25_7[6] , \nOut25_7[5] , \nOut25_7[4] , 
        \nOut25_7[3] , \nOut25_7[2] , \nOut25_7[1] , \nOut25_7[0] }), 
        .SouthIn({\nOut25_9[7] , \nOut25_9[6] , \nOut25_9[5] , \nOut25_9[4] , 
        \nOut25_9[3] , \nOut25_9[2] , \nOut25_9[1] , \nOut25_9[0] }), .EastIn(
        {\nOut26_8[7] , \nOut26_8[6] , \nOut26_8[5] , \nOut26_8[4] , 
        \nOut26_8[3] , \nOut26_8[2] , \nOut26_8[1] , \nOut26_8[0] }), .WestIn(
        {\nOut24_8[7] , \nOut24_8[6] , \nOut24_8[5] , \nOut24_8[4] , 
        \nOut24_8[3] , \nOut24_8[2] , \nOut24_8[1] , \nOut24_8[0] }), .Out({
        \nOut25_8[7] , \nOut25_8[6] , \nOut25_8[5] , \nOut25_8[4] , 
        \nOut25_8[3] , \nOut25_8[2] , \nOut25_8[1] , \nOut25_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_998 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut999[7] , \nScanOut999[6] , 
        \nScanOut999[5] , \nScanOut999[4] , \nScanOut999[3] , \nScanOut999[2] , 
        \nScanOut999[1] , \nScanOut999[0] }), .ScanOut({\nScanOut998[7] , 
        \nScanOut998[6] , \nScanOut998[5] , \nScanOut998[4] , \nScanOut998[3] , 
        \nScanOut998[2] , \nScanOut998[1] , \nScanOut998[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut31_6[7] , \nOut31_6[6] , 
        \nOut31_6[5] , \nOut31_6[4] , \nOut31_6[3] , \nOut31_6[2] , 
        \nOut31_6[1] , \nOut31_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_167 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut168[7] , \nScanOut168[6] , 
        \nScanOut168[5] , \nScanOut168[4] , \nScanOut168[3] , \nScanOut168[2] , 
        \nScanOut168[1] , \nScanOut168[0] }), .ScanOut({\nScanOut167[7] , 
        \nScanOut167[6] , \nScanOut167[5] , \nScanOut167[4] , \nScanOut167[3] , 
        \nScanOut167[2] , \nScanOut167[1] , \nScanOut167[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_6[7] , \nOut5_6[6] , \nOut5_6[5] , \nOut5_6[4] , \nOut5_6[3] , 
        \nOut5_6[2] , \nOut5_6[1] , \nOut5_6[0] }), .SouthIn({\nOut5_8[7] , 
        \nOut5_8[6] , \nOut5_8[5] , \nOut5_8[4] , \nOut5_8[3] , \nOut5_8[2] , 
        \nOut5_8[1] , \nOut5_8[0] }), .EastIn({\nOut6_7[7] , \nOut6_7[6] , 
        \nOut6_7[5] , \nOut6_7[4] , \nOut6_7[3] , \nOut6_7[2] , \nOut6_7[1] , 
        \nOut6_7[0] }), .WestIn({\nOut4_7[7] , \nOut4_7[6] , \nOut4_7[5] , 
        \nOut4_7[4] , \nOut4_7[3] , \nOut4_7[2] , \nOut4_7[1] , \nOut4_7[0] }), 
        .Out({\nOut5_7[7] , \nOut5_7[6] , \nOut5_7[5] , \nOut5_7[4] , 
        \nOut5_7[3] , \nOut5_7[2] , \nOut5_7[1] , \nOut5_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_257 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut258[7] , \nScanOut258[6] , 
        \nScanOut258[5] , \nScanOut258[4] , \nScanOut258[3] , \nScanOut258[2] , 
        \nScanOut258[1] , \nScanOut258[0] }), .ScanOut({\nScanOut257[7] , 
        \nScanOut257[6] , \nScanOut257[5] , \nScanOut257[4] , \nScanOut257[3] , 
        \nScanOut257[2] , \nScanOut257[1] , \nScanOut257[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_0[7] , \nOut8_0[6] , \nOut8_0[5] , \nOut8_0[4] , \nOut8_0[3] , 
        \nOut8_0[2] , \nOut8_0[1] , \nOut8_0[0] }), .SouthIn({\nOut8_2[7] , 
        \nOut8_2[6] , \nOut8_2[5] , \nOut8_2[4] , \nOut8_2[3] , \nOut8_2[2] , 
        \nOut8_2[1] , \nOut8_2[0] }), .EastIn({\nOut9_1[7] , \nOut9_1[6] , 
        \nOut9_1[5] , \nOut9_1[4] , \nOut9_1[3] , \nOut9_1[2] , \nOut9_1[1] , 
        \nOut9_1[0] }), .WestIn({\nOut7_1[7] , \nOut7_1[6] , \nOut7_1[5] , 
        \nOut7_1[4] , \nOut7_1[3] , \nOut7_1[2] , \nOut7_1[1] , \nOut7_1[0] }), 
        .Out({\nOut8_1[7] , \nOut8_1[6] , \nOut8_1[5] , \nOut8_1[4] , 
        \nOut8_1[3] , \nOut8_1[2] , \nOut8_1[1] , \nOut8_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_270 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut271[7] , \nScanOut271[6] , 
        \nScanOut271[5] , \nScanOut271[4] , \nScanOut271[3] , \nScanOut271[2] , 
        \nScanOut271[1] , \nScanOut271[0] }), .ScanOut({\nScanOut270[7] , 
        \nScanOut270[6] , \nScanOut270[5] , \nScanOut270[4] , \nScanOut270[3] , 
        \nScanOut270[2] , \nScanOut270[1] , \nScanOut270[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }), 
        .SouthIn({\nOut8_15[7] , \nOut8_15[6] , \nOut8_15[5] , \nOut8_15[4] , 
        \nOut8_15[3] , \nOut8_15[2] , \nOut8_15[1] , \nOut8_15[0] }), .EastIn(
        {\nOut9_14[7] , \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , 
        \nOut9_14[3] , \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }), .WestIn(
        {\nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }), .Out({
        \nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_751 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut752[7] , \nScanOut752[6] , 
        \nScanOut752[5] , \nScanOut752[4] , \nScanOut752[3] , \nScanOut752[2] , 
        \nScanOut752[1] , \nScanOut752[0] }), .ScanOut({\nScanOut751[7] , 
        \nScanOut751[6] , \nScanOut751[5] , \nScanOut751[4] , \nScanOut751[3] , 
        \nScanOut751[2] , \nScanOut751[1] , \nScanOut751[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_14[7] , \nOut23_14[6] , \nOut23_14[5] , \nOut23_14[4] , 
        \nOut23_14[3] , \nOut23_14[2] , \nOut23_14[1] , \nOut23_14[0] }), 
        .SouthIn({\nOut23_16[7] , \nOut23_16[6] , \nOut23_16[5] , 
        \nOut23_16[4] , \nOut23_16[3] , \nOut23_16[2] , \nOut23_16[1] , 
        \nOut23_16[0] }), .EastIn({\nOut24_15[7] , \nOut24_15[6] , 
        \nOut24_15[5] , \nOut24_15[4] , \nOut24_15[3] , \nOut24_15[2] , 
        \nOut24_15[1] , \nOut24_15[0] }), .WestIn({\nOut22_15[7] , 
        \nOut22_15[6] , \nOut22_15[5] , \nOut22_15[4] , \nOut22_15[3] , 
        \nOut22_15[2] , \nOut22_15[1] , \nOut22_15[0] }), .Out({\nOut23_15[7] , 
        \nOut23_15[6] , \nOut23_15[5] , \nOut23_15[4] , \nOut23_15[3] , 
        \nOut23_15[2] , \nOut23_15[1] , \nOut23_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_446 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut447[7] , \nScanOut447[6] , 
        \nScanOut447[5] , \nScanOut447[4] , \nScanOut447[3] , \nScanOut447[2] , 
        \nScanOut447[1] , \nScanOut447[0] }), .ScanOut({\nScanOut446[7] , 
        \nScanOut446[6] , \nScanOut446[5] , \nScanOut446[4] , \nScanOut446[3] , 
        \nScanOut446[2] , \nScanOut446[1] , \nScanOut446[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_29[7] , \nOut13_29[6] , \nOut13_29[5] , \nOut13_29[4] , 
        \nOut13_29[3] , \nOut13_29[2] , \nOut13_29[1] , \nOut13_29[0] }), 
        .SouthIn({\nOut13_31[7] , \nOut13_31[6] , \nOut13_31[5] , 
        \nOut13_31[4] , \nOut13_31[3] , \nOut13_31[2] , \nOut13_31[1] , 
        \nOut13_31[0] }), .EastIn({\nOut14_30[7] , \nOut14_30[6] , 
        \nOut14_30[5] , \nOut14_30[4] , \nOut14_30[3] , \nOut14_30[2] , 
        \nOut14_30[1] , \nOut14_30[0] }), .WestIn({\nOut12_30[7] , 
        \nOut12_30[6] , \nOut12_30[5] , \nOut12_30[4] , \nOut12_30[3] , 
        \nOut12_30[2] , \nOut12_30[1] , \nOut12_30[0] }), .Out({\nOut13_30[7] , 
        \nOut13_30[6] , \nOut13_30[5] , \nOut13_30[4] , \nOut13_30[3] , 
        \nOut13_30[2] , \nOut13_30[1] , \nOut13_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_461 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut462[7] , \nScanOut462[6] , 
        \nScanOut462[5] , \nScanOut462[4] , \nScanOut462[3] , \nScanOut462[2] , 
        \nScanOut462[1] , \nScanOut462[0] }), .ScanOut({\nScanOut461[7] , 
        \nScanOut461[6] , \nScanOut461[5] , \nScanOut461[4] , \nScanOut461[3] , 
        \nScanOut461[2] , \nScanOut461[1] , \nScanOut461[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_12[7] , \nOut14_12[6] , \nOut14_12[5] , \nOut14_12[4] , 
        \nOut14_12[3] , \nOut14_12[2] , \nOut14_12[1] , \nOut14_12[0] }), 
        .SouthIn({\nOut14_14[7] , \nOut14_14[6] , \nOut14_14[5] , 
        \nOut14_14[4] , \nOut14_14[3] , \nOut14_14[2] , \nOut14_14[1] , 
        \nOut14_14[0] }), .EastIn({\nOut15_13[7] , \nOut15_13[6] , 
        \nOut15_13[5] , \nOut15_13[4] , \nOut15_13[3] , \nOut15_13[2] , 
        \nOut15_13[1] , \nOut15_13[0] }), .WestIn({\nOut13_13[7] , 
        \nOut13_13[6] , \nOut13_13[5] , \nOut13_13[4] , \nOut13_13[3] , 
        \nOut13_13[2] , \nOut13_13[1] , \nOut13_13[0] }), .Out({\nOut14_13[7] , 
        \nOut14_13[6] , \nOut14_13[5] , \nOut14_13[4] , \nOut14_13[3] , 
        \nOut14_13[2] , \nOut14_13[1] , \nOut14_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_813 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut814[7] , \nScanOut814[6] , 
        \nScanOut814[5] , \nScanOut814[4] , \nScanOut814[3] , \nScanOut814[2] , 
        \nScanOut814[1] , \nScanOut814[0] }), .ScanOut({\nScanOut813[7] , 
        \nScanOut813[6] , \nScanOut813[5] , \nScanOut813[4] , \nScanOut813[3] , 
        \nScanOut813[2] , \nScanOut813[1] , \nScanOut813[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_12[7] , \nOut25_12[6] , \nOut25_12[5] , \nOut25_12[4] , 
        \nOut25_12[3] , \nOut25_12[2] , \nOut25_12[1] , \nOut25_12[0] }), 
        .SouthIn({\nOut25_14[7] , \nOut25_14[6] , \nOut25_14[5] , 
        \nOut25_14[4] , \nOut25_14[3] , \nOut25_14[2] , \nOut25_14[1] , 
        \nOut25_14[0] }), .EastIn({\nOut26_13[7] , \nOut26_13[6] , 
        \nOut26_13[5] , \nOut26_13[4] , \nOut26_13[3] , \nOut26_13[2] , 
        \nOut26_13[1] , \nOut26_13[0] }), .WestIn({\nOut24_13[7] , 
        \nOut24_13[6] , \nOut24_13[5] , \nOut24_13[4] , \nOut24_13[3] , 
        \nOut24_13[2] , \nOut24_13[1] , \nOut24_13[0] }), .Out({\nOut25_13[7] , 
        \nOut25_13[6] , \nOut25_13[5] , \nOut25_13[4] , \nOut25_13[3] , 
        \nOut25_13[2] , \nOut25_13[1] , \nOut25_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_983 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut984[7] , \nScanOut984[6] , 
        \nScanOut984[5] , \nScanOut984[4] , \nScanOut984[3] , \nScanOut984[2] , 
        \nScanOut984[1] , \nScanOut984[0] }), .ScanOut({\nScanOut983[7] , 
        \nScanOut983[6] , \nScanOut983[5] , \nScanOut983[4] , \nScanOut983[3] , 
        \nScanOut983[2] , \nScanOut983[1] , \nScanOut983[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_22[7] , \nOut30_22[6] , \nOut30_22[5] , \nOut30_22[4] , 
        \nOut30_22[3] , \nOut30_22[2] , \nOut30_22[1] , \nOut30_22[0] }), 
        .SouthIn({\nOut30_24[7] , \nOut30_24[6] , \nOut30_24[5] , 
        \nOut30_24[4] , \nOut30_24[3] , \nOut30_24[2] , \nOut30_24[1] , 
        \nOut30_24[0] }), .EastIn({\nOut31_23[7] , \nOut31_23[6] , 
        \nOut31_23[5] , \nOut31_23[4] , \nOut31_23[3] , \nOut31_23[2] , 
        \nOut31_23[1] , \nOut31_23[0] }), .WestIn({\nOut29_23[7] , 
        \nOut29_23[6] , \nOut29_23[5] , \nOut29_23[4] , \nOut29_23[3] , 
        \nOut29_23[2] , \nOut29_23[1] , \nOut29_23[0] }), .Out({\nOut30_23[7] , 
        \nOut30_23[6] , \nOut30_23[5] , \nOut30_23[4] , \nOut30_23[3] , 
        \nOut30_23[2] , \nOut30_23[1] , \nOut30_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_776 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut777[7] , \nScanOut777[6] , 
        \nScanOut777[5] , \nScanOut777[4] , \nScanOut777[3] , \nScanOut777[2] , 
        \nScanOut777[1] , \nScanOut777[0] }), .ScanOut({\nScanOut776[7] , 
        \nScanOut776[6] , \nScanOut776[5] , \nScanOut776[4] , \nScanOut776[3] , 
        \nScanOut776[2] , \nScanOut776[1] , \nScanOut776[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_7[7] , \nOut24_7[6] , \nOut24_7[5] , \nOut24_7[4] , 
        \nOut24_7[3] , \nOut24_7[2] , \nOut24_7[1] , \nOut24_7[0] }), 
        .SouthIn({\nOut24_9[7] , \nOut24_9[6] , \nOut24_9[5] , \nOut24_9[4] , 
        \nOut24_9[3] , \nOut24_9[2] , \nOut24_9[1] , \nOut24_9[0] }), .EastIn(
        {\nOut25_8[7] , \nOut25_8[6] , \nOut25_8[5] , \nOut25_8[4] , 
        \nOut25_8[3] , \nOut25_8[2] , \nOut25_8[1] , \nOut25_8[0] }), .WestIn(
        {\nOut23_8[7] , \nOut23_8[6] , \nOut23_8[5] , \nOut23_8[4] , 
        \nOut23_8[3] , \nOut23_8[2] , \nOut23_8[1] , \nOut23_8[0] }), .Out({
        \nOut24_8[7] , \nOut24_8[6] , \nOut24_8[5] , \nOut24_8[4] , 
        \nOut24_8[3] , \nOut24_8[2] , \nOut24_8[1] , \nOut24_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_834 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut835[7] , \nScanOut835[6] , 
        \nScanOut835[5] , \nScanOut835[4] , \nScanOut835[3] , \nScanOut835[2] , 
        \nScanOut835[1] , \nScanOut835[0] }), .ScanOut({\nScanOut834[7] , 
        \nScanOut834[6] , \nScanOut834[5] , \nScanOut834[4] , \nScanOut834[3] , 
        \nScanOut834[2] , \nScanOut834[1] , \nScanOut834[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_1[7] , \nOut26_1[6] , \nOut26_1[5] , \nOut26_1[4] , 
        \nOut26_1[3] , \nOut26_1[2] , \nOut26_1[1] , \nOut26_1[0] }), 
        .SouthIn({\nOut26_3[7] , \nOut26_3[6] , \nOut26_3[5] , \nOut26_3[4] , 
        \nOut26_3[3] , \nOut26_3[2] , \nOut26_3[1] , \nOut26_3[0] }), .EastIn(
        {\nOut27_2[7] , \nOut27_2[6] , \nOut27_2[5] , \nOut27_2[4] , 
        \nOut27_2[3] , \nOut27_2[2] , \nOut27_2[1] , \nOut27_2[0] }), .WestIn(
        {\nOut25_2[7] , \nOut25_2[6] , \nOut25_2[5] , \nOut25_2[4] , 
        \nOut25_2[3] , \nOut25_2[2] , \nOut25_2[1] , \nOut25_2[0] }), .Out({
        \nOut26_2[7] , \nOut26_2[6] , \nOut26_2[5] , \nOut26_2[4] , 
        \nOut26_2[3] , \nOut26_2[2] , \nOut26_2[1] , \nOut26_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_898 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut899[7] , \nScanOut899[6] , 
        \nScanOut899[5] , \nScanOut899[4] , \nScanOut899[3] , \nScanOut899[2] , 
        \nScanOut899[1] , \nScanOut899[0] }), .ScanOut({\nScanOut898[7] , 
        \nScanOut898[6] , \nScanOut898[5] , \nScanOut898[4] , \nScanOut898[3] , 
        \nScanOut898[2] , \nScanOut898[1] , \nScanOut898[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_1[7] , \nOut28_1[6] , \nOut28_1[5] , \nOut28_1[4] , 
        \nOut28_1[3] , \nOut28_1[2] , \nOut28_1[1] , \nOut28_1[0] }), 
        .SouthIn({\nOut28_3[7] , \nOut28_3[6] , \nOut28_3[5] , \nOut28_3[4] , 
        \nOut28_3[3] , \nOut28_3[2] , \nOut28_3[1] , \nOut28_3[0] }), .EastIn(
        {\nOut29_2[7] , \nOut29_2[6] , \nOut29_2[5] , \nOut29_2[4] , 
        \nOut29_2[3] , \nOut29_2[2] , \nOut29_2[1] , \nOut29_2[0] }), .WestIn(
        {\nOut27_2[7] , \nOut27_2[6] , \nOut27_2[5] , \nOut27_2[4] , 
        \nOut27_2[3] , \nOut27_2[2] , \nOut27_2[1] , \nOut27_2[0] }), .Out({
        \nOut28_2[7] , \nOut28_2[6] , \nOut28_2[5] , \nOut28_2[4] , 
        \nOut28_2[3] , \nOut28_2[2] , \nOut28_2[1] , \nOut28_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_908 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut909[7] , \nScanOut909[6] , 
        \nScanOut909[5] , \nScanOut909[4] , \nScanOut909[3] , \nScanOut909[2] , 
        \nScanOut909[1] , \nScanOut909[0] }), .ScanOut({\nScanOut908[7] , 
        \nScanOut908[6] , \nScanOut908[5] , \nScanOut908[4] , \nScanOut908[3] , 
        \nScanOut908[2] , \nScanOut908[1] , \nScanOut908[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_11[7] , \nOut28_11[6] , \nOut28_11[5] , \nOut28_11[4] , 
        \nOut28_11[3] , \nOut28_11[2] , \nOut28_11[1] , \nOut28_11[0] }), 
        .SouthIn({\nOut28_13[7] , \nOut28_13[6] , \nOut28_13[5] , 
        \nOut28_13[4] , \nOut28_13[3] , \nOut28_13[2] , \nOut28_13[1] , 
        \nOut28_13[0] }), .EastIn({\nOut29_12[7] , \nOut29_12[6] , 
        \nOut29_12[5] , \nOut29_12[4] , \nOut29_12[3] , \nOut29_12[2] , 
        \nOut29_12[1] , \nOut29_12[0] }), .WestIn({\nOut27_12[7] , 
        \nOut27_12[6] , \nOut27_12[5] , \nOut27_12[4] , \nOut27_12[3] , 
        \nOut27_12[2] , \nOut27_12[1] , \nOut27_12[0] }), .Out({\nOut28_12[7] , 
        \nOut28_12[6] , \nOut28_12[5] , \nOut28_12[4] , \nOut28_12[3] , 
        \nOut28_12[2] , \nOut28_12[1] , \nOut28_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_322 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut323[7] , \nScanOut323[6] , 
        \nScanOut323[5] , \nScanOut323[4] , \nScanOut323[3] , \nScanOut323[2] , 
        \nScanOut323[1] , \nScanOut323[0] }), .ScanOut({\nScanOut322[7] , 
        \nScanOut322[6] , \nScanOut322[5] , \nScanOut322[4] , \nScanOut322[3] , 
        \nScanOut322[2] , \nScanOut322[1] , \nScanOut322[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_1[7] , \nOut10_1[6] , \nOut10_1[5] , \nOut10_1[4] , 
        \nOut10_1[3] , \nOut10_1[2] , \nOut10_1[1] , \nOut10_1[0] }), 
        .SouthIn({\nOut10_3[7] , \nOut10_3[6] , \nOut10_3[5] , \nOut10_3[4] , 
        \nOut10_3[3] , \nOut10_3[2] , \nOut10_3[1] , \nOut10_3[0] }), .EastIn(
        {\nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }), .WestIn(
        {\nOut9_2[7] , \nOut9_2[6] , \nOut9_2[5] , \nOut9_2[4] , \nOut9_2[3] , 
        \nOut9_2[2] , \nOut9_2[1] , \nOut9_2[0] }), .Out({\nOut10_2[7] , 
        \nOut10_2[6] , \nOut10_2[5] , \nOut10_2[4] , \nOut10_2[3] , 
        \nOut10_2[2] , \nOut10_2[1] , \nOut10_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_533 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut534[7] , \nScanOut534[6] , 
        \nScanOut534[5] , \nScanOut534[4] , \nScanOut534[3] , \nScanOut534[2] , 
        \nScanOut534[1] , \nScanOut534[0] }), .ScanOut({\nScanOut533[7] , 
        \nScanOut533[6] , \nScanOut533[5] , \nScanOut533[4] , \nScanOut533[3] , 
        \nScanOut533[2] , \nScanOut533[1] , \nScanOut533[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_20[7] , \nOut16_20[6] , \nOut16_20[5] , \nOut16_20[4] , 
        \nOut16_20[3] , \nOut16_20[2] , \nOut16_20[1] , \nOut16_20[0] }), 
        .SouthIn({\nOut16_22[7] , \nOut16_22[6] , \nOut16_22[5] , 
        \nOut16_22[4] , \nOut16_22[3] , \nOut16_22[2] , \nOut16_22[1] , 
        \nOut16_22[0] }), .EastIn({\nOut17_21[7] , \nOut17_21[6] , 
        \nOut17_21[5] , \nOut17_21[4] , \nOut17_21[3] , \nOut17_21[2] , 
        \nOut17_21[1] , \nOut17_21[0] }), .WestIn({\nOut15_21[7] , 
        \nOut15_21[6] , \nOut15_21[5] , \nOut15_21[4] , \nOut15_21[3] , 
        \nOut15_21[2] , \nOut15_21[1] , \nOut15_21[0] }), .Out({\nOut16_21[7] , 
        \nOut16_21[6] , \nOut16_21[5] , \nOut16_21[4] , \nOut16_21[3] , 
        \nOut16_21[2] , \nOut16_21[1] , \nOut16_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_941 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut942[7] , \nScanOut942[6] , 
        \nScanOut942[5] , \nScanOut942[4] , \nScanOut942[3] , \nScanOut942[2] , 
        \nScanOut942[1] , \nScanOut942[0] }), .ScanOut({\nScanOut941[7] , 
        \nScanOut941[6] , \nScanOut941[5] , \nScanOut941[4] , \nScanOut941[3] , 
        \nScanOut941[2] , \nScanOut941[1] , \nScanOut941[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_12[7] , \nOut29_12[6] , \nOut29_12[5] , \nOut29_12[4] , 
        \nOut29_12[3] , \nOut29_12[2] , \nOut29_12[1] , \nOut29_12[0] }), 
        .SouthIn({\nOut29_14[7] , \nOut29_14[6] , \nOut29_14[5] , 
        \nOut29_14[4] , \nOut29_14[3] , \nOut29_14[2] , \nOut29_14[1] , 
        \nOut29_14[0] }), .EastIn({\nOut30_13[7] , \nOut30_13[6] , 
        \nOut30_13[5] , \nOut30_13[4] , \nOut30_13[3] , \nOut30_13[2] , 
        \nOut30_13[1] , \nOut30_13[0] }), .WestIn({\nOut28_13[7] , 
        \nOut28_13[6] , \nOut28_13[5] , \nOut28_13[4] , \nOut28_13[3] , 
        \nOut28_13[2] , \nOut28_13[1] , \nOut28_13[0] }), .Out({\nOut29_13[7] , 
        \nOut29_13[6] , \nOut29_13[5] , \nOut29_13[4] , \nOut29_13[3] , 
        \nOut29_13[2] , \nOut29_13[1] , \nOut29_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_18 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut19[7] , \nScanOut19[6] , 
        \nScanOut19[5] , \nScanOut19[4] , \nScanOut19[3] , \nScanOut19[2] , 
        \nScanOut19[1] , \nScanOut19[0] }), .ScanOut({\nScanOut18[7] , 
        \nScanOut18[6] , \nScanOut18[5] , \nScanOut18[4] , \nScanOut18[3] , 
        \nScanOut18[2] , \nScanOut18[1] , \nScanOut18[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_18[7] , \nOut0_18[6] , 
        \nOut0_18[5] , \nOut0_18[4] , \nOut0_18[3] , \nOut0_18[2] , 
        \nOut0_18[1] , \nOut0_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_23 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut24[7] , \nScanOut24[6] , 
        \nScanOut24[5] , \nScanOut24[4] , \nScanOut24[3] , \nScanOut24[2] , 
        \nScanOut24[1] , \nScanOut24[0] }), .ScanOut({\nScanOut23[7] , 
        \nScanOut23[6] , \nScanOut23[5] , \nScanOut23[4] , \nScanOut23[3] , 
        \nScanOut23[2] , \nScanOut23[1] , \nScanOut23[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_23[7] , \nOut0_23[6] , 
        \nOut0_23[5] , \nOut0_23[4] , \nOut0_23[3] , \nOut0_23[2] , 
        \nOut0_23[1] , \nOut0_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_31 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut32[7] , \nScanOut32[6] , 
        \nScanOut32[5] , \nScanOut32[4] , \nScanOut32[3] , \nScanOut32[2] , 
        \nScanOut32[1] , \nScanOut32[0] }), .ScanOut({\nScanOut31[7] , 
        \nScanOut31[6] , \nScanOut31[5] , \nScanOut31[4] , \nScanOut31[3] , 
        \nScanOut31[2] , \nScanOut31[1] , \nScanOut31[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_182 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut183[7] , \nScanOut183[6] , 
        \nScanOut183[5] , \nScanOut183[4] , \nScanOut183[3] , \nScanOut183[2] , 
        \nScanOut183[1] , \nScanOut183[0] }), .ScanOut({\nScanOut182[7] , 
        \nScanOut182[6] , \nScanOut182[5] , \nScanOut182[4] , \nScanOut182[3] , 
        \nScanOut182[2] , \nScanOut182[1] , \nScanOut182[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_21[7] , \nOut5_21[6] , \nOut5_21[5] , \nOut5_21[4] , 
        \nOut5_21[3] , \nOut5_21[2] , \nOut5_21[1] , \nOut5_21[0] }), 
        .SouthIn({\nOut5_23[7] , \nOut5_23[6] , \nOut5_23[5] , \nOut5_23[4] , 
        \nOut5_23[3] , \nOut5_23[2] , \nOut5_23[1] , \nOut5_23[0] }), .EastIn(
        {\nOut6_22[7] , \nOut6_22[6] , \nOut6_22[5] , \nOut6_22[4] , 
        \nOut6_22[3] , \nOut6_22[2] , \nOut6_22[1] , \nOut6_22[0] }), .WestIn(
        {\nOut4_22[7] , \nOut4_22[6] , \nOut4_22[5] , \nOut4_22[4] , 
        \nOut4_22[3] , \nOut4_22[2] , \nOut4_22[1] , \nOut4_22[0] }), .Out({
        \nOut5_22[7] , \nOut5_22[6] , \nOut5_22[5] , \nOut5_22[4] , 
        \nOut5_22[3] , \nOut5_22[2] , \nOut5_22[1] , \nOut5_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_603 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut604[7] , \nScanOut604[6] , 
        \nScanOut604[5] , \nScanOut604[4] , \nScanOut604[3] , \nScanOut604[2] , 
        \nScanOut604[1] , \nScanOut604[0] }), .ScanOut({\nScanOut603[7] , 
        \nScanOut603[6] , \nScanOut603[5] , \nScanOut603[4] , \nScanOut603[3] , 
        \nScanOut603[2] , \nScanOut603[1] , \nScanOut603[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_26[7] , \nOut18_26[6] , \nOut18_26[5] , \nOut18_26[4] , 
        \nOut18_26[3] , \nOut18_26[2] , \nOut18_26[1] , \nOut18_26[0] }), 
        .SouthIn({\nOut18_28[7] , \nOut18_28[6] , \nOut18_28[5] , 
        \nOut18_28[4] , \nOut18_28[3] , \nOut18_28[2] , \nOut18_28[1] , 
        \nOut18_28[0] }), .EastIn({\nOut19_27[7] , \nOut19_27[6] , 
        \nOut19_27[5] , \nOut19_27[4] , \nOut19_27[3] , \nOut19_27[2] , 
        \nOut19_27[1] , \nOut19_27[0] }), .WestIn({\nOut17_27[7] , 
        \nOut17_27[6] , \nOut17_27[5] , \nOut17_27[4] , \nOut17_27[3] , 
        \nOut17_27[2] , \nOut17_27[1] , \nOut17_27[0] }), .Out({\nOut18_27[7] , 
        \nOut18_27[6] , \nOut18_27[5] , \nOut18_27[4] , \nOut18_27[3] , 
        \nOut18_27[2] , \nOut18_27[1] , \nOut18_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_793 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut794[7] , \nScanOut794[6] , 
        \nScanOut794[5] , \nScanOut794[4] , \nScanOut794[3] , \nScanOut794[2] , 
        \nScanOut794[1] , \nScanOut794[0] }), .ScanOut({\nScanOut793[7] , 
        \nScanOut793[6] , \nScanOut793[5] , \nScanOut793[4] , \nScanOut793[3] , 
        \nScanOut793[2] , \nScanOut793[1] , \nScanOut793[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_24[7] , \nOut24_24[6] , \nOut24_24[5] , \nOut24_24[4] , 
        \nOut24_24[3] , \nOut24_24[2] , \nOut24_24[1] , \nOut24_24[0] }), 
        .SouthIn({\nOut24_26[7] , \nOut24_26[6] , \nOut24_26[5] , 
        \nOut24_26[4] , \nOut24_26[3] , \nOut24_26[2] , \nOut24_26[1] , 
        \nOut24_26[0] }), .EastIn({\nOut25_25[7] , \nOut25_25[6] , 
        \nOut25_25[5] , \nOut25_25[4] , \nOut25_25[3] , \nOut25_25[2] , 
        \nOut25_25[1] , \nOut25_25[0] }), .WestIn({\nOut23_25[7] , 
        \nOut23_25[6] , \nOut23_25[5] , \nOut23_25[4] , \nOut23_25[3] , 
        \nOut23_25[2] , \nOut23_25[1] , \nOut23_25[0] }), .Out({\nOut24_25[7] , 
        \nOut24_25[6] , \nOut24_25[5] , \nOut24_25[4] , \nOut24_25[3] , 
        \nOut24_25[2] , \nOut24_25[1] , \nOut24_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_109 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut110[7] , \nScanOut110[6] , 
        \nScanOut110[5] , \nScanOut110[4] , \nScanOut110[3] , \nScanOut110[2] , 
        \nScanOut110[1] , \nScanOut110[0] }), .ScanOut({\nScanOut109[7] , 
        \nScanOut109[6] , \nScanOut109[5] , \nScanOut109[4] , \nScanOut109[3] , 
        \nScanOut109[2] , \nScanOut109[1] , \nScanOut109[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }), 
        .SouthIn({\nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }), .EastIn(
        {\nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }), .WestIn(
        {\nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), .Out({
        \nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_239 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut240[7] , \nScanOut240[6] , 
        \nScanOut240[5] , \nScanOut240[4] , \nScanOut240[3] , \nScanOut240[2] , 
        \nScanOut240[1] , \nScanOut240[0] }), .ScanOut({\nScanOut239[7] , 
        \nScanOut239[6] , \nScanOut239[5] , \nScanOut239[4] , \nScanOut239[3] , 
        \nScanOut239[2] , \nScanOut239[1] , \nScanOut239[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }), 
        .SouthIn({\nOut7_16[7] , \nOut7_16[6] , \nOut7_16[5] , \nOut7_16[4] , 
        \nOut7_16[3] , \nOut7_16[2] , \nOut7_16[1] , \nOut7_16[0] }), .EastIn(
        {\nOut8_15[7] , \nOut8_15[6] , \nOut8_15[5] , \nOut8_15[4] , 
        \nOut8_15[3] , \nOut8_15[2] , \nOut8_15[1] , \nOut8_15[0] }), .WestIn(
        {\nOut6_15[7] , \nOut6_15[6] , \nOut6_15[5] , \nOut6_15[4] , 
        \nOut6_15[3] , \nOut6_15[2] , \nOut6_15[1] , \nOut6_15[0] }), .Out({
        \nOut7_15[7] , \nOut7_15[6] , \nOut7_15[5] , \nOut7_15[4] , 
        \nOut7_15[3] , \nOut7_15[2] , \nOut7_15[1] , \nOut7_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_295 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut296[7] , \nScanOut296[6] , 
        \nScanOut296[5] , \nScanOut296[4] , \nScanOut296[3] , \nScanOut296[2] , 
        \nScanOut296[1] , \nScanOut296[0] }), .ScanOut({\nScanOut295[7] , 
        \nScanOut295[6] , \nScanOut295[5] , \nScanOut295[4] , \nScanOut295[3] , 
        \nScanOut295[2] , \nScanOut295[1] , \nScanOut295[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_6[7] , \nOut9_6[6] , \nOut9_6[5] , \nOut9_6[4] , \nOut9_6[3] , 
        \nOut9_6[2] , \nOut9_6[1] , \nOut9_6[0] }), .SouthIn({\nOut9_8[7] , 
        \nOut9_8[6] , \nOut9_8[5] , \nOut9_8[4] , \nOut9_8[3] , \nOut9_8[2] , 
        \nOut9_8[1] , \nOut9_8[0] }), .EastIn({\nOut10_7[7] , \nOut10_7[6] , 
        \nOut10_7[5] , \nOut10_7[4] , \nOut10_7[3] , \nOut10_7[2] , 
        \nOut10_7[1] , \nOut10_7[0] }), .WestIn({\nOut8_7[7] , \nOut8_7[6] , 
        \nOut8_7[5] , \nOut8_7[4] , \nOut8_7[3] , \nOut8_7[2] , \nOut8_7[1] , 
        \nOut8_7[0] }), .Out({\nOut9_7[7] , \nOut9_7[6] , \nOut9_7[5] , 
        \nOut9_7[4] , \nOut9_7[3] , \nOut9_7[2] , \nOut9_7[1] , \nOut9_7[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_305 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut306[7] , \nScanOut306[6] , 
        \nScanOut306[5] , \nScanOut306[4] , \nScanOut306[3] , \nScanOut306[2] , 
        \nScanOut306[1] , \nScanOut306[0] }), .ScanOut({\nScanOut305[7] , 
        \nScanOut305[6] , \nScanOut305[5] , \nScanOut305[4] , \nScanOut305[3] , 
        \nScanOut305[2] , \nScanOut305[1] , \nScanOut305[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_16[7] , \nOut9_16[6] , \nOut9_16[5] , \nOut9_16[4] , 
        \nOut9_16[3] , \nOut9_16[2] , \nOut9_16[1] , \nOut9_16[0] }), 
        .SouthIn({\nOut9_18[7] , \nOut9_18[6] , \nOut9_18[5] , \nOut9_18[4] , 
        \nOut9_18[3] , \nOut9_18[2] , \nOut9_18[1] , \nOut9_18[0] }), .EastIn(
        {\nOut10_17[7] , \nOut10_17[6] , \nOut10_17[5] , \nOut10_17[4] , 
        \nOut10_17[3] , \nOut10_17[2] , \nOut10_17[1] , \nOut10_17[0] }), 
        .WestIn({\nOut8_17[7] , \nOut8_17[6] , \nOut8_17[5] , \nOut8_17[4] , 
        \nOut8_17[3] , \nOut8_17[2] , \nOut8_17[1] , \nOut8_17[0] }), .Out({
        \nOut9_17[7] , \nOut9_17[6] , \nOut9_17[5] , \nOut9_17[4] , 
        \nOut9_17[3] , \nOut9_17[2] , \nOut9_17[1] , \nOut9_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_484 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut485[7] , \nScanOut485[6] , 
        \nScanOut485[5] , \nScanOut485[4] , \nScanOut485[3] , \nScanOut485[2] , 
        \nScanOut485[1] , \nScanOut485[0] }), .ScanOut({\nScanOut484[7] , 
        \nScanOut484[6] , \nScanOut484[5] , \nScanOut484[4] , \nScanOut484[3] , 
        \nScanOut484[2] , \nScanOut484[1] , \nScanOut484[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_3[7] , \nOut15_3[6] , \nOut15_3[5] , \nOut15_3[4] , 
        \nOut15_3[3] , \nOut15_3[2] , \nOut15_3[1] , \nOut15_3[0] }), 
        .SouthIn({\nOut15_5[7] , \nOut15_5[6] , \nOut15_5[5] , \nOut15_5[4] , 
        \nOut15_5[3] , \nOut15_5[2] , \nOut15_5[1] , \nOut15_5[0] }), .EastIn(
        {\nOut16_4[7] , \nOut16_4[6] , \nOut16_4[5] , \nOut16_4[4] , 
        \nOut16_4[3] , \nOut16_4[2] , \nOut16_4[1] , \nOut16_4[0] }), .WestIn(
        {\nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }), .Out({
        \nOut15_4[7] , \nOut15_4[6] , \nOut15_4[5] , \nOut15_4[4] , 
        \nOut15_4[3] , \nOut15_4[2] , \nOut15_4[1] , \nOut15_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_624 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut625[7] , \nScanOut625[6] , 
        \nScanOut625[5] , \nScanOut625[4] , \nScanOut625[3] , \nScanOut625[2] , 
        \nScanOut625[1] , \nScanOut625[0] }), .ScanOut({\nScanOut624[7] , 
        \nScanOut624[6] , \nScanOut624[5] , \nScanOut624[4] , \nScanOut624[3] , 
        \nScanOut624[2] , \nScanOut624[1] , \nScanOut624[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_15[7] , \nOut19_15[6] , \nOut19_15[5] , \nOut19_15[4] , 
        \nOut19_15[3] , \nOut19_15[2] , \nOut19_15[1] , \nOut19_15[0] }), 
        .SouthIn({\nOut19_17[7] , \nOut19_17[6] , \nOut19_17[5] , 
        \nOut19_17[4] , \nOut19_17[3] , \nOut19_17[2] , \nOut19_17[1] , 
        \nOut19_17[0] }), .EastIn({\nOut20_16[7] , \nOut20_16[6] , 
        \nOut20_16[5] , \nOut20_16[4] , \nOut20_16[3] , \nOut20_16[2] , 
        \nOut20_16[1] , \nOut20_16[0] }), .WestIn({\nOut18_16[7] , 
        \nOut18_16[6] , \nOut18_16[5] , \nOut18_16[4] , \nOut18_16[3] , 
        \nOut18_16[2] , \nOut18_16[1] , \nOut18_16[0] }), .Out({\nOut19_16[7] , 
        \nOut19_16[6] , \nOut19_16[5] , \nOut19_16[4] , \nOut19_16[3] , 
        \nOut19_16[2] , \nOut19_16[1] , \nOut19_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_514 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut515[7] , \nScanOut515[6] , 
        \nScanOut515[5] , \nScanOut515[4] , \nScanOut515[3] , \nScanOut515[2] , 
        \nScanOut515[1] , \nScanOut515[0] }), .ScanOut({\nScanOut514[7] , 
        \nScanOut514[6] , \nScanOut514[5] , \nScanOut514[4] , \nScanOut514[3] , 
        \nScanOut514[2] , \nScanOut514[1] , \nScanOut514[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_1[7] , \nOut16_1[6] , \nOut16_1[5] , \nOut16_1[4] , 
        \nOut16_1[3] , \nOut16_1[2] , \nOut16_1[1] , \nOut16_1[0] }), 
        .SouthIn({\nOut16_3[7] , \nOut16_3[6] , \nOut16_3[5] , \nOut16_3[4] , 
        \nOut16_3[3] , \nOut16_3[2] , \nOut16_3[1] , \nOut16_3[0] }), .EastIn(
        {\nOut17_2[7] , \nOut17_2[6] , \nOut17_2[5] , \nOut17_2[4] , 
        \nOut17_2[3] , \nOut17_2[2] , \nOut17_2[1] , \nOut17_2[0] }), .WestIn(
        {\nOut15_2[7] , \nOut15_2[6] , \nOut15_2[5] , \nOut15_2[4] , 
        \nOut15_2[3] , \nOut15_2[2] , \nOut15_2[1] , \nOut15_2[0] }), .Out({
        \nOut16_2[7] , \nOut16_2[6] , \nOut16_2[5] , \nOut16_2[4] , 
        \nOut16_2[3] , \nOut16_2[2] , \nOut16_2[1] , \nOut16_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_966 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut967[7] , \nScanOut967[6] , 
        \nScanOut967[5] , \nScanOut967[4] , \nScanOut967[3] , \nScanOut967[2] , 
        \nScanOut967[1] , \nScanOut967[0] }), .ScanOut({\nScanOut966[7] , 
        \nScanOut966[6] , \nScanOut966[5] , \nScanOut966[4] , \nScanOut966[3] , 
        \nScanOut966[2] , \nScanOut966[1] , \nScanOut966[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_5[7] , \nOut30_5[6] , \nOut30_5[5] , \nOut30_5[4] , 
        \nOut30_5[3] , \nOut30_5[2] , \nOut30_5[1] , \nOut30_5[0] }), 
        .SouthIn({\nOut30_7[7] , \nOut30_7[6] , \nOut30_7[5] , \nOut30_7[4] , 
        \nOut30_7[3] , \nOut30_7[2] , \nOut30_7[1] , \nOut30_7[0] }), .EastIn(
        {\nOut31_6[7] , \nOut31_6[6] , \nOut31_6[5] , \nOut31_6[4] , 
        \nOut31_6[3] , \nOut31_6[2] , \nOut31_6[1] , \nOut31_6[0] }), .WestIn(
        {\nOut29_6[7] , \nOut29_6[6] , \nOut29_6[5] , \nOut29_6[4] , 
        \nOut29_6[3] , \nOut29_6[2] , \nOut29_6[1] , \nOut29_6[0] }), .Out({
        \nOut30_6[7] , \nOut30_6[6] , \nOut30_6[5] , \nOut30_6[4] , 
        \nOut30_6[3] , \nOut30_6[2] , \nOut30_6[1] , \nOut30_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_428 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut429[7] , \nScanOut429[6] , 
        \nScanOut429[5] , \nScanOut429[4] , \nScanOut429[3] , \nScanOut429[2] , 
        \nScanOut429[1] , \nScanOut429[0] }), .ScanOut({\nScanOut428[7] , 
        \nScanOut428[6] , \nScanOut428[5] , \nScanOut428[4] , \nScanOut428[3] , 
        \nScanOut428[2] , \nScanOut428[1] , \nScanOut428[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_11[7] , \nOut13_11[6] , \nOut13_11[5] , \nOut13_11[4] , 
        \nOut13_11[3] , \nOut13_11[2] , \nOut13_11[1] , \nOut13_11[0] }), 
        .SouthIn({\nOut13_13[7] , \nOut13_13[6] , \nOut13_13[5] , 
        \nOut13_13[4] , \nOut13_13[3] , \nOut13_13[2] , \nOut13_13[1] , 
        \nOut13_13[0] }), .EastIn({\nOut14_12[7] , \nOut14_12[6] , 
        \nOut14_12[5] , \nOut14_12[4] , \nOut14_12[3] , \nOut14_12[2] , 
        \nOut14_12[1] , \nOut14_12[0] }), .WestIn({\nOut12_12[7] , 
        \nOut12_12[6] , \nOut12_12[5] , \nOut12_12[4] , \nOut12_12[3] , 
        \nOut12_12[2] , \nOut12_12[1] , \nOut12_12[0] }), .Out({\nOut13_12[7] , 
        \nOut13_12[6] , \nOut13_12[5] , \nOut13_12[4] , \nOut13_12[3] , 
        \nOut13_12[2] , \nOut13_12[1] , \nOut13_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_190 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut191[7] , \nScanOut191[6] , 
        \nScanOut191[5] , \nScanOut191[4] , \nScanOut191[3] , \nScanOut191[2] , 
        \nScanOut191[1] , \nScanOut191[0] }), .ScanOut({\nScanOut190[7] , 
        \nScanOut190[6] , \nScanOut190[5] , \nScanOut190[4] , \nScanOut190[3] , 
        \nScanOut190[2] , \nScanOut190[1] , \nScanOut190[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_29[7] , \nOut5_29[6] , \nOut5_29[5] , \nOut5_29[4] , 
        \nOut5_29[3] , \nOut5_29[2] , \nOut5_29[1] , \nOut5_29[0] }), 
        .SouthIn({\nOut5_31[7] , \nOut5_31[6] , \nOut5_31[5] , \nOut5_31[4] , 
        \nOut5_31[3] , \nOut5_31[2] , \nOut5_31[1] , \nOut5_31[0] }), .EastIn(
        {\nOut6_30[7] , \nOut6_30[6] , \nOut6_30[5] , \nOut6_30[4] , 
        \nOut6_30[3] , \nOut6_30[2] , \nOut6_30[1] , \nOut6_30[0] }), .WestIn(
        {\nOut4_30[7] , \nOut4_30[6] , \nOut4_30[5] , \nOut4_30[4] , 
        \nOut4_30[3] , \nOut4_30[2] , \nOut4_30[1] , \nOut4_30[0] }), .Out({
        \nOut5_30[7] , \nOut5_30[6] , \nOut5_30[5] , \nOut5_30[4] , 
        \nOut5_30[3] , \nOut5_30[2] , \nOut5_30[1] , \nOut5_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_330 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut331[7] , \nScanOut331[6] , 
        \nScanOut331[5] , \nScanOut331[4] , \nScanOut331[3] , \nScanOut331[2] , 
        \nScanOut331[1] , \nScanOut331[0] }), .ScanOut({\nScanOut330[7] , 
        \nScanOut330[6] , \nScanOut330[5] , \nScanOut330[4] , \nScanOut330[3] , 
        \nScanOut330[2] , \nScanOut330[1] , \nScanOut330[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_9[7] , \nOut10_9[6] , \nOut10_9[5] , \nOut10_9[4] , 
        \nOut10_9[3] , \nOut10_9[2] , \nOut10_9[1] , \nOut10_9[0] }), 
        .SouthIn({\nOut10_11[7] , \nOut10_11[6] , \nOut10_11[5] , 
        \nOut10_11[4] , \nOut10_11[3] , \nOut10_11[2] , \nOut10_11[1] , 
        \nOut10_11[0] }), .EastIn({\nOut11_10[7] , \nOut11_10[6] , 
        \nOut11_10[5] , \nOut11_10[4] , \nOut11_10[3] , \nOut11_10[2] , 
        \nOut11_10[1] , \nOut11_10[0] }), .WestIn({\nOut9_10[7] , 
        \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , \nOut9_10[3] , 
        \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }), .Out({\nOut10_10[7] , 
        \nOut10_10[6] , \nOut10_10[5] , \nOut10_10[4] , \nOut10_10[3] , 
        \nOut10_10[2] , \nOut10_10[1] , \nOut10_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_688 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut689[7] , \nScanOut689[6] , 
        \nScanOut689[5] , \nScanOut689[4] , \nScanOut689[3] , \nScanOut689[2] , 
        \nScanOut689[1] , \nScanOut689[0] }), .ScanOut({\nScanOut688[7] , 
        \nScanOut688[6] , \nScanOut688[5] , \nScanOut688[4] , \nScanOut688[3] , 
        \nScanOut688[2] , \nScanOut688[1] , \nScanOut688[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_15[7] , \nOut21_15[6] , \nOut21_15[5] , \nOut21_15[4] , 
        \nOut21_15[3] , \nOut21_15[2] , \nOut21_15[1] , \nOut21_15[0] }), 
        .SouthIn({\nOut21_17[7] , \nOut21_17[6] , \nOut21_17[5] , 
        \nOut21_17[4] , \nOut21_17[3] , \nOut21_17[2] , \nOut21_17[1] , 
        \nOut21_17[0] }), .EastIn({\nOut22_16[7] , \nOut22_16[6] , 
        \nOut22_16[5] , \nOut22_16[4] , \nOut22_16[3] , \nOut22_16[2] , 
        \nOut22_16[1] , \nOut22_16[0] }), .WestIn({\nOut20_16[7] , 
        \nOut20_16[6] , \nOut20_16[5] , \nOut20_16[4] , \nOut20_16[3] , 
        \nOut20_16[2] , \nOut20_16[1] , \nOut20_16[0] }), .Out({\nOut21_16[7] , 
        \nOut21_16[6] , \nOut21_16[5] , \nOut21_16[4] , \nOut21_16[3] , 
        \nOut21_16[2] , \nOut21_16[1] , \nOut21_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_718 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut719[7] , \nScanOut719[6] , 
        \nScanOut719[5] , \nScanOut719[4] , \nScanOut719[3] , \nScanOut719[2] , 
        \nScanOut719[1] , \nScanOut719[0] }), .ScanOut({\nScanOut718[7] , 
        \nScanOut718[6] , \nScanOut718[5] , \nScanOut718[4] , \nScanOut718[3] , 
        \nScanOut718[2] , \nScanOut718[1] , \nScanOut718[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_13[7] , \nOut22_13[6] , \nOut22_13[5] , \nOut22_13[4] , 
        \nOut22_13[3] , \nOut22_13[2] , \nOut22_13[1] , \nOut22_13[0] }), 
        .SouthIn({\nOut22_15[7] , \nOut22_15[6] , \nOut22_15[5] , 
        \nOut22_15[4] , \nOut22_15[3] , \nOut22_15[2] , \nOut22_15[1] , 
        \nOut22_15[0] }), .EastIn({\nOut23_14[7] , \nOut23_14[6] , 
        \nOut23_14[5] , \nOut23_14[4] , \nOut23_14[3] , \nOut23_14[2] , 
        \nOut23_14[1] , \nOut23_14[0] }), .WestIn({\nOut21_14[7] , 
        \nOut21_14[6] , \nOut21_14[5] , \nOut21_14[4] , \nOut21_14[3] , 
        \nOut21_14[2] , \nOut21_14[1] , \nOut21_14[0] }), .Out({\nOut22_14[7] , 
        \nOut22_14[6] , \nOut22_14[5] , \nOut22_14[4] , \nOut22_14[3] , 
        \nOut22_14[2] , \nOut22_14[1] , \nOut22_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_848 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut849[7] , \nScanOut849[6] , 
        \nScanOut849[5] , \nScanOut849[4] , \nScanOut849[3] , \nScanOut849[2] , 
        \nScanOut849[1] , \nScanOut849[0] }), .ScanOut({\nScanOut848[7] , 
        \nScanOut848[6] , \nScanOut848[5] , \nScanOut848[4] , \nScanOut848[3] , 
        \nScanOut848[2] , \nScanOut848[1] , \nScanOut848[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_15[7] , \nOut26_15[6] , \nOut26_15[5] , \nOut26_15[4] , 
        \nOut26_15[3] , \nOut26_15[2] , \nOut26_15[1] , \nOut26_15[0] }), 
        .SouthIn({\nOut26_17[7] , \nOut26_17[6] , \nOut26_17[5] , 
        \nOut26_17[4] , \nOut26_17[3] , \nOut26_17[2] , \nOut26_17[1] , 
        \nOut26_17[0] }), .EastIn({\nOut27_16[7] , \nOut27_16[6] , 
        \nOut27_16[5] , \nOut27_16[4] , \nOut27_16[3] , \nOut27_16[2] , 
        \nOut27_16[1] , \nOut27_16[0] }), .WestIn({\nOut25_16[7] , 
        \nOut25_16[6] , \nOut25_16[5] , \nOut25_16[4] , \nOut25_16[3] , 
        \nOut25_16[2] , \nOut25_16[1] , \nOut25_16[0] }), .Out({\nOut26_16[7] , 
        \nOut26_16[6] , \nOut26_16[5] , \nOut26_16[4] , \nOut26_16[3] , 
        \nOut26_16[2] , \nOut26_16[1] , \nOut26_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_953 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut954[7] , \nScanOut954[6] , 
        \nScanOut954[5] , \nScanOut954[4] , \nScanOut954[3] , \nScanOut954[2] , 
        \nScanOut954[1] , \nScanOut954[0] }), .ScanOut({\nScanOut953[7] , 
        \nScanOut953[6] , \nScanOut953[5] , \nScanOut953[4] , \nScanOut953[3] , 
        \nScanOut953[2] , \nScanOut953[1] , \nScanOut953[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_24[7] , \nOut29_24[6] , \nOut29_24[5] , \nOut29_24[4] , 
        \nOut29_24[3] , \nOut29_24[2] , \nOut29_24[1] , \nOut29_24[0] }), 
        .SouthIn({\nOut29_26[7] , \nOut29_26[6] , \nOut29_26[5] , 
        \nOut29_26[4] , \nOut29_26[3] , \nOut29_26[2] , \nOut29_26[1] , 
        \nOut29_26[0] }), .EastIn({\nOut30_25[7] , \nOut30_25[6] , 
        \nOut30_25[5] , \nOut30_25[4] , \nOut30_25[3] , \nOut30_25[2] , 
        \nOut30_25[1] , \nOut30_25[0] }), .WestIn({\nOut28_25[7] , 
        \nOut28_25[6] , \nOut28_25[5] , \nOut28_25[4] , \nOut28_25[3] , 
        \nOut28_25[2] , \nOut28_25[1] , \nOut28_25[0] }), .Out({\nOut29_25[7] , 
        \nOut29_25[6] , \nOut29_25[5] , \nOut29_25[4] , \nOut29_25[3] , 
        \nOut29_25[2] , \nOut29_25[1] , \nOut29_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_521 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut522[7] , \nScanOut522[6] , 
        \nScanOut522[5] , \nScanOut522[4] , \nScanOut522[3] , \nScanOut522[2] , 
        \nScanOut522[1] , \nScanOut522[0] }), .ScanOut({\nScanOut521[7] , 
        \nScanOut521[6] , \nScanOut521[5] , \nScanOut521[4] , \nScanOut521[3] , 
        \nScanOut521[2] , \nScanOut521[1] , \nScanOut521[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_8[7] , \nOut16_8[6] , \nOut16_8[5] , \nOut16_8[4] , 
        \nOut16_8[3] , \nOut16_8[2] , \nOut16_8[1] , \nOut16_8[0] }), 
        .SouthIn({\nOut16_10[7] , \nOut16_10[6] , \nOut16_10[5] , 
        \nOut16_10[4] , \nOut16_10[3] , \nOut16_10[2] , \nOut16_10[1] , 
        \nOut16_10[0] }), .EastIn({\nOut17_9[7] , \nOut17_9[6] , \nOut17_9[5] , 
        \nOut17_9[4] , \nOut17_9[3] , \nOut17_9[2] , \nOut17_9[1] , 
        \nOut17_9[0] }), .WestIn({\nOut15_9[7] , \nOut15_9[6] , \nOut15_9[5] , 
        \nOut15_9[4] , \nOut15_9[3] , \nOut15_9[2] , \nOut15_9[1] , 
        \nOut15_9[0] }), .Out({\nOut16_9[7] , \nOut16_9[6] , \nOut16_9[5] , 
        \nOut16_9[4] , \nOut16_9[3] , \nOut16_9[2] , \nOut16_9[1] , 
        \nOut16_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_781 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut782[7] , \nScanOut782[6] , 
        \nScanOut782[5] , \nScanOut782[4] , \nScanOut782[3] , \nScanOut782[2] , 
        \nScanOut782[1] , \nScanOut782[0] }), .ScanOut({\nScanOut781[7] , 
        \nScanOut781[6] , \nScanOut781[5] , \nScanOut781[4] , \nScanOut781[3] , 
        \nScanOut781[2] , \nScanOut781[1] , \nScanOut781[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_12[7] , \nOut24_12[6] , \nOut24_12[5] , \nOut24_12[4] , 
        \nOut24_12[3] , \nOut24_12[2] , \nOut24_12[1] , \nOut24_12[0] }), 
        .SouthIn({\nOut24_14[7] , \nOut24_14[6] , \nOut24_14[5] , 
        \nOut24_14[4] , \nOut24_14[3] , \nOut24_14[2] , \nOut24_14[1] , 
        \nOut24_14[0] }), .EastIn({\nOut25_13[7] , \nOut25_13[6] , 
        \nOut25_13[5] , \nOut25_13[4] , \nOut25_13[3] , \nOut25_13[2] , 
        \nOut25_13[1] , \nOut25_13[0] }), .WestIn({\nOut23_13[7] , 
        \nOut23_13[6] , \nOut23_13[5] , \nOut23_13[4] , \nOut23_13[3] , 
        \nOut23_13[2] , \nOut23_13[1] , \nOut23_13[0] }), .Out({\nOut24_13[7] , 
        \nOut24_13[6] , \nOut24_13[5] , \nOut24_13[4] , \nOut24_13[3] , 
        \nOut24_13[2] , \nOut24_13[1] , \nOut24_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_611 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut612[7] , \nScanOut612[6] , 
        \nScanOut612[5] , \nScanOut612[4] , \nScanOut612[3] , \nScanOut612[2] , 
        \nScanOut612[1] , \nScanOut612[0] }), .ScanOut({\nScanOut611[7] , 
        \nScanOut611[6] , \nScanOut611[5] , \nScanOut611[4] , \nScanOut611[3] , 
        \nScanOut611[2] , \nScanOut611[1] , \nScanOut611[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_2[7] , \nOut19_2[6] , \nOut19_2[5] , \nOut19_2[4] , 
        \nOut19_2[3] , \nOut19_2[2] , \nOut19_2[1] , \nOut19_2[0] }), 
        .SouthIn({\nOut19_4[7] , \nOut19_4[6] , \nOut19_4[5] , \nOut19_4[4] , 
        \nOut19_4[3] , \nOut19_4[2] , \nOut19_4[1] , \nOut19_4[0] }), .EastIn(
        {\nOut20_3[7] , \nOut20_3[6] , \nOut20_3[5] , \nOut20_3[4] , 
        \nOut20_3[3] , \nOut20_3[2] , \nOut20_3[1] , \nOut20_3[0] }), .WestIn(
        {\nOut18_3[7] , \nOut18_3[6] , \nOut18_3[5] , \nOut18_3[4] , 
        \nOut18_3[3] , \nOut18_3[2] , \nOut18_3[1] , \nOut18_3[0] }), .Out({
        \nOut19_3[7] , \nOut19_3[6] , \nOut19_3[5] , \nOut19_3[4] , 
        \nOut19_3[3] , \nOut19_3[2] , \nOut19_3[1] , \nOut19_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_38 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut39[7] , \nScanOut39[6] , 
        \nScanOut39[5] , \nScanOut39[4] , \nScanOut39[3] , \nScanOut39[2] , 
        \nScanOut39[1] , \nScanOut39[0] }), .ScanOut({\nScanOut38[7] , 
        \nScanOut38[6] , \nScanOut38[5] , \nScanOut38[4] , \nScanOut38[3] , 
        \nScanOut38[2] , \nScanOut38[1] , \nScanOut38[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , \nOut1_5[4] , \nOut1_5[3] , 
        \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }), .SouthIn({\nOut1_7[7] , 
        \nOut1_7[6] , \nOut1_7[5] , \nOut1_7[4] , \nOut1_7[3] , \nOut1_7[2] , 
        \nOut1_7[1] , \nOut1_7[0] }), .EastIn({\nOut2_6[7] , \nOut2_6[6] , 
        \nOut2_6[5] , \nOut2_6[4] , \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , 
        \nOut2_6[0] }), .WestIn({\nOut0_6[7] , \nOut0_6[6] , \nOut0_6[5] , 
        \nOut0_6[4] , \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , \nOut0_6[0] }), 
        .Out({\nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , \nOut1_6[4] , 
        \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_56 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut57[7] , \nScanOut57[6] , 
        \nScanOut57[5] , \nScanOut57[4] , \nScanOut57[3] , \nScanOut57[2] , 
        \nScanOut57[1] , \nScanOut57[0] }), .ScanOut({\nScanOut56[7] , 
        \nScanOut56[6] , \nScanOut56[5] , \nScanOut56[4] , \nScanOut56[3] , 
        \nScanOut56[2] , \nScanOut56[1] , \nScanOut56[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_23[7] , \nOut1_23[6] , \nOut1_23[5] , \nOut1_23[4] , 
        \nOut1_23[3] , \nOut1_23[2] , \nOut1_23[1] , \nOut1_23[0] }), 
        .SouthIn({\nOut1_25[7] , \nOut1_25[6] , \nOut1_25[5] , \nOut1_25[4] , 
        \nOut1_25[3] , \nOut1_25[2] , \nOut1_25[1] , \nOut1_25[0] }), .EastIn(
        {\nOut2_24[7] , \nOut2_24[6] , \nOut2_24[5] , \nOut2_24[4] , 
        \nOut2_24[3] , \nOut2_24[2] , \nOut2_24[1] , \nOut2_24[0] }), .WestIn(
        {\nOut0_24[7] , \nOut0_24[6] , \nOut0_24[5] , \nOut0_24[4] , 
        \nOut0_24[3] , \nOut0_24[2] , \nOut0_24[1] , \nOut0_24[0] }), .Out({
        \nOut1_24[7] , \nOut1_24[6] , \nOut1_24[5] , \nOut1_24[4] , 
        \nOut1_24[3] , \nOut1_24[2] , \nOut1_24[1] , \nOut1_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_71 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut72[7] , \nScanOut72[6] , 
        \nScanOut72[5] , \nScanOut72[4] , \nScanOut72[3] , \nScanOut72[2] , 
        \nScanOut72[1] , \nScanOut72[0] }), .ScanOut({\nScanOut71[7] , 
        \nScanOut71[6] , \nScanOut71[5] , \nScanOut71[4] , \nScanOut71[3] , 
        \nScanOut71[2] , \nScanOut71[1] , \nScanOut71[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_6[7] , \nOut2_6[6] , \nOut2_6[5] , \nOut2_6[4] , \nOut2_6[3] , 
        \nOut2_6[2] , \nOut2_6[1] , \nOut2_6[0] }), .SouthIn({\nOut2_8[7] , 
        \nOut2_8[6] , \nOut2_8[5] , \nOut2_8[4] , \nOut2_8[3] , \nOut2_8[2] , 
        \nOut2_8[1] , \nOut2_8[0] }), .EastIn({\nOut3_7[7] , \nOut3_7[6] , 
        \nOut3_7[5] , \nOut3_7[4] , \nOut3_7[3] , \nOut3_7[2] , \nOut3_7[1] , 
        \nOut3_7[0] }), .WestIn({\nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , 
        \nOut1_7[4] , \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }), 
        .Out({\nOut2_7[7] , \nOut2_7[6] , \nOut2_7[5] , \nOut2_7[4] , 
        \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , \nOut2_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_149 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut150[7] , \nScanOut150[6] , 
        \nScanOut150[5] , \nScanOut150[4] , \nScanOut150[3] , \nScanOut150[2] , 
        \nScanOut150[1] , \nScanOut150[0] }), .ScanOut({\nScanOut149[7] , 
        \nScanOut149[6] , \nScanOut149[5] , \nScanOut149[4] , \nScanOut149[3] , 
        \nScanOut149[2] , \nScanOut149[1] , \nScanOut149[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_20[7] , \nOut4_20[6] , \nOut4_20[5] , \nOut4_20[4] , 
        \nOut4_20[3] , \nOut4_20[2] , \nOut4_20[1] , \nOut4_20[0] }), 
        .SouthIn({\nOut4_22[7] , \nOut4_22[6] , \nOut4_22[5] , \nOut4_22[4] , 
        \nOut4_22[3] , \nOut4_22[2] , \nOut4_22[1] , \nOut4_22[0] }), .EastIn(
        {\nOut5_21[7] , \nOut5_21[6] , \nOut5_21[5] , \nOut5_21[4] , 
        \nOut5_21[3] , \nOut5_21[2] , \nOut5_21[1] , \nOut5_21[0] }), .WestIn(
        {\nOut3_21[7] , \nOut3_21[6] , \nOut3_21[5] , \nOut3_21[4] , 
        \nOut3_21[3] , \nOut3_21[2] , \nOut3_21[1] , \nOut3_21[0] }), .Out({
        \nOut4_21[7] , \nOut4_21[6] , \nOut4_21[5] , \nOut4_21[4] , 
        \nOut4_21[3] , \nOut4_21[2] , \nOut4_21[1] , \nOut4_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_152 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut153[7] , \nScanOut153[6] , 
        \nScanOut153[5] , \nScanOut153[4] , \nScanOut153[3] , \nScanOut153[2] , 
        \nScanOut153[1] , \nScanOut153[0] }), .ScanOut({\nScanOut152[7] , 
        \nScanOut152[6] , \nScanOut152[5] , \nScanOut152[4] , \nScanOut152[3] , 
        \nScanOut152[2] , \nScanOut152[1] , \nScanOut152[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_23[7] , \nOut4_23[6] , \nOut4_23[5] , \nOut4_23[4] , 
        \nOut4_23[3] , \nOut4_23[2] , \nOut4_23[1] , \nOut4_23[0] }), 
        .SouthIn({\nOut4_25[7] , \nOut4_25[6] , \nOut4_25[5] , \nOut4_25[4] , 
        \nOut4_25[3] , \nOut4_25[2] , \nOut4_25[1] , \nOut4_25[0] }), .EastIn(
        {\nOut5_24[7] , \nOut5_24[6] , \nOut5_24[5] , \nOut5_24[4] , 
        \nOut5_24[3] , \nOut5_24[2] , \nOut5_24[1] , \nOut5_24[0] }), .WestIn(
        {\nOut3_24[7] , \nOut3_24[6] , \nOut3_24[5] , \nOut3_24[4] , 
        \nOut3_24[3] , \nOut3_24[2] , \nOut3_24[1] , \nOut3_24[0] }), .Out({
        \nOut4_24[7] , \nOut4_24[6] , \nOut4_24[5] , \nOut4_24[4] , 
        \nOut4_24[3] , \nOut4_24[2] , \nOut4_24[1] , \nOut4_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_287 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut288[7] , \nScanOut288[6] , 
        \nScanOut288[5] , \nScanOut288[4] , \nScanOut288[3] , \nScanOut288[2] , 
        \nScanOut288[1] , \nScanOut288[0] }), .ScanOut({\nScanOut287[7] , 
        \nScanOut287[6] , \nScanOut287[5] , \nScanOut287[4] , \nScanOut287[3] , 
        \nScanOut287[2] , \nScanOut287[1] , \nScanOut287[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut8_31[7] , \nOut8_31[6] , 
        \nOut8_31[5] , \nOut8_31[4] , \nOut8_31[3] , \nOut8_31[2] , 
        \nOut8_31[1] , \nOut8_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_506 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut507[7] , \nScanOut507[6] , 
        \nScanOut507[5] , \nScanOut507[4] , \nScanOut507[3] , \nScanOut507[2] , 
        \nScanOut507[1] , \nScanOut507[0] }), .ScanOut({\nScanOut506[7] , 
        \nScanOut506[6] , \nScanOut506[5] , \nScanOut506[4] , \nScanOut506[3] , 
        \nScanOut506[2] , \nScanOut506[1] , \nScanOut506[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_25[7] , \nOut15_25[6] , \nOut15_25[5] , \nOut15_25[4] , 
        \nOut15_25[3] , \nOut15_25[2] , \nOut15_25[1] , \nOut15_25[0] }), 
        .SouthIn({\nOut15_27[7] , \nOut15_27[6] , \nOut15_27[5] , 
        \nOut15_27[4] , \nOut15_27[3] , \nOut15_27[2] , \nOut15_27[1] , 
        \nOut15_27[0] }), .EastIn({\nOut16_26[7] , \nOut16_26[6] , 
        \nOut16_26[5] , \nOut16_26[4] , \nOut16_26[3] , \nOut16_26[2] , 
        \nOut16_26[1] , \nOut16_26[0] }), .WestIn({\nOut14_26[7] , 
        \nOut14_26[6] , \nOut14_26[5] , \nOut14_26[4] , \nOut14_26[3] , 
        \nOut14_26[2] , \nOut14_26[1] , \nOut14_26[0] }), .Out({\nOut15_26[7] , 
        \nOut15_26[6] , \nOut15_26[5] , \nOut15_26[4] , \nOut15_26[3] , 
        \nOut15_26[2] , \nOut15_26[1] , \nOut15_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_636 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut637[7] , \nScanOut637[6] , 
        \nScanOut637[5] , \nScanOut637[4] , \nScanOut637[3] , \nScanOut637[2] , 
        \nScanOut637[1] , \nScanOut637[0] }), .ScanOut({\nScanOut636[7] , 
        \nScanOut636[6] , \nScanOut636[5] , \nScanOut636[4] , \nScanOut636[3] , 
        \nScanOut636[2] , \nScanOut636[1] , \nScanOut636[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_27[7] , \nOut19_27[6] , \nOut19_27[5] , \nOut19_27[4] , 
        \nOut19_27[3] , \nOut19_27[2] , \nOut19_27[1] , \nOut19_27[0] }), 
        .SouthIn({\nOut19_29[7] , \nOut19_29[6] , \nOut19_29[5] , 
        \nOut19_29[4] , \nOut19_29[3] , \nOut19_29[2] , \nOut19_29[1] , 
        \nOut19_29[0] }), .EastIn({\nOut20_28[7] , \nOut20_28[6] , 
        \nOut20_28[5] , \nOut20_28[4] , \nOut20_28[3] , \nOut20_28[2] , 
        \nOut20_28[1] , \nOut20_28[0] }), .WestIn({\nOut18_28[7] , 
        \nOut18_28[6] , \nOut18_28[5] , \nOut18_28[4] , \nOut18_28[3] , 
        \nOut18_28[2] , \nOut18_28[1] , \nOut18_28[0] }), .Out({\nOut19_28[7] , 
        \nOut19_28[6] , \nOut19_28[5] , \nOut19_28[4] , \nOut19_28[3] , 
        \nOut19_28[2] , \nOut19_28[1] , \nOut19_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_974 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut975[7] , \nScanOut975[6] , 
        \nScanOut975[5] , \nScanOut975[4] , \nScanOut975[3] , \nScanOut975[2] , 
        \nScanOut975[1] , \nScanOut975[0] }), .ScanOut({\nScanOut974[7] , 
        \nScanOut974[6] , \nScanOut974[5] , \nScanOut974[4] , \nScanOut974[3] , 
        \nScanOut974[2] , \nScanOut974[1] , \nScanOut974[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_13[7] , \nOut30_13[6] , \nOut30_13[5] , \nOut30_13[4] , 
        \nOut30_13[3] , \nOut30_13[2] , \nOut30_13[1] , \nOut30_13[0] }), 
        .SouthIn({\nOut30_15[7] , \nOut30_15[6] , \nOut30_15[5] , 
        \nOut30_15[4] , \nOut30_15[3] , \nOut30_15[2] , \nOut30_15[1] , 
        \nOut30_15[0] }), .EastIn({\nOut31_14[7] , \nOut31_14[6] , 
        \nOut31_14[5] , \nOut31_14[4] , \nOut31_14[3] , \nOut31_14[2] , 
        \nOut31_14[1] , \nOut31_14[0] }), .WestIn({\nOut29_14[7] , 
        \nOut29_14[6] , \nOut29_14[5] , \nOut29_14[4] , \nOut29_14[3] , 
        \nOut29_14[2] , \nOut29_14[1] , \nOut29_14[0] }), .Out({\nOut30_14[7] , 
        \nOut30_14[6] , \nOut30_14[5] , \nOut30_14[4] , \nOut30_14[3] , 
        \nOut30_14[2] , \nOut30_14[1] , \nOut30_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_317 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut318[7] , \nScanOut318[6] , 
        \nScanOut318[5] , \nScanOut318[4] , \nScanOut318[3] , \nScanOut318[2] , 
        \nScanOut318[1] , \nScanOut318[0] }), .ScanOut({\nScanOut317[7] , 
        \nScanOut317[6] , \nScanOut317[5] , \nScanOut317[4] , \nScanOut317[3] , 
        \nScanOut317[2] , \nScanOut317[1] , \nScanOut317[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_28[7] , \nOut9_28[6] , \nOut9_28[5] , \nOut9_28[4] , 
        \nOut9_28[3] , \nOut9_28[2] , \nOut9_28[1] , \nOut9_28[0] }), 
        .SouthIn({\nOut9_30[7] , \nOut9_30[6] , \nOut9_30[5] , \nOut9_30[4] , 
        \nOut9_30[3] , \nOut9_30[2] , \nOut9_30[1] , \nOut9_30[0] }), .EastIn(
        {\nOut10_29[7] , \nOut10_29[6] , \nOut10_29[5] , \nOut10_29[4] , 
        \nOut10_29[3] , \nOut10_29[2] , \nOut10_29[1] , \nOut10_29[0] }), 
        .WestIn({\nOut8_29[7] , \nOut8_29[6] , \nOut8_29[5] , \nOut8_29[4] , 
        \nOut8_29[3] , \nOut8_29[2] , \nOut8_29[1] , \nOut8_29[0] }), .Out({
        \nOut9_29[7] , \nOut9_29[6] , \nOut9_29[5] , \nOut9_29[4] , 
        \nOut9_29[3] , \nOut9_29[2] , \nOut9_29[1] , \nOut9_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_496 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut497[7] , \nScanOut497[6] , 
        \nScanOut497[5] , \nScanOut497[4] , \nScanOut497[3] , \nScanOut497[2] , 
        \nScanOut497[1] , \nScanOut497[0] }), .ScanOut({\nScanOut496[7] , 
        \nScanOut496[6] , \nScanOut496[5] , \nScanOut496[4] , \nScanOut496[3] , 
        \nScanOut496[2] , \nScanOut496[1] , \nScanOut496[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_15[7] , \nOut15_15[6] , \nOut15_15[5] , \nOut15_15[4] , 
        \nOut15_15[3] , \nOut15_15[2] , \nOut15_15[1] , \nOut15_15[0] }), 
        .SouthIn({\nOut15_17[7] , \nOut15_17[6] , \nOut15_17[5] , 
        \nOut15_17[4] , \nOut15_17[3] , \nOut15_17[2] , \nOut15_17[1] , 
        \nOut15_17[0] }), .EastIn({\nOut16_16[7] , \nOut16_16[6] , 
        \nOut16_16[5] , \nOut16_16[4] , \nOut16_16[3] , \nOut16_16[2] , 
        \nOut16_16[1] , \nOut16_16[0] }), .WestIn({\nOut14_16[7] , 
        \nOut14_16[6] , \nOut14_16[5] , \nOut14_16[4] , \nOut14_16[3] , 
        \nOut14_16[2] , \nOut14_16[1] , \nOut14_16[0] }), .Out({\nOut15_16[7] , 
        \nOut15_16[6] , \nOut15_16[5] , \nOut15_16[4] , \nOut15_16[3] , 
        \nOut15_16[2] , \nOut15_16[1] , \nOut15_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_379 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut380[7] , \nScanOut380[6] , 
        \nScanOut380[5] , \nScanOut380[4] , \nScanOut380[3] , \nScanOut380[2] , 
        \nScanOut380[1] , \nScanOut380[0] }), .ScanOut({\nScanOut379[7] , 
        \nScanOut379[6] , \nScanOut379[5] , \nScanOut379[4] , \nScanOut379[3] , 
        \nScanOut379[2] , \nScanOut379[1] , \nScanOut379[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_26[7] , \nOut11_26[6] , \nOut11_26[5] , \nOut11_26[4] , 
        \nOut11_26[3] , \nOut11_26[2] , \nOut11_26[1] , \nOut11_26[0] }), 
        .SouthIn({\nOut11_28[7] , \nOut11_28[6] , \nOut11_28[5] , 
        \nOut11_28[4] , \nOut11_28[3] , \nOut11_28[2] , \nOut11_28[1] , 
        \nOut11_28[0] }), .EastIn({\nOut12_27[7] , \nOut12_27[6] , 
        \nOut12_27[5] , \nOut12_27[4] , \nOut12_27[3] , \nOut12_27[2] , 
        \nOut12_27[1] , \nOut12_27[0] }), .WestIn({\nOut10_27[7] , 
        \nOut10_27[6] , \nOut10_27[5] , \nOut10_27[4] , \nOut10_27[3] , 
        \nOut10_27[2] , \nOut10_27[1] , \nOut10_27[0] }), .Out({\nOut11_27[7] , 
        \nOut11_27[6] , \nOut11_27[5] , \nOut11_27[4] , \nOut11_27[3] , 
        \nOut11_27[2] , \nOut11_27[1] , \nOut11_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_658 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut659[7] , \nScanOut659[6] , 
        \nScanOut659[5] , \nScanOut659[4] , \nScanOut659[3] , \nScanOut659[2] , 
        \nScanOut659[1] , \nScanOut659[0] }), .ScanOut({\nScanOut658[7] , 
        \nScanOut658[6] , \nScanOut658[5] , \nScanOut658[4] , \nScanOut658[3] , 
        \nScanOut658[2] , \nScanOut658[1] , \nScanOut658[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_17[7] , \nOut20_17[6] , \nOut20_17[5] , \nOut20_17[4] , 
        \nOut20_17[3] , \nOut20_17[2] , \nOut20_17[1] , \nOut20_17[0] }), 
        .SouthIn({\nOut20_19[7] , \nOut20_19[6] , \nOut20_19[5] , 
        \nOut20_19[4] , \nOut20_19[3] , \nOut20_19[2] , \nOut20_19[1] , 
        \nOut20_19[0] }), .EastIn({\nOut21_18[7] , \nOut21_18[6] , 
        \nOut21_18[5] , \nOut21_18[4] , \nOut21_18[3] , \nOut21_18[2] , 
        \nOut21_18[1] , \nOut21_18[0] }), .WestIn({\nOut19_18[7] , 
        \nOut19_18[6] , \nOut19_18[5] , \nOut19_18[4] , \nOut19_18[3] , 
        \nOut19_18[2] , \nOut19_18[1] , \nOut19_18[0] }), .Out({\nOut20_18[7] , 
        \nOut20_18[6] , \nOut20_18[5] , \nOut20_18[4] , \nOut20_18[3] , 
        \nOut20_18[2] , \nOut20_18[1] , \nOut20_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_568 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut569[7] , \nScanOut569[6] , 
        \nScanOut569[5] , \nScanOut569[4] , \nScanOut569[3] , \nScanOut569[2] , 
        \nScanOut569[1] , \nScanOut569[0] }), .ScanOut({\nScanOut568[7] , 
        \nScanOut568[6] , \nScanOut568[5] , \nScanOut568[4] , \nScanOut568[3] , 
        \nScanOut568[2] , \nScanOut568[1] , \nScanOut568[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_23[7] , \nOut17_23[6] , \nOut17_23[5] , \nOut17_23[4] , 
        \nOut17_23[3] , \nOut17_23[2] , \nOut17_23[1] , \nOut17_23[0] }), 
        .SouthIn({\nOut17_25[7] , \nOut17_25[6] , \nOut17_25[5] , 
        \nOut17_25[4] , \nOut17_25[3] , \nOut17_25[2] , \nOut17_25[1] , 
        \nOut17_25[0] }), .EastIn({\nOut18_24[7] , \nOut18_24[6] , 
        \nOut18_24[5] , \nOut18_24[4] , \nOut18_24[3] , \nOut18_24[2] , 
        \nOut18_24[1] , \nOut18_24[0] }), .WestIn({\nOut16_24[7] , 
        \nOut16_24[6] , \nOut16_24[5] , \nOut16_24[4] , \nOut16_24[3] , 
        \nOut16_24[2] , \nOut16_24[1] , \nOut16_24[0] }), .Out({\nOut17_24[7] , 
        \nOut17_24[6] , \nOut17_24[5] , \nOut17_24[4] , \nOut17_24[3] , 
        \nOut17_24[2] , \nOut17_24[1] , \nOut17_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_743 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut744[7] , \nScanOut744[6] , 
        \nScanOut744[5] , \nScanOut744[4] , \nScanOut744[3] , \nScanOut744[2] , 
        \nScanOut744[1] , \nScanOut744[0] }), .ScanOut({\nScanOut743[7] , 
        \nScanOut743[6] , \nScanOut743[5] , \nScanOut743[4] , \nScanOut743[3] , 
        \nScanOut743[2] , \nScanOut743[1] , \nScanOut743[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_6[7] , \nOut23_6[6] , \nOut23_6[5] , \nOut23_6[4] , 
        \nOut23_6[3] , \nOut23_6[2] , \nOut23_6[1] , \nOut23_6[0] }), 
        .SouthIn({\nOut23_8[7] , \nOut23_8[6] , \nOut23_8[5] , \nOut23_8[4] , 
        \nOut23_8[3] , \nOut23_8[2] , \nOut23_8[1] , \nOut23_8[0] }), .EastIn(
        {\nOut24_7[7] , \nOut24_7[6] , \nOut24_7[5] , \nOut24_7[4] , 
        \nOut24_7[3] , \nOut24_7[2] , \nOut24_7[1] , \nOut24_7[0] }), .WestIn(
        {\nOut22_7[7] , \nOut22_7[6] , \nOut22_7[5] , \nOut22_7[4] , 
        \nOut22_7[3] , \nOut22_7[2] , \nOut22_7[1] , \nOut22_7[0] }), .Out({
        \nOut23_7[7] , \nOut23_7[6] , \nOut23_7[5] , \nOut23_7[4] , 
        \nOut23_7[3] , \nOut23_7[2] , \nOut23_7[1] , \nOut23_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_175 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut176[7] , \nScanOut176[6] , 
        \nScanOut176[5] , \nScanOut176[4] , \nScanOut176[3] , \nScanOut176[2] , 
        \nScanOut176[1] , \nScanOut176[0] }), .ScanOut({\nScanOut175[7] , 
        \nScanOut175[6] , \nScanOut175[5] , \nScanOut175[4] , \nScanOut175[3] , 
        \nScanOut175[2] , \nScanOut175[1] , \nScanOut175[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }), 
        .SouthIn({\nOut5_16[7] , \nOut5_16[6] , \nOut5_16[5] , \nOut5_16[4] , 
        \nOut5_16[3] , \nOut5_16[2] , \nOut5_16[1] , \nOut5_16[0] }), .EastIn(
        {\nOut6_15[7] , \nOut6_15[6] , \nOut6_15[5] , \nOut6_15[4] , 
        \nOut6_15[3] , \nOut6_15[2] , \nOut6_15[1] , \nOut6_15[0] }), .WestIn(
        {\nOut4_15[7] , \nOut4_15[6] , \nOut4_15[5] , \nOut4_15[4] , 
        \nOut4_15[3] , \nOut4_15[2] , \nOut4_15[1] , \nOut4_15[0] }), .Out({
        \nOut5_15[7] , \nOut5_15[6] , \nOut5_15[5] , \nOut5_15[4] , 
        \nOut5_15[3] , \nOut5_15[2] , \nOut5_15[1] , \nOut5_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_245 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut246[7] , \nScanOut246[6] , 
        \nScanOut246[5] , \nScanOut246[4] , \nScanOut246[3] , \nScanOut246[2] , 
        \nScanOut246[1] , \nScanOut246[0] }), .ScanOut({\nScanOut245[7] , 
        \nScanOut245[6] , \nScanOut245[5] , \nScanOut245[4] , \nScanOut245[3] , 
        \nScanOut245[2] , \nScanOut245[1] , \nScanOut245[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_20[7] , \nOut7_20[6] , \nOut7_20[5] , \nOut7_20[4] , 
        \nOut7_20[3] , \nOut7_20[2] , \nOut7_20[1] , \nOut7_20[0] }), 
        .SouthIn({\nOut7_22[7] , \nOut7_22[6] , \nOut7_22[5] , \nOut7_22[4] , 
        \nOut7_22[3] , \nOut7_22[2] , \nOut7_22[1] , \nOut7_22[0] }), .EastIn(
        {\nOut8_21[7] , \nOut8_21[6] , \nOut8_21[5] , \nOut8_21[4] , 
        \nOut8_21[3] , \nOut8_21[2] , \nOut8_21[1] , \nOut8_21[0] }), .WestIn(
        {\nOut6_21[7] , \nOut6_21[6] , \nOut6_21[5] , \nOut6_21[4] , 
        \nOut6_21[3] , \nOut6_21[2] , \nOut6_21[1] , \nOut6_21[0] }), .Out({
        \nOut7_21[7] , \nOut7_21[6] , \nOut7_21[5] , \nOut7_21[4] , 
        \nOut7_21[3] , \nOut7_21[2] , \nOut7_21[1] , \nOut7_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_262 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut263[7] , \nScanOut263[6] , 
        \nScanOut263[5] , \nScanOut263[4] , \nScanOut263[3] , \nScanOut263[2] , 
        \nScanOut263[1] , \nScanOut263[0] }), .ScanOut({\nScanOut262[7] , 
        \nScanOut262[6] , \nScanOut262[5] , \nScanOut262[4] , \nScanOut262[3] , 
        \nScanOut262[2] , \nScanOut262[1] , \nScanOut262[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_5[7] , \nOut8_5[6] , \nOut8_5[5] , \nOut8_5[4] , \nOut8_5[3] , 
        \nOut8_5[2] , \nOut8_5[1] , \nOut8_5[0] }), .SouthIn({\nOut8_7[7] , 
        \nOut8_7[6] , \nOut8_7[5] , \nOut8_7[4] , \nOut8_7[3] , \nOut8_7[2] , 
        \nOut8_7[1] , \nOut8_7[0] }), .EastIn({\nOut9_6[7] , \nOut9_6[6] , 
        \nOut9_6[5] , \nOut9_6[4] , \nOut9_6[3] , \nOut9_6[2] , \nOut9_6[1] , 
        \nOut9_6[0] }), .WestIn({\nOut7_6[7] , \nOut7_6[6] , \nOut7_6[5] , 
        \nOut7_6[4] , \nOut7_6[3] , \nOut7_6[2] , \nOut7_6[1] , \nOut7_6[0] }), 
        .Out({\nOut8_6[7] , \nOut8_6[6] , \nOut8_6[5] , \nOut8_6[4] , 
        \nOut8_6[3] , \nOut8_6[2] , \nOut8_6[1] , \nOut8_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_473 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut474[7] , \nScanOut474[6] , 
        \nScanOut474[5] , \nScanOut474[4] , \nScanOut474[3] , \nScanOut474[2] , 
        \nScanOut474[1] , \nScanOut474[0] }), .ScanOut({\nScanOut473[7] , 
        \nScanOut473[6] , \nScanOut473[5] , \nScanOut473[4] , \nScanOut473[3] , 
        \nScanOut473[2] , \nScanOut473[1] , \nScanOut473[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_24[7] , \nOut14_24[6] , \nOut14_24[5] , \nOut14_24[4] , 
        \nOut14_24[3] , \nOut14_24[2] , \nOut14_24[1] , \nOut14_24[0] }), 
        .SouthIn({\nOut14_26[7] , \nOut14_26[6] , \nOut14_26[5] , 
        \nOut14_26[4] , \nOut14_26[3] , \nOut14_26[2] , \nOut14_26[1] , 
        \nOut14_26[0] }), .EastIn({\nOut15_25[7] , \nOut15_25[6] , 
        \nOut15_25[5] , \nOut15_25[4] , \nOut15_25[3] , \nOut15_25[2] , 
        \nOut15_25[1] , \nOut15_25[0] }), .WestIn({\nOut13_25[7] , 
        \nOut13_25[6] , \nOut13_25[5] , \nOut13_25[4] , \nOut13_25[3] , 
        \nOut13_25[2] , \nOut13_25[1] , \nOut13_25[0] }), .Out({\nOut14_25[7] , 
        \nOut14_25[6] , \nOut14_25[5] , \nOut14_25[4] , \nOut14_25[3] , 
        \nOut14_25[2] , \nOut14_25[1] , \nOut14_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_801 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut802[7] , \nScanOut802[6] , 
        \nScanOut802[5] , \nScanOut802[4] , \nScanOut802[3] , \nScanOut802[2] , 
        \nScanOut802[1] , \nScanOut802[0] }), .ScanOut({\nScanOut801[7] , 
        \nScanOut801[6] , \nScanOut801[5] , \nScanOut801[4] , \nScanOut801[3] , 
        \nScanOut801[2] , \nScanOut801[1] , \nScanOut801[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_0[7] , \nOut25_0[6] , \nOut25_0[5] , \nOut25_0[4] , 
        \nOut25_0[3] , \nOut25_0[2] , \nOut25_0[1] , \nOut25_0[0] }), 
        .SouthIn({\nOut25_2[7] , \nOut25_2[6] , \nOut25_2[5] , \nOut25_2[4] , 
        \nOut25_2[3] , \nOut25_2[2] , \nOut25_2[1] , \nOut25_2[0] }), .EastIn(
        {\nOut26_1[7] , \nOut26_1[6] , \nOut26_1[5] , \nOut26_1[4] , 
        \nOut26_1[3] , \nOut26_1[2] , \nOut26_1[1] , \nOut26_1[0] }), .WestIn(
        {\nOut24_1[7] , \nOut24_1[6] , \nOut24_1[5] , \nOut24_1[4] , 
        \nOut24_1[3] , \nOut24_1[2] , \nOut24_1[1] , \nOut24_1[0] }), .Out({
        \nOut25_1[7] , \nOut25_1[6] , \nOut25_1[5] , \nOut25_1[4] , 
        \nOut25_1[3] , \nOut25_1[2] , \nOut25_1[1] , \nOut25_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_991 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut992[7] , \nScanOut992[6] , 
        \nScanOut992[5] , \nScanOut992[4] , \nScanOut992[3] , \nScanOut992[2] , 
        \nScanOut992[1] , \nScanOut992[0] }), .ScanOut({\nScanOut991[7] , 
        \nScanOut991[6] , \nScanOut991[5] , \nScanOut991[4] , \nScanOut991[3] , 
        \nScanOut991[2] , \nScanOut991[1] , \nScanOut991[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut30_31[7] , \nOut30_31[6] , 
        \nOut30_31[5] , \nOut30_31[4] , \nOut30_31[3] , \nOut30_31[2] , 
        \nOut30_31[1] , \nOut30_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_826 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut827[7] , \nScanOut827[6] , 
        \nScanOut827[5] , \nScanOut827[4] , \nScanOut827[3] , \nScanOut827[2] , 
        \nScanOut827[1] , \nScanOut827[0] }), .ScanOut({\nScanOut826[7] , 
        \nScanOut826[6] , \nScanOut826[5] , \nScanOut826[4] , \nScanOut826[3] , 
        \nScanOut826[2] , \nScanOut826[1] , \nScanOut826[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_25[7] , \nOut25_25[6] , \nOut25_25[5] , \nOut25_25[4] , 
        \nOut25_25[3] , \nOut25_25[2] , \nOut25_25[1] , \nOut25_25[0] }), 
        .SouthIn({\nOut25_27[7] , \nOut25_27[6] , \nOut25_27[5] , 
        \nOut25_27[4] , \nOut25_27[3] , \nOut25_27[2] , \nOut25_27[1] , 
        \nOut25_27[0] }), .EastIn({\nOut26_26[7] , \nOut26_26[6] , 
        \nOut26_26[5] , \nOut26_26[4] , \nOut26_26[3] , \nOut26_26[2] , 
        \nOut26_26[1] , \nOut26_26[0] }), .WestIn({\nOut24_26[7] , 
        \nOut24_26[6] , \nOut24_26[5] , \nOut24_26[4] , \nOut24_26[3] , 
        \nOut24_26[2] , \nOut24_26[1] , \nOut24_26[0] }), .Out({\nOut25_26[7] , 
        \nOut25_26[6] , \nOut25_26[5] , \nOut25_26[4] , \nOut25_26[3] , 
        \nOut25_26[2] , \nOut25_26[1] , \nOut25_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_454 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut455[7] , \nScanOut455[6] , 
        \nScanOut455[5] , \nScanOut455[4] , \nScanOut455[3] , \nScanOut455[2] , 
        \nScanOut455[1] , \nScanOut455[0] }), .ScanOut({\nScanOut454[7] , 
        \nScanOut454[6] , \nScanOut454[5] , \nScanOut454[4] , \nScanOut454[3] , 
        \nScanOut454[2] , \nScanOut454[1] , \nScanOut454[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }), 
        .SouthIn({\nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }), .EastIn(
        {\nOut15_6[7] , \nOut15_6[6] , \nOut15_6[5] , \nOut15_6[4] , 
        \nOut15_6[3] , \nOut15_6[2] , \nOut15_6[1] , \nOut15_6[0] }), .WestIn(
        {\nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }), .Out({
        \nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_279 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut280[7] , \nScanOut280[6] , 
        \nScanOut280[5] , \nScanOut280[4] , \nScanOut280[3] , \nScanOut280[2] , 
        \nScanOut280[1] , \nScanOut280[0] }), .ScanOut({\nScanOut279[7] , 
        \nScanOut279[6] , \nScanOut279[5] , \nScanOut279[4] , \nScanOut279[3] , 
        \nScanOut279[2] , \nScanOut279[1] , \nScanOut279[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_22[7] , \nOut8_22[6] , \nOut8_22[5] , \nOut8_22[4] , 
        \nOut8_22[3] , \nOut8_22[2] , \nOut8_22[1] , \nOut8_22[0] }), 
        .SouthIn({\nOut8_24[7] , \nOut8_24[6] , \nOut8_24[5] , \nOut8_24[4] , 
        \nOut8_24[3] , \nOut8_24[2] , \nOut8_24[1] , \nOut8_24[0] }), .EastIn(
        {\nOut9_23[7] , \nOut9_23[6] , \nOut9_23[5] , \nOut9_23[4] , 
        \nOut9_23[3] , \nOut9_23[2] , \nOut9_23[1] , \nOut9_23[0] }), .WestIn(
        {\nOut7_23[7] , \nOut7_23[6] , \nOut7_23[5] , \nOut7_23[4] , 
        \nOut7_23[3] , \nOut7_23[2] , \nOut7_23[1] , \nOut7_23[0] }), .Out({
        \nOut8_23[7] , \nOut8_23[6] , \nOut8_23[5] , \nOut8_23[4] , 
        \nOut8_23[3] , \nOut8_23[2] , \nOut8_23[1] , \nOut8_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_468 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut469[7] , \nScanOut469[6] , 
        \nScanOut469[5] , \nScanOut469[4] , \nScanOut469[3] , \nScanOut469[2] , 
        \nScanOut469[1] , \nScanOut469[0] }), .ScanOut({\nScanOut468[7] , 
        \nScanOut468[6] , \nScanOut468[5] , \nScanOut468[4] , \nScanOut468[3] , 
        \nScanOut468[2] , \nScanOut468[1] , \nScanOut468[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_19[7] , \nOut14_19[6] , \nOut14_19[5] , \nOut14_19[4] , 
        \nOut14_19[3] , \nOut14_19[2] , \nOut14_19[1] , \nOut14_19[0] }), 
        .SouthIn({\nOut14_21[7] , \nOut14_21[6] , \nOut14_21[5] , 
        \nOut14_21[4] , \nOut14_21[3] , \nOut14_21[2] , \nOut14_21[1] , 
        \nOut14_21[0] }), .EastIn({\nOut15_20[7] , \nOut15_20[6] , 
        \nOut15_20[5] , \nOut15_20[4] , \nOut15_20[3] , \nOut15_20[2] , 
        \nOut15_20[1] , \nOut15_20[0] }), .WestIn({\nOut13_20[7] , 
        \nOut13_20[6] , \nOut13_20[5] , \nOut13_20[4] , \nOut13_20[3] , 
        \nOut13_20[2] , \nOut13_20[1] , \nOut13_20[0] }), .Out({\nOut14_20[7] , 
        \nOut14_20[6] , \nOut14_20[5] , \nOut14_20[4] , \nOut14_20[3] , 
        \nOut14_20[2] , \nOut14_20[1] , \nOut14_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_764 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut765[7] , \nScanOut765[6] , 
        \nScanOut765[5] , \nScanOut765[4] , \nScanOut765[3] , \nScanOut765[2] , 
        \nScanOut765[1] , \nScanOut765[0] }), .ScanOut({\nScanOut764[7] , 
        \nScanOut764[6] , \nScanOut764[5] , \nScanOut764[4] , \nScanOut764[3] , 
        \nScanOut764[2] , \nScanOut764[1] , \nScanOut764[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_27[7] , \nOut23_27[6] , \nOut23_27[5] , \nOut23_27[4] , 
        \nOut23_27[3] , \nOut23_27[2] , \nOut23_27[1] , \nOut23_27[0] }), 
        .SouthIn({\nOut23_29[7] , \nOut23_29[6] , \nOut23_29[5] , 
        \nOut23_29[4] , \nOut23_29[3] , \nOut23_29[2] , \nOut23_29[1] , 
        \nOut23_29[0] }), .EastIn({\nOut24_28[7] , \nOut24_28[6] , 
        \nOut24_28[5] , \nOut24_28[4] , \nOut24_28[3] , \nOut24_28[2] , 
        \nOut24_28[1] , \nOut24_28[0] }), .WestIn({\nOut22_28[7] , 
        \nOut22_28[6] , \nOut22_28[5] , \nOut22_28[4] , \nOut22_28[3] , 
        \nOut22_28[2] , \nOut22_28[1] , \nOut22_28[0] }), .Out({\nOut23_28[7] , 
        \nOut23_28[6] , \nOut23_28[5] , \nOut23_28[4] , \nOut23_28[3] , 
        \nOut23_28[2] , \nOut23_28[1] , \nOut23_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_758 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut759[7] , \nScanOut759[6] , 
        \nScanOut759[5] , \nScanOut759[4] , \nScanOut759[3] , \nScanOut759[2] , 
        \nScanOut759[1] , \nScanOut759[0] }), .ScanOut({\nScanOut758[7] , 
        \nScanOut758[6] , \nScanOut758[5] , \nScanOut758[4] , \nScanOut758[3] , 
        \nScanOut758[2] , \nScanOut758[1] , \nScanOut758[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_21[7] , \nOut23_21[6] , \nOut23_21[5] , \nOut23_21[4] , 
        \nOut23_21[3] , \nOut23_21[2] , \nOut23_21[1] , \nOut23_21[0] }), 
        .SouthIn({\nOut23_23[7] , \nOut23_23[6] , \nOut23_23[5] , 
        \nOut23_23[4] , \nOut23_23[3] , \nOut23_23[2] , \nOut23_23[1] , 
        \nOut23_23[0] }), .EastIn({\nOut24_22[7] , \nOut24_22[6] , 
        \nOut24_22[5] , \nOut24_22[4] , \nOut24_22[3] , \nOut24_22[2] , 
        \nOut24_22[1] , \nOut24_22[0] }), .WestIn({\nOut22_22[7] , 
        \nOut22_22[6] , \nOut22_22[5] , \nOut22_22[4] , \nOut22_22[3] , 
        \nOut22_22[2] , \nOut22_22[1] , \nOut22_22[0] }), .Out({\nOut23_22[7] , 
        \nOut23_22[6] , \nOut23_22[5] , \nOut23_22[4] , \nOut23_22[3] , 
        \nOut23_22[2] , \nOut23_22[1] , \nOut23_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_664 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut665[7] , \nScanOut665[6] , 
        \nScanOut665[5] , \nScanOut665[4] , \nScanOut665[3] , \nScanOut665[2] , 
        \nScanOut665[1] , \nScanOut665[0] }), .ScanOut({\nScanOut664[7] , 
        \nScanOut664[6] , \nScanOut664[5] , \nScanOut664[4] , \nScanOut664[3] , 
        \nScanOut664[2] , \nScanOut664[1] , \nScanOut664[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_23[7] , \nOut20_23[6] , \nOut20_23[5] , \nOut20_23[4] , 
        \nOut20_23[3] , \nOut20_23[2] , \nOut20_23[1] , \nOut20_23[0] }), 
        .SouthIn({\nOut20_25[7] , \nOut20_25[6] , \nOut20_25[5] , 
        \nOut20_25[4] , \nOut20_25[3] , \nOut20_25[2] , \nOut20_25[1] , 
        \nOut20_25[0] }), .EastIn({\nOut21_24[7] , \nOut21_24[6] , 
        \nOut21_24[5] , \nOut21_24[4] , \nOut21_24[3] , \nOut21_24[2] , 
        \nOut21_24[1] , \nOut21_24[0] }), .WestIn({\nOut19_24[7] , 
        \nOut19_24[6] , \nOut19_24[5] , \nOut19_24[4] , \nOut19_24[3] , 
        \nOut19_24[2] , \nOut19_24[1] , \nOut19_24[0] }), .Out({\nOut20_24[7] , 
        \nOut20_24[6] , \nOut20_24[5] , \nOut20_24[4] , \nOut20_24[3] , 
        \nOut20_24[2] , \nOut20_24[1] , \nOut20_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_345 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut346[7] , \nScanOut346[6] , 
        \nScanOut346[5] , \nScanOut346[4] , \nScanOut346[3] , \nScanOut346[2] , 
        \nScanOut346[1] , \nScanOut346[0] }), .ScanOut({\nScanOut345[7] , 
        \nScanOut345[6] , \nScanOut345[5] , \nScanOut345[4] , \nScanOut345[3] , 
        \nScanOut345[2] , \nScanOut345[1] , \nScanOut345[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_24[7] , \nOut10_24[6] , \nOut10_24[5] , \nOut10_24[4] , 
        \nOut10_24[3] , \nOut10_24[2] , \nOut10_24[1] , \nOut10_24[0] }), 
        .SouthIn({\nOut10_26[7] , \nOut10_26[6] , \nOut10_26[5] , 
        \nOut10_26[4] , \nOut10_26[3] , \nOut10_26[2] , \nOut10_26[1] , 
        \nOut10_26[0] }), .EastIn({\nOut11_25[7] , \nOut11_25[6] , 
        \nOut11_25[5] , \nOut11_25[4] , \nOut11_25[3] , \nOut11_25[2] , 
        \nOut11_25[1] , \nOut11_25[0] }), .WestIn({\nOut9_25[7] , 
        \nOut9_25[6] , \nOut9_25[5] , \nOut9_25[4] , \nOut9_25[3] , 
        \nOut9_25[2] , \nOut9_25[1] , \nOut9_25[0] }), .Out({\nOut10_25[7] , 
        \nOut10_25[6] , \nOut10_25[5] , \nOut10_25[4] , \nOut10_25[3] , 
        \nOut10_25[2] , \nOut10_25[1] , \nOut10_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_554 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut555[7] , \nScanOut555[6] , 
        \nScanOut555[5] , \nScanOut555[4] , \nScanOut555[3] , \nScanOut555[2] , 
        \nScanOut555[1] , \nScanOut555[0] }), .ScanOut({\nScanOut554[7] , 
        \nScanOut554[6] , \nScanOut554[5] , \nScanOut554[4] , \nScanOut554[3] , 
        \nScanOut554[2] , \nScanOut554[1] , \nScanOut554[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_9[7] , \nOut17_9[6] , \nOut17_9[5] , \nOut17_9[4] , 
        \nOut17_9[3] , \nOut17_9[2] , \nOut17_9[1] , \nOut17_9[0] }), 
        .SouthIn({\nOut17_11[7] , \nOut17_11[6] , \nOut17_11[5] , 
        \nOut17_11[4] , \nOut17_11[3] , \nOut17_11[2] , \nOut17_11[1] , 
        \nOut17_11[0] }), .EastIn({\nOut18_10[7] , \nOut18_10[6] , 
        \nOut18_10[5] , \nOut18_10[4] , \nOut18_10[3] , \nOut18_10[2] , 
        \nOut18_10[1] , \nOut18_10[0] }), .WestIn({\nOut16_10[7] , 
        \nOut16_10[6] , \nOut16_10[5] , \nOut16_10[4] , \nOut16_10[3] , 
        \nOut16_10[2] , \nOut16_10[1] , \nOut16_10[0] }), .Out({\nOut17_10[7] , 
        \nOut17_10[6] , \nOut17_10[5] , \nOut17_10[4] , \nOut17_10[3] , 
        \nOut17_10[2] , \nOut17_10[1] , \nOut17_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_926 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut927[7] , \nScanOut927[6] , 
        \nScanOut927[5] , \nScanOut927[4] , \nScanOut927[3] , \nScanOut927[2] , 
        \nScanOut927[1] , \nScanOut927[0] }), .ScanOut({\nScanOut926[7] , 
        \nScanOut926[6] , \nScanOut926[5] , \nScanOut926[4] , \nScanOut926[3] , 
        \nScanOut926[2] , \nScanOut926[1] , \nScanOut926[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_29[7] , \nOut28_29[6] , \nOut28_29[5] , \nOut28_29[4] , 
        \nOut28_29[3] , \nOut28_29[2] , \nOut28_29[1] , \nOut28_29[0] }), 
        .SouthIn({\nOut28_31[7] , \nOut28_31[6] , \nOut28_31[5] , 
        \nOut28_31[4] , \nOut28_31[3] , \nOut28_31[2] , \nOut28_31[1] , 
        \nOut28_31[0] }), .EastIn({\nOut29_30[7] , \nOut29_30[6] , 
        \nOut29_30[5] , \nOut29_30[4] , \nOut29_30[3] , \nOut29_30[2] , 
        \nOut29_30[1] , \nOut29_30[0] }), .WestIn({\nOut27_30[7] , 
        \nOut27_30[6] , \nOut27_30[5] , \nOut27_30[4] , \nOut27_30[3] , 
        \nOut27_30[2] , \nOut27_30[1] , \nOut27_30[0] }), .Out({\nOut28_30[7] , 
        \nOut28_30[6] , \nOut28_30[5] , \nOut28_30[4] , \nOut28_30[3] , 
        \nOut28_30[2] , \nOut28_30[1] , \nOut28_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_362 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut363[7] , \nScanOut363[6] , 
        \nScanOut363[5] , \nScanOut363[4] , \nScanOut363[3] , \nScanOut363[2] , 
        \nScanOut363[1] , \nScanOut363[0] }), .ScanOut({\nScanOut362[7] , 
        \nScanOut362[6] , \nScanOut362[5] , \nScanOut362[4] , \nScanOut362[3] , 
        \nScanOut362[2] , \nScanOut362[1] , \nScanOut362[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , \nOut11_9[4] , 
        \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , \nOut11_9[0] }), 
        .SouthIn({\nOut11_11[7] , \nOut11_11[6] , \nOut11_11[5] , 
        \nOut11_11[4] , \nOut11_11[3] , \nOut11_11[2] , \nOut11_11[1] , 
        \nOut11_11[0] }), .EastIn({\nOut12_10[7] , \nOut12_10[6] , 
        \nOut12_10[5] , \nOut12_10[4] , \nOut12_10[3] , \nOut12_10[2] , 
        \nOut12_10[1] , \nOut12_10[0] }), .WestIn({\nOut10_10[7] , 
        \nOut10_10[6] , \nOut10_10[5] , \nOut10_10[4] , \nOut10_10[3] , 
        \nOut10_10[2] , \nOut10_10[1] , \nOut10_10[0] }), .Out({\nOut11_10[7] , 
        \nOut11_10[6] , \nOut11_10[5] , \nOut11_10[4] , \nOut11_10[3] , 
        \nOut11_10[2] , \nOut11_10[1] , \nOut11_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_891 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut892[7] , \nScanOut892[6] , 
        \nScanOut892[5] , \nScanOut892[4] , \nScanOut892[3] , \nScanOut892[2] , 
        \nScanOut892[1] , \nScanOut892[0] }), .ScanOut({\nScanOut891[7] , 
        \nScanOut891[6] , \nScanOut891[5] , \nScanOut891[4] , \nScanOut891[3] , 
        \nScanOut891[2] , \nScanOut891[1] , \nScanOut891[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_26[7] , \nOut27_26[6] , \nOut27_26[5] , \nOut27_26[4] , 
        \nOut27_26[3] , \nOut27_26[2] , \nOut27_26[1] , \nOut27_26[0] }), 
        .SouthIn({\nOut27_28[7] , \nOut27_28[6] , \nOut27_28[5] , 
        \nOut27_28[4] , \nOut27_28[3] , \nOut27_28[2] , \nOut27_28[1] , 
        \nOut27_28[0] }), .EastIn({\nOut28_27[7] , \nOut28_27[6] , 
        \nOut28_27[5] , \nOut28_27[4] , \nOut28_27[3] , \nOut28_27[2] , 
        \nOut28_27[1] , \nOut28_27[0] }), .WestIn({\nOut26_27[7] , 
        \nOut26_27[6] , \nOut26_27[5] , \nOut26_27[4] , \nOut26_27[3] , 
        \nOut26_27[2] , \nOut26_27[1] , \nOut26_27[0] }), .Out({\nOut27_27[7] , 
        \nOut27_27[6] , \nOut27_27[5] , \nOut27_27[4] , \nOut27_27[3] , 
        \nOut27_27[2] , \nOut27_27[1] , \nOut27_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_901 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut902[7] , \nScanOut902[6] , 
        \nScanOut902[5] , \nScanOut902[4] , \nScanOut902[3] , \nScanOut902[2] , 
        \nScanOut902[1] , \nScanOut902[0] }), .ScanOut({\nScanOut901[7] , 
        \nScanOut901[6] , \nScanOut901[5] , \nScanOut901[4] , \nScanOut901[3] , 
        \nScanOut901[2] , \nScanOut901[1] , \nScanOut901[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_4[7] , \nOut28_4[6] , \nOut28_4[5] , \nOut28_4[4] , 
        \nOut28_4[3] , \nOut28_4[2] , \nOut28_4[1] , \nOut28_4[0] }), 
        .SouthIn({\nOut28_6[7] , \nOut28_6[6] , \nOut28_6[5] , \nOut28_6[4] , 
        \nOut28_6[3] , \nOut28_6[2] , \nOut28_6[1] , \nOut28_6[0] }), .EastIn(
        {\nOut29_5[7] , \nOut29_5[6] , \nOut29_5[5] , \nOut29_5[4] , 
        \nOut29_5[3] , \nOut29_5[2] , \nOut29_5[1] , \nOut29_5[0] }), .WestIn(
        {\nOut27_5[7] , \nOut27_5[6] , \nOut27_5[5] , \nOut27_5[4] , 
        \nOut27_5[3] , \nOut27_5[2] , \nOut27_5[1] , \nOut27_5[0] }), .Out({
        \nOut28_5[7] , \nOut28_5[6] , \nOut28_5[5] , \nOut28_5[4] , 
        \nOut28_5[3] , \nOut28_5[2] , \nOut28_5[1] , \nOut28_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_573 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut574[7] , \nScanOut574[6] , 
        \nScanOut574[5] , \nScanOut574[4] , \nScanOut574[3] , \nScanOut574[2] , 
        \nScanOut574[1] , \nScanOut574[0] }), .ScanOut({\nScanOut573[7] , 
        \nScanOut573[6] , \nScanOut573[5] , \nScanOut573[4] , \nScanOut573[3] , 
        \nScanOut573[2] , \nScanOut573[1] , \nScanOut573[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_28[7] , \nOut17_28[6] , \nOut17_28[5] , \nOut17_28[4] , 
        \nOut17_28[3] , \nOut17_28[2] , \nOut17_28[1] , \nOut17_28[0] }), 
        .SouthIn({\nOut17_30[7] , \nOut17_30[6] , \nOut17_30[5] , 
        \nOut17_30[4] , \nOut17_30[3] , \nOut17_30[2] , \nOut17_30[1] , 
        \nOut17_30[0] }), .EastIn({\nOut18_29[7] , \nOut18_29[6] , 
        \nOut18_29[5] , \nOut18_29[4] , \nOut18_29[3] , \nOut18_29[2] , 
        \nOut18_29[1] , \nOut18_29[0] }), .WestIn({\nOut16_29[7] , 
        \nOut16_29[6] , \nOut16_29[5] , \nOut16_29[4] , \nOut16_29[3] , 
        \nOut16_29[2] , \nOut16_29[1] , \nOut16_29[0] }), .Out({\nOut17_29[7] , 
        \nOut17_29[6] , \nOut17_29[5] , \nOut17_29[4] , \nOut17_29[3] , 
        \nOut17_29[2] , \nOut17_29[1] , \nOut17_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_643 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut644[7] , \nScanOut644[6] , 
        \nScanOut644[5] , \nScanOut644[4] , \nScanOut644[3] , \nScanOut644[2] , 
        \nScanOut644[1] , \nScanOut644[0] }), .ScanOut({\nScanOut643[7] , 
        \nScanOut643[6] , \nScanOut643[5] , \nScanOut643[4] , \nScanOut643[3] , 
        \nScanOut643[2] , \nScanOut643[1] , \nScanOut643[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_2[7] , \nOut20_2[6] , \nOut20_2[5] , \nOut20_2[4] , 
        \nOut20_2[3] , \nOut20_2[2] , \nOut20_2[1] , \nOut20_2[0] }), 
        .SouthIn({\nOut20_4[7] , \nOut20_4[6] , \nOut20_4[5] , \nOut20_4[4] , 
        \nOut20_4[3] , \nOut20_4[2] , \nOut20_4[1] , \nOut20_4[0] }), .EastIn(
        {\nOut21_3[7] , \nOut21_3[6] , \nOut21_3[5] , \nOut21_3[4] , 
        \nOut21_3[3] , \nOut21_3[2] , \nOut21_3[1] , \nOut21_3[0] }), .WestIn(
        {\nOut19_3[7] , \nOut19_3[6] , \nOut19_3[5] , \nOut19_3[4] , 
        \nOut19_3[3] , \nOut19_3[2] , \nOut19_3[1] , \nOut19_3[0] }), .Out({
        \nOut20_3[7] , \nOut20_3[6] , \nOut20_3[5] , \nOut20_3[4] , 
        \nOut20_3[3] , \nOut20_3[2] , \nOut20_3[1] , \nOut20_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_94 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut95[7] , \nScanOut95[6] , 
        \nScanOut95[5] , \nScanOut95[4] , \nScanOut95[3] , \nScanOut95[2] , 
        \nScanOut95[1] , \nScanOut95[0] }), .ScanOut({\nScanOut94[7] , 
        \nScanOut94[6] , \nScanOut94[5] , \nScanOut94[4] , \nScanOut94[3] , 
        \nScanOut94[2] , \nScanOut94[1] , \nScanOut94[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_29[7] , \nOut2_29[6] , \nOut2_29[5] , \nOut2_29[4] , 
        \nOut2_29[3] , \nOut2_29[2] , \nOut2_29[1] , \nOut2_29[0] }), 
        .SouthIn({\nOut2_31[7] , \nOut2_31[6] , \nOut2_31[5] , \nOut2_31[4] , 
        \nOut2_31[3] , \nOut2_31[2] , \nOut2_31[1] , \nOut2_31[0] }), .EastIn(
        {\nOut3_30[7] , \nOut3_30[6] , \nOut3_30[5] , \nOut3_30[4] , 
        \nOut3_30[3] , \nOut3_30[2] , \nOut3_30[1] , \nOut3_30[0] }), .WestIn(
        {\nOut1_30[7] , \nOut1_30[6] , \nOut1_30[5] , \nOut1_30[4] , 
        \nOut1_30[3] , \nOut1_30[2] , \nOut1_30[1] , \nOut1_30[0] }), .Out({
        \nOut2_30[7] , \nOut2_30[6] , \nOut2_30[5] , \nOut2_30[4] , 
        \nOut2_30[3] , \nOut2_30[2] , \nOut2_30[1] , \nOut2_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_127 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut128[7] , \nScanOut128[6] , 
        \nScanOut128[5] , \nScanOut128[4] , \nScanOut128[3] , \nScanOut128[2] , 
        \nScanOut128[1] , \nScanOut128[0] }), .ScanOut({\nScanOut127[7] , 
        \nScanOut127[6] , \nScanOut127[5] , \nScanOut127[4] , \nScanOut127[3] , 
        \nScanOut127[2] , \nScanOut127[1] , \nScanOut127[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut3_31[7] , \nOut3_31[6] , 
        \nOut3_31[5] , \nOut3_31[4] , \nOut3_31[3] , \nOut3_31[2] , 
        \nOut3_31[1] , \nOut3_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_217 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut218[7] , \nScanOut218[6] , 
        \nScanOut218[5] , \nScanOut218[4] , \nScanOut218[3] , \nScanOut218[2] , 
        \nScanOut218[1] , \nScanOut218[0] }), .ScanOut({\nScanOut217[7] , 
        \nScanOut217[6] , \nScanOut217[5] , \nScanOut217[4] , \nScanOut217[3] , 
        \nScanOut217[2] , \nScanOut217[1] , \nScanOut217[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_24[7] , \nOut6_24[6] , \nOut6_24[5] , \nOut6_24[4] , 
        \nOut6_24[3] , \nOut6_24[2] , \nOut6_24[1] , \nOut6_24[0] }), 
        .SouthIn({\nOut6_26[7] , \nOut6_26[6] , \nOut6_26[5] , \nOut6_26[4] , 
        \nOut6_26[3] , \nOut6_26[2] , \nOut6_26[1] , \nOut6_26[0] }), .EastIn(
        {\nOut7_25[7] , \nOut7_25[6] , \nOut7_25[5] , \nOut7_25[4] , 
        \nOut7_25[3] , \nOut7_25[2] , \nOut7_25[1] , \nOut7_25[0] }), .WestIn(
        {\nOut5_25[7] , \nOut5_25[6] , \nOut5_25[5] , \nOut5_25[4] , 
        \nOut5_25[3] , \nOut5_25[2] , \nOut5_25[1] , \nOut5_25[0] }), .Out({
        \nOut6_25[7] , \nOut6_25[6] , \nOut6_25[5] , \nOut6_25[4] , 
        \nOut6_25[3] , \nOut6_25[2] , \nOut6_25[1] , \nOut6_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_596 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut597[7] , \nScanOut597[6] , 
        \nScanOut597[5] , \nScanOut597[4] , \nScanOut597[3] , \nScanOut597[2] , 
        \nScanOut597[1] , \nScanOut597[0] }), .ScanOut({\nScanOut596[7] , 
        \nScanOut596[6] , \nScanOut596[5] , \nScanOut596[4] , \nScanOut596[3] , 
        \nScanOut596[2] , \nScanOut596[1] , \nScanOut596[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_19[7] , \nOut18_19[6] , \nOut18_19[5] , \nOut18_19[4] , 
        \nOut18_19[3] , \nOut18_19[2] , \nOut18_19[1] , \nOut18_19[0] }), 
        .SouthIn({\nOut18_21[7] , \nOut18_21[6] , \nOut18_21[5] , 
        \nOut18_21[4] , \nOut18_21[3] , \nOut18_21[2] , \nOut18_21[1] , 
        \nOut18_21[0] }), .EastIn({\nOut19_20[7] , \nOut19_20[6] , 
        \nOut19_20[5] , \nOut19_20[4] , \nOut19_20[3] , \nOut19_20[2] , 
        \nOut19_20[1] , \nOut19_20[0] }), .WestIn({\nOut17_20[7] , 
        \nOut17_20[6] , \nOut17_20[5] , \nOut17_20[4] , \nOut17_20[3] , 
        \nOut17_20[2] , \nOut17_20[1] , \nOut17_20[0] }), .Out({\nOut18_20[7] , 
        \nOut18_20[6] , \nOut18_20[5] , \nOut18_20[4] , \nOut18_20[3] , 
        \nOut18_20[2] , \nOut18_20[1] , \nOut18_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_874 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut875[7] , \nScanOut875[6] , 
        \nScanOut875[5] , \nScanOut875[4] , \nScanOut875[3] , \nScanOut875[2] , 
        \nScanOut875[1] , \nScanOut875[0] }), .ScanOut({\nScanOut874[7] , 
        \nScanOut874[6] , \nScanOut874[5] , \nScanOut874[4] , \nScanOut874[3] , 
        \nScanOut874[2] , \nScanOut874[1] , \nScanOut874[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_9[7] , \nOut27_9[6] , \nOut27_9[5] , \nOut27_9[4] , 
        \nOut27_9[3] , \nOut27_9[2] , \nOut27_9[1] , \nOut27_9[0] }), 
        .SouthIn({\nOut27_11[7] , \nOut27_11[6] , \nOut27_11[5] , 
        \nOut27_11[4] , \nOut27_11[3] , \nOut27_11[2] , \nOut27_11[1] , 
        \nOut27_11[0] }), .EastIn({\nOut28_10[7] , \nOut28_10[6] , 
        \nOut28_10[5] , \nOut28_10[4] , \nOut28_10[3] , \nOut28_10[2] , 
        \nOut28_10[1] , \nOut28_10[0] }), .WestIn({\nOut26_10[7] , 
        \nOut26_10[6] , \nOut26_10[5] , \nOut26_10[4] , \nOut26_10[3] , 
        \nOut26_10[2] , \nOut26_10[1] , \nOut26_10[0] }), .Out({\nOut27_10[7] , 
        \nOut27_10[6] , \nOut27_10[5] , \nOut27_10[4] , \nOut27_10[3] , 
        \nOut27_10[2] , \nOut27_10[1] , \nOut27_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_948 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut949[7] , \nScanOut949[6] , 
        \nScanOut949[5] , \nScanOut949[4] , \nScanOut949[3] , \nScanOut949[2] , 
        \nScanOut949[1] , \nScanOut949[0] }), .ScanOut({\nScanOut948[7] , 
        \nScanOut948[6] , \nScanOut948[5] , \nScanOut948[4] , \nScanOut948[3] , 
        \nScanOut948[2] , \nScanOut948[1] , \nScanOut948[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_19[7] , \nOut29_19[6] , \nOut29_19[5] , \nOut29_19[4] , 
        \nOut29_19[3] , \nOut29_19[2] , \nOut29_19[1] , \nOut29_19[0] }), 
        .SouthIn({\nOut29_21[7] , \nOut29_21[6] , \nOut29_21[5] , 
        \nOut29_21[4] , \nOut29_21[3] , \nOut29_21[2] , \nOut29_21[1] , 
        \nOut29_21[0] }), .EastIn({\nOut30_20[7] , \nOut30_20[6] , 
        \nOut30_20[5] , \nOut30_20[4] , \nOut30_20[3] , \nOut30_20[2] , 
        \nOut30_20[1] , \nOut30_20[0] }), .WestIn({\nOut28_20[7] , 
        \nOut28_20[6] , \nOut28_20[5] , \nOut28_20[4] , \nOut28_20[3] , 
        \nOut28_20[2] , \nOut28_20[1] , \nOut28_20[0] }), .Out({\nOut29_20[7] , 
        \nOut29_20[6] , \nOut29_20[5] , \nOut29_20[4] , \nOut29_20[3] , 
        \nOut29_20[2] , \nOut29_20[1] , \nOut29_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_387 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut388[7] , \nScanOut388[6] , 
        \nScanOut388[5] , \nScanOut388[4] , \nScanOut388[3] , \nScanOut388[2] , 
        \nScanOut388[1] , \nScanOut388[0] }), .ScanOut({\nScanOut387[7] , 
        \nScanOut387[6] , \nScanOut387[5] , \nScanOut387[4] , \nScanOut387[3] , 
        \nScanOut387[2] , \nScanOut387[1] , \nScanOut387[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }), 
        .SouthIn({\nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }), .EastIn(
        {\nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }), .WestIn(
        {\nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }), .Out({
        \nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_406 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut407[7] , \nScanOut407[6] , 
        \nScanOut407[5] , \nScanOut407[4] , \nScanOut407[3] , \nScanOut407[2] , 
        \nScanOut407[1] , \nScanOut407[0] }), .ScanOut({\nScanOut406[7] , 
        \nScanOut406[6] , \nScanOut406[5] , \nScanOut406[4] , \nScanOut406[3] , 
        \nScanOut406[2] , \nScanOut406[1] , \nScanOut406[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_21[7] , \nOut12_21[6] , \nOut12_21[5] , \nOut12_21[4] , 
        \nOut12_21[3] , \nOut12_21[2] , \nOut12_21[1] , \nOut12_21[0] }), 
        .SouthIn({\nOut12_23[7] , \nOut12_23[6] , \nOut12_23[5] , 
        \nOut12_23[4] , \nOut12_23[3] , \nOut12_23[2] , \nOut12_23[1] , 
        \nOut12_23[0] }), .EastIn({\nOut13_22[7] , \nOut13_22[6] , 
        \nOut13_22[5] , \nOut13_22[4] , \nOut13_22[3] , \nOut13_22[2] , 
        \nOut13_22[1] , \nOut13_22[0] }), .WestIn({\nOut11_22[7] , 
        \nOut11_22[6] , \nOut11_22[5] , \nOut11_22[4] , \nOut11_22[3] , 
        \nOut11_22[2] , \nOut11_22[1] , \nOut11_22[0] }), .Out({\nOut12_22[7] , 
        \nOut12_22[6] , \nOut12_22[5] , \nOut12_22[4] , \nOut12_22[3] , 
        \nOut12_22[2] , \nOut12_22[1] , \nOut12_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_736 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut737[7] , \nScanOut737[6] , 
        \nScanOut737[5] , \nScanOut737[4] , \nScanOut737[3] , \nScanOut737[2] , 
        \nScanOut737[1] , \nScanOut737[0] }), .ScanOut({\nScanOut736[7] , 
        \nScanOut736[6] , \nScanOut736[5] , \nScanOut736[4] , \nScanOut736[3] , 
        \nScanOut736[2] , \nScanOut736[1] , \nScanOut736[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut23_0[7] , \nOut23_0[6] , 
        \nOut23_0[5] , \nOut23_0[4] , \nOut23_0[3] , \nOut23_0[2] , 
        \nOut23_0[1] , \nOut23_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_100 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut101[7] , \nScanOut101[6] , 
        \nScanOut101[5] , \nScanOut101[4] , \nScanOut101[3] , \nScanOut101[2] , 
        \nScanOut101[1] , \nScanOut101[0] }), .ScanOut({\nScanOut100[7] , 
        \nScanOut100[6] , \nScanOut100[5] , \nScanOut100[4] , \nScanOut100[3] , 
        \nScanOut100[2] , \nScanOut100[1] , \nScanOut100[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_3[7] , \nOut3_3[6] , \nOut3_3[5] , \nOut3_3[4] , \nOut3_3[3] , 
        \nOut3_3[2] , \nOut3_3[1] , \nOut3_3[0] }), .SouthIn({\nOut3_5[7] , 
        \nOut3_5[6] , \nOut3_5[5] , \nOut3_5[4] , \nOut3_5[3] , \nOut3_5[2] , 
        \nOut3_5[1] , \nOut3_5[0] }), .EastIn({\nOut4_4[7] , \nOut4_4[6] , 
        \nOut4_4[5] , \nOut4_4[4] , \nOut4_4[3] , \nOut4_4[2] , \nOut4_4[1] , 
        \nOut4_4[0] }), .WestIn({\nOut2_4[7] , \nOut2_4[6] , \nOut2_4[5] , 
        \nOut2_4[4] , \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , \nOut2_4[0] }), 
        .Out({\nOut3_4[7] , \nOut3_4[6] , \nOut3_4[5] , \nOut3_4[4] , 
        \nOut3_4[3] , \nOut3_4[2] , \nOut3_4[1] , \nOut3_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_711 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut712[7] , \nScanOut712[6] , 
        \nScanOut712[5] , \nScanOut712[4] , \nScanOut712[3] , \nScanOut712[2] , 
        \nScanOut712[1] , \nScanOut712[0] }), .ScanOut({\nScanOut711[7] , 
        \nScanOut711[6] , \nScanOut711[5] , \nScanOut711[4] , \nScanOut711[3] , 
        \nScanOut711[2] , \nScanOut711[1] , \nScanOut711[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_6[7] , \nOut22_6[6] , \nOut22_6[5] , \nOut22_6[4] , 
        \nOut22_6[3] , \nOut22_6[2] , \nOut22_6[1] , \nOut22_6[0] }), 
        .SouthIn({\nOut22_8[7] , \nOut22_8[6] , \nOut22_8[5] , \nOut22_8[4] , 
        \nOut22_8[3] , \nOut22_8[2] , \nOut22_8[1] , \nOut22_8[0] }), .EastIn(
        {\nOut23_7[7] , \nOut23_7[6] , \nOut23_7[5] , \nOut23_7[4] , 
        \nOut23_7[3] , \nOut23_7[2] , \nOut23_7[1] , \nOut23_7[0] }), .WestIn(
        {\nOut21_7[7] , \nOut21_7[6] , \nOut21_7[5] , \nOut21_7[4] , 
        \nOut21_7[3] , \nOut21_7[2] , \nOut21_7[1] , \nOut21_7[0] }), .Out({
        \nOut22_7[7] , \nOut22_7[6] , \nOut22_7[5] , \nOut22_7[4] , 
        \nOut22_7[3] , \nOut22_7[2] , \nOut22_7[1] , \nOut22_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_230 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut231[7] , \nScanOut231[6] , 
        \nScanOut231[5] , \nScanOut231[4] , \nScanOut231[3] , \nScanOut231[2] , 
        \nScanOut231[1] , \nScanOut231[0] }), .ScanOut({\nScanOut230[7] , 
        \nScanOut230[6] , \nScanOut230[5] , \nScanOut230[4] , \nScanOut230[3] , 
        \nScanOut230[2] , \nScanOut230[1] , \nScanOut230[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_5[7] , \nOut7_5[6] , \nOut7_5[5] , \nOut7_5[4] , \nOut7_5[3] , 
        \nOut7_5[2] , \nOut7_5[1] , \nOut7_5[0] }), .SouthIn({\nOut7_7[7] , 
        \nOut7_7[6] , \nOut7_7[5] , \nOut7_7[4] , \nOut7_7[3] , \nOut7_7[2] , 
        \nOut7_7[1] , \nOut7_7[0] }), .EastIn({\nOut8_6[7] , \nOut8_6[6] , 
        \nOut8_6[5] , \nOut8_6[4] , \nOut8_6[3] , \nOut8_6[2] , \nOut8_6[1] , 
        \nOut8_6[0] }), .WestIn({\nOut6_6[7] , \nOut6_6[6] , \nOut6_6[5] , 
        \nOut6_6[4] , \nOut6_6[3] , \nOut6_6[2] , \nOut6_6[1] , \nOut6_6[0] }), 
        .Out({\nOut7_6[7] , \nOut7_6[6] , \nOut7_6[5] , \nOut7_6[4] , 
        \nOut7_6[3] , \nOut7_6[2] , \nOut7_6[1] , \nOut7_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_421 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut422[7] , \nScanOut422[6] , 
        \nScanOut422[5] , \nScanOut422[4] , \nScanOut422[3] , \nScanOut422[2] , 
        \nScanOut422[1] , \nScanOut422[0] }), .ScanOut({\nScanOut421[7] , 
        \nScanOut421[6] , \nScanOut421[5] , \nScanOut421[4] , \nScanOut421[3] , 
        \nScanOut421[2] , \nScanOut421[1] , \nScanOut421[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }), 
        .SouthIn({\nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }), .EastIn(
        {\nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }), .WestIn(
        {\nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }), .Out({
        \nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_681 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut682[7] , \nScanOut682[6] , 
        \nScanOut682[5] , \nScanOut682[4] , \nScanOut682[3] , \nScanOut682[2] , 
        \nScanOut682[1] , \nScanOut682[0] }), .ScanOut({\nScanOut681[7] , 
        \nScanOut681[6] , \nScanOut681[5] , \nScanOut681[4] , \nScanOut681[3] , 
        \nScanOut681[2] , \nScanOut681[1] , \nScanOut681[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_8[7] , \nOut21_8[6] , \nOut21_8[5] , \nOut21_8[4] , 
        \nOut21_8[3] , \nOut21_8[2] , \nOut21_8[1] , \nOut21_8[0] }), 
        .SouthIn({\nOut21_10[7] , \nOut21_10[6] , \nOut21_10[5] , 
        \nOut21_10[4] , \nOut21_10[3] , \nOut21_10[2] , \nOut21_10[1] , 
        \nOut21_10[0] }), .EastIn({\nOut22_9[7] , \nOut22_9[6] , \nOut22_9[5] , 
        \nOut22_9[4] , \nOut22_9[3] , \nOut22_9[2] , \nOut22_9[1] , 
        \nOut22_9[0] }), .WestIn({\nOut20_9[7] , \nOut20_9[6] , \nOut20_9[5] , 
        \nOut20_9[4] , \nOut20_9[3] , \nOut20_9[2] , \nOut20_9[1] , 
        \nOut20_9[0] }), .Out({\nOut21_9[7] , \nOut21_9[6] , \nOut21_9[5] , 
        \nOut21_9[4] , \nOut21_9[3] , \nOut21_9[2] , \nOut21_9[1] , 
        \nOut21_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_853 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut854[7] , \nScanOut854[6] , 
        \nScanOut854[5] , \nScanOut854[4] , \nScanOut854[3] , \nScanOut854[2] , 
        \nScanOut854[1] , \nScanOut854[0] }), .ScanOut({\nScanOut853[7] , 
        \nScanOut853[6] , \nScanOut853[5] , \nScanOut853[4] , \nScanOut853[3] , 
        \nScanOut853[2] , \nScanOut853[1] , \nScanOut853[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_20[7] , \nOut26_20[6] , \nOut26_20[5] , \nOut26_20[4] , 
        \nOut26_20[3] , \nOut26_20[2] , \nOut26_20[1] , \nOut26_20[0] }), 
        .SouthIn({\nOut26_22[7] , \nOut26_22[6] , \nOut26_22[5] , 
        \nOut26_22[4] , \nOut26_22[3] , \nOut26_22[2] , \nOut26_22[1] , 
        \nOut26_22[0] }), .EastIn({\nOut27_21[7] , \nOut27_21[6] , 
        \nOut27_21[5] , \nOut27_21[4] , \nOut27_21[3] , \nOut27_21[2] , 
        \nOut27_21[1] , \nOut27_21[0] }), .WestIn({\nOut25_21[7] , 
        \nOut25_21[6] , \nOut25_21[5] , \nOut25_21[4] , \nOut25_21[3] , 
        \nOut25_21[2] , \nOut25_21[1] , \nOut25_21[0] }), .Out({\nOut26_21[7] , 
        \nOut26_21[6] , \nOut26_21[5] , \nOut26_21[4] , \nOut26_21[3] , 
        \nOut26_21[2] , \nOut26_21[1] , \nOut26_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1017 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1018[7] , \nScanOut1018[6] , 
        \nScanOut1018[5] , \nScanOut1018[4] , \nScanOut1018[3] , 
        \nScanOut1018[2] , \nScanOut1018[1] , \nScanOut1018[0] }), .ScanOut({
        \nScanOut1017[7] , \nScanOut1017[6] , \nScanOut1017[5] , 
        \nScanOut1017[4] , \nScanOut1017[3] , \nScanOut1017[2] , 
        \nScanOut1017[1] , \nScanOut1017[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_25[7] , \nOut31_25[6] , \nOut31_25[5] , 
        \nOut31_25[4] , \nOut31_25[3] , \nOut31_25[2] , \nOut31_25[1] , 
        \nOut31_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_24 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut25[7] , \nScanOut25[6] , 
        \nScanOut25[5] , \nScanOut25[4] , \nScanOut25[3] , \nScanOut25[2] , 
        \nScanOut25[1] , \nScanOut25[0] }), .ScanOut({\nScanOut24[7] , 
        \nScanOut24[6] , \nScanOut24[5] , \nScanOut24[4] , \nScanOut24[3] , 
        \nScanOut24[2] , \nScanOut24[1] , \nScanOut24[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_24[7] , \nOut0_24[6] , 
        \nOut0_24[5] , \nOut0_24[4] , \nOut0_24[3] , \nOut0_24[2] , 
        \nOut0_24[1] , \nOut0_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_51 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut52[7] , \nScanOut52[6] , 
        \nScanOut52[5] , \nScanOut52[4] , \nScanOut52[3] , \nScanOut52[2] , 
        \nScanOut52[1] , \nScanOut52[0] }), .ScanOut({\nScanOut51[7] , 
        \nScanOut51[6] , \nScanOut51[5] , \nScanOut51[4] , \nScanOut51[3] , 
        \nScanOut51[2] , \nScanOut51[1] , \nScanOut51[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_18[7] , \nOut1_18[6] , \nOut1_18[5] , \nOut1_18[4] , 
        \nOut1_18[3] , \nOut1_18[2] , \nOut1_18[1] , \nOut1_18[0] }), 
        .SouthIn({\nOut1_20[7] , \nOut1_20[6] , \nOut1_20[5] , \nOut1_20[4] , 
        \nOut1_20[3] , \nOut1_20[2] , \nOut1_20[1] , \nOut1_20[0] }), .EastIn(
        {\nOut2_19[7] , \nOut2_19[6] , \nOut2_19[5] , \nOut2_19[4] , 
        \nOut2_19[3] , \nOut2_19[2] , \nOut2_19[1] , \nOut2_19[0] }), .WestIn(
        {\nOut0_19[7] , \nOut0_19[6] , \nOut0_19[5] , \nOut0_19[4] , 
        \nOut0_19[3] , \nOut0_19[2] , \nOut0_19[1] , \nOut0_19[0] }), .Out({
        \nOut1_19[7] , \nOut1_19[6] , \nOut1_19[5] , \nOut1_19[4] , 
        \nOut1_19[3] , \nOut1_19[2] , \nOut1_19[1] , \nOut1_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_93 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut94[7] , \nScanOut94[6] , 
        \nScanOut94[5] , \nScanOut94[4] , \nScanOut94[3] , \nScanOut94[2] , 
        \nScanOut94[1] , \nScanOut94[0] }), .ScanOut({\nScanOut93[7] , 
        \nScanOut93[6] , \nScanOut93[5] , \nScanOut93[4] , \nScanOut93[3] , 
        \nScanOut93[2] , \nScanOut93[1] , \nScanOut93[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_28[7] , \nOut2_28[6] , \nOut2_28[5] , \nOut2_28[4] , 
        \nOut2_28[3] , \nOut2_28[2] , \nOut2_28[1] , \nOut2_28[0] }), 
        .SouthIn({\nOut2_30[7] , \nOut2_30[6] , \nOut2_30[5] , \nOut2_30[4] , 
        \nOut2_30[3] , \nOut2_30[2] , \nOut2_30[1] , \nOut2_30[0] }), .EastIn(
        {\nOut3_29[7] , \nOut3_29[6] , \nOut3_29[5] , \nOut3_29[4] , 
        \nOut3_29[3] , \nOut3_29[2] , \nOut3_29[1] , \nOut3_29[0] }), .WestIn(
        {\nOut1_29[7] , \nOut1_29[6] , \nOut1_29[5] , \nOut1_29[4] , 
        \nOut1_29[3] , \nOut1_29[2] , \nOut1_29[1] , \nOut1_29[0] }), .Out({
        \nOut2_29[7] , \nOut2_29[6] , \nOut2_29[5] , \nOut2_29[4] , 
        \nOut2_29[3] , \nOut2_29[2] , \nOut2_29[1] , \nOut2_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_107 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut108[7] , \nScanOut108[6] , 
        \nScanOut108[5] , \nScanOut108[4] , \nScanOut108[3] , \nScanOut108[2] , 
        \nScanOut108[1] , \nScanOut108[0] }), .ScanOut({\nScanOut107[7] , 
        \nScanOut107[6] , \nScanOut107[5] , \nScanOut107[4] , \nScanOut107[3] , 
        \nScanOut107[2] , \nScanOut107[1] , \nScanOut107[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_10[7] , \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , 
        \nOut3_10[3] , \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }), 
        .SouthIn({\nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }), .EastIn(
        {\nOut4_11[7] , \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , 
        \nOut4_11[3] , \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }), .WestIn(
        {\nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), .Out({
        \nOut3_11[7] , \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , 
        \nOut3_11[3] , \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_237 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut238[7] , \nScanOut238[6] , 
        \nScanOut238[5] , \nScanOut238[4] , \nScanOut238[3] , \nScanOut238[2] , 
        \nScanOut238[1] , \nScanOut238[0] }), .ScanOut({\nScanOut237[7] , 
        \nScanOut237[6] , \nScanOut237[5] , \nScanOut237[4] , \nScanOut237[3] , 
        \nScanOut237[2] , \nScanOut237[1] , \nScanOut237[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }), 
        .SouthIn({\nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }), .EastIn(
        {\nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }), .WestIn(
        {\nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }), .Out({
        \nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_968 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut969[7] , \nScanOut969[6] , 
        \nScanOut969[5] , \nScanOut969[4] , \nScanOut969[3] , \nScanOut969[2] , 
        \nScanOut969[1] , \nScanOut969[0] }), .ScanOut({\nScanOut968[7] , 
        \nScanOut968[6] , \nScanOut968[5] , \nScanOut968[4] , \nScanOut968[3] , 
        \nScanOut968[2] , \nScanOut968[1] , \nScanOut968[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_7[7] , \nOut30_7[6] , \nOut30_7[5] , \nOut30_7[4] , 
        \nOut30_7[3] , \nOut30_7[2] , \nOut30_7[1] , \nOut30_7[0] }), 
        .SouthIn({\nOut30_9[7] , \nOut30_9[6] , \nOut30_9[5] , \nOut30_9[4] , 
        \nOut30_9[3] , \nOut30_9[2] , \nOut30_9[1] , \nOut30_9[0] }), .EastIn(
        {\nOut31_8[7] , \nOut31_8[6] , \nOut31_8[5] , \nOut31_8[4] , 
        \nOut31_8[3] , \nOut31_8[2] , \nOut31_8[1] , \nOut31_8[0] }), .WestIn(
        {\nOut29_8[7] , \nOut29_8[6] , \nOut29_8[5] , \nOut29_8[4] , 
        \nOut29_8[3] , \nOut29_8[2] , \nOut29_8[1] , \nOut29_8[0] }), .Out({
        \nOut30_8[7] , \nOut30_8[6] , \nOut30_8[5] , \nOut30_8[4] , 
        \nOut30_8[3] , \nOut30_8[2] , \nOut30_8[1] , \nOut30_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_426 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut427[7] , \nScanOut427[6] , 
        \nScanOut427[5] , \nScanOut427[4] , \nScanOut427[3] , \nScanOut427[2] , 
        \nScanOut427[1] , \nScanOut427[0] }), .ScanOut({\nScanOut426[7] , 
        \nScanOut426[6] , \nScanOut426[5] , \nScanOut426[4] , \nScanOut426[3] , 
        \nScanOut426[2] , \nScanOut426[1] , \nScanOut426[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , \nOut13_9[4] , 
        \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , \nOut13_9[0] }), 
        .SouthIn({\nOut13_11[7] , \nOut13_11[6] , \nOut13_11[5] , 
        \nOut13_11[4] , \nOut13_11[3] , \nOut13_11[2] , \nOut13_11[1] , 
        \nOut13_11[0] }), .EastIn({\nOut14_10[7] , \nOut14_10[6] , 
        \nOut14_10[5] , \nOut14_10[4] , \nOut14_10[3] , \nOut14_10[2] , 
        \nOut14_10[1] , \nOut14_10[0] }), .WestIn({\nOut12_10[7] , 
        \nOut12_10[6] , \nOut12_10[5] , \nOut12_10[4] , \nOut12_10[3] , 
        \nOut12_10[2] , \nOut12_10[1] , \nOut12_10[0] }), .Out({\nOut13_10[7] , 
        \nOut13_10[6] , \nOut13_10[5] , \nOut13_10[4] , \nOut13_10[3] , 
        \nOut13_10[2] , \nOut13_10[1] , \nOut13_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_686 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut687[7] , \nScanOut687[6] , 
        \nScanOut687[5] , \nScanOut687[4] , \nScanOut687[3] , \nScanOut687[2] , 
        \nScanOut687[1] , \nScanOut687[0] }), .ScanOut({\nScanOut686[7] , 
        \nScanOut686[6] , \nScanOut686[5] , \nScanOut686[4] , \nScanOut686[3] , 
        \nScanOut686[2] , \nScanOut686[1] , \nScanOut686[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_13[7] , \nOut21_13[6] , \nOut21_13[5] , \nOut21_13[4] , 
        \nOut21_13[3] , \nOut21_13[2] , \nOut21_13[1] , \nOut21_13[0] }), 
        .SouthIn({\nOut21_15[7] , \nOut21_15[6] , \nOut21_15[5] , 
        \nOut21_15[4] , \nOut21_15[3] , \nOut21_15[2] , \nOut21_15[1] , 
        \nOut21_15[0] }), .EastIn({\nOut22_14[7] , \nOut22_14[6] , 
        \nOut22_14[5] , \nOut22_14[4] , \nOut22_14[3] , \nOut22_14[2] , 
        \nOut22_14[1] , \nOut22_14[0] }), .WestIn({\nOut20_14[7] , 
        \nOut20_14[6] , \nOut20_14[5] , \nOut20_14[4] , \nOut20_14[3] , 
        \nOut20_14[2] , \nOut20_14[1] , \nOut20_14[0] }), .Out({\nOut21_14[7] , 
        \nOut21_14[6] , \nOut21_14[5] , \nOut21_14[4] , \nOut21_14[3] , 
        \nOut21_14[2] , \nOut21_14[1] , \nOut21_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_854 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut855[7] , \nScanOut855[6] , 
        \nScanOut855[5] , \nScanOut855[4] , \nScanOut855[3] , \nScanOut855[2] , 
        \nScanOut855[1] , \nScanOut855[0] }), .ScanOut({\nScanOut854[7] , 
        \nScanOut854[6] , \nScanOut854[5] , \nScanOut854[4] , \nScanOut854[3] , 
        \nScanOut854[2] , \nScanOut854[1] , \nScanOut854[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_21[7] , \nOut26_21[6] , \nOut26_21[5] , \nOut26_21[4] , 
        \nOut26_21[3] , \nOut26_21[2] , \nOut26_21[1] , \nOut26_21[0] }), 
        .SouthIn({\nOut26_23[7] , \nOut26_23[6] , \nOut26_23[5] , 
        \nOut26_23[4] , \nOut26_23[3] , \nOut26_23[2] , \nOut26_23[1] , 
        \nOut26_23[0] }), .EastIn({\nOut27_22[7] , \nOut27_22[6] , 
        \nOut27_22[5] , \nOut27_22[4] , \nOut27_22[3] , \nOut27_22[2] , 
        \nOut27_22[1] , \nOut27_22[0] }), .WestIn({\nOut25_22[7] , 
        \nOut25_22[6] , \nOut25_22[5] , \nOut25_22[4] , \nOut25_22[3] , 
        \nOut25_22[2] , \nOut25_22[1] , \nOut25_22[0] }), .Out({\nOut26_22[7] , 
        \nOut26_22[6] , \nOut26_22[5] , \nOut26_22[4] , \nOut26_22[3] , 
        \nOut26_22[2] , \nOut26_22[1] , \nOut26_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1010 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1011[7] , \nScanOut1011[6] , 
        \nScanOut1011[5] , \nScanOut1011[4] , \nScanOut1011[3] , 
        \nScanOut1011[2] , \nScanOut1011[1] , \nScanOut1011[0] }), .ScanOut({
        \nScanOut1010[7] , \nScanOut1010[6] , \nScanOut1010[5] , 
        \nScanOut1010[4] , \nScanOut1010[3] , \nScanOut1010[2] , 
        \nScanOut1010[1] , \nScanOut1010[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_18[7] , \nOut31_18[6] , \nOut31_18[5] , 
        \nOut31_18[4] , \nOut31_18[3] , \nOut31_18[2] , \nOut31_18[1] , 
        \nOut31_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_716 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut717[7] , \nScanOut717[6] , 
        \nScanOut717[5] , \nScanOut717[4] , \nScanOut717[3] , \nScanOut717[2] , 
        \nScanOut717[1] , \nScanOut717[0] }), .ScanOut({\nScanOut716[7] , 
        \nScanOut716[6] , \nScanOut716[5] , \nScanOut716[4] , \nScanOut716[3] , 
        \nScanOut716[2] , \nScanOut716[1] , \nScanOut716[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_11[7] , \nOut22_11[6] , \nOut22_11[5] , \nOut22_11[4] , 
        \nOut22_11[3] , \nOut22_11[2] , \nOut22_11[1] , \nOut22_11[0] }), 
        .SouthIn({\nOut22_13[7] , \nOut22_13[6] , \nOut22_13[5] , 
        \nOut22_13[4] , \nOut22_13[3] , \nOut22_13[2] , \nOut22_13[1] , 
        \nOut22_13[0] }), .EastIn({\nOut23_12[7] , \nOut23_12[6] , 
        \nOut23_12[5] , \nOut23_12[4] , \nOut23_12[3] , \nOut23_12[2] , 
        \nOut23_12[1] , \nOut23_12[0] }), .WestIn({\nOut21_12[7] , 
        \nOut21_12[6] , \nOut21_12[5] , \nOut21_12[4] , \nOut21_12[3] , 
        \nOut21_12[2] , \nOut21_12[1] , \nOut21_12[0] }), .Out({\nOut22_12[7] , 
        \nOut22_12[6] , \nOut22_12[5] , \nOut22_12[4] , \nOut22_12[3] , 
        \nOut22_12[2] , \nOut22_12[1] , \nOut22_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_120 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut121[7] , \nScanOut121[6] , 
        \nScanOut121[5] , \nScanOut121[4] , \nScanOut121[3] , \nScanOut121[2] , 
        \nScanOut121[1] , \nScanOut121[0] }), .ScanOut({\nScanOut120[7] , 
        \nScanOut120[6] , \nScanOut120[5] , \nScanOut120[4] , \nScanOut120[3] , 
        \nScanOut120[2] , \nScanOut120[1] , \nScanOut120[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_23[7] , \nOut3_23[6] , \nOut3_23[5] , \nOut3_23[4] , 
        \nOut3_23[3] , \nOut3_23[2] , \nOut3_23[1] , \nOut3_23[0] }), 
        .SouthIn({\nOut3_25[7] , \nOut3_25[6] , \nOut3_25[5] , \nOut3_25[4] , 
        \nOut3_25[3] , \nOut3_25[2] , \nOut3_25[1] , \nOut3_25[0] }), .EastIn(
        {\nOut4_24[7] , \nOut4_24[6] , \nOut4_24[5] , \nOut4_24[4] , 
        \nOut4_24[3] , \nOut4_24[2] , \nOut4_24[1] , \nOut4_24[0] }), .WestIn(
        {\nOut2_24[7] , \nOut2_24[6] , \nOut2_24[5] , \nOut2_24[4] , 
        \nOut2_24[3] , \nOut2_24[2] , \nOut2_24[1] , \nOut2_24[0] }), .Out({
        \nOut3_24[7] , \nOut3_24[6] , \nOut3_24[5] , \nOut3_24[4] , 
        \nOut3_24[3] , \nOut3_24[2] , \nOut3_24[1] , \nOut3_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_731 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut732[7] , \nScanOut732[6] , 
        \nScanOut732[5] , \nScanOut732[4] , \nScanOut732[3] , \nScanOut732[2] , 
        \nScanOut732[1] , \nScanOut732[0] }), .ScanOut({\nScanOut731[7] , 
        \nScanOut731[6] , \nScanOut731[5] , \nScanOut731[4] , \nScanOut731[3] , 
        \nScanOut731[2] , \nScanOut731[1] , \nScanOut731[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_26[7] , \nOut22_26[6] , \nOut22_26[5] , \nOut22_26[4] , 
        \nOut22_26[3] , \nOut22_26[2] , \nOut22_26[1] , \nOut22_26[0] }), 
        .SouthIn({\nOut22_28[7] , \nOut22_28[6] , \nOut22_28[5] , 
        \nOut22_28[4] , \nOut22_28[3] , \nOut22_28[2] , \nOut22_28[1] , 
        \nOut22_28[0] }), .EastIn({\nOut23_27[7] , \nOut23_27[6] , 
        \nOut23_27[5] , \nOut23_27[4] , \nOut23_27[3] , \nOut23_27[2] , 
        \nOut23_27[1] , \nOut23_27[0] }), .WestIn({\nOut21_27[7] , 
        \nOut21_27[6] , \nOut21_27[5] , \nOut21_27[4] , \nOut21_27[3] , 
        \nOut21_27[2] , \nOut21_27[1] , \nOut21_27[0] }), .Out({\nOut22_27[7] , 
        \nOut22_27[6] , \nOut22_27[5] , \nOut22_27[4] , \nOut22_27[3] , 
        \nOut22_27[2] , \nOut22_27[1] , \nOut22_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_169 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut170[7] , \nScanOut170[6] , 
        \nScanOut170[5] , \nScanOut170[4] , \nScanOut170[3] , \nScanOut170[2] , 
        \nScanOut170[1] , \nScanOut170[0] }), .ScanOut({\nScanOut169[7] , 
        \nScanOut169[6] , \nScanOut169[5] , \nScanOut169[4] , \nScanOut169[3] , 
        \nScanOut169[2] , \nScanOut169[1] , \nScanOut169[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_8[7] , \nOut5_8[6] , \nOut5_8[5] , \nOut5_8[4] , \nOut5_8[3] , 
        \nOut5_8[2] , \nOut5_8[1] , \nOut5_8[0] }), .SouthIn({\nOut5_10[7] , 
        \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , \nOut5_10[3] , 
        \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }), .EastIn({\nOut6_9[7] , 
        \nOut6_9[6] , \nOut6_9[5] , \nOut6_9[4] , \nOut6_9[3] , \nOut6_9[2] , 
        \nOut6_9[1] , \nOut6_9[0] }), .WestIn({\nOut4_9[7] , \nOut4_9[6] , 
        \nOut4_9[5] , \nOut4_9[4] , \nOut4_9[3] , \nOut4_9[2] , \nOut4_9[1] , 
        \nOut4_9[0] }), .Out({\nOut5_9[7] , \nOut5_9[6] , \nOut5_9[5] , 
        \nOut5_9[4] , \nOut5_9[3] , \nOut5_9[2] , \nOut5_9[1] , \nOut5_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_210 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut211[7] , \nScanOut211[6] , 
        \nScanOut211[5] , \nScanOut211[4] , \nScanOut211[3] , \nScanOut211[2] , 
        \nScanOut211[1] , \nScanOut211[0] }), .ScanOut({\nScanOut210[7] , 
        \nScanOut210[6] , \nScanOut210[5] , \nScanOut210[4] , \nScanOut210[3] , 
        \nScanOut210[2] , \nScanOut210[1] , \nScanOut210[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_17[7] , \nOut6_17[6] , \nOut6_17[5] , \nOut6_17[4] , 
        \nOut6_17[3] , \nOut6_17[2] , \nOut6_17[1] , \nOut6_17[0] }), 
        .SouthIn({\nOut6_19[7] , \nOut6_19[6] , \nOut6_19[5] , \nOut6_19[4] , 
        \nOut6_19[3] , \nOut6_19[2] , \nOut6_19[1] , \nOut6_19[0] }), .EastIn(
        {\nOut7_18[7] , \nOut7_18[6] , \nOut7_18[5] , \nOut7_18[4] , 
        \nOut7_18[3] , \nOut7_18[2] , \nOut7_18[1] , \nOut7_18[0] }), .WestIn(
        {\nOut5_18[7] , \nOut5_18[6] , \nOut5_18[5] , \nOut5_18[4] , 
        \nOut5_18[3] , \nOut5_18[2] , \nOut5_18[1] , \nOut5_18[0] }), .Out({
        \nOut6_18[7] , \nOut6_18[6] , \nOut6_18[5] , \nOut6_18[4] , 
        \nOut6_18[3] , \nOut6_18[2] , \nOut6_18[1] , \nOut6_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_380 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut381[7] , \nScanOut381[6] , 
        \nScanOut381[5] , \nScanOut381[4] , \nScanOut381[3] , \nScanOut381[2] , 
        \nScanOut381[1] , \nScanOut381[0] }), .ScanOut({\nScanOut380[7] , 
        \nScanOut380[6] , \nScanOut380[5] , \nScanOut380[4] , \nScanOut380[3] , 
        \nScanOut380[2] , \nScanOut380[1] , \nScanOut380[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_27[7] , \nOut11_27[6] , \nOut11_27[5] , \nOut11_27[4] , 
        \nOut11_27[3] , \nOut11_27[2] , \nOut11_27[1] , \nOut11_27[0] }), 
        .SouthIn({\nOut11_29[7] , \nOut11_29[6] , \nOut11_29[5] , 
        \nOut11_29[4] , \nOut11_29[3] , \nOut11_29[2] , \nOut11_29[1] , 
        \nOut11_29[0] }), .EastIn({\nOut12_28[7] , \nOut12_28[6] , 
        \nOut12_28[5] , \nOut12_28[4] , \nOut12_28[3] , \nOut12_28[2] , 
        \nOut12_28[1] , \nOut12_28[0] }), .WestIn({\nOut10_28[7] , 
        \nOut10_28[6] , \nOut10_28[5] , \nOut10_28[4] , \nOut10_28[3] , 
        \nOut10_28[2] , \nOut10_28[1] , \nOut10_28[0] }), .Out({\nOut11_28[7] , 
        \nOut11_28[6] , \nOut11_28[5] , \nOut11_28[4] , \nOut11_28[3] , 
        \nOut11_28[2] , \nOut11_28[1] , \nOut11_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_401 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut402[7] , \nScanOut402[6] , 
        \nScanOut402[5] , \nScanOut402[4] , \nScanOut402[3] , \nScanOut402[2] , 
        \nScanOut402[1] , \nScanOut402[0] }), .ScanOut({\nScanOut401[7] , 
        \nScanOut401[6] , \nScanOut401[5] , \nScanOut401[4] , \nScanOut401[3] , 
        \nScanOut401[2] , \nScanOut401[1] , \nScanOut401[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_16[7] , \nOut12_16[6] , \nOut12_16[5] , \nOut12_16[4] , 
        \nOut12_16[3] , \nOut12_16[2] , \nOut12_16[1] , \nOut12_16[0] }), 
        .SouthIn({\nOut12_18[7] , \nOut12_18[6] , \nOut12_18[5] , 
        \nOut12_18[4] , \nOut12_18[3] , \nOut12_18[2] , \nOut12_18[1] , 
        \nOut12_18[0] }), .EastIn({\nOut13_17[7] , \nOut13_17[6] , 
        \nOut13_17[5] , \nOut13_17[4] , \nOut13_17[3] , \nOut13_17[2] , 
        \nOut13_17[1] , \nOut13_17[0] }), .WestIn({\nOut11_17[7] , 
        \nOut11_17[6] , \nOut11_17[5] , \nOut11_17[4] , \nOut11_17[3] , 
        \nOut11_17[2] , \nOut11_17[1] , \nOut11_17[0] }), .Out({\nOut12_17[7] , 
        \nOut12_17[6] , \nOut12_17[5] , \nOut12_17[4] , \nOut12_17[3] , 
        \nOut12_17[2] , \nOut12_17[1] , \nOut12_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_259 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut260[7] , \nScanOut260[6] , 
        \nScanOut260[5] , \nScanOut260[4] , \nScanOut260[3] , \nScanOut260[2] , 
        \nScanOut260[1] , \nScanOut260[0] }), .ScanOut({\nScanOut259[7] , 
        \nScanOut259[6] , \nScanOut259[5] , \nScanOut259[4] , \nScanOut259[3] , 
        \nScanOut259[2] , \nScanOut259[1] , \nScanOut259[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_2[7] , \nOut8_2[6] , \nOut8_2[5] , \nOut8_2[4] , \nOut8_2[3] , 
        \nOut8_2[2] , \nOut8_2[1] , \nOut8_2[0] }), .SouthIn({\nOut8_4[7] , 
        \nOut8_4[6] , \nOut8_4[5] , \nOut8_4[4] , \nOut8_4[3] , \nOut8_4[2] , 
        \nOut8_4[1] , \nOut8_4[0] }), .EastIn({\nOut9_3[7] , \nOut9_3[6] , 
        \nOut9_3[5] , \nOut9_3[4] , \nOut9_3[3] , \nOut9_3[2] , \nOut9_3[1] , 
        \nOut9_3[0] }), .WestIn({\nOut7_3[7] , \nOut7_3[6] , \nOut7_3[5] , 
        \nOut7_3[4] , \nOut7_3[3] , \nOut7_3[2] , \nOut7_3[1] , \nOut7_3[0] }), 
        .Out({\nOut8_3[7] , \nOut8_3[6] , \nOut8_3[5] , \nOut8_3[4] , 
        \nOut8_3[3] , \nOut8_3[2] , \nOut8_3[1] , \nOut8_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_448 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut449[7] , \nScanOut449[6] , 
        \nScanOut449[5] , \nScanOut449[4] , \nScanOut449[3] , \nScanOut449[2] , 
        \nScanOut449[1] , \nScanOut449[0] }), .ScanOut({\nScanOut448[7] , 
        \nScanOut448[6] , \nScanOut448[5] , \nScanOut448[4] , \nScanOut448[3] , 
        \nScanOut448[2] , \nScanOut448[1] , \nScanOut448[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut14_0[7] , \nOut14_0[6] , 
        \nOut14_0[5] , \nOut14_0[4] , \nOut14_0[3] , \nOut14_0[2] , 
        \nOut14_0[1] , \nOut14_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_591 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut592[7] , \nScanOut592[6] , 
        \nScanOut592[5] , \nScanOut592[4] , \nScanOut592[3] , \nScanOut592[2] , 
        \nScanOut592[1] , \nScanOut592[0] }), .ScanOut({\nScanOut591[7] , 
        \nScanOut591[6] , \nScanOut591[5] , \nScanOut591[4] , \nScanOut591[3] , 
        \nScanOut591[2] , \nScanOut591[1] , \nScanOut591[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_14[7] , \nOut18_14[6] , \nOut18_14[5] , \nOut18_14[4] , 
        \nOut18_14[3] , \nOut18_14[2] , \nOut18_14[1] , \nOut18_14[0] }), 
        .SouthIn({\nOut18_16[7] , \nOut18_16[6] , \nOut18_16[5] , 
        \nOut18_16[4] , \nOut18_16[3] , \nOut18_16[2] , \nOut18_16[1] , 
        \nOut18_16[0] }), .EastIn({\nOut19_15[7] , \nOut19_15[6] , 
        \nOut19_15[5] , \nOut19_15[4] , \nOut19_15[3] , \nOut19_15[2] , 
        \nOut19_15[1] , \nOut19_15[0] }), .WestIn({\nOut17_15[7] , 
        \nOut17_15[6] , \nOut17_15[5] , \nOut17_15[4] , \nOut17_15[3] , 
        \nOut17_15[2] , \nOut17_15[1] , \nOut17_15[0] }), .Out({\nOut18_15[7] , 
        \nOut18_15[6] , \nOut18_15[5] , \nOut18_15[4] , \nOut18_15[3] , 
        \nOut18_15[2] , \nOut18_15[1] , \nOut18_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_873 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut874[7] , \nScanOut874[6] , 
        \nScanOut874[5] , \nScanOut874[4] , \nScanOut874[3] , \nScanOut874[2] , 
        \nScanOut874[1] , \nScanOut874[0] }), .ScanOut({\nScanOut873[7] , 
        \nScanOut873[6] , \nScanOut873[5] , \nScanOut873[4] , \nScanOut873[3] , 
        \nScanOut873[2] , \nScanOut873[1] , \nScanOut873[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_8[7] , \nOut27_8[6] , \nOut27_8[5] , \nOut27_8[4] , 
        \nOut27_8[3] , \nOut27_8[2] , \nOut27_8[1] , \nOut27_8[0] }), 
        .SouthIn({\nOut27_10[7] , \nOut27_10[6] , \nOut27_10[5] , 
        \nOut27_10[4] , \nOut27_10[3] , \nOut27_10[2] , \nOut27_10[1] , 
        \nOut27_10[0] }), .EastIn({\nOut28_9[7] , \nOut28_9[6] , \nOut28_9[5] , 
        \nOut28_9[4] , \nOut28_9[3] , \nOut28_9[2] , \nOut28_9[1] , 
        \nOut28_9[0] }), .WestIn({\nOut26_9[7] , \nOut26_9[6] , \nOut26_9[5] , 
        \nOut26_9[4] , \nOut26_9[3] , \nOut26_9[2] , \nOut26_9[1] , 
        \nOut26_9[0] }), .Out({\nOut27_9[7] , \nOut27_9[6] , \nOut27_9[5] , 
        \nOut27_9[4] , \nOut27_9[3] , \nOut27_9[2] , \nOut27_9[1] , 
        \nOut27_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_778 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut779[7] , \nScanOut779[6] , 
        \nScanOut779[5] , \nScanOut779[4] , \nScanOut779[3] , \nScanOut779[2] , 
        \nScanOut779[1] , \nScanOut779[0] }), .ScanOut({\nScanOut778[7] , 
        \nScanOut778[6] , \nScanOut778[5] , \nScanOut778[4] , \nScanOut778[3] , 
        \nScanOut778[2] , \nScanOut778[1] , \nScanOut778[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_9[7] , \nOut24_9[6] , \nOut24_9[5] , \nOut24_9[4] , 
        \nOut24_9[3] , \nOut24_9[2] , \nOut24_9[1] , \nOut24_9[0] }), 
        .SouthIn({\nOut24_11[7] , \nOut24_11[6] , \nOut24_11[5] , 
        \nOut24_11[4] , \nOut24_11[3] , \nOut24_11[2] , \nOut24_11[1] , 
        \nOut24_11[0] }), .EastIn({\nOut25_10[7] , \nOut25_10[6] , 
        \nOut25_10[5] , \nOut25_10[4] , \nOut25_10[3] , \nOut25_10[2] , 
        \nOut25_10[1] , \nOut25_10[0] }), .WestIn({\nOut23_10[7] , 
        \nOut23_10[6] , \nOut23_10[5] , \nOut23_10[4] , \nOut23_10[3] , 
        \nOut23_10[2] , \nOut23_10[1] , \nOut23_10[0] }), .Out({\nOut24_10[7] , 
        \nOut24_10[6] , \nOut24_10[5] , \nOut24_10[4] , \nOut24_10[3] , 
        \nOut24_10[2] , \nOut24_10[1] , \nOut24_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_76 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut77[7] , \nScanOut77[6] , 
        \nScanOut77[5] , \nScanOut77[4] , \nScanOut77[3] , \nScanOut77[2] , 
        \nScanOut77[1] , \nScanOut77[0] }), .ScanOut({\nScanOut76[7] , 
        \nScanOut76[6] , \nScanOut76[5] , \nScanOut76[4] , \nScanOut76[3] , 
        \nScanOut76[2] , \nScanOut76[1] , \nScanOut76[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), 
        .SouthIn({\nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), .EastIn(
        {\nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }), .WestIn(
        {\nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), .Out({
        \nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_342 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut343[7] , \nScanOut343[6] , 
        \nScanOut343[5] , \nScanOut343[4] , \nScanOut343[3] , \nScanOut343[2] , 
        \nScanOut343[1] , \nScanOut343[0] }), .ScanOut({\nScanOut342[7] , 
        \nScanOut342[6] , \nScanOut342[5] , \nScanOut342[4] , \nScanOut342[3] , 
        \nScanOut342[2] , \nScanOut342[1] , \nScanOut342[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_21[7] , \nOut10_21[6] , \nOut10_21[5] , \nOut10_21[4] , 
        \nOut10_21[3] , \nOut10_21[2] , \nOut10_21[1] , \nOut10_21[0] }), 
        .SouthIn({\nOut10_23[7] , \nOut10_23[6] , \nOut10_23[5] , 
        \nOut10_23[4] , \nOut10_23[3] , \nOut10_23[2] , \nOut10_23[1] , 
        \nOut10_23[0] }), .EastIn({\nOut11_22[7] , \nOut11_22[6] , 
        \nOut11_22[5] , \nOut11_22[4] , \nOut11_22[3] , \nOut11_22[2] , 
        \nOut11_22[1] , \nOut11_22[0] }), .WestIn({\nOut9_22[7] , 
        \nOut9_22[6] , \nOut9_22[5] , \nOut9_22[4] , \nOut9_22[3] , 
        \nOut9_22[2] , \nOut9_22[1] , \nOut9_22[0] }), .Out({\nOut10_22[7] , 
        \nOut10_22[6] , \nOut10_22[5] , \nOut10_22[4] , \nOut10_22[3] , 
        \nOut10_22[2] , \nOut10_22[1] , \nOut10_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_365 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut366[7] , \nScanOut366[6] , 
        \nScanOut366[5] , \nScanOut366[4] , \nScanOut366[3] , \nScanOut366[2] , 
        \nScanOut366[1] , \nScanOut366[0] }), .ScanOut({\nScanOut365[7] , 
        \nScanOut365[6] , \nScanOut365[5] , \nScanOut365[4] , \nScanOut365[3] , 
        \nScanOut365[2] , \nScanOut365[1] , \nScanOut365[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_12[7] , \nOut11_12[6] , \nOut11_12[5] , \nOut11_12[4] , 
        \nOut11_12[3] , \nOut11_12[2] , \nOut11_12[1] , \nOut11_12[0] }), 
        .SouthIn({\nOut11_14[7] , \nOut11_14[6] , \nOut11_14[5] , 
        \nOut11_14[4] , \nOut11_14[3] , \nOut11_14[2] , \nOut11_14[1] , 
        \nOut11_14[0] }), .EastIn({\nOut12_13[7] , \nOut12_13[6] , 
        \nOut12_13[5] , \nOut12_13[4] , \nOut12_13[3] , \nOut12_13[2] , 
        \nOut12_13[1] , \nOut12_13[0] }), .WestIn({\nOut10_13[7] , 
        \nOut10_13[6] , \nOut10_13[5] , \nOut10_13[4] , \nOut10_13[3] , 
        \nOut10_13[2] , \nOut10_13[1] , \nOut10_13[0] }), .Out({\nOut11_13[7] , 
        \nOut11_13[6] , \nOut11_13[5] , \nOut11_13[4] , \nOut11_13[3] , 
        \nOut11_13[2] , \nOut11_13[1] , \nOut11_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_574 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut575[7] , \nScanOut575[6] , 
        \nScanOut575[5] , \nScanOut575[4] , \nScanOut575[3] , \nScanOut575[2] , 
        \nScanOut575[1] , \nScanOut575[0] }), .ScanOut({\nScanOut574[7] , 
        \nScanOut574[6] , \nScanOut574[5] , \nScanOut574[4] , \nScanOut574[3] , 
        \nScanOut574[2] , \nScanOut574[1] , \nScanOut574[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_29[7] , \nOut17_29[6] , \nOut17_29[5] , \nOut17_29[4] , 
        \nOut17_29[3] , \nOut17_29[2] , \nOut17_29[1] , \nOut17_29[0] }), 
        .SouthIn({\nOut17_31[7] , \nOut17_31[6] , \nOut17_31[5] , 
        \nOut17_31[4] , \nOut17_31[3] , \nOut17_31[2] , \nOut17_31[1] , 
        \nOut17_31[0] }), .EastIn({\nOut18_30[7] , \nOut18_30[6] , 
        \nOut18_30[5] , \nOut18_30[4] , \nOut18_30[3] , \nOut18_30[2] , 
        \nOut18_30[1] , \nOut18_30[0] }), .WestIn({\nOut16_30[7] , 
        \nOut16_30[6] , \nOut16_30[5] , \nOut16_30[4] , \nOut16_30[3] , 
        \nOut16_30[2] , \nOut16_30[1] , \nOut16_30[0] }), .Out({\nOut17_30[7] , 
        \nOut17_30[6] , \nOut17_30[5] , \nOut17_30[4] , \nOut17_30[3] , 
        \nOut17_30[2] , \nOut17_30[1] , \nOut17_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_644 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut645[7] , \nScanOut645[6] , 
        \nScanOut645[5] , \nScanOut645[4] , \nScanOut645[3] , \nScanOut645[2] , 
        \nScanOut645[1] , \nScanOut645[0] }), .ScanOut({\nScanOut644[7] , 
        \nScanOut644[6] , \nScanOut644[5] , \nScanOut644[4] , \nScanOut644[3] , 
        \nScanOut644[2] , \nScanOut644[1] , \nScanOut644[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_3[7] , \nOut20_3[6] , \nOut20_3[5] , \nOut20_3[4] , 
        \nOut20_3[3] , \nOut20_3[2] , \nOut20_3[1] , \nOut20_3[0] }), 
        .SouthIn({\nOut20_5[7] , \nOut20_5[6] , \nOut20_5[5] , \nOut20_5[4] , 
        \nOut20_5[3] , \nOut20_5[2] , \nOut20_5[1] , \nOut20_5[0] }), .EastIn(
        {\nOut21_4[7] , \nOut21_4[6] , \nOut21_4[5] , \nOut21_4[4] , 
        \nOut21_4[3] , \nOut21_4[2] , \nOut21_4[1] , \nOut21_4[0] }), .WestIn(
        {\nOut19_4[7] , \nOut19_4[6] , \nOut19_4[5] , \nOut19_4[4] , 
        \nOut19_4[3] , \nOut19_4[2] , \nOut19_4[1] , \nOut19_4[0] }), .Out({
        \nOut20_4[7] , \nOut20_4[6] , \nOut20_4[5] , \nOut20_4[4] , 
        \nOut20_4[3] , \nOut20_4[2] , \nOut20_4[1] , \nOut20_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_896 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut897[7] , \nScanOut897[6] , 
        \nScanOut897[5] , \nScanOut897[4] , \nScanOut897[3] , \nScanOut897[2] , 
        \nScanOut897[1] , \nScanOut897[0] }), .ScanOut({\nScanOut896[7] , 
        \nScanOut896[6] , \nScanOut896[5] , \nScanOut896[4] , \nScanOut896[3] , 
        \nScanOut896[2] , \nScanOut896[1] , \nScanOut896[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut28_0[7] , \nOut28_0[6] , 
        \nOut28_0[5] , \nOut28_0[4] , \nOut28_0[3] , \nOut28_0[2] , 
        \nOut28_0[1] , \nOut28_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_906 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut907[7] , \nScanOut907[6] , 
        \nScanOut907[5] , \nScanOut907[4] , \nScanOut907[3] , \nScanOut907[2] , 
        \nScanOut907[1] , \nScanOut907[0] }), .ScanOut({\nScanOut906[7] , 
        \nScanOut906[6] , \nScanOut906[5] , \nScanOut906[4] , \nScanOut906[3] , 
        \nScanOut906[2] , \nScanOut906[1] , \nScanOut906[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_9[7] , \nOut28_9[6] , \nOut28_9[5] , \nOut28_9[4] , 
        \nOut28_9[3] , \nOut28_9[2] , \nOut28_9[1] , \nOut28_9[0] }), 
        .SouthIn({\nOut28_11[7] , \nOut28_11[6] , \nOut28_11[5] , 
        \nOut28_11[4] , \nOut28_11[3] , \nOut28_11[2] , \nOut28_11[1] , 
        \nOut28_11[0] }), .EastIn({\nOut29_10[7] , \nOut29_10[6] , 
        \nOut29_10[5] , \nOut29_10[4] , \nOut29_10[3] , \nOut29_10[2] , 
        \nOut29_10[1] , \nOut29_10[0] }), .WestIn({\nOut27_10[7] , 
        \nOut27_10[6] , \nOut27_10[5] , \nOut27_10[4] , \nOut27_10[3] , 
        \nOut27_10[2] , \nOut27_10[1] , \nOut27_10[0] }), .Out({\nOut28_10[7] , 
        \nOut28_10[6] , \nOut28_10[5] , \nOut28_10[4] , \nOut28_10[3] , 
        \nOut28_10[2] , \nOut28_10[1] , \nOut28_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_553 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut554[7] , \nScanOut554[6] , 
        \nScanOut554[5] , \nScanOut554[4] , \nScanOut554[3] , \nScanOut554[2] , 
        \nScanOut554[1] , \nScanOut554[0] }), .ScanOut({\nScanOut553[7] , 
        \nScanOut553[6] , \nScanOut553[5] , \nScanOut553[4] , \nScanOut553[3] , 
        \nScanOut553[2] , \nScanOut553[1] , \nScanOut553[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_8[7] , \nOut17_8[6] , \nOut17_8[5] , \nOut17_8[4] , 
        \nOut17_8[3] , \nOut17_8[2] , \nOut17_8[1] , \nOut17_8[0] }), 
        .SouthIn({\nOut17_10[7] , \nOut17_10[6] , \nOut17_10[5] , 
        \nOut17_10[4] , \nOut17_10[3] , \nOut17_10[2] , \nOut17_10[1] , 
        \nOut17_10[0] }), .EastIn({\nOut18_9[7] , \nOut18_9[6] , \nOut18_9[5] , 
        \nOut18_9[4] , \nOut18_9[3] , \nOut18_9[2] , \nOut18_9[1] , 
        \nOut18_9[0] }), .WestIn({\nOut16_9[7] , \nOut16_9[6] , \nOut16_9[5] , 
        \nOut16_9[4] , \nOut16_9[3] , \nOut16_9[2] , \nOut16_9[1] , 
        \nOut16_9[0] }), .Out({\nOut17_9[7] , \nOut17_9[6] , \nOut17_9[5] , 
        \nOut17_9[4] , \nOut17_9[3] , \nOut17_9[2] , \nOut17_9[1] , 
        \nOut17_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_921 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut922[7] , \nScanOut922[6] , 
        \nScanOut922[5] , \nScanOut922[4] , \nScanOut922[3] , \nScanOut922[2] , 
        \nScanOut922[1] , \nScanOut922[0] }), .ScanOut({\nScanOut921[7] , 
        \nScanOut921[6] , \nScanOut921[5] , \nScanOut921[4] , \nScanOut921[3] , 
        \nScanOut921[2] , \nScanOut921[1] , \nScanOut921[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_24[7] , \nOut28_24[6] , \nOut28_24[5] , \nOut28_24[4] , 
        \nOut28_24[3] , \nOut28_24[2] , \nOut28_24[1] , \nOut28_24[0] }), 
        .SouthIn({\nOut28_26[7] , \nOut28_26[6] , \nOut28_26[5] , 
        \nOut28_26[4] , \nOut28_26[3] , \nOut28_26[2] , \nOut28_26[1] , 
        \nOut28_26[0] }), .EastIn({\nOut29_25[7] , \nOut29_25[6] , 
        \nOut29_25[5] , \nOut29_25[4] , \nOut29_25[3] , \nOut29_25[2] , 
        \nOut29_25[1] , \nOut29_25[0] }), .WestIn({\nOut27_25[7] , 
        \nOut27_25[6] , \nOut27_25[5] , \nOut27_25[4] , \nOut27_25[3] , 
        \nOut27_25[2] , \nOut27_25[1] , \nOut27_25[0] }), .Out({\nOut28_25[7] , 
        \nOut28_25[6] , \nOut28_25[5] , \nOut28_25[4] , \nOut28_25[3] , 
        \nOut28_25[2] , \nOut28_25[1] , \nOut28_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_88 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut89[7] , \nScanOut89[6] , 
        \nScanOut89[5] , \nScanOut89[4] , \nScanOut89[3] , \nScanOut89[2] , 
        \nScanOut89[1] , \nScanOut89[0] }), .ScanOut({\nScanOut88[7] , 
        \nScanOut88[6] , \nScanOut88[5] , \nScanOut88[4] , \nScanOut88[3] , 
        \nScanOut88[2] , \nScanOut88[1] , \nScanOut88[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_23[7] , \nOut2_23[6] , \nOut2_23[5] , \nOut2_23[4] , 
        \nOut2_23[3] , \nOut2_23[2] , \nOut2_23[1] , \nOut2_23[0] }), 
        .SouthIn({\nOut2_25[7] , \nOut2_25[6] , \nOut2_25[5] , \nOut2_25[4] , 
        \nOut2_25[3] , \nOut2_25[2] , \nOut2_25[1] , \nOut2_25[0] }), .EastIn(
        {\nOut3_24[7] , \nOut3_24[6] , \nOut3_24[5] , \nOut3_24[4] , 
        \nOut3_24[3] , \nOut3_24[2] , \nOut3_24[1] , \nOut3_24[0] }), .WestIn(
        {\nOut1_24[7] , \nOut1_24[6] , \nOut1_24[5] , \nOut1_24[4] , 
        \nOut1_24[3] , \nOut1_24[2] , \nOut1_24[1] , \nOut1_24[0] }), .Out({
        \nOut2_24[7] , \nOut2_24[6] , \nOut2_24[5] , \nOut2_24[4] , 
        \nOut2_24[3] , \nOut2_24[2] , \nOut2_24[1] , \nOut2_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_155 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut156[7] , \nScanOut156[6] , 
        \nScanOut156[5] , \nScanOut156[4] , \nScanOut156[3] , \nScanOut156[2] , 
        \nScanOut156[1] , \nScanOut156[0] }), .ScanOut({\nScanOut155[7] , 
        \nScanOut155[6] , \nScanOut155[5] , \nScanOut155[4] , \nScanOut155[3] , 
        \nScanOut155[2] , \nScanOut155[1] , \nScanOut155[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_26[7] , \nOut4_26[6] , \nOut4_26[5] , \nOut4_26[4] , 
        \nOut4_26[3] , \nOut4_26[2] , \nOut4_26[1] , \nOut4_26[0] }), 
        .SouthIn({\nOut4_28[7] , \nOut4_28[6] , \nOut4_28[5] , \nOut4_28[4] , 
        \nOut4_28[3] , \nOut4_28[2] , \nOut4_28[1] , \nOut4_28[0] }), .EastIn(
        {\nOut5_27[7] , \nOut5_27[6] , \nOut5_27[5] , \nOut5_27[4] , 
        \nOut5_27[3] , \nOut5_27[2] , \nOut5_27[1] , \nOut5_27[0] }), .WestIn(
        {\nOut3_27[7] , \nOut3_27[6] , \nOut3_27[5] , \nOut3_27[4] , 
        \nOut3_27[3] , \nOut3_27[2] , \nOut3_27[1] , \nOut3_27[0] }), .Out({
        \nOut4_27[7] , \nOut4_27[6] , \nOut4_27[5] , \nOut4_27[4] , 
        \nOut4_27[3] , \nOut4_27[2] , \nOut4_27[1] , \nOut4_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_172 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut173[7] , \nScanOut173[6] , 
        \nScanOut173[5] , \nScanOut173[4] , \nScanOut173[3] , \nScanOut173[2] , 
        \nScanOut173[1] , \nScanOut173[0] }), .ScanOut({\nScanOut172[7] , 
        \nScanOut172[6] , \nScanOut172[5] , \nScanOut172[4] , \nScanOut172[3] , 
        \nScanOut172[2] , \nScanOut172[1] , \nScanOut172[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_11[7] , \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , 
        \nOut5_11[3] , \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }), 
        .SouthIn({\nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }), .EastIn(
        {\nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }), .WestIn(
        {\nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }), .Out({
        \nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_359 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut360[7] , \nScanOut360[6] , 
        \nScanOut360[5] , \nScanOut360[4] , \nScanOut360[3] , \nScanOut360[2] , 
        \nScanOut360[1] , \nScanOut360[0] }), .ScanOut({\nScanOut359[7] , 
        \nScanOut359[6] , \nScanOut359[5] , \nScanOut359[4] , \nScanOut359[3] , 
        \nScanOut359[2] , \nScanOut359[1] , \nScanOut359[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }), 
        .SouthIn({\nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }), .EastIn(
        {\nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }), .WestIn(
        {\nOut10_7[7] , \nOut10_7[6] , \nOut10_7[5] , \nOut10_7[4] , 
        \nOut10_7[3] , \nOut10_7[2] , \nOut10_7[1] , \nOut10_7[0] }), .Out({
        \nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_663 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut664[7] , \nScanOut664[6] , 
        \nScanOut664[5] , \nScanOut664[4] , \nScanOut664[3] , \nScanOut664[2] , 
        \nScanOut664[1] , \nScanOut664[0] }), .ScanOut({\nScanOut663[7] , 
        \nScanOut663[6] , \nScanOut663[5] , \nScanOut663[4] , \nScanOut663[3] , 
        \nScanOut663[2] , \nScanOut663[1] , \nScanOut663[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_22[7] , \nOut20_22[6] , \nOut20_22[5] , \nOut20_22[4] , 
        \nOut20_22[3] , \nOut20_22[2] , \nOut20_22[1] , \nOut20_22[0] }), 
        .SouthIn({\nOut20_24[7] , \nOut20_24[6] , \nOut20_24[5] , 
        \nOut20_24[4] , \nOut20_24[3] , \nOut20_24[2] , \nOut20_24[1] , 
        \nOut20_24[0] }), .EastIn({\nOut21_23[7] , \nOut21_23[6] , 
        \nOut21_23[5] , \nOut21_23[4] , \nOut21_23[3] , \nOut21_23[2] , 
        \nOut21_23[1] , \nOut21_23[0] }), .WestIn({\nOut19_23[7] , 
        \nOut19_23[6] , \nOut19_23[5] , \nOut19_23[4] , \nOut19_23[3] , 
        \nOut19_23[2] , \nOut19_23[1] , \nOut19_23[0] }), .Out({\nOut20_23[7] , 
        \nOut20_23[6] , \nOut20_23[5] , \nOut20_23[4] , \nOut20_23[3] , 
        \nOut20_23[2] , \nOut20_23[1] , \nOut20_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_678 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut679[7] , \nScanOut679[6] , 
        \nScanOut679[5] , \nScanOut679[4] , \nScanOut679[3] , \nScanOut679[2] , 
        \nScanOut679[1] , \nScanOut679[0] }), .ScanOut({\nScanOut678[7] , 
        \nScanOut678[6] , \nScanOut678[5] , \nScanOut678[4] , \nScanOut678[3] , 
        \nScanOut678[2] , \nScanOut678[1] , \nScanOut678[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_5[7] , \nOut21_5[6] , \nOut21_5[5] , \nOut21_5[4] , 
        \nOut21_5[3] , \nOut21_5[2] , \nOut21_5[1] , \nOut21_5[0] }), 
        .SouthIn({\nOut21_7[7] , \nOut21_7[6] , \nOut21_7[5] , \nOut21_7[4] , 
        \nOut21_7[3] , \nOut21_7[2] , \nOut21_7[1] , \nOut21_7[0] }), .EastIn(
        {\nOut22_6[7] , \nOut22_6[6] , \nOut22_6[5] , \nOut22_6[4] , 
        \nOut22_6[3] , \nOut22_6[2] , \nOut22_6[1] , \nOut22_6[0] }), .WestIn(
        {\nOut20_6[7] , \nOut20_6[6] , \nOut20_6[5] , \nOut20_6[4] , 
        \nOut20_6[3] , \nOut20_6[2] , \nOut20_6[1] , \nOut20_6[0] }), .Out({
        \nOut21_6[7] , \nOut21_6[6] , \nOut21_6[5] , \nOut21_6[4] , 
        \nOut21_6[3] , \nOut21_6[2] , \nOut21_6[1] , \nOut21_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_548 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut549[7] , \nScanOut549[6] , 
        \nScanOut549[5] , \nScanOut549[4] , \nScanOut549[3] , \nScanOut549[2] , 
        \nScanOut549[1] , \nScanOut549[0] }), .ScanOut({\nScanOut548[7] , 
        \nScanOut548[6] , \nScanOut548[5] , \nScanOut548[4] , \nScanOut548[3] , 
        \nScanOut548[2] , \nScanOut548[1] , \nScanOut548[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_3[7] , \nOut17_3[6] , \nOut17_3[5] , \nOut17_3[4] , 
        \nOut17_3[3] , \nOut17_3[2] , \nOut17_3[1] , \nOut17_3[0] }), 
        .SouthIn({\nOut17_5[7] , \nOut17_5[6] , \nOut17_5[5] , \nOut17_5[4] , 
        \nOut17_5[3] , \nOut17_5[2] , \nOut17_5[1] , \nOut17_5[0] }), .EastIn(
        {\nOut18_4[7] , \nOut18_4[6] , \nOut18_4[5] , \nOut18_4[4] , 
        \nOut18_4[3] , \nOut18_4[2] , \nOut18_4[1] , \nOut18_4[0] }), .WestIn(
        {\nOut16_4[7] , \nOut16_4[6] , \nOut16_4[5] , \nOut16_4[4] , 
        \nOut16_4[3] , \nOut16_4[2] , \nOut16_4[1] , \nOut16_4[0] }), .Out({
        \nOut17_4[7] , \nOut17_4[6] , \nOut17_4[5] , \nOut17_4[4] , 
        \nOut17_4[3] , \nOut17_4[2] , \nOut17_4[1] , \nOut17_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_763 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut764[7] , \nScanOut764[6] , 
        \nScanOut764[5] , \nScanOut764[4] , \nScanOut764[3] , \nScanOut764[2] , 
        \nScanOut764[1] , \nScanOut764[0] }), .ScanOut({\nScanOut763[7] , 
        \nScanOut763[6] , \nScanOut763[5] , \nScanOut763[4] , \nScanOut763[3] , 
        \nScanOut763[2] , \nScanOut763[1] , \nScanOut763[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_26[7] , \nOut23_26[6] , \nOut23_26[5] , \nOut23_26[4] , 
        \nOut23_26[3] , \nOut23_26[2] , \nOut23_26[1] , \nOut23_26[0] }), 
        .SouthIn({\nOut23_28[7] , \nOut23_28[6] , \nOut23_28[5] , 
        \nOut23_28[4] , \nOut23_28[3] , \nOut23_28[2] , \nOut23_28[1] , 
        \nOut23_28[0] }), .EastIn({\nOut24_27[7] , \nOut24_27[6] , 
        \nOut24_27[5] , \nOut24_27[4] , \nOut24_27[3] , \nOut24_27[2] , 
        \nOut24_27[1] , \nOut24_27[0] }), .WestIn({\nOut22_27[7] , 
        \nOut22_27[6] , \nOut22_27[5] , \nOut22_27[4] , \nOut22_27[3] , 
        \nOut22_27[2] , \nOut22_27[1] , \nOut22_27[0] }), .Out({\nOut23_27[7] , 
        \nOut23_27[6] , \nOut23_27[5] , \nOut23_27[4] , \nOut23_27[3] , 
        \nOut23_27[2] , \nOut23_27[1] , \nOut23_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_242 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut243[7] , \nScanOut243[6] , 
        \nScanOut243[5] , \nScanOut243[4] , \nScanOut243[3] , \nScanOut243[2] , 
        \nScanOut243[1] , \nScanOut243[0] }), .ScanOut({\nScanOut242[7] , 
        \nScanOut242[6] , \nScanOut242[5] , \nScanOut242[4] , \nScanOut242[3] , 
        \nScanOut242[2] , \nScanOut242[1] , \nScanOut242[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_17[7] , \nOut7_17[6] , \nOut7_17[5] , \nOut7_17[4] , 
        \nOut7_17[3] , \nOut7_17[2] , \nOut7_17[1] , \nOut7_17[0] }), 
        .SouthIn({\nOut7_19[7] , \nOut7_19[6] , \nOut7_19[5] , \nOut7_19[4] , 
        \nOut7_19[3] , \nOut7_19[2] , \nOut7_19[1] , \nOut7_19[0] }), .EastIn(
        {\nOut8_18[7] , \nOut8_18[6] , \nOut8_18[5] , \nOut8_18[4] , 
        \nOut8_18[3] , \nOut8_18[2] , \nOut8_18[1] , \nOut8_18[0] }), .WestIn(
        {\nOut6_18[7] , \nOut6_18[6] , \nOut6_18[5] , \nOut6_18[4] , 
        \nOut6_18[3] , \nOut6_18[2] , \nOut6_18[1] , \nOut6_18[0] }), .Out({
        \nOut7_18[7] , \nOut7_18[6] , \nOut7_18[5] , \nOut7_18[4] , 
        \nOut7_18[3] , \nOut7_18[2] , \nOut7_18[1] , \nOut7_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_453 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut454[7] , \nScanOut454[6] , 
        \nScanOut454[5] , \nScanOut454[4] , \nScanOut454[3] , \nScanOut454[2] , 
        \nScanOut454[1] , \nScanOut454[0] }), .ScanOut({\nScanOut453[7] , 
        \nScanOut453[6] , \nScanOut453[5] , \nScanOut453[4] , \nScanOut453[3] , 
        \nScanOut453[2] , \nScanOut453[1] , \nScanOut453[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }), 
        .SouthIn({\nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }), .EastIn(
        {\nOut15_5[7] , \nOut15_5[6] , \nOut15_5[5] , \nOut15_5[4] , 
        \nOut15_5[3] , \nOut15_5[2] , \nOut15_5[1] , \nOut15_5[0] }), .WestIn(
        {\nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }), .Out({
        \nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_265 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut266[7] , \nScanOut266[6] , 
        \nScanOut266[5] , \nScanOut266[4] , \nScanOut266[3] , \nScanOut266[2] , 
        \nScanOut266[1] , \nScanOut266[0] }), .ScanOut({\nScanOut265[7] , 
        \nScanOut265[6] , \nScanOut265[5] , \nScanOut265[4] , \nScanOut265[3] , 
        \nScanOut265[2] , \nScanOut265[1] , \nScanOut265[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_8[7] , \nOut8_8[6] , \nOut8_8[5] , \nOut8_8[4] , \nOut8_8[3] , 
        \nOut8_8[2] , \nOut8_8[1] , \nOut8_8[0] }), .SouthIn({\nOut8_10[7] , 
        \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , \nOut8_10[3] , 
        \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }), .EastIn({\nOut9_9[7] , 
        \nOut9_9[6] , \nOut9_9[5] , \nOut9_9[4] , \nOut9_9[3] , \nOut9_9[2] , 
        \nOut9_9[1] , \nOut9_9[0] }), .WestIn({\nOut7_9[7] , \nOut7_9[6] , 
        \nOut7_9[5] , \nOut7_9[4] , \nOut7_9[3] , \nOut7_9[2] , \nOut7_9[1] , 
        \nOut7_9[0] }), .Out({\nOut8_9[7] , \nOut8_9[6] , \nOut8_9[5] , 
        \nOut8_9[4] , \nOut8_9[3] , \nOut8_9[2] , \nOut8_9[1] , \nOut8_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_821 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut822[7] , \nScanOut822[6] , 
        \nScanOut822[5] , \nScanOut822[4] , \nScanOut822[3] , \nScanOut822[2] , 
        \nScanOut822[1] , \nScanOut822[0] }), .ScanOut({\nScanOut821[7] , 
        \nScanOut821[6] , \nScanOut821[5] , \nScanOut821[4] , \nScanOut821[3] , 
        \nScanOut821[2] , \nScanOut821[1] , \nScanOut821[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_20[7] , \nOut25_20[6] , \nOut25_20[5] , \nOut25_20[4] , 
        \nOut25_20[3] , \nOut25_20[2] , \nOut25_20[1] , \nOut25_20[0] }), 
        .SouthIn({\nOut25_22[7] , \nOut25_22[6] , \nOut25_22[5] , 
        \nOut25_22[4] , \nOut25_22[3] , \nOut25_22[2] , \nOut25_22[1] , 
        \nOut25_22[0] }), .EastIn({\nOut26_21[7] , \nOut26_21[6] , 
        \nOut26_21[5] , \nOut26_21[4] , \nOut26_21[3] , \nOut26_21[2] , 
        \nOut26_21[1] , \nOut26_21[0] }), .WestIn({\nOut24_21[7] , 
        \nOut24_21[6] , \nOut24_21[5] , \nOut24_21[4] , \nOut24_21[3] , 
        \nOut24_21[2] , \nOut24_21[1] , \nOut24_21[0] }), .Out({\nOut25_21[7] , 
        \nOut25_21[6] , \nOut25_21[5] , \nOut25_21[4] , \nOut25_21[3] , 
        \nOut25_21[2] , \nOut25_21[1] , \nOut25_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_474 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut475[7] , \nScanOut475[6] , 
        \nScanOut475[5] , \nScanOut475[4] , \nScanOut475[3] , \nScanOut475[2] , 
        \nScanOut475[1] , \nScanOut475[0] }), .ScanOut({\nScanOut474[7] , 
        \nScanOut474[6] , \nScanOut474[5] , \nScanOut474[4] , \nScanOut474[3] , 
        \nScanOut474[2] , \nScanOut474[1] , \nScanOut474[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_25[7] , \nOut14_25[6] , \nOut14_25[5] , \nOut14_25[4] , 
        \nOut14_25[3] , \nOut14_25[2] , \nOut14_25[1] , \nOut14_25[0] }), 
        .SouthIn({\nOut14_27[7] , \nOut14_27[6] , \nOut14_27[5] , 
        \nOut14_27[4] , \nOut14_27[3] , \nOut14_27[2] , \nOut14_27[1] , 
        \nOut14_27[0] }), .EastIn({\nOut15_26[7] , \nOut15_26[6] , 
        \nOut15_26[5] , \nOut15_26[4] , \nOut15_26[3] , \nOut15_26[2] , 
        \nOut15_26[1] , \nOut15_26[0] }), .WestIn({\nOut13_26[7] , 
        \nOut13_26[6] , \nOut13_26[5] , \nOut13_26[4] , \nOut13_26[3] , 
        \nOut13_26[2] , \nOut13_26[1] , \nOut13_26[0] }), .Out({\nOut14_26[7] , 
        \nOut14_26[6] , \nOut14_26[5] , \nOut14_26[4] , \nOut14_26[3] , 
        \nOut14_26[2] , \nOut14_26[1] , \nOut14_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_806 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut807[7] , \nScanOut807[6] , 
        \nScanOut807[5] , \nScanOut807[4] , \nScanOut807[3] , \nScanOut807[2] , 
        \nScanOut807[1] , \nScanOut807[0] }), .ScanOut({\nScanOut806[7] , 
        \nScanOut806[6] , \nScanOut806[5] , \nScanOut806[4] , \nScanOut806[3] , 
        \nScanOut806[2] , \nScanOut806[1] , \nScanOut806[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_5[7] , \nOut25_5[6] , \nOut25_5[5] , \nOut25_5[4] , 
        \nOut25_5[3] , \nOut25_5[2] , \nOut25_5[1] , \nOut25_5[0] }), 
        .SouthIn({\nOut25_7[7] , \nOut25_7[6] , \nOut25_7[5] , \nOut25_7[4] , 
        \nOut25_7[3] , \nOut25_7[2] , \nOut25_7[1] , \nOut25_7[0] }), .EastIn(
        {\nOut26_6[7] , \nOut26_6[6] , \nOut26_6[5] , \nOut26_6[4] , 
        \nOut26_6[3] , \nOut26_6[2] , \nOut26_6[1] , \nOut26_6[0] }), .WestIn(
        {\nOut24_6[7] , \nOut24_6[6] , \nOut24_6[5] , \nOut24_6[4] , 
        \nOut24_6[3] , \nOut24_6[2] , \nOut24_6[1] , \nOut24_6[0] }), .Out({
        \nOut25_6[7] , \nOut25_6[6] , \nOut25_6[5] , \nOut25_6[4] , 
        \nOut25_6[3] , \nOut25_6[2] , \nOut25_6[1] , \nOut25_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_996 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut997[7] , \nScanOut997[6] , 
        \nScanOut997[5] , \nScanOut997[4] , \nScanOut997[3] , \nScanOut997[2] , 
        \nScanOut997[1] , \nScanOut997[0] }), .ScanOut({\nScanOut996[7] , 
        \nScanOut996[6] , \nScanOut996[5] , \nScanOut996[4] , \nScanOut996[3] , 
        \nScanOut996[2] , \nScanOut996[1] , \nScanOut996[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut31_4[7] , \nOut31_4[6] , 
        \nOut31_4[5] , \nOut31_4[4] , \nOut31_4[3] , \nOut31_4[2] , 
        \nOut31_4[1] , \nOut31_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_744 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut745[7] , \nScanOut745[6] , 
        \nScanOut745[5] , \nScanOut745[4] , \nScanOut745[3] , \nScanOut745[2] , 
        \nScanOut745[1] , \nScanOut745[0] }), .ScanOut({\nScanOut744[7] , 
        \nScanOut744[6] , \nScanOut744[5] , \nScanOut744[4] , \nScanOut744[3] , 
        \nScanOut744[2] , \nScanOut744[1] , \nScanOut744[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_7[7] , \nOut23_7[6] , \nOut23_7[5] , \nOut23_7[4] , 
        \nOut23_7[3] , \nOut23_7[2] , \nOut23_7[1] , \nOut23_7[0] }), 
        .SouthIn({\nOut23_9[7] , \nOut23_9[6] , \nOut23_9[5] , \nOut23_9[4] , 
        \nOut23_9[3] , \nOut23_9[2] , \nOut23_9[1] , \nOut23_9[0] }), .EastIn(
        {\nOut24_8[7] , \nOut24_8[6] , \nOut24_8[5] , \nOut24_8[4] , 
        \nOut24_8[3] , \nOut24_8[2] , \nOut24_8[1] , \nOut24_8[0] }), .WestIn(
        {\nOut22_8[7] , \nOut22_8[6] , \nOut22_8[5] , \nOut22_8[4] , 
        \nOut22_8[3] , \nOut22_8[2] , \nOut22_8[1] , \nOut22_8[0] }), .Out({
        \nOut23_8[7] , \nOut23_8[6] , \nOut23_8[5] , \nOut23_8[4] , 
        \nOut23_8[3] , \nOut23_8[2] , \nOut23_8[1] , \nOut23_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_868 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut869[7] , \nScanOut869[6] , 
        \nScanOut869[5] , \nScanOut869[4] , \nScanOut869[3] , \nScanOut869[2] , 
        \nScanOut869[1] , \nScanOut869[0] }), .ScanOut({\nScanOut868[7] , 
        \nScanOut868[6] , \nScanOut868[5] , \nScanOut868[4] , \nScanOut868[3] , 
        \nScanOut868[2] , \nScanOut868[1] , \nScanOut868[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_3[7] , \nOut27_3[6] , \nOut27_3[5] , \nOut27_3[4] , 
        \nOut27_3[3] , \nOut27_3[2] , \nOut27_3[1] , \nOut27_3[0] }), 
        .SouthIn({\nOut27_5[7] , \nOut27_5[6] , \nOut27_5[5] , \nOut27_5[4] , 
        \nOut27_5[3] , \nOut27_5[2] , \nOut27_5[1] , \nOut27_5[0] }), .EastIn(
        {\nOut28_4[7] , \nOut28_4[6] , \nOut28_4[5] , \nOut28_4[4] , 
        \nOut28_4[3] , \nOut28_4[2] , \nOut28_4[1] , \nOut28_4[0] }), .WestIn(
        {\nOut26_4[7] , \nOut26_4[6] , \nOut26_4[5] , \nOut26_4[4] , 
        \nOut26_4[3] , \nOut26_4[2] , \nOut26_4[1] , \nOut26_4[0] }), .Out({
        \nOut27_4[7] , \nOut27_4[6] , \nOut27_4[5] , \nOut27_4[4] , 
        \nOut27_4[3] , \nOut27_4[2] , \nOut27_4[1] , \nOut27_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_280 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut281[7] , \nScanOut281[6] , 
        \nScanOut281[5] , \nScanOut281[4] , \nScanOut281[3] , \nScanOut281[2] , 
        \nScanOut281[1] , \nScanOut281[0] }), .ScanOut({\nScanOut280[7] , 
        \nScanOut280[6] , \nScanOut280[5] , \nScanOut280[4] , \nScanOut280[3] , 
        \nScanOut280[2] , \nScanOut280[1] , \nScanOut280[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_23[7] , \nOut8_23[6] , \nOut8_23[5] , \nOut8_23[4] , 
        \nOut8_23[3] , \nOut8_23[2] , \nOut8_23[1] , \nOut8_23[0] }), 
        .SouthIn({\nOut8_25[7] , \nOut8_25[6] , \nOut8_25[5] , \nOut8_25[4] , 
        \nOut8_25[3] , \nOut8_25[2] , \nOut8_25[1] , \nOut8_25[0] }), .EastIn(
        {\nOut9_24[7] , \nOut9_24[6] , \nOut9_24[5] , \nOut9_24[4] , 
        \nOut9_24[3] , \nOut9_24[2] , \nOut9_24[1] , \nOut9_24[0] }), .WestIn(
        {\nOut7_24[7] , \nOut7_24[6] , \nOut7_24[5] , \nOut7_24[4] , 
        \nOut7_24[3] , \nOut7_24[2] , \nOut7_24[1] , \nOut7_24[0] }), .Out({
        \nOut8_24[7] , \nOut8_24[6] , \nOut8_24[5] , \nOut8_24[4] , 
        \nOut8_24[3] , \nOut8_24[2] , \nOut8_24[1] , \nOut8_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_310 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut311[7] , \nScanOut311[6] , 
        \nScanOut311[5] , \nScanOut311[4] , \nScanOut311[3] , \nScanOut311[2] , 
        \nScanOut311[1] , \nScanOut311[0] }), .ScanOut({\nScanOut310[7] , 
        \nScanOut310[6] , \nScanOut310[5] , \nScanOut310[4] , \nScanOut310[3] , 
        \nScanOut310[2] , \nScanOut310[1] , \nScanOut310[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_21[7] , \nOut9_21[6] , \nOut9_21[5] , \nOut9_21[4] , 
        \nOut9_21[3] , \nOut9_21[2] , \nOut9_21[1] , \nOut9_21[0] }), 
        .SouthIn({\nOut9_23[7] , \nOut9_23[6] , \nOut9_23[5] , \nOut9_23[4] , 
        \nOut9_23[3] , \nOut9_23[2] , \nOut9_23[1] , \nOut9_23[0] }), .EastIn(
        {\nOut10_22[7] , \nOut10_22[6] , \nOut10_22[5] , \nOut10_22[4] , 
        \nOut10_22[3] , \nOut10_22[2] , \nOut10_22[1] , \nOut10_22[0] }), 
        .WestIn({\nOut8_22[7] , \nOut8_22[6] , \nOut8_22[5] , \nOut8_22[4] , 
        \nOut8_22[3] , \nOut8_22[2] , \nOut8_22[1] , \nOut8_22[0] }), .Out({
        \nOut9_22[7] , \nOut9_22[6] , \nOut9_22[5] , \nOut9_22[4] , 
        \nOut9_22[3] , \nOut9_22[2] , \nOut9_22[1] , \nOut9_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_491 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut492[7] , \nScanOut492[6] , 
        \nScanOut492[5] , \nScanOut492[4] , \nScanOut492[3] , \nScanOut492[2] , 
        \nScanOut492[1] , \nScanOut492[0] }), .ScanOut({\nScanOut491[7] , 
        \nScanOut491[6] , \nScanOut491[5] , \nScanOut491[4] , \nScanOut491[3] , 
        \nScanOut491[2] , \nScanOut491[1] , \nScanOut491[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_10[7] , \nOut15_10[6] , \nOut15_10[5] , \nOut15_10[4] , 
        \nOut15_10[3] , \nOut15_10[2] , \nOut15_10[1] , \nOut15_10[0] }), 
        .SouthIn({\nOut15_12[7] , \nOut15_12[6] , \nOut15_12[5] , 
        \nOut15_12[4] , \nOut15_12[3] , \nOut15_12[2] , \nOut15_12[1] , 
        \nOut15_12[0] }), .EastIn({\nOut16_11[7] , \nOut16_11[6] , 
        \nOut16_11[5] , \nOut16_11[4] , \nOut16_11[3] , \nOut16_11[2] , 
        \nOut16_11[1] , \nOut16_11[0] }), .WestIn({\nOut14_11[7] , 
        \nOut14_11[6] , \nOut14_11[5] , \nOut14_11[4] , \nOut14_11[3] , 
        \nOut14_11[2] , \nOut14_11[1] , \nOut14_11[0] }), .Out({\nOut15_11[7] , 
        \nOut15_11[6] , \nOut15_11[5] , \nOut15_11[4] , \nOut15_11[3] , 
        \nOut15_11[2] , \nOut15_11[1] , \nOut15_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_501 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut502[7] , \nScanOut502[6] , 
        \nScanOut502[5] , \nScanOut502[4] , \nScanOut502[3] , \nScanOut502[2] , 
        \nScanOut502[1] , \nScanOut502[0] }), .ScanOut({\nScanOut501[7] , 
        \nScanOut501[6] , \nScanOut501[5] , \nScanOut501[4] , \nScanOut501[3] , 
        \nScanOut501[2] , \nScanOut501[1] , \nScanOut501[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_20[7] , \nOut15_20[6] , \nOut15_20[5] , \nOut15_20[4] , 
        \nOut15_20[3] , \nOut15_20[2] , \nOut15_20[1] , \nOut15_20[0] }), 
        .SouthIn({\nOut15_22[7] , \nOut15_22[6] , \nOut15_22[5] , 
        \nOut15_22[4] , \nOut15_22[3] , \nOut15_22[2] , \nOut15_22[1] , 
        \nOut15_22[0] }), .EastIn({\nOut16_21[7] , \nOut16_21[6] , 
        \nOut16_21[5] , \nOut16_21[4] , \nOut16_21[3] , \nOut16_21[2] , 
        \nOut16_21[1] , \nOut16_21[0] }), .WestIn({\nOut14_21[7] , 
        \nOut14_21[6] , \nOut14_21[5] , \nOut14_21[4] , \nOut14_21[3] , 
        \nOut14_21[2] , \nOut14_21[1] , \nOut14_21[0] }), .Out({\nOut15_21[7] , 
        \nOut15_21[6] , \nOut15_21[5] , \nOut15_21[4] , \nOut15_21[3] , 
        \nOut15_21[2] , \nOut15_21[1] , \nOut15_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_631 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut632[7] , \nScanOut632[6] , 
        \nScanOut632[5] , \nScanOut632[4] , \nScanOut632[3] , \nScanOut632[2] , 
        \nScanOut632[1] , \nScanOut632[0] }), .ScanOut({\nScanOut631[7] , 
        \nScanOut631[6] , \nScanOut631[5] , \nScanOut631[4] , \nScanOut631[3] , 
        \nScanOut631[2] , \nScanOut631[1] , \nScanOut631[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_22[7] , \nOut19_22[6] , \nOut19_22[5] , \nOut19_22[4] , 
        \nOut19_22[3] , \nOut19_22[2] , \nOut19_22[1] , \nOut19_22[0] }), 
        .SouthIn({\nOut19_24[7] , \nOut19_24[6] , \nOut19_24[5] , 
        \nOut19_24[4] , \nOut19_24[3] , \nOut19_24[2] , \nOut19_24[1] , 
        \nOut19_24[0] }), .EastIn({\nOut20_23[7] , \nOut20_23[6] , 
        \nOut20_23[5] , \nOut20_23[4] , \nOut20_23[3] , \nOut20_23[2] , 
        \nOut20_23[1] , \nOut20_23[0] }), .WestIn({\nOut18_23[7] , 
        \nOut18_23[6] , \nOut18_23[5] , \nOut18_23[4] , \nOut18_23[3] , 
        \nOut18_23[2] , \nOut18_23[1] , \nOut18_23[0] }), .Out({\nOut19_23[7] , 
        \nOut19_23[6] , \nOut19_23[5] , \nOut19_23[4] , \nOut19_23[3] , 
        \nOut19_23[2] , \nOut19_23[1] , \nOut19_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_973 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut974[7] , \nScanOut974[6] , 
        \nScanOut974[5] , \nScanOut974[4] , \nScanOut974[3] , \nScanOut974[2] , 
        \nScanOut974[1] , \nScanOut974[0] }), .ScanOut({\nScanOut973[7] , 
        \nScanOut973[6] , \nScanOut973[5] , \nScanOut973[4] , \nScanOut973[3] , 
        \nScanOut973[2] , \nScanOut973[1] , \nScanOut973[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_12[7] , \nOut30_12[6] , \nOut30_12[5] , \nOut30_12[4] , 
        \nOut30_12[3] , \nOut30_12[2] , \nOut30_12[1] , \nOut30_12[0] }), 
        .SouthIn({\nOut30_14[7] , \nOut30_14[6] , \nOut30_14[5] , 
        \nOut30_14[4] , \nOut30_14[3] , \nOut30_14[2] , \nOut30_14[1] , 
        \nOut30_14[0] }), .EastIn({\nOut31_13[7] , \nOut31_13[6] , 
        \nOut31_13[5] , \nOut31_13[4] , \nOut31_13[3] , \nOut31_13[2] , 
        \nOut31_13[1] , \nOut31_13[0] }), .WestIn({\nOut29_13[7] , 
        \nOut29_13[6] , \nOut29_13[5] , \nOut29_13[4] , \nOut29_13[3] , 
        \nOut29_13[2] , \nOut29_13[1] , \nOut29_13[0] }), .Out({\nOut30_13[7] , 
        \nOut30_13[6] , \nOut30_13[5] , \nOut30_13[4] , \nOut30_13[3] , 
        \nOut30_13[2] , \nOut30_13[1] , \nOut30_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_36 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut37[7] , \nScanOut37[6] , 
        \nScanOut37[5] , \nScanOut37[4] , \nScanOut37[3] , \nScanOut37[2] , 
        \nScanOut37[1] , \nScanOut37[0] }), .ScanOut({\nScanOut36[7] , 
        \nScanOut36[6] , \nScanOut36[5] , \nScanOut36[4] , \nScanOut36[3] , 
        \nScanOut36[2] , \nScanOut36[1] , \nScanOut36[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , \nOut1_3[3] , 
        \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }), .SouthIn({\nOut1_5[7] , 
        \nOut1_5[6] , \nOut1_5[5] , \nOut1_5[4] , \nOut1_5[3] , \nOut1_5[2] , 
        \nOut1_5[1] , \nOut1_5[0] }), .EastIn({\nOut2_4[7] , \nOut2_4[6] , 
        \nOut2_4[5] , \nOut2_4[4] , \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , 
        \nOut2_4[0] }), .WestIn({\nOut0_4[7] , \nOut0_4[6] , \nOut0_4[5] , 
        \nOut0_4[4] , \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , \nOut0_4[0] }), 
        .Out({\nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , \nOut1_4[4] , 
        \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_197 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut198[7] , \nScanOut198[6] , 
        \nScanOut198[5] , \nScanOut198[4] , \nScanOut198[3] , \nScanOut198[2] , 
        \nScanOut198[1] , \nScanOut198[0] }), .ScanOut({\nScanOut197[7] , 
        \nScanOut197[6] , \nScanOut197[5] , \nScanOut197[4] , \nScanOut197[3] , 
        \nScanOut197[2] , \nScanOut197[1] , \nScanOut197[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_4[7] , \nOut6_4[6] , \nOut6_4[5] , \nOut6_4[4] , \nOut6_4[3] , 
        \nOut6_4[2] , \nOut6_4[1] , \nOut6_4[0] }), .SouthIn({\nOut6_6[7] , 
        \nOut6_6[6] , \nOut6_6[5] , \nOut6_6[4] , \nOut6_6[3] , \nOut6_6[2] , 
        \nOut6_6[1] , \nOut6_6[0] }), .EastIn({\nOut7_5[7] , \nOut7_5[6] , 
        \nOut7_5[5] , \nOut7_5[4] , \nOut7_5[3] , \nOut7_5[2] , \nOut7_5[1] , 
        \nOut7_5[0] }), .WestIn({\nOut5_5[7] , \nOut5_5[6] , \nOut5_5[5] , 
        \nOut5_5[4] , \nOut5_5[3] , \nOut5_5[2] , \nOut5_5[1] , \nOut5_5[0] }), 
        .Out({\nOut6_5[7] , \nOut6_5[6] , \nOut6_5[5] , \nOut6_5[4] , 
        \nOut6_5[3] , \nOut6_5[2] , \nOut6_5[1] , \nOut6_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_616 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut617[7] , \nScanOut617[6] , 
        \nScanOut617[5] , \nScanOut617[4] , \nScanOut617[3] , \nScanOut617[2] , 
        \nScanOut617[1] , \nScanOut617[0] }), .ScanOut({\nScanOut616[7] , 
        \nScanOut616[6] , \nScanOut616[5] , \nScanOut616[4] , \nScanOut616[3] , 
        \nScanOut616[2] , \nScanOut616[1] , \nScanOut616[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_7[7] , \nOut19_7[6] , \nOut19_7[5] , \nOut19_7[4] , 
        \nOut19_7[3] , \nOut19_7[2] , \nOut19_7[1] , \nOut19_7[0] }), 
        .SouthIn({\nOut19_9[7] , \nOut19_9[6] , \nOut19_9[5] , \nOut19_9[4] , 
        \nOut19_9[3] , \nOut19_9[2] , \nOut19_9[1] , \nOut19_9[0] }), .EastIn(
        {\nOut20_8[7] , \nOut20_8[6] , \nOut20_8[5] , \nOut20_8[4] , 
        \nOut20_8[3] , \nOut20_8[2] , \nOut20_8[1] , \nOut20_8[0] }), .WestIn(
        {\nOut18_8[7] , \nOut18_8[6] , \nOut18_8[5] , \nOut18_8[4] , 
        \nOut18_8[3] , \nOut18_8[2] , \nOut18_8[1] , \nOut18_8[0] }), .Out({
        \nOut19_8[7] , \nOut19_8[6] , \nOut19_8[5] , \nOut19_8[4] , 
        \nOut19_8[3] , \nOut19_8[2] , \nOut19_8[1] , \nOut19_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_292 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut293[7] , \nScanOut293[6] , 
        \nScanOut293[5] , \nScanOut293[4] , \nScanOut293[3] , \nScanOut293[2] , 
        \nScanOut293[1] , \nScanOut293[0] }), .ScanOut({\nScanOut292[7] , 
        \nScanOut292[6] , \nScanOut292[5] , \nScanOut292[4] , \nScanOut292[3] , 
        \nScanOut292[2] , \nScanOut292[1] , \nScanOut292[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_3[7] , \nOut9_3[6] , \nOut9_3[5] , \nOut9_3[4] , \nOut9_3[3] , 
        \nOut9_3[2] , \nOut9_3[1] , \nOut9_3[0] }), .SouthIn({\nOut9_5[7] , 
        \nOut9_5[6] , \nOut9_5[5] , \nOut9_5[4] , \nOut9_5[3] , \nOut9_5[2] , 
        \nOut9_5[1] , \nOut9_5[0] }), .EastIn({\nOut10_4[7] , \nOut10_4[6] , 
        \nOut10_4[5] , \nOut10_4[4] , \nOut10_4[3] , \nOut10_4[2] , 
        \nOut10_4[1] , \nOut10_4[0] }), .WestIn({\nOut8_4[7] , \nOut8_4[6] , 
        \nOut8_4[5] , \nOut8_4[4] , \nOut8_4[3] , \nOut8_4[2] , \nOut8_4[1] , 
        \nOut8_4[0] }), .Out({\nOut9_4[7] , \nOut9_4[6] , \nOut9_4[5] , 
        \nOut9_4[4] , \nOut9_4[3] , \nOut9_4[2] , \nOut9_4[1] , \nOut9_4[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_337 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut338[7] , \nScanOut338[6] , 
        \nScanOut338[5] , \nScanOut338[4] , \nScanOut338[3] , \nScanOut338[2] , 
        \nScanOut338[1] , \nScanOut338[0] }), .ScanOut({\nScanOut337[7] , 
        \nScanOut337[6] , \nScanOut337[5] , \nScanOut337[4] , \nScanOut337[3] , 
        \nScanOut337[2] , \nScanOut337[1] , \nScanOut337[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_16[7] , \nOut10_16[6] , \nOut10_16[5] , \nOut10_16[4] , 
        \nOut10_16[3] , \nOut10_16[2] , \nOut10_16[1] , \nOut10_16[0] }), 
        .SouthIn({\nOut10_18[7] , \nOut10_18[6] , \nOut10_18[5] , 
        \nOut10_18[4] , \nOut10_18[3] , \nOut10_18[2] , \nOut10_18[1] , 
        \nOut10_18[0] }), .EastIn({\nOut11_17[7] , \nOut11_17[6] , 
        \nOut11_17[5] , \nOut11_17[4] , \nOut11_17[3] , \nOut11_17[2] , 
        \nOut11_17[1] , \nOut11_17[0] }), .WestIn({\nOut9_17[7] , 
        \nOut9_17[6] , \nOut9_17[5] , \nOut9_17[4] , \nOut9_17[3] , 
        \nOut9_17[2] , \nOut9_17[1] , \nOut9_17[0] }), .Out({\nOut10_17[7] , 
        \nOut10_17[6] , \nOut10_17[5] , \nOut10_17[4] , \nOut10_17[3] , 
        \nOut10_17[2] , \nOut10_17[1] , \nOut10_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_526 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut527[7] , \nScanOut527[6] , 
        \nScanOut527[5] , \nScanOut527[4] , \nScanOut527[3] , \nScanOut527[2] , 
        \nScanOut527[1] , \nScanOut527[0] }), .ScanOut({\nScanOut526[7] , 
        \nScanOut526[6] , \nScanOut526[5] , \nScanOut526[4] , \nScanOut526[3] , 
        \nScanOut526[2] , \nScanOut526[1] , \nScanOut526[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_13[7] , \nOut16_13[6] , \nOut16_13[5] , \nOut16_13[4] , 
        \nOut16_13[3] , \nOut16_13[2] , \nOut16_13[1] , \nOut16_13[0] }), 
        .SouthIn({\nOut16_15[7] , \nOut16_15[6] , \nOut16_15[5] , 
        \nOut16_15[4] , \nOut16_15[3] , \nOut16_15[2] , \nOut16_15[1] , 
        \nOut16_15[0] }), .EastIn({\nOut17_14[7] , \nOut17_14[6] , 
        \nOut17_14[5] , \nOut17_14[4] , \nOut17_14[3] , \nOut17_14[2] , 
        \nOut17_14[1] , \nOut17_14[0] }), .WestIn({\nOut15_14[7] , 
        \nOut15_14[6] , \nOut15_14[5] , \nOut15_14[4] , \nOut15_14[3] , 
        \nOut15_14[2] , \nOut15_14[1] , \nOut15_14[0] }), .Out({\nOut16_14[7] , 
        \nOut16_14[6] , \nOut16_14[5] , \nOut16_14[4] , \nOut16_14[3] , 
        \nOut16_14[2] , \nOut16_14[1] , \nOut16_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_786 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut787[7] , \nScanOut787[6] , 
        \nScanOut787[5] , \nScanOut787[4] , \nScanOut787[3] , \nScanOut787[2] , 
        \nScanOut787[1] , \nScanOut787[0] }), .ScanOut({\nScanOut786[7] , 
        \nScanOut786[6] , \nScanOut786[5] , \nScanOut786[4] , \nScanOut786[3] , 
        \nScanOut786[2] , \nScanOut786[1] , \nScanOut786[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_17[7] , \nOut24_17[6] , \nOut24_17[5] , \nOut24_17[4] , 
        \nOut24_17[3] , \nOut24_17[2] , \nOut24_17[1] , \nOut24_17[0] }), 
        .SouthIn({\nOut24_19[7] , \nOut24_19[6] , \nOut24_19[5] , 
        \nOut24_19[4] , \nOut24_19[3] , \nOut24_19[2] , \nOut24_19[1] , 
        \nOut24_19[0] }), .EastIn({\nOut25_18[7] , \nOut25_18[6] , 
        \nOut25_18[5] , \nOut25_18[4] , \nOut25_18[3] , \nOut25_18[2] , 
        \nOut25_18[1] , \nOut25_18[0] }), .WestIn({\nOut23_18[7] , 
        \nOut23_18[6] , \nOut23_18[5] , \nOut23_18[4] , \nOut23_18[3] , 
        \nOut23_18[2] , \nOut23_18[1] , \nOut23_18[0] }), .Out({\nOut24_18[7] , 
        \nOut24_18[6] , \nOut24_18[5] , \nOut24_18[4] , \nOut24_18[3] , 
        \nOut24_18[2] , \nOut24_18[1] , \nOut24_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_954 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut955[7] , \nScanOut955[6] , 
        \nScanOut955[5] , \nScanOut955[4] , \nScanOut955[3] , \nScanOut955[2] , 
        \nScanOut955[1] , \nScanOut955[0] }), .ScanOut({\nScanOut954[7] , 
        \nScanOut954[6] , \nScanOut954[5] , \nScanOut954[4] , \nScanOut954[3] , 
        \nScanOut954[2] , \nScanOut954[1] , \nScanOut954[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_25[7] , \nOut29_25[6] , \nOut29_25[5] , \nOut29_25[4] , 
        \nOut29_25[3] , \nOut29_25[2] , \nOut29_25[1] , \nOut29_25[0] }), 
        .SouthIn({\nOut29_27[7] , \nOut29_27[6] , \nOut29_27[5] , 
        \nOut29_27[4] , \nOut29_27[3] , \nOut29_27[2] , \nOut29_27[1] , 
        \nOut29_27[0] }), .EastIn({\nOut30_26[7] , \nOut30_26[6] , 
        \nOut30_26[5] , \nOut30_26[4] , \nOut30_26[3] , \nOut30_26[2] , 
        \nOut30_26[1] , \nOut30_26[0] }), .WestIn({\nOut28_26[7] , 
        \nOut28_26[6] , \nOut28_26[5] , \nOut28_26[4] , \nOut28_26[3] , 
        \nOut28_26[2] , \nOut28_26[1] , \nOut28_26[0] }), .Out({\nOut29_26[7] , 
        \nOut29_26[6] , \nOut29_26[5] , \nOut29_26[4] , \nOut29_26[3] , 
        \nOut29_26[2] , \nOut29_26[1] , \nOut29_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_961 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut962[7] , \nScanOut962[6] , 
        \nScanOut962[5] , \nScanOut962[4] , \nScanOut962[3] , \nScanOut962[2] , 
        \nScanOut962[1] , \nScanOut962[0] }), .ScanOut({\nScanOut961[7] , 
        \nScanOut961[6] , \nScanOut961[5] , \nScanOut961[4] , \nScanOut961[3] , 
        \nScanOut961[2] , \nScanOut961[1] , \nScanOut961[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_0[7] , \nOut30_0[6] , \nOut30_0[5] , \nOut30_0[4] , 
        \nOut30_0[3] , \nOut30_0[2] , \nOut30_0[1] , \nOut30_0[0] }), 
        .SouthIn({\nOut30_2[7] , \nOut30_2[6] , \nOut30_2[5] , \nOut30_2[4] , 
        \nOut30_2[3] , \nOut30_2[2] , \nOut30_2[1] , \nOut30_2[0] }), .EastIn(
        {\nOut31_1[7] , \nOut31_1[6] , \nOut31_1[5] , \nOut31_1[4] , 
        \nOut31_1[3] , \nOut31_1[2] , \nOut31_1[1] , \nOut31_1[0] }), .WestIn(
        {\nOut29_1[7] , \nOut29_1[6] , \nOut29_1[5] , \nOut29_1[4] , 
        \nOut29_1[3] , \nOut29_1[2] , \nOut29_1[1] , \nOut29_1[0] }), .Out({
        \nOut30_1[7] , \nOut30_1[6] , \nOut30_1[5] , \nOut30_1[4] , 
        \nOut30_1[3] , \nOut30_1[2] , \nOut30_1[1] , \nOut30_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_302 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut303[7] , \nScanOut303[6] , 
        \nScanOut303[5] , \nScanOut303[4] , \nScanOut303[3] , \nScanOut303[2] , 
        \nScanOut303[1] , \nScanOut303[0] }), .ScanOut({\nScanOut302[7] , 
        \nScanOut302[6] , \nScanOut302[5] , \nScanOut302[4] , \nScanOut302[3] , 
        \nScanOut302[2] , \nScanOut302[1] , \nScanOut302[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_13[7] , \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , 
        \nOut9_13[3] , \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }), 
        .SouthIn({\nOut9_15[7] , \nOut9_15[6] , \nOut9_15[5] , \nOut9_15[4] , 
        \nOut9_15[3] , \nOut9_15[2] , \nOut9_15[1] , \nOut9_15[0] }), .EastIn(
        {\nOut10_14[7] , \nOut10_14[6] , \nOut10_14[5] , \nOut10_14[4] , 
        \nOut10_14[3] , \nOut10_14[2] , \nOut10_14[1] , \nOut10_14[0] }), 
        .WestIn({\nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }), .Out({
        \nOut9_14[7] , \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , 
        \nOut9_14[3] , \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_513 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut514[7] , \nScanOut514[6] , 
        \nScanOut514[5] , \nScanOut514[4] , \nScanOut514[3] , \nScanOut514[2] , 
        \nScanOut514[1] , \nScanOut514[0] }), .ScanOut({\nScanOut513[7] , 
        \nScanOut513[6] , \nScanOut513[5] , \nScanOut513[4] , \nScanOut513[3] , 
        \nScanOut513[2] , \nScanOut513[1] , \nScanOut513[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_0[7] , \nOut16_0[6] , \nOut16_0[5] , \nOut16_0[4] , 
        \nOut16_0[3] , \nOut16_0[2] , \nOut16_0[1] , \nOut16_0[0] }), 
        .SouthIn({\nOut16_2[7] , \nOut16_2[6] , \nOut16_2[5] , \nOut16_2[4] , 
        \nOut16_2[3] , \nOut16_2[2] , \nOut16_2[1] , \nOut16_2[0] }), .EastIn(
        {\nOut17_1[7] , \nOut17_1[6] , \nOut17_1[5] , \nOut17_1[4] , 
        \nOut17_1[3] , \nOut17_1[2] , \nOut17_1[1] , \nOut17_1[0] }), .WestIn(
        {\nOut15_1[7] , \nOut15_1[6] , \nOut15_1[5] , \nOut15_1[4] , 
        \nOut15_1[3] , \nOut15_1[2] , \nOut15_1[1] , \nOut15_1[0] }), .Out({
        \nOut16_1[7] , \nOut16_1[6] , \nOut16_1[5] , \nOut16_1[4] , 
        \nOut16_1[3] , \nOut16_1[2] , \nOut16_1[1] , \nOut16_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_483 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut484[7] , \nScanOut484[6] , 
        \nScanOut484[5] , \nScanOut484[4] , \nScanOut484[3] , \nScanOut484[2] , 
        \nScanOut484[1] , \nScanOut484[0] }), .ScanOut({\nScanOut483[7] , 
        \nScanOut483[6] , \nScanOut483[5] , \nScanOut483[4] , \nScanOut483[3] , 
        \nScanOut483[2] , \nScanOut483[1] , \nScanOut483[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_2[7] , \nOut15_2[6] , \nOut15_2[5] , \nOut15_2[4] , 
        \nOut15_2[3] , \nOut15_2[2] , \nOut15_2[1] , \nOut15_2[0] }), 
        .SouthIn({\nOut15_4[7] , \nOut15_4[6] , \nOut15_4[5] , \nOut15_4[4] , 
        \nOut15_4[3] , \nOut15_4[2] , \nOut15_4[1] , \nOut15_4[0] }), .EastIn(
        {\nOut16_3[7] , \nOut16_3[6] , \nOut16_3[5] , \nOut16_3[4] , 
        \nOut16_3[3] , \nOut16_3[2] , \nOut16_3[1] , \nOut16_3[0] }), .WestIn(
        {\nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }), .Out({
        \nOut15_3[7] , \nOut15_3[6] , \nOut15_3[5] , \nOut15_3[4] , 
        \nOut15_3[3] , \nOut15_3[2] , \nOut15_3[1] , \nOut15_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_623 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut624[7] , \nScanOut624[6] , 
        \nScanOut624[5] , \nScanOut624[4] , \nScanOut624[3] , \nScanOut624[2] , 
        \nScanOut624[1] , \nScanOut624[0] }), .ScanOut({\nScanOut623[7] , 
        \nScanOut623[6] , \nScanOut623[5] , \nScanOut623[4] , \nScanOut623[3] , 
        \nScanOut623[2] , \nScanOut623[1] , \nScanOut623[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_14[7] , \nOut19_14[6] , \nOut19_14[5] , \nOut19_14[4] , 
        \nOut19_14[3] , \nOut19_14[2] , \nOut19_14[1] , \nOut19_14[0] }), 
        .SouthIn({\nOut19_16[7] , \nOut19_16[6] , \nOut19_16[5] , 
        \nOut19_16[4] , \nOut19_16[3] , \nOut19_16[2] , \nOut19_16[1] , 
        \nOut19_16[0] }), .EastIn({\nOut20_15[7] , \nOut20_15[6] , 
        \nOut20_15[5] , \nOut20_15[4] , \nOut20_15[3] , \nOut20_15[2] , 
        \nOut20_15[1] , \nOut20_15[0] }), .WestIn({\nOut18_15[7] , 
        \nOut18_15[6] , \nOut18_15[5] , \nOut18_15[4] , \nOut18_15[3] , 
        \nOut18_15[2] , \nOut18_15[1] , \nOut18_15[0] }), .Out({\nOut19_15[7] , 
        \nOut19_15[6] , \nOut19_15[5] , \nOut19_15[4] , \nOut19_15[3] , 
        \nOut19_15[2] , \nOut19_15[1] , \nOut19_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_185 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut186[7] , \nScanOut186[6] , 
        \nScanOut186[5] , \nScanOut186[4] , \nScanOut186[3] , \nScanOut186[2] , 
        \nScanOut186[1] , \nScanOut186[0] }), .ScanOut({\nScanOut185[7] , 
        \nScanOut185[6] , \nScanOut185[5] , \nScanOut185[4] , \nScanOut185[3] , 
        \nScanOut185[2] , \nScanOut185[1] , \nScanOut185[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_24[7] , \nOut5_24[6] , \nOut5_24[5] , \nOut5_24[4] , 
        \nOut5_24[3] , \nOut5_24[2] , \nOut5_24[1] , \nOut5_24[0] }), 
        .SouthIn({\nOut5_26[7] , \nOut5_26[6] , \nOut5_26[5] , \nOut5_26[4] , 
        \nOut5_26[3] , \nOut5_26[2] , \nOut5_26[1] , \nOut5_26[0] }), .EastIn(
        {\nOut6_25[7] , \nOut6_25[6] , \nOut6_25[5] , \nOut6_25[4] , 
        \nOut6_25[3] , \nOut6_25[2] , \nOut6_25[1] , \nOut6_25[0] }), .WestIn(
        {\nOut4_25[7] , \nOut4_25[6] , \nOut4_25[5] , \nOut4_25[4] , 
        \nOut4_25[3] , \nOut4_25[2] , \nOut4_25[1] , \nOut4_25[0] }), .Out({
        \nOut5_25[7] , \nOut5_25[6] , \nOut5_25[5] , \nOut5_25[4] , 
        \nOut5_25[3] , \nOut5_25[2] , \nOut5_25[1] , \nOut5_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_604 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut605[7] , \nScanOut605[6] , 
        \nScanOut605[5] , \nScanOut605[4] , \nScanOut605[3] , \nScanOut605[2] , 
        \nScanOut605[1] , \nScanOut605[0] }), .ScanOut({\nScanOut604[7] , 
        \nScanOut604[6] , \nScanOut604[5] , \nScanOut604[4] , \nScanOut604[3] , 
        \nScanOut604[2] , \nScanOut604[1] , \nScanOut604[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_27[7] , \nOut18_27[6] , \nOut18_27[5] , \nOut18_27[4] , 
        \nOut18_27[3] , \nOut18_27[2] , \nOut18_27[1] , \nOut18_27[0] }), 
        .SouthIn({\nOut18_29[7] , \nOut18_29[6] , \nOut18_29[5] , 
        \nOut18_29[4] , \nOut18_29[3] , \nOut18_29[2] , \nOut18_29[1] , 
        \nOut18_29[0] }), .EastIn({\nOut19_28[7] , \nOut19_28[6] , 
        \nOut19_28[5] , \nOut19_28[4] , \nOut19_28[3] , \nOut19_28[2] , 
        \nOut19_28[1] , \nOut19_28[0] }), .WestIn({\nOut17_28[7] , 
        \nOut17_28[6] , \nOut17_28[5] , \nOut17_28[4] , \nOut17_28[3] , 
        \nOut17_28[2] , \nOut17_28[1] , \nOut17_28[0] }), .Out({\nOut18_28[7] , 
        \nOut18_28[6] , \nOut18_28[5] , \nOut18_28[4] , \nOut18_28[3] , 
        \nOut18_28[2] , \nOut18_28[1] , \nOut18_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_794 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut795[7] , \nScanOut795[6] , 
        \nScanOut795[5] , \nScanOut795[4] , \nScanOut795[3] , \nScanOut795[2] , 
        \nScanOut795[1] , \nScanOut795[0] }), .ScanOut({\nScanOut794[7] , 
        \nScanOut794[6] , \nScanOut794[5] , \nScanOut794[4] , \nScanOut794[3] , 
        \nScanOut794[2] , \nScanOut794[1] , \nScanOut794[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_25[7] , \nOut24_25[6] , \nOut24_25[5] , \nOut24_25[4] , 
        \nOut24_25[3] , \nOut24_25[2] , \nOut24_25[1] , \nOut24_25[0] }), 
        .SouthIn({\nOut24_27[7] , \nOut24_27[6] , \nOut24_27[5] , 
        \nOut24_27[4] , \nOut24_27[3] , \nOut24_27[2] , \nOut24_27[1] , 
        \nOut24_27[0] }), .EastIn({\nOut25_26[7] , \nOut25_26[6] , 
        \nOut25_26[5] , \nOut25_26[4] , \nOut25_26[3] , \nOut25_26[2] , 
        \nOut25_26[1] , \nOut25_26[0] }), .WestIn({\nOut23_26[7] , 
        \nOut23_26[6] , \nOut23_26[5] , \nOut23_26[4] , \nOut23_26[3] , 
        \nOut23_26[2] , \nOut23_26[1] , \nOut23_26[0] }), .Out({\nOut24_26[7] , 
        \nOut24_26[6] , \nOut24_26[5] , \nOut24_26[4] , \nOut24_26[3] , 
        \nOut24_26[2] , \nOut24_26[1] , \nOut24_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_43 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut44[7] , \nScanOut44[6] , 
        \nScanOut44[5] , \nScanOut44[4] , \nScanOut44[3] , \nScanOut44[2] , 
        \nScanOut44[1] , \nScanOut44[0] }), .ScanOut({\nScanOut43[7] , 
        \nScanOut43[6] , \nScanOut43[5] , \nScanOut43[4] , \nScanOut43[3] , 
        \nScanOut43[2] , \nScanOut43[1] , \nScanOut43[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_10[7] , \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , 
        \nOut1_10[3] , \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), 
        .SouthIn({\nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), .EastIn(
        {\nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), .WestIn(
        {\nOut0_11[7] , \nOut0_11[6] , \nOut0_11[5] , \nOut0_11[4] , 
        \nOut0_11[3] , \nOut0_11[2] , \nOut0_11[1] , \nOut0_11[0] }), .Out({
        \nOut1_11[7] , \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , 
        \nOut1_11[3] , \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_58 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut59[7] , \nScanOut59[6] , 
        \nScanOut59[5] , \nScanOut59[4] , \nScanOut59[3] , \nScanOut59[2] , 
        \nScanOut59[1] , \nScanOut59[0] }), .ScanOut({\nScanOut58[7] , 
        \nScanOut58[6] , \nScanOut58[5] , \nScanOut58[4] , \nScanOut58[3] , 
        \nScanOut58[2] , \nScanOut58[1] , \nScanOut58[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_25[7] , \nOut1_25[6] , \nOut1_25[5] , \nOut1_25[4] , 
        \nOut1_25[3] , \nOut1_25[2] , \nOut1_25[1] , \nOut1_25[0] }), 
        .SouthIn({\nOut1_27[7] , \nOut1_27[6] , \nOut1_27[5] , \nOut1_27[4] , 
        \nOut1_27[3] , \nOut1_27[2] , \nOut1_27[1] , \nOut1_27[0] }), .EastIn(
        {\nOut2_26[7] , \nOut2_26[6] , \nOut2_26[5] , \nOut2_26[4] , 
        \nOut2_26[3] , \nOut2_26[2] , \nOut2_26[1] , \nOut2_26[0] }), .WestIn(
        {\nOut0_26[7] , \nOut0_26[6] , \nOut0_26[5] , \nOut0_26[4] , 
        \nOut0_26[3] , \nOut0_26[2] , \nOut0_26[1] , \nOut0_26[0] }), .Out({
        \nOut1_26[7] , \nOut1_26[6] , \nOut1_26[5] , \nOut1_26[4] , 
        \nOut1_26[3] , \nOut1_26[2] , \nOut1_26[1] , \nOut1_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_129 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut130[7] , \nScanOut130[6] , 
        \nScanOut130[5] , \nScanOut130[4] , \nScanOut130[3] , \nScanOut130[2] , 
        \nScanOut130[1] , \nScanOut130[0] }), .ScanOut({\nScanOut129[7] , 
        \nScanOut129[6] , \nScanOut129[5] , \nScanOut129[4] , \nScanOut129[3] , 
        \nScanOut129[2] , \nScanOut129[1] , \nScanOut129[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_0[7] , \nOut4_0[6] , \nOut4_0[5] , \nOut4_0[4] , \nOut4_0[3] , 
        \nOut4_0[2] , \nOut4_0[1] , \nOut4_0[0] }), .SouthIn({\nOut4_2[7] , 
        \nOut4_2[6] , \nOut4_2[5] , \nOut4_2[4] , \nOut4_2[3] , \nOut4_2[2] , 
        \nOut4_2[1] , \nOut4_2[0] }), .EastIn({\nOut5_1[7] , \nOut5_1[6] , 
        \nOut5_1[5] , \nOut5_1[4] , \nOut5_1[3] , \nOut5_1[2] , \nOut5_1[1] , 
        \nOut5_1[0] }), .WestIn({\nOut3_1[7] , \nOut3_1[6] , \nOut3_1[5] , 
        \nOut3_1[4] , \nOut3_1[3] , \nOut3_1[2] , \nOut3_1[1] , \nOut3_1[0] }), 
        .Out({\nOut4_1[7] , \nOut4_1[6] , \nOut4_1[5] , \nOut4_1[4] , 
        \nOut4_1[3] , \nOut4_1[2] , \nOut4_1[1] , \nOut4_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_219 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut220[7] , \nScanOut220[6] , 
        \nScanOut220[5] , \nScanOut220[4] , \nScanOut220[3] , \nScanOut220[2] , 
        \nScanOut220[1] , \nScanOut220[0] }), .ScanOut({\nScanOut219[7] , 
        \nScanOut219[6] , \nScanOut219[5] , \nScanOut219[4] , \nScanOut219[3] , 
        \nScanOut219[2] , \nScanOut219[1] , \nScanOut219[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_26[7] , \nOut6_26[6] , \nOut6_26[5] , \nOut6_26[4] , 
        \nOut6_26[3] , \nOut6_26[2] , \nOut6_26[1] , \nOut6_26[0] }), 
        .SouthIn({\nOut6_28[7] , \nOut6_28[6] , \nOut6_28[5] , \nOut6_28[4] , 
        \nOut6_28[3] , \nOut6_28[2] , \nOut6_28[1] , \nOut6_28[0] }), .EastIn(
        {\nOut7_27[7] , \nOut7_27[6] , \nOut7_27[5] , \nOut7_27[4] , 
        \nOut7_27[3] , \nOut7_27[2] , \nOut7_27[1] , \nOut7_27[0] }), .WestIn(
        {\nOut5_27[7] , \nOut5_27[6] , \nOut5_27[5] , \nOut5_27[4] , 
        \nOut5_27[3] , \nOut5_27[2] , \nOut5_27[1] , \nOut5_27[0] }), .Out({
        \nOut6_27[7] , \nOut6_27[6] , \nOut6_27[5] , \nOut6_27[4] , 
        \nOut6_27[3] , \nOut6_27[2] , \nOut6_27[1] , \nOut6_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_325 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut326[7] , \nScanOut326[6] , 
        \nScanOut326[5] , \nScanOut326[4] , \nScanOut326[3] , \nScanOut326[2] , 
        \nScanOut326[1] , \nScanOut326[0] }), .ScanOut({\nScanOut325[7] , 
        \nScanOut325[6] , \nScanOut325[5] , \nScanOut325[4] , \nScanOut325[3] , 
        \nScanOut325[2] , \nScanOut325[1] , \nScanOut325[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_4[7] , \nOut10_4[6] , \nOut10_4[5] , \nOut10_4[4] , 
        \nOut10_4[3] , \nOut10_4[2] , \nOut10_4[1] , \nOut10_4[0] }), 
        .SouthIn({\nOut10_6[7] , \nOut10_6[6] , \nOut10_6[5] , \nOut10_6[4] , 
        \nOut10_6[3] , \nOut10_6[2] , \nOut10_6[1] , \nOut10_6[0] }), .EastIn(
        {\nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }), .WestIn(
        {\nOut9_5[7] , \nOut9_5[6] , \nOut9_5[5] , \nOut9_5[4] , \nOut9_5[3] , 
        \nOut9_5[2] , \nOut9_5[1] , \nOut9_5[0] }), .Out({\nOut10_5[7] , 
        \nOut10_5[6] , \nOut10_5[5] , \nOut10_5[4] , \nOut10_5[3] , 
        \nOut10_5[2] , \nOut10_5[1] , \nOut10_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_946 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut947[7] , \nScanOut947[6] , 
        \nScanOut947[5] , \nScanOut947[4] , \nScanOut947[3] , \nScanOut947[2] , 
        \nScanOut947[1] , \nScanOut947[0] }), .ScanOut({\nScanOut946[7] , 
        \nScanOut946[6] , \nScanOut946[5] , \nScanOut946[4] , \nScanOut946[3] , 
        \nScanOut946[2] , \nScanOut946[1] , \nScanOut946[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_17[7] , \nOut29_17[6] , \nOut29_17[5] , \nOut29_17[4] , 
        \nOut29_17[3] , \nOut29_17[2] , \nOut29_17[1] , \nOut29_17[0] }), 
        .SouthIn({\nOut29_19[7] , \nOut29_19[6] , \nOut29_19[5] , 
        \nOut29_19[4] , \nOut29_19[3] , \nOut29_19[2] , \nOut29_19[1] , 
        \nOut29_19[0] }), .EastIn({\nOut30_18[7] , \nOut30_18[6] , 
        \nOut30_18[5] , \nOut30_18[4] , \nOut30_18[3] , \nOut30_18[2] , 
        \nOut30_18[1] , \nOut30_18[0] }), .WestIn({\nOut28_18[7] , 
        \nOut28_18[6] , \nOut28_18[5] , \nOut28_18[4] , \nOut28_18[3] , 
        \nOut28_18[2] , \nOut28_18[1] , \nOut28_18[0] }), .Out({\nOut29_18[7] , 
        \nOut29_18[6] , \nOut29_18[5] , \nOut29_18[4] , \nOut29_18[3] , 
        \nOut29_18[2] , \nOut29_18[1] , \nOut29_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_534 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut535[7] , \nScanOut535[6] , 
        \nScanOut535[5] , \nScanOut535[4] , \nScanOut535[3] , \nScanOut535[2] , 
        \nScanOut535[1] , \nScanOut535[0] }), .ScanOut({\nScanOut534[7] , 
        \nScanOut534[6] , \nScanOut534[5] , \nScanOut534[4] , \nScanOut534[3] , 
        \nScanOut534[2] , \nScanOut534[1] , \nScanOut534[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_21[7] , \nOut16_21[6] , \nOut16_21[5] , \nOut16_21[4] , 
        \nOut16_21[3] , \nOut16_21[2] , \nOut16_21[1] , \nOut16_21[0] }), 
        .SouthIn({\nOut16_23[7] , \nOut16_23[6] , \nOut16_23[5] , 
        \nOut16_23[4] , \nOut16_23[3] , \nOut16_23[2] , \nOut16_23[1] , 
        \nOut16_23[0] }), .EastIn({\nOut17_22[7] , \nOut17_22[6] , 
        \nOut17_22[5] , \nOut17_22[4] , \nOut17_22[3] , \nOut17_22[2] , 
        \nOut17_22[1] , \nOut17_22[0] }), .WestIn({\nOut15_22[7] , 
        \nOut15_22[6] , \nOut15_22[5] , \nOut15_22[4] , \nOut15_22[3] , 
        \nOut15_22[2] , \nOut15_22[1] , \nOut15_22[0] }), .Out({\nOut16_22[7] , 
        \nOut16_22[6] , \nOut16_22[5] , \nOut16_22[4] , \nOut16_22[3] , 
        \nOut16_22[2] , \nOut16_22[1] , \nOut16_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_389 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut390[7] , \nScanOut390[6] , 
        \nScanOut390[5] , \nScanOut390[4] , \nScanOut390[3] , \nScanOut390[2] , 
        \nScanOut390[1] , \nScanOut390[0] }), .ScanOut({\nScanOut389[7] , 
        \nScanOut389[6] , \nScanOut389[5] , \nScanOut389[4] , \nScanOut389[3] , 
        \nScanOut389[2] , \nScanOut389[1] , \nScanOut389[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }), 
        .SouthIn({\nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }), .EastIn(
        {\nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }), .WestIn(
        {\nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }), .Out({
        \nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_598 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut599[7] , \nScanOut599[6] , 
        \nScanOut599[5] , \nScanOut599[4] , \nScanOut599[3] , \nScanOut599[2] , 
        \nScanOut599[1] , \nScanOut599[0] }), .ScanOut({\nScanOut598[7] , 
        \nScanOut598[6] , \nScanOut598[5] , \nScanOut598[4] , \nScanOut598[3] , 
        \nScanOut598[2] , \nScanOut598[1] , \nScanOut598[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_21[7] , \nOut18_21[6] , \nOut18_21[5] , \nOut18_21[4] , 
        \nOut18_21[3] , \nOut18_21[2] , \nOut18_21[1] , \nOut18_21[0] }), 
        .SouthIn({\nOut18_23[7] , \nOut18_23[6] , \nOut18_23[5] , 
        \nOut18_23[4] , \nOut18_23[3] , \nOut18_23[2] , \nOut18_23[1] , 
        \nOut18_23[0] }), .EastIn({\nOut19_22[7] , \nOut19_22[6] , 
        \nOut19_22[5] , \nOut19_22[4] , \nOut19_22[3] , \nOut19_22[2] , 
        \nOut19_22[1] , \nOut19_22[0] }), .WestIn({\nOut17_22[7] , 
        \nOut17_22[6] , \nOut17_22[5] , \nOut17_22[4] , \nOut17_22[3] , 
        \nOut17_22[2] , \nOut17_22[1] , \nOut17_22[0] }), .Out({\nOut18_22[7] , 
        \nOut18_22[6] , \nOut18_22[5] , \nOut18_22[4] , \nOut18_22[3] , 
        \nOut18_22[2] , \nOut18_22[1] , \nOut18_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_408 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut409[7] , \nScanOut409[6] , 
        \nScanOut409[5] , \nScanOut409[4] , \nScanOut409[3] , \nScanOut409[2] , 
        \nScanOut409[1] , \nScanOut409[0] }), .ScanOut({\nScanOut408[7] , 
        \nScanOut408[6] , \nScanOut408[5] , \nScanOut408[4] , \nScanOut408[3] , 
        \nScanOut408[2] , \nScanOut408[1] , \nScanOut408[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_23[7] , \nOut12_23[6] , \nOut12_23[5] , \nOut12_23[4] , 
        \nOut12_23[3] , \nOut12_23[2] , \nOut12_23[1] , \nOut12_23[0] }), 
        .SouthIn({\nOut12_25[7] , \nOut12_25[6] , \nOut12_25[5] , 
        \nOut12_25[4] , \nOut12_25[3] , \nOut12_25[2] , \nOut12_25[1] , 
        \nOut12_25[0] }), .EastIn({\nOut13_24[7] , \nOut13_24[6] , 
        \nOut13_24[5] , \nOut13_24[4] , \nOut13_24[3] , \nOut13_24[2] , 
        \nOut13_24[1] , \nOut13_24[0] }), .WestIn({\nOut11_24[7] , 
        \nOut11_24[6] , \nOut11_24[5] , \nOut11_24[4] , \nOut11_24[3] , 
        \nOut11_24[2] , \nOut11_24[1] , \nOut11_24[0] }), .Out({\nOut12_24[7] , 
        \nOut12_24[6] , \nOut12_24[5] , \nOut12_24[4] , \nOut12_24[3] , 
        \nOut12_24[2] , \nOut12_24[1] , \nOut12_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_147 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut148[7] , \nScanOut148[6] , 
        \nScanOut148[5] , \nScanOut148[4] , \nScanOut148[3] , \nScanOut148[2] , 
        \nScanOut148[1] , \nScanOut148[0] }), .ScanOut({\nScanOut147[7] , 
        \nScanOut147[6] , \nScanOut147[5] , \nScanOut147[4] , \nScanOut147[3] , 
        \nScanOut147[2] , \nScanOut147[1] , \nScanOut147[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_18[7] , \nOut4_18[6] , \nOut4_18[5] , \nOut4_18[4] , 
        \nOut4_18[3] , \nOut4_18[2] , \nOut4_18[1] , \nOut4_18[0] }), 
        .SouthIn({\nOut4_20[7] , \nOut4_20[6] , \nOut4_20[5] , \nOut4_20[4] , 
        \nOut4_20[3] , \nOut4_20[2] , \nOut4_20[1] , \nOut4_20[0] }), .EastIn(
        {\nOut5_19[7] , \nOut5_19[6] , \nOut5_19[5] , \nOut5_19[4] , 
        \nOut5_19[3] , \nOut5_19[2] , \nOut5_19[1] , \nOut5_19[0] }), .WestIn(
        {\nOut3_19[7] , \nOut3_19[6] , \nOut3_19[5] , \nOut3_19[4] , 
        \nOut3_19[3] , \nOut3_19[2] , \nOut3_19[1] , \nOut3_19[0] }), .Out({
        \nOut4_19[7] , \nOut4_19[6] , \nOut4_19[5] , \nOut4_19[4] , 
        \nOut4_19[3] , \nOut4_19[2] , \nOut4_19[1] , \nOut4_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_160 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut161[7] , \nScanOut161[6] , 
        \nScanOut161[5] , \nScanOut161[4] , \nScanOut161[3] , \nScanOut161[2] , 
        \nScanOut161[1] , \nScanOut161[0] }), .ScanOut({\nScanOut160[7] , 
        \nScanOut160[6] , \nScanOut160[5] , \nScanOut160[4] , \nScanOut160[3] , 
        \nScanOut160[2] , \nScanOut160[1] , \nScanOut160[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut5_0[7] , \nOut5_0[6] , 
        \nOut5_0[5] , \nOut5_0[4] , \nOut5_0[3] , \nOut5_0[2] , \nOut5_0[1] , 
        \nOut5_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_738 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut739[7] , \nScanOut739[6] , 
        \nScanOut739[5] , \nScanOut739[4] , \nScanOut739[3] , \nScanOut739[2] , 
        \nScanOut739[1] , \nScanOut739[0] }), .ScanOut({\nScanOut738[7] , 
        \nScanOut738[6] , \nScanOut738[5] , \nScanOut738[4] , \nScanOut738[3] , 
        \nScanOut738[2] , \nScanOut738[1] , \nScanOut738[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_1[7] , \nOut23_1[6] , \nOut23_1[5] , \nOut23_1[4] , 
        \nOut23_1[3] , \nOut23_1[2] , \nOut23_1[1] , \nOut23_1[0] }), 
        .SouthIn({\nOut23_3[7] , \nOut23_3[6] , \nOut23_3[5] , \nOut23_3[4] , 
        \nOut23_3[3] , \nOut23_3[2] , \nOut23_3[1] , \nOut23_3[0] }), .EastIn(
        {\nOut24_2[7] , \nOut24_2[6] , \nOut24_2[5] , \nOut24_2[4] , 
        \nOut24_2[3] , \nOut24_2[2] , \nOut24_2[1] , \nOut24_2[0] }), .WestIn(
        {\nOut22_2[7] , \nOut22_2[6] , \nOut22_2[5] , \nOut22_2[4] , 
        \nOut22_2[3] , \nOut22_2[2] , \nOut22_2[1] , \nOut22_2[0] }), .Out({
        \nOut23_2[7] , \nOut23_2[6] , \nOut23_2[5] , \nOut23_2[4] , 
        \nOut23_2[3] , \nOut23_2[2] , \nOut23_2[1] , \nOut23_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1019 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1020[7] , \nScanOut1020[6] , 
        \nScanOut1020[5] , \nScanOut1020[4] , \nScanOut1020[3] , 
        \nScanOut1020[2] , \nScanOut1020[1] , \nScanOut1020[0] }), .ScanOut({
        \nScanOut1019[7] , \nScanOut1019[6] , \nScanOut1019[5] , 
        \nScanOut1019[4] , \nScanOut1019[3] , \nScanOut1019[2] , 
        \nScanOut1019[1] , \nScanOut1019[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_27[7] , \nOut31_27[6] , \nOut31_27[5] , 
        \nOut31_27[4] , \nOut31_27[3] , \nOut31_27[2] , \nOut31_27[1] , 
        \nOut31_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_250 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut251[7] , \nScanOut251[6] , 
        \nScanOut251[5] , \nScanOut251[4] , \nScanOut251[3] , \nScanOut251[2] , 
        \nScanOut251[1] , \nScanOut251[0] }), .ScanOut({\nScanOut250[7] , 
        \nScanOut250[6] , \nScanOut250[5] , \nScanOut250[4] , \nScanOut250[3] , 
        \nScanOut250[2] , \nScanOut250[1] , \nScanOut250[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_25[7] , \nOut7_25[6] , \nOut7_25[5] , \nOut7_25[4] , 
        \nOut7_25[3] , \nOut7_25[2] , \nOut7_25[1] , \nOut7_25[0] }), 
        .SouthIn({\nOut7_27[7] , \nOut7_27[6] , \nOut7_27[5] , \nOut7_27[4] , 
        \nOut7_27[3] , \nOut7_27[2] , \nOut7_27[1] , \nOut7_27[0] }), .EastIn(
        {\nOut8_26[7] , \nOut8_26[6] , \nOut8_26[5] , \nOut8_26[4] , 
        \nOut8_26[3] , \nOut8_26[2] , \nOut8_26[1] , \nOut8_26[0] }), .WestIn(
        {\nOut6_26[7] , \nOut6_26[6] , \nOut6_26[5] , \nOut6_26[4] , 
        \nOut6_26[3] , \nOut6_26[2] , \nOut6_26[1] , \nOut6_26[0] }), .Out({
        \nOut7_26[7] , \nOut7_26[6] , \nOut7_26[5] , \nOut7_26[4] , 
        \nOut7_26[3] , \nOut7_26[2] , \nOut7_26[1] , \nOut7_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_771 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut772[7] , \nScanOut772[6] , 
        \nScanOut772[5] , \nScanOut772[4] , \nScanOut772[3] , \nScanOut772[2] , 
        \nScanOut772[1] , \nScanOut772[0] }), .ScanOut({\nScanOut771[7] , 
        \nScanOut771[6] , \nScanOut771[5] , \nScanOut771[4] , \nScanOut771[3] , 
        \nScanOut771[2] , \nScanOut771[1] , \nScanOut771[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_2[7] , \nOut24_2[6] , \nOut24_2[5] , \nOut24_2[4] , 
        \nOut24_2[3] , \nOut24_2[2] , \nOut24_2[1] , \nOut24_2[0] }), 
        .SouthIn({\nOut24_4[7] , \nOut24_4[6] , \nOut24_4[5] , \nOut24_4[4] , 
        \nOut24_4[3] , \nOut24_4[2] , \nOut24_4[1] , \nOut24_4[0] }), .EastIn(
        {\nOut25_3[7] , \nOut25_3[6] , \nOut25_3[5] , \nOut25_3[4] , 
        \nOut25_3[3] , \nOut25_3[2] , \nOut25_3[1] , \nOut25_3[0] }), .WestIn(
        {\nOut23_3[7] , \nOut23_3[6] , \nOut23_3[5] , \nOut23_3[4] , 
        \nOut23_3[3] , \nOut23_3[2] , \nOut23_3[1] , \nOut23_3[0] }), .Out({
        \nOut24_3[7] , \nOut24_3[6] , \nOut24_3[5] , \nOut24_3[4] , 
        \nOut24_3[3] , \nOut24_3[2] , \nOut24_3[1] , \nOut24_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_833 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut834[7] , \nScanOut834[6] , 
        \nScanOut834[5] , \nScanOut834[4] , \nScanOut834[3] , \nScanOut834[2] , 
        \nScanOut834[1] , \nScanOut834[0] }), .ScanOut({\nScanOut833[7] , 
        \nScanOut833[6] , \nScanOut833[5] , \nScanOut833[4] , \nScanOut833[3] , 
        \nScanOut833[2] , \nScanOut833[1] , \nScanOut833[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_0[7] , \nOut26_0[6] , \nOut26_0[5] , \nOut26_0[4] , 
        \nOut26_0[3] , \nOut26_0[2] , \nOut26_0[1] , \nOut26_0[0] }), 
        .SouthIn({\nOut26_2[7] , \nOut26_2[6] , \nOut26_2[5] , \nOut26_2[4] , 
        \nOut26_2[3] , \nOut26_2[2] , \nOut26_2[1] , \nOut26_2[0] }), .EastIn(
        {\nOut27_1[7] , \nOut27_1[6] , \nOut27_1[5] , \nOut27_1[4] , 
        \nOut27_1[3] , \nOut27_1[2] , \nOut27_1[1] , \nOut27_1[0] }), .WestIn(
        {\nOut25_1[7] , \nOut25_1[6] , \nOut25_1[5] , \nOut25_1[4] , 
        \nOut25_1[3] , \nOut25_1[2] , \nOut25_1[1] , \nOut25_1[0] }), .Out({
        \nOut26_1[7] , \nOut26_1[6] , \nOut26_1[5] , \nOut26_1[4] , 
        \nOut26_1[3] , \nOut26_1[2] , \nOut26_1[1] , \nOut26_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_277 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut278[7] , \nScanOut278[6] , 
        \nScanOut278[5] , \nScanOut278[4] , \nScanOut278[3] , \nScanOut278[2] , 
        \nScanOut278[1] , \nScanOut278[0] }), .ScanOut({\nScanOut277[7] , 
        \nScanOut277[6] , \nScanOut277[5] , \nScanOut277[4] , \nScanOut277[3] , 
        \nScanOut277[2] , \nScanOut277[1] , \nScanOut277[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_20[7] , \nOut8_20[6] , \nOut8_20[5] , \nOut8_20[4] , 
        \nOut8_20[3] , \nOut8_20[2] , \nOut8_20[1] , \nOut8_20[0] }), 
        .SouthIn({\nOut8_22[7] , \nOut8_22[6] , \nOut8_22[5] , \nOut8_22[4] , 
        \nOut8_22[3] , \nOut8_22[2] , \nOut8_22[1] , \nOut8_22[0] }), .EastIn(
        {\nOut9_21[7] , \nOut9_21[6] , \nOut9_21[5] , \nOut9_21[4] , 
        \nOut9_21[3] , \nOut9_21[2] , \nOut9_21[1] , \nOut9_21[0] }), .WestIn(
        {\nOut7_21[7] , \nOut7_21[6] , \nOut7_21[5] , \nOut7_21[4] , 
        \nOut7_21[3] , \nOut7_21[2] , \nOut7_21[1] , \nOut7_21[0] }), .Out({
        \nOut8_21[7] , \nOut8_21[6] , \nOut8_21[5] , \nOut8_21[4] , 
        \nOut8_21[3] , \nOut8_21[2] , \nOut8_21[1] , \nOut8_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_441 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut442[7] , \nScanOut442[6] , 
        \nScanOut442[5] , \nScanOut442[4] , \nScanOut442[3] , \nScanOut442[2] , 
        \nScanOut442[1] , \nScanOut442[0] }), .ScanOut({\nScanOut441[7] , 
        \nScanOut441[6] , \nScanOut441[5] , \nScanOut441[4] , \nScanOut441[3] , 
        \nScanOut441[2] , \nScanOut441[1] , \nScanOut441[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_24[7] , \nOut13_24[6] , \nOut13_24[5] , \nOut13_24[4] , 
        \nOut13_24[3] , \nOut13_24[2] , \nOut13_24[1] , \nOut13_24[0] }), 
        .SouthIn({\nOut13_26[7] , \nOut13_26[6] , \nOut13_26[5] , 
        \nOut13_26[4] , \nOut13_26[3] , \nOut13_26[2] , \nOut13_26[1] , 
        \nOut13_26[0] }), .EastIn({\nOut14_25[7] , \nOut14_25[6] , 
        \nOut14_25[5] , \nOut14_25[4] , \nOut14_25[3] , \nOut14_25[2] , 
        \nOut14_25[1] , \nOut14_25[0] }), .WestIn({\nOut12_25[7] , 
        \nOut12_25[6] , \nOut12_25[5] , \nOut12_25[4] , \nOut12_25[3] , 
        \nOut12_25[2] , \nOut12_25[1] , \nOut12_25[0] }), .Out({\nOut13_25[7] , 
        \nOut13_25[6] , \nOut13_25[5] , \nOut13_25[4] , \nOut13_25[3] , 
        \nOut13_25[2] , \nOut13_25[1] , \nOut13_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_466 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut467[7] , \nScanOut467[6] , 
        \nScanOut467[5] , \nScanOut467[4] , \nScanOut467[3] , \nScanOut467[2] , 
        \nScanOut467[1] , \nScanOut467[0] }), .ScanOut({\nScanOut466[7] , 
        \nScanOut466[6] , \nScanOut466[5] , \nScanOut466[4] , \nScanOut466[3] , 
        \nScanOut466[2] , \nScanOut466[1] , \nScanOut466[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_17[7] , \nOut14_17[6] , \nOut14_17[5] , \nOut14_17[4] , 
        \nOut14_17[3] , \nOut14_17[2] , \nOut14_17[1] , \nOut14_17[0] }), 
        .SouthIn({\nOut14_19[7] , \nOut14_19[6] , \nOut14_19[5] , 
        \nOut14_19[4] , \nOut14_19[3] , \nOut14_19[2] , \nOut14_19[1] , 
        \nOut14_19[0] }), .EastIn({\nOut15_18[7] , \nOut15_18[6] , 
        \nOut15_18[5] , \nOut15_18[4] , \nOut15_18[3] , \nOut15_18[2] , 
        \nOut15_18[1] , \nOut15_18[0] }), .WestIn({\nOut13_18[7] , 
        \nOut13_18[6] , \nOut13_18[5] , \nOut13_18[4] , \nOut13_18[3] , 
        \nOut13_18[2] , \nOut13_18[1] , \nOut13_18[0] }), .Out({\nOut14_18[7] , 
        \nOut14_18[6] , \nOut14_18[5] , \nOut14_18[4] , \nOut14_18[3] , 
        \nOut14_18[2] , \nOut14_18[1] , \nOut14_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_814 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut815[7] , \nScanOut815[6] , 
        \nScanOut815[5] , \nScanOut815[4] , \nScanOut815[3] , \nScanOut815[2] , 
        \nScanOut815[1] , \nScanOut815[0] }), .ScanOut({\nScanOut814[7] , 
        \nScanOut814[6] , \nScanOut814[5] , \nScanOut814[4] , \nScanOut814[3] , 
        \nScanOut814[2] , \nScanOut814[1] , \nScanOut814[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_13[7] , \nOut25_13[6] , \nOut25_13[5] , \nOut25_13[4] , 
        \nOut25_13[3] , \nOut25_13[2] , \nOut25_13[1] , \nOut25_13[0] }), 
        .SouthIn({\nOut25_15[7] , \nOut25_15[6] , \nOut25_15[5] , 
        \nOut25_15[4] , \nOut25_15[3] , \nOut25_15[2] , \nOut25_15[1] , 
        \nOut25_15[0] }), .EastIn({\nOut26_14[7] , \nOut26_14[6] , 
        \nOut26_14[5] , \nOut26_14[4] , \nOut26_14[3] , \nOut26_14[2] , 
        \nOut26_14[1] , \nOut26_14[0] }), .WestIn({\nOut24_14[7] , 
        \nOut24_14[6] , \nOut24_14[5] , \nOut24_14[4] , \nOut24_14[3] , 
        \nOut24_14[2] , \nOut24_14[1] , \nOut24_14[0] }), .Out({\nOut25_14[7] , 
        \nOut25_14[6] , \nOut25_14[5] , \nOut25_14[4] , \nOut25_14[3] , 
        \nOut25_14[2] , \nOut25_14[1] , \nOut25_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_984 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut985[7] , \nScanOut985[6] , 
        \nScanOut985[5] , \nScanOut985[4] , \nScanOut985[3] , \nScanOut985[2] , 
        \nScanOut985[1] , \nScanOut985[0] }), .ScanOut({\nScanOut984[7] , 
        \nScanOut984[6] , \nScanOut984[5] , \nScanOut984[4] , \nScanOut984[3] , 
        \nScanOut984[2] , \nScanOut984[1] , \nScanOut984[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_23[7] , \nOut30_23[6] , \nOut30_23[5] , \nOut30_23[4] , 
        \nOut30_23[3] , \nOut30_23[2] , \nOut30_23[1] , \nOut30_23[0] }), 
        .SouthIn({\nOut30_25[7] , \nOut30_25[6] , \nOut30_25[5] , 
        \nOut30_25[4] , \nOut30_25[3] , \nOut30_25[2] , \nOut30_25[1] , 
        \nOut30_25[0] }), .EastIn({\nOut31_24[7] , \nOut31_24[6] , 
        \nOut31_24[5] , \nOut31_24[4] , \nOut31_24[3] , \nOut31_24[2] , 
        \nOut31_24[1] , \nOut31_24[0] }), .WestIn({\nOut29_24[7] , 
        \nOut29_24[6] , \nOut29_24[5] , \nOut29_24[4] , \nOut29_24[3] , 
        \nOut29_24[2] , \nOut29_24[1] , \nOut29_24[0] }), .Out({\nOut30_24[7] , 
        \nOut30_24[6] , \nOut30_24[5] , \nOut30_24[4] , \nOut30_24[3] , 
        \nOut30_24[2] , \nOut30_24[1] , \nOut30_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_756 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut757[7] , \nScanOut757[6] , 
        \nScanOut757[5] , \nScanOut757[4] , \nScanOut757[3] , \nScanOut757[2] , 
        \nScanOut757[1] , \nScanOut757[0] }), .ScanOut({\nScanOut756[7] , 
        \nScanOut756[6] , \nScanOut756[5] , \nScanOut756[4] , \nScanOut756[3] , 
        \nScanOut756[2] , \nScanOut756[1] , \nScanOut756[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_19[7] , \nOut23_19[6] , \nOut23_19[5] , \nOut23_19[4] , 
        \nOut23_19[3] , \nOut23_19[2] , \nOut23_19[1] , \nOut23_19[0] }), 
        .SouthIn({\nOut23_21[7] , \nOut23_21[6] , \nOut23_21[5] , 
        \nOut23_21[4] , \nOut23_21[3] , \nOut23_21[2] , \nOut23_21[1] , 
        \nOut23_21[0] }), .EastIn({\nOut24_20[7] , \nOut24_20[6] , 
        \nOut24_20[5] , \nOut24_20[4] , \nOut24_20[3] , \nOut24_20[2] , 
        \nOut24_20[1] , \nOut24_20[0] }), .WestIn({\nOut22_20[7] , 
        \nOut22_20[6] , \nOut22_20[5] , \nOut22_20[4] , \nOut22_20[3] , 
        \nOut22_20[2] , \nOut22_20[1] , \nOut22_20[0] }), .Out({\nOut23_20[7] , 
        \nOut23_20[6] , \nOut23_20[5] , \nOut23_20[4] , \nOut23_20[3] , 
        \nOut23_20[2] , \nOut23_20[1] , \nOut23_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_928 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut929[7] , \nScanOut929[6] , 
        \nScanOut929[5] , \nScanOut929[4] , \nScanOut929[3] , \nScanOut929[2] , 
        \nScanOut929[1] , \nScanOut929[0] }), .ScanOut({\nScanOut928[7] , 
        \nScanOut928[6] , \nScanOut928[5] , \nScanOut928[4] , \nScanOut928[3] , 
        \nScanOut928[2] , \nScanOut928[1] , \nScanOut928[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut29_0[7] , \nOut29_0[6] , 
        \nOut29_0[5] , \nOut29_0[4] , \nOut29_0[3] , \nOut29_0[2] , 
        \nOut29_0[1] , \nOut29_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_656 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut657[7] , \nScanOut657[6] , 
        \nScanOut657[5] , \nScanOut657[4] , \nScanOut657[3] , \nScanOut657[2] , 
        \nScanOut657[1] , \nScanOut657[0] }), .ScanOut({\nScanOut656[7] , 
        \nScanOut656[6] , \nScanOut656[5] , \nScanOut656[4] , \nScanOut656[3] , 
        \nScanOut656[2] , \nScanOut656[1] , \nScanOut656[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_15[7] , \nOut20_15[6] , \nOut20_15[5] , \nOut20_15[4] , 
        \nOut20_15[3] , \nOut20_15[2] , \nOut20_15[1] , \nOut20_15[0] }), 
        .SouthIn({\nOut20_17[7] , \nOut20_17[6] , \nOut20_17[5] , 
        \nOut20_17[4] , \nOut20_17[3] , \nOut20_17[2] , \nOut20_17[1] , 
        \nOut20_17[0] }), .EastIn({\nOut21_16[7] , \nOut21_16[6] , 
        \nOut21_16[5] , \nOut21_16[4] , \nOut21_16[3] , \nOut21_16[2] , 
        \nOut21_16[1] , \nOut21_16[0] }), .WestIn({\nOut19_16[7] , 
        \nOut19_16[6] , \nOut19_16[5] , \nOut19_16[4] , \nOut19_16[3] , 
        \nOut19_16[2] , \nOut19_16[1] , \nOut19_16[0] }), .Out({\nOut20_16[7] , 
        \nOut20_16[6] , \nOut20_16[5] , \nOut20_16[4] , \nOut20_16[3] , 
        \nOut20_16[2] , \nOut20_16[1] , \nOut20_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_7 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut8[7] , \nScanOut8[6] , 
        \nScanOut8[5] , \nScanOut8[4] , \nScanOut8[3] , \nScanOut8[2] , 
        \nScanOut8[1] , \nScanOut8[0] }), .ScanOut({\nScanOut7[7] , 
        \nScanOut7[6] , \nScanOut7[5] , \nScanOut7[4] , \nScanOut7[3] , 
        \nScanOut7[2] , \nScanOut7[1] , \nScanOut7[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_7[7] , \nOut0_7[6] , 
        \nOut0_7[5] , \nOut0_7[4] , \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , 
        \nOut0_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_26 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut27[7] , \nScanOut27[6] , 
        \nScanOut27[5] , \nScanOut27[4] , \nScanOut27[3] , \nScanOut27[2] , 
        \nScanOut27[1] , \nScanOut27[0] }), .ScanOut({\nScanOut26[7] , 
        \nScanOut26[6] , \nScanOut26[5] , \nScanOut26[4] , \nScanOut26[3] , 
        \nScanOut26[2] , \nScanOut26[1] , \nScanOut26[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_26[7] , \nOut0_26[6] , 
        \nOut0_26[5] , \nOut0_26[4] , \nOut0_26[3] , \nOut0_26[2] , 
        \nOut0_26[1] , \nOut0_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_64 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut65[7] , \nScanOut65[6] , 
        \nScanOut65[5] , \nScanOut65[4] , \nScanOut65[3] , \nScanOut65[2] , 
        \nScanOut65[1] , \nScanOut65[0] }), .ScanOut({\nScanOut64[7] , 
        \nScanOut64[6] , \nScanOut64[5] , \nScanOut64[4] , \nScanOut64[3] , 
        \nScanOut64[2] , \nScanOut64[1] , \nScanOut64[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut2_0[7] , \nOut2_0[6] , 
        \nOut2_0[5] , \nOut2_0[4] , \nOut2_0[3] , \nOut2_0[2] , \nOut2_0[1] , 
        \nOut2_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_350 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut351[7] , \nScanOut351[6] , 
        \nScanOut351[5] , \nScanOut351[4] , \nScanOut351[3] , \nScanOut351[2] , 
        \nScanOut351[1] , \nScanOut351[0] }), .ScanOut({\nScanOut350[7] , 
        \nScanOut350[6] , \nScanOut350[5] , \nScanOut350[4] , \nScanOut350[3] , 
        \nScanOut350[2] , \nScanOut350[1] , \nScanOut350[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_29[7] , \nOut10_29[6] , \nOut10_29[5] , \nOut10_29[4] , 
        \nOut10_29[3] , \nOut10_29[2] , \nOut10_29[1] , \nOut10_29[0] }), 
        .SouthIn({\nOut10_31[7] , \nOut10_31[6] , \nOut10_31[5] , 
        \nOut10_31[4] , \nOut10_31[3] , \nOut10_31[2] , \nOut10_31[1] , 
        \nOut10_31[0] }), .EastIn({\nOut11_30[7] , \nOut11_30[6] , 
        \nOut11_30[5] , \nOut11_30[4] , \nOut11_30[3] , \nOut11_30[2] , 
        \nOut11_30[1] , \nOut11_30[0] }), .WestIn({\nOut9_30[7] , 
        \nOut9_30[6] , \nOut9_30[5] , \nOut9_30[4] , \nOut9_30[3] , 
        \nOut9_30[2] , \nOut9_30[1] , \nOut9_30[0] }), .Out({\nOut10_30[7] , 
        \nOut10_30[6] , \nOut10_30[5] , \nOut10_30[4] , \nOut10_30[3] , 
        \nOut10_30[2] , \nOut10_30[1] , \nOut10_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_377 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut378[7] , \nScanOut378[6] , 
        \nScanOut378[5] , \nScanOut378[4] , \nScanOut378[3] , \nScanOut378[2] , 
        \nScanOut378[1] , \nScanOut378[0] }), .ScanOut({\nScanOut377[7] , 
        \nScanOut377[6] , \nScanOut377[5] , \nScanOut377[4] , \nScanOut377[3] , 
        \nScanOut377[2] , \nScanOut377[1] , \nScanOut377[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_24[7] , \nOut11_24[6] , \nOut11_24[5] , \nOut11_24[4] , 
        \nOut11_24[3] , \nOut11_24[2] , \nOut11_24[1] , \nOut11_24[0] }), 
        .SouthIn({\nOut11_26[7] , \nOut11_26[6] , \nOut11_26[5] , 
        \nOut11_26[4] , \nOut11_26[3] , \nOut11_26[2] , \nOut11_26[1] , 
        \nOut11_26[0] }), .EastIn({\nOut12_25[7] , \nOut12_25[6] , 
        \nOut12_25[5] , \nOut12_25[4] , \nOut12_25[3] , \nOut12_25[2] , 
        \nOut12_25[1] , \nOut12_25[0] }), .WestIn({\nOut10_25[7] , 
        \nOut10_25[6] , \nOut10_25[5] , \nOut10_25[4] , \nOut10_25[3] , 
        \nOut10_25[2] , \nOut10_25[1] , \nOut10_25[0] }), .Out({\nOut11_25[7] , 
        \nOut11_25[6] , \nOut11_25[5] , \nOut11_25[4] , \nOut11_25[3] , 
        \nOut11_25[2] , \nOut11_25[1] , \nOut11_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_884 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut885[7] , \nScanOut885[6] , 
        \nScanOut885[5] , \nScanOut885[4] , \nScanOut885[3] , \nScanOut885[2] , 
        \nScanOut885[1] , \nScanOut885[0] }), .ScanOut({\nScanOut884[7] , 
        \nScanOut884[6] , \nScanOut884[5] , \nScanOut884[4] , \nScanOut884[3] , 
        \nScanOut884[2] , \nScanOut884[1] , \nScanOut884[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_19[7] , \nOut27_19[6] , \nOut27_19[5] , \nOut27_19[4] , 
        \nOut27_19[3] , \nOut27_19[2] , \nOut27_19[1] , \nOut27_19[0] }), 
        .SouthIn({\nOut27_21[7] , \nOut27_21[6] , \nOut27_21[5] , 
        \nOut27_21[4] , \nOut27_21[3] , \nOut27_21[2] , \nOut27_21[1] , 
        \nOut27_21[0] }), .EastIn({\nOut28_20[7] , \nOut28_20[6] , 
        \nOut28_20[5] , \nOut28_20[4] , \nOut28_20[3] , \nOut28_20[2] , 
        \nOut28_20[1] , \nOut28_20[0] }), .WestIn({\nOut26_20[7] , 
        \nOut26_20[6] , \nOut26_20[5] , \nOut26_20[4] , \nOut26_20[3] , 
        \nOut26_20[2] , \nOut26_20[1] , \nOut26_20[0] }), .Out({\nOut27_20[7] , 
        \nOut27_20[6] , \nOut27_20[5] , \nOut27_20[4] , \nOut27_20[3] , 
        \nOut27_20[2] , \nOut27_20[1] , \nOut27_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_914 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut915[7] , \nScanOut915[6] , 
        \nScanOut915[5] , \nScanOut915[4] , \nScanOut915[3] , \nScanOut915[2] , 
        \nScanOut915[1] , \nScanOut915[0] }), .ScanOut({\nScanOut914[7] , 
        \nScanOut914[6] , \nScanOut914[5] , \nScanOut914[4] , \nScanOut914[3] , 
        \nScanOut914[2] , \nScanOut914[1] , \nScanOut914[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_17[7] , \nOut28_17[6] , \nOut28_17[5] , \nOut28_17[4] , 
        \nOut28_17[3] , \nOut28_17[2] , \nOut28_17[1] , \nOut28_17[0] }), 
        .SouthIn({\nOut28_19[7] , \nOut28_19[6] , \nOut28_19[5] , 
        \nOut28_19[4] , \nOut28_19[3] , \nOut28_19[2] , \nOut28_19[1] , 
        \nOut28_19[0] }), .EastIn({\nOut29_18[7] , \nOut29_18[6] , 
        \nOut29_18[5] , \nOut29_18[4] , \nOut29_18[3] , \nOut29_18[2] , 
        \nOut29_18[1] , \nOut29_18[0] }), .WestIn({\nOut27_18[7] , 
        \nOut27_18[6] , \nOut27_18[5] , \nOut27_18[4] , \nOut27_18[3] , 
        \nOut27_18[2] , \nOut27_18[1] , \nOut27_18[0] }), .Out({\nOut28_18[7] , 
        \nOut28_18[6] , \nOut28_18[5] , \nOut28_18[4] , \nOut28_18[3] , 
        \nOut28_18[2] , \nOut28_18[1] , \nOut28_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_541 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut542[7] , \nScanOut542[6] , 
        \nScanOut542[5] , \nScanOut542[4] , \nScanOut542[3] , \nScanOut542[2] , 
        \nScanOut542[1] , \nScanOut542[0] }), .ScanOut({\nScanOut541[7] , 
        \nScanOut541[6] , \nScanOut541[5] , \nScanOut541[4] , \nScanOut541[3] , 
        \nScanOut541[2] , \nScanOut541[1] , \nScanOut541[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_28[7] , \nOut16_28[6] , \nOut16_28[5] , \nOut16_28[4] , 
        \nOut16_28[3] , \nOut16_28[2] , \nOut16_28[1] , \nOut16_28[0] }), 
        .SouthIn({\nOut16_30[7] , \nOut16_30[6] , \nOut16_30[5] , 
        \nOut16_30[4] , \nOut16_30[3] , \nOut16_30[2] , \nOut16_30[1] , 
        \nOut16_30[0] }), .EastIn({\nOut17_29[7] , \nOut17_29[6] , 
        \nOut17_29[5] , \nOut17_29[4] , \nOut17_29[3] , \nOut17_29[2] , 
        \nOut17_29[1] , \nOut17_29[0] }), .WestIn({\nOut15_29[7] , 
        \nOut15_29[6] , \nOut15_29[5] , \nOut15_29[4] , \nOut15_29[3] , 
        \nOut15_29[2] , \nOut15_29[1] , \nOut15_29[0] }), .Out({\nOut16_29[7] , 
        \nOut16_29[6] , \nOut16_29[5] , \nOut16_29[4] , \nOut16_29[3] , 
        \nOut16_29[2] , \nOut16_29[1] , \nOut16_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_566 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut567[7] , \nScanOut567[6] , 
        \nScanOut567[5] , \nScanOut567[4] , \nScanOut567[3] , \nScanOut567[2] , 
        \nScanOut567[1] , \nScanOut567[0] }), .ScanOut({\nScanOut566[7] , 
        \nScanOut566[6] , \nScanOut566[5] , \nScanOut566[4] , \nScanOut566[3] , 
        \nScanOut566[2] , \nScanOut566[1] , \nScanOut566[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_21[7] , \nOut17_21[6] , \nOut17_21[5] , \nOut17_21[4] , 
        \nOut17_21[3] , \nOut17_21[2] , \nOut17_21[1] , \nOut17_21[0] }), 
        .SouthIn({\nOut17_23[7] , \nOut17_23[6] , \nOut17_23[5] , 
        \nOut17_23[4] , \nOut17_23[3] , \nOut17_23[2] , \nOut17_23[1] , 
        \nOut17_23[0] }), .EastIn({\nOut18_22[7] , \nOut18_22[6] , 
        \nOut18_22[5] , \nOut18_22[4] , \nOut18_22[3] , \nOut18_22[2] , 
        \nOut18_22[1] , \nOut18_22[0] }), .WestIn({\nOut16_22[7] , 
        \nOut16_22[6] , \nOut16_22[5] , \nOut16_22[4] , \nOut16_22[3] , 
        \nOut16_22[2] , \nOut16_22[1] , \nOut16_22[0] }), .Out({\nOut17_22[7] , 
        \nOut17_22[6] , \nOut17_22[5] , \nOut17_22[4] , \nOut17_22[3] , 
        \nOut17_22[2] , \nOut17_22[1] , \nOut17_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_933 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut934[7] , \nScanOut934[6] , 
        \nScanOut934[5] , \nScanOut934[4] , \nScanOut934[3] , \nScanOut934[2] , 
        \nScanOut934[1] , \nScanOut934[0] }), .ScanOut({\nScanOut933[7] , 
        \nScanOut933[6] , \nScanOut933[5] , \nScanOut933[4] , \nScanOut933[3] , 
        \nScanOut933[2] , \nScanOut933[1] , \nScanOut933[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_4[7] , \nOut29_4[6] , \nOut29_4[5] , \nOut29_4[4] , 
        \nOut29_4[3] , \nOut29_4[2] , \nOut29_4[1] , \nOut29_4[0] }), 
        .SouthIn({\nOut29_6[7] , \nOut29_6[6] , \nOut29_6[5] , \nOut29_6[4] , 
        \nOut29_6[3] , \nOut29_6[2] , \nOut29_6[1] , \nOut29_6[0] }), .EastIn(
        {\nOut30_5[7] , \nOut30_5[6] , \nOut30_5[5] , \nOut30_5[4] , 
        \nOut30_5[3] , \nOut30_5[2] , \nOut30_5[1] , \nOut30_5[0] }), .WestIn(
        {\nOut28_5[7] , \nOut28_5[6] , \nOut28_5[5] , \nOut28_5[4] , 
        \nOut28_5[3] , \nOut28_5[2] , \nOut28_5[1] , \nOut28_5[0] }), .Out({
        \nOut29_5[7] , \nOut29_5[6] , \nOut29_5[5] , \nOut29_5[4] , 
        \nOut29_5[3] , \nOut29_5[2] , \nOut29_5[1] , \nOut29_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_81 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut82[7] , \nScanOut82[6] , 
        \nScanOut82[5] , \nScanOut82[4] , \nScanOut82[3] , \nScanOut82[2] , 
        \nScanOut82[1] , \nScanOut82[0] }), .ScanOut({\nScanOut81[7] , 
        \nScanOut81[6] , \nScanOut81[5] , \nScanOut81[4] , \nScanOut81[3] , 
        \nScanOut81[2] , \nScanOut81[1] , \nScanOut81[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_16[7] , \nOut2_16[6] , \nOut2_16[5] , \nOut2_16[4] , 
        \nOut2_16[3] , \nOut2_16[2] , \nOut2_16[1] , \nOut2_16[0] }), 
        .SouthIn({\nOut2_18[7] , \nOut2_18[6] , \nOut2_18[5] , \nOut2_18[4] , 
        \nOut2_18[3] , \nOut2_18[2] , \nOut2_18[1] , \nOut2_18[0] }), .EastIn(
        {\nOut3_17[7] , \nOut3_17[6] , \nOut3_17[5] , \nOut3_17[4] , 
        \nOut3_17[3] , \nOut3_17[2] , \nOut3_17[1] , \nOut3_17[0] }), .WestIn(
        {\nOut1_17[7] , \nOut1_17[6] , \nOut1_17[5] , \nOut1_17[4] , 
        \nOut1_17[3] , \nOut1_17[2] , \nOut1_17[1] , \nOut1_17[0] }), .Out({
        \nOut2_17[7] , \nOut2_17[6] , \nOut2_17[5] , \nOut2_17[4] , 
        \nOut2_17[3] , \nOut2_17[2] , \nOut2_17[1] , \nOut2_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_115 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut116[7] , \nScanOut116[6] , 
        \nScanOut116[5] , \nScanOut116[4] , \nScanOut116[3] , \nScanOut116[2] , 
        \nScanOut116[1] , \nScanOut116[0] }), .ScanOut({\nScanOut115[7] , 
        \nScanOut115[6] , \nScanOut115[5] , \nScanOut115[4] , \nScanOut115[3] , 
        \nScanOut115[2] , \nScanOut115[1] , \nScanOut115[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_18[7] , \nOut3_18[6] , \nOut3_18[5] , \nOut3_18[4] , 
        \nOut3_18[3] , \nOut3_18[2] , \nOut3_18[1] , \nOut3_18[0] }), 
        .SouthIn({\nOut3_20[7] , \nOut3_20[6] , \nOut3_20[5] , \nOut3_20[4] , 
        \nOut3_20[3] , \nOut3_20[2] , \nOut3_20[1] , \nOut3_20[0] }), .EastIn(
        {\nOut4_19[7] , \nOut4_19[6] , \nOut4_19[5] , \nOut4_19[4] , 
        \nOut4_19[3] , \nOut4_19[2] , \nOut4_19[1] , \nOut4_19[0] }), .WestIn(
        {\nOut2_19[7] , \nOut2_19[6] , \nOut2_19[5] , \nOut2_19[4] , 
        \nOut2_19[3] , \nOut2_19[2] , \nOut2_19[1] , \nOut2_19[0] }), .Out({
        \nOut3_19[7] , \nOut3_19[6] , \nOut3_19[5] , \nOut3_19[4] , 
        \nOut3_19[3] , \nOut3_19[2] , \nOut3_19[1] , \nOut3_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_225 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut226[7] , \nScanOut226[6] , 
        \nScanOut226[5] , \nScanOut226[4] , \nScanOut226[3] , \nScanOut226[2] , 
        \nScanOut226[1] , \nScanOut226[0] }), .ScanOut({\nScanOut225[7] , 
        \nScanOut225[6] , \nScanOut225[5] , \nScanOut225[4] , \nScanOut225[3] , 
        \nScanOut225[2] , \nScanOut225[1] , \nScanOut225[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_0[7] , \nOut7_0[6] , \nOut7_0[5] , \nOut7_0[4] , \nOut7_0[3] , 
        \nOut7_0[2] , \nOut7_0[1] , \nOut7_0[0] }), .SouthIn({\nOut7_2[7] , 
        \nOut7_2[6] , \nOut7_2[5] , \nOut7_2[4] , \nOut7_2[3] , \nOut7_2[2] , 
        \nOut7_2[1] , \nOut7_2[0] }), .EastIn({\nOut8_1[7] , \nOut8_1[6] , 
        \nOut8_1[5] , \nOut8_1[4] , \nOut8_1[3] , \nOut8_1[2] , \nOut8_1[1] , 
        \nOut8_1[0] }), .WestIn({\nOut6_1[7] , \nOut6_1[6] , \nOut6_1[5] , 
        \nOut6_1[4] , \nOut6_1[3] , \nOut6_1[2] , \nOut6_1[1] , \nOut6_1[0] }), 
        .Out({\nOut7_1[7] , \nOut7_1[6] , \nOut7_1[5] , \nOut7_1[4] , 
        \nOut7_1[3] , \nOut7_1[2] , \nOut7_1[1] , \nOut7_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_434 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut435[7] , \nScanOut435[6] , 
        \nScanOut435[5] , \nScanOut435[4] , \nScanOut435[3] , \nScanOut435[2] , 
        \nScanOut435[1] , \nScanOut435[0] }), .ScanOut({\nScanOut434[7] , 
        \nScanOut434[6] , \nScanOut434[5] , \nScanOut434[4] , \nScanOut434[3] , 
        \nScanOut434[2] , \nScanOut434[1] , \nScanOut434[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_17[7] , \nOut13_17[6] , \nOut13_17[5] , \nOut13_17[4] , 
        \nOut13_17[3] , \nOut13_17[2] , \nOut13_17[1] , \nOut13_17[0] }), 
        .SouthIn({\nOut13_19[7] , \nOut13_19[6] , \nOut13_19[5] , 
        \nOut13_19[4] , \nOut13_19[3] , \nOut13_19[2] , \nOut13_19[1] , 
        \nOut13_19[0] }), .EastIn({\nOut14_18[7] , \nOut14_18[6] , 
        \nOut14_18[5] , \nOut14_18[4] , \nOut14_18[3] , \nOut14_18[2] , 
        \nOut14_18[1] , \nOut14_18[0] }), .WestIn({\nOut12_18[7] , 
        \nOut12_18[6] , \nOut12_18[5] , \nOut12_18[4] , \nOut12_18[3] , 
        \nOut12_18[2] , \nOut12_18[1] , \nOut12_18[0] }), .Out({\nOut13_18[7] , 
        \nOut13_18[6] , \nOut13_18[5] , \nOut13_18[4] , \nOut13_18[3] , 
        \nOut13_18[2] , \nOut13_18[1] , \nOut13_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_671 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut672[7] , \nScanOut672[6] , 
        \nScanOut672[5] , \nScanOut672[4] , \nScanOut672[3] , \nScanOut672[2] , 
        \nScanOut672[1] , \nScanOut672[0] }), .ScanOut({\nScanOut671[7] , 
        \nScanOut671[6] , \nScanOut671[5] , \nScanOut671[4] , \nScanOut671[3] , 
        \nScanOut671[2] , \nScanOut671[1] , \nScanOut671[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut20_31[7] , \nOut20_31[6] , 
        \nOut20_31[5] , \nOut20_31[4] , \nOut20_31[3] , \nOut20_31[2] , 
        \nOut20_31[1] , \nOut20_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_828 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut829[7] , \nScanOut829[6] , 
        \nScanOut829[5] , \nScanOut829[4] , \nScanOut829[3] , \nScanOut829[2] , 
        \nScanOut829[1] , \nScanOut829[0] }), .ScanOut({\nScanOut828[7] , 
        \nScanOut828[6] , \nScanOut828[5] , \nScanOut828[4] , \nScanOut828[3] , 
        \nScanOut828[2] , \nScanOut828[1] , \nScanOut828[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_27[7] , \nOut25_27[6] , \nOut25_27[5] , \nOut25_27[4] , 
        \nOut25_27[3] , \nOut25_27[2] , \nOut25_27[1] , \nOut25_27[0] }), 
        .SouthIn({\nOut25_29[7] , \nOut25_29[6] , \nOut25_29[5] , 
        \nOut25_29[4] , \nOut25_29[3] , \nOut25_29[2] , \nOut25_29[1] , 
        \nOut25_29[0] }), .EastIn({\nOut26_28[7] , \nOut26_28[6] , 
        \nOut26_28[5] , \nOut26_28[4] , \nOut26_28[3] , \nOut26_28[2] , 
        \nOut26_28[1] , \nOut26_28[0] }), .WestIn({\nOut24_28[7] , 
        \nOut24_28[6] , \nOut24_28[5] , \nOut24_28[4] , \nOut24_28[3] , 
        \nOut24_28[2] , \nOut24_28[1] , \nOut24_28[0] }), .Out({\nOut25_28[7] , 
        \nOut25_28[6] , \nOut25_28[5] , \nOut25_28[4] , \nOut25_28[3] , 
        \nOut25_28[2] , \nOut25_28[1] , \nOut25_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_846 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut847[7] , \nScanOut847[6] , 
        \nScanOut847[5] , \nScanOut847[4] , \nScanOut847[3] , \nScanOut847[2] , 
        \nScanOut847[1] , \nScanOut847[0] }), .ScanOut({\nScanOut846[7] , 
        \nScanOut846[6] , \nScanOut846[5] , \nScanOut846[4] , \nScanOut846[3] , 
        \nScanOut846[2] , \nScanOut846[1] , \nScanOut846[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_13[7] , \nOut26_13[6] , \nOut26_13[5] , \nOut26_13[4] , 
        \nOut26_13[3] , \nOut26_13[2] , \nOut26_13[1] , \nOut26_13[0] }), 
        .SouthIn({\nOut26_15[7] , \nOut26_15[6] , \nOut26_15[5] , 
        \nOut26_15[4] , \nOut26_15[3] , \nOut26_15[2] , \nOut26_15[1] , 
        \nOut26_15[0] }), .EastIn({\nOut27_14[7] , \nOut27_14[6] , 
        \nOut27_14[5] , \nOut27_14[4] , \nOut27_14[3] , \nOut27_14[2] , 
        \nOut27_14[1] , \nOut27_14[0] }), .WestIn({\nOut25_14[7] , 
        \nOut25_14[6] , \nOut25_14[5] , \nOut25_14[4] , \nOut25_14[3] , 
        \nOut25_14[2] , \nOut25_14[1] , \nOut25_14[0] }), .Out({\nOut26_14[7] , 
        \nOut26_14[6] , \nOut26_14[5] , \nOut26_14[4] , \nOut26_14[3] , 
        \nOut26_14[2] , \nOut26_14[1] , \nOut26_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_694 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut695[7] , \nScanOut695[6] , 
        \nScanOut695[5] , \nScanOut695[4] , \nScanOut695[3] , \nScanOut695[2] , 
        \nScanOut695[1] , \nScanOut695[0] }), .ScanOut({\nScanOut694[7] , 
        \nScanOut694[6] , \nScanOut694[5] , \nScanOut694[4] , \nScanOut694[3] , 
        \nScanOut694[2] , \nScanOut694[1] , \nScanOut694[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_21[7] , \nOut21_21[6] , \nOut21_21[5] , \nOut21_21[4] , 
        \nOut21_21[3] , \nOut21_21[2] , \nOut21_21[1] , \nOut21_21[0] }), 
        .SouthIn({\nOut21_23[7] , \nOut21_23[6] , \nOut21_23[5] , 
        \nOut21_23[4] , \nOut21_23[3] , \nOut21_23[2] , \nOut21_23[1] , 
        \nOut21_23[0] }), .EastIn({\nOut22_22[7] , \nOut22_22[6] , 
        \nOut22_22[5] , \nOut22_22[4] , \nOut22_22[3] , \nOut22_22[2] , 
        \nOut22_22[1] , \nOut22_22[0] }), .WestIn({\nOut20_22[7] , 
        \nOut20_22[6] , \nOut20_22[5] , \nOut20_22[4] , \nOut20_22[3] , 
        \nOut20_22[2] , \nOut20_22[1] , \nOut20_22[0] }), .Out({\nOut21_22[7] , 
        \nOut21_22[6] , \nOut21_22[5] , \nOut21_22[4] , \nOut21_22[3] , 
        \nOut21_22[2] , \nOut21_22[1] , \nOut21_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_704 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut705[7] , \nScanOut705[6] , 
        \nScanOut705[5] , \nScanOut705[4] , \nScanOut705[3] , \nScanOut705[2] , 
        \nScanOut705[1] , \nScanOut705[0] }), .ScanOut({\nScanOut704[7] , 
        \nScanOut704[6] , \nScanOut704[5] , \nScanOut704[4] , \nScanOut704[3] , 
        \nScanOut704[2] , \nScanOut704[1] , \nScanOut704[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut22_0[7] , \nOut22_0[6] , 
        \nOut22_0[5] , \nOut22_0[4] , \nOut22_0[3] , \nOut22_0[2] , 
        \nOut22_0[1] , \nOut22_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1002 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1003[7] , \nScanOut1003[6] , 
        \nScanOut1003[5] , \nScanOut1003[4] , \nScanOut1003[3] , 
        \nScanOut1003[2] , \nScanOut1003[1] , \nScanOut1003[0] }), .ScanOut({
        \nScanOut1002[7] , \nScanOut1002[6] , \nScanOut1002[5] , 
        \nScanOut1002[4] , \nScanOut1002[3] , \nScanOut1002[2] , 
        \nScanOut1002[1] , \nScanOut1002[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_10[7] , \nOut31_10[6] , \nOut31_10[5] , 
        \nOut31_10[4] , \nOut31_10[3] , \nOut31_10[2] , \nOut31_10[1] , 
        \nOut31_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_132 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut133[7] , \nScanOut133[6] , 
        \nScanOut133[5] , \nScanOut133[4] , \nScanOut133[3] , \nScanOut133[2] , 
        \nScanOut133[1] , \nScanOut133[0] }), .ScanOut({\nScanOut132[7] , 
        \nScanOut132[6] , \nScanOut132[5] , \nScanOut132[4] , \nScanOut132[3] , 
        \nScanOut132[2] , \nScanOut132[1] , \nScanOut132[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_3[7] , \nOut4_3[6] , \nOut4_3[5] , \nOut4_3[4] , \nOut4_3[3] , 
        \nOut4_3[2] , \nOut4_3[1] , \nOut4_3[0] }), .SouthIn({\nOut4_5[7] , 
        \nOut4_5[6] , \nOut4_5[5] , \nOut4_5[4] , \nOut4_5[3] , \nOut4_5[2] , 
        \nOut4_5[1] , \nOut4_5[0] }), .EastIn({\nOut5_4[7] , \nOut5_4[6] , 
        \nOut5_4[5] , \nOut5_4[4] , \nOut5_4[3] , \nOut5_4[2] , \nOut5_4[1] , 
        \nOut5_4[0] }), .WestIn({\nOut3_4[7] , \nOut3_4[6] , \nOut3_4[5] , 
        \nOut3_4[4] , \nOut3_4[3] , \nOut3_4[2] , \nOut3_4[1] , \nOut3_4[0] }), 
        .Out({\nOut4_4[7] , \nOut4_4[6] , \nOut4_4[5] , \nOut4_4[4] , 
        \nOut4_4[3] , \nOut4_4[2] , \nOut4_4[1] , \nOut4_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_195 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut196[7] , \nScanOut196[6] , 
        \nScanOut196[5] , \nScanOut196[4] , \nScanOut196[3] , \nScanOut196[2] , 
        \nScanOut196[1] , \nScanOut196[0] }), .ScanOut({\nScanOut195[7] , 
        \nScanOut195[6] , \nScanOut195[5] , \nScanOut195[4] , \nScanOut195[3] , 
        \nScanOut195[2] , \nScanOut195[1] , \nScanOut195[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_2[7] , \nOut6_2[6] , \nOut6_2[5] , \nOut6_2[4] , \nOut6_2[3] , 
        \nOut6_2[2] , \nOut6_2[1] , \nOut6_2[0] }), .SouthIn({\nOut6_4[7] , 
        \nOut6_4[6] , \nOut6_4[5] , \nOut6_4[4] , \nOut6_4[3] , \nOut6_4[2] , 
        \nOut6_4[1] , \nOut6_4[0] }), .EastIn({\nOut7_3[7] , \nOut7_3[6] , 
        \nOut7_3[5] , \nOut7_3[4] , \nOut7_3[3] , \nOut7_3[2] , \nOut7_3[1] , 
        \nOut7_3[0] }), .WestIn({\nOut5_3[7] , \nOut5_3[6] , \nOut5_3[5] , 
        \nOut5_3[4] , \nOut5_3[3] , \nOut5_3[2] , \nOut5_3[1] , \nOut5_3[0] }), 
        .Out({\nOut6_3[7] , \nOut6_3[6] , \nOut6_3[5] , \nOut6_3[4] , 
        \nOut6_3[3] , \nOut6_3[2] , \nOut6_3[1] , \nOut6_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_202 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut203[7] , \nScanOut203[6] , 
        \nScanOut203[5] , \nScanOut203[4] , \nScanOut203[3] , \nScanOut203[2] , 
        \nScanOut203[1] , \nScanOut203[0] }), .ScanOut({\nScanOut202[7] , 
        \nScanOut202[6] , \nScanOut202[5] , \nScanOut202[4] , \nScanOut202[3] , 
        \nScanOut202[2] , \nScanOut202[1] , \nScanOut202[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_9[7] , \nOut6_9[6] , \nOut6_9[5] , \nOut6_9[4] , \nOut6_9[3] , 
        \nOut6_9[2] , \nOut6_9[1] , \nOut6_9[0] }), .SouthIn({\nOut6_11[7] , 
        \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , \nOut6_11[3] , 
        \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }), .EastIn({\nOut7_10[7] , 
        \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , \nOut7_10[3] , 
        \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }), .WestIn({\nOut5_10[7] , 
        \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , \nOut5_10[3] , 
        \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }), .Out({\nOut6_10[7] , 
        \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , \nOut6_10[3] , 
        \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_723 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut724[7] , \nScanOut724[6] , 
        \nScanOut724[5] , \nScanOut724[4] , \nScanOut724[3] , \nScanOut724[2] , 
        \nScanOut724[1] , \nScanOut724[0] }), .ScanOut({\nScanOut723[7] , 
        \nScanOut723[6] , \nScanOut723[5] , \nScanOut723[4] , \nScanOut723[3] , 
        \nScanOut723[2] , \nScanOut723[1] , \nScanOut723[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_18[7] , \nOut22_18[6] , \nOut22_18[5] , \nOut22_18[4] , 
        \nOut22_18[3] , \nOut22_18[2] , \nOut22_18[1] , \nOut22_18[0] }), 
        .SouthIn({\nOut22_20[7] , \nOut22_20[6] , \nOut22_20[5] , 
        \nOut22_20[4] , \nOut22_20[3] , \nOut22_20[2] , \nOut22_20[1] , 
        \nOut22_20[0] }), .EastIn({\nOut23_19[7] , \nOut23_19[6] , 
        \nOut23_19[5] , \nOut23_19[4] , \nOut23_19[3] , \nOut23_19[2] , 
        \nOut23_19[1] , \nOut23_19[0] }), .WestIn({\nOut21_19[7] , 
        \nOut21_19[6] , \nOut21_19[5] , \nOut21_19[4] , \nOut21_19[3] , 
        \nOut21_19[2] , \nOut21_19[1] , \nOut21_19[0] }), .Out({\nOut22_19[7] , 
        \nOut22_19[6] , \nOut22_19[5] , \nOut22_19[4] , \nOut22_19[3] , 
        \nOut22_19[2] , \nOut22_19[1] , \nOut22_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_861 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut862[7] , \nScanOut862[6] , 
        \nScanOut862[5] , \nScanOut862[4] , \nScanOut862[3] , \nScanOut862[2] , 
        \nScanOut862[1] , \nScanOut862[0] }), .ScanOut({\nScanOut861[7] , 
        \nScanOut861[6] , \nScanOut861[5] , \nScanOut861[4] , \nScanOut861[3] , 
        \nScanOut861[2] , \nScanOut861[1] , \nScanOut861[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_28[7] , \nOut26_28[6] , \nOut26_28[5] , \nOut26_28[4] , 
        \nOut26_28[3] , \nOut26_28[2] , \nOut26_28[1] , \nOut26_28[0] }), 
        .SouthIn({\nOut26_30[7] , \nOut26_30[6] , \nOut26_30[5] , 
        \nOut26_30[4] , \nOut26_30[3] , \nOut26_30[2] , \nOut26_30[1] , 
        \nOut26_30[0] }), .EastIn({\nOut27_29[7] , \nOut27_29[6] , 
        \nOut27_29[5] , \nOut27_29[4] , \nOut27_29[3] , \nOut27_29[2] , 
        \nOut27_29[1] , \nOut27_29[0] }), .WestIn({\nOut25_29[7] , 
        \nOut25_29[6] , \nOut25_29[5] , \nOut25_29[4] , \nOut25_29[3] , 
        \nOut25_29[2] , \nOut25_29[1] , \nOut25_29[0] }), .Out({\nOut26_29[7] , 
        \nOut26_29[6] , \nOut26_29[5] , \nOut26_29[4] , \nOut26_29[3] , 
        \nOut26_29[2] , \nOut26_29[1] , \nOut26_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_289 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut290[7] , \nScanOut290[6] , 
        \nScanOut290[5] , \nScanOut290[4] , \nScanOut290[3] , \nScanOut290[2] , 
        \nScanOut290[1] , \nScanOut290[0] }), .ScanOut({\nScanOut289[7] , 
        \nScanOut289[6] , \nScanOut289[5] , \nScanOut289[4] , \nScanOut289[3] , 
        \nScanOut289[2] , \nScanOut289[1] , \nScanOut289[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_0[7] , \nOut9_0[6] , \nOut9_0[5] , \nOut9_0[4] , \nOut9_0[3] , 
        \nOut9_0[2] , \nOut9_0[1] , \nOut9_0[0] }), .SouthIn({\nOut9_2[7] , 
        \nOut9_2[6] , \nOut9_2[5] , \nOut9_2[4] , \nOut9_2[3] , \nOut9_2[2] , 
        \nOut9_2[1] , \nOut9_2[0] }), .EastIn({\nOut10_1[7] , \nOut10_1[6] , 
        \nOut10_1[5] , \nOut10_1[4] , \nOut10_1[3] , \nOut10_1[2] , 
        \nOut10_1[1] , \nOut10_1[0] }), .WestIn({\nOut8_1[7] , \nOut8_1[6] , 
        \nOut8_1[5] , \nOut8_1[4] , \nOut8_1[3] , \nOut8_1[2] , \nOut8_1[1] , 
        \nOut8_1[0] }), .Out({\nOut9_1[7] , \nOut9_1[6] , \nOut9_1[5] , 
        \nOut9_1[4] , \nOut9_1[3] , \nOut9_1[2] , \nOut9_1[1] , \nOut9_1[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_392 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut393[7] , \nScanOut393[6] , 
        \nScanOut393[5] , \nScanOut393[4] , \nScanOut393[3] , \nScanOut393[2] , 
        \nScanOut393[1] , \nScanOut393[0] }), .ScanOut({\nScanOut392[7] , 
        \nScanOut392[6] , \nScanOut392[5] , \nScanOut392[4] , \nScanOut392[3] , 
        \nScanOut392[2] , \nScanOut392[1] , \nScanOut392[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }), 
        .SouthIn({\nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , \nOut12_9[4] , 
        \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , \nOut12_9[0] }), .EastIn(
        {\nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }), .WestIn(
        {\nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }), .Out({
        \nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_583 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut584[7] , \nScanOut584[6] , 
        \nScanOut584[5] , \nScanOut584[4] , \nScanOut584[3] , \nScanOut584[2] , 
        \nScanOut584[1] , \nScanOut584[0] }), .ScanOut({\nScanOut583[7] , 
        \nScanOut583[6] , \nScanOut583[5] , \nScanOut583[4] , \nScanOut583[3] , 
        \nScanOut583[2] , \nScanOut583[1] , \nScanOut583[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_6[7] , \nOut18_6[6] , \nOut18_6[5] , \nOut18_6[4] , 
        \nOut18_6[3] , \nOut18_6[2] , \nOut18_6[1] , \nOut18_6[0] }), 
        .SouthIn({\nOut18_8[7] , \nOut18_8[6] , \nOut18_8[5] , \nOut18_8[4] , 
        \nOut18_8[3] , \nOut18_8[2] , \nOut18_8[1] , \nOut18_8[0] }), .EastIn(
        {\nOut19_7[7] , \nOut19_7[6] , \nOut19_7[5] , \nOut19_7[4] , 
        \nOut19_7[3] , \nOut19_7[2] , \nOut19_7[1] , \nOut19_7[0] }), .WestIn(
        {\nOut17_7[7] , \nOut17_7[6] , \nOut17_7[5] , \nOut17_7[4] , 
        \nOut17_7[3] , \nOut17_7[2] , \nOut17_7[1] , \nOut17_7[0] }), .Out({
        \nOut18_7[7] , \nOut18_7[6] , \nOut18_7[5] , \nOut18_7[4] , 
        \nOut18_7[3] , \nOut18_7[2] , \nOut18_7[1] , \nOut18_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_413 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut414[7] , \nScanOut414[6] , 
        \nScanOut414[5] , \nScanOut414[4] , \nScanOut414[3] , \nScanOut414[2] , 
        \nScanOut414[1] , \nScanOut414[0] }), .ScanOut({\nScanOut413[7] , 
        \nScanOut413[6] , \nScanOut413[5] , \nScanOut413[4] , \nScanOut413[3] , 
        \nScanOut413[2] , \nScanOut413[1] , \nScanOut413[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_28[7] , \nOut12_28[6] , \nOut12_28[5] , \nOut12_28[4] , 
        \nOut12_28[3] , \nOut12_28[2] , \nOut12_28[1] , \nOut12_28[0] }), 
        .SouthIn({\nOut12_30[7] , \nOut12_30[6] , \nOut12_30[5] , 
        \nOut12_30[4] , \nOut12_30[3] , \nOut12_30[2] , \nOut12_30[1] , 
        \nOut12_30[0] }), .EastIn({\nOut13_29[7] , \nOut13_29[6] , 
        \nOut13_29[5] , \nOut13_29[4] , \nOut13_29[3] , \nOut13_29[2] , 
        \nOut13_29[1] , \nOut13_29[0] }), .WestIn({\nOut11_29[7] , 
        \nOut11_29[6] , \nOut11_29[5] , \nOut11_29[4] , \nOut11_29[3] , 
        \nOut11_29[2] , \nOut11_29[1] , \nOut11_29[0] }), .Out({\nOut12_29[7] , 
        \nOut12_29[6] , \nOut12_29[5] , \nOut12_29[4] , \nOut12_29[3] , 
        \nOut12_29[2] , \nOut12_29[1] , \nOut12_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_638 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut639[7] , \nScanOut639[6] , 
        \nScanOut639[5] , \nScanOut639[4] , \nScanOut639[3] , \nScanOut639[2] , 
        \nScanOut639[1] , \nScanOut639[0] }), .ScanOut({\nScanOut638[7] , 
        \nScanOut638[6] , \nScanOut638[5] , \nScanOut638[4] , \nScanOut638[3] , 
        \nScanOut638[2] , \nScanOut638[1] , \nScanOut638[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_29[7] , \nOut19_29[6] , \nOut19_29[5] , \nOut19_29[4] , 
        \nOut19_29[3] , \nOut19_29[2] , \nOut19_29[1] , \nOut19_29[0] }), 
        .SouthIn({\nOut19_31[7] , \nOut19_31[6] , \nOut19_31[5] , 
        \nOut19_31[4] , \nOut19_31[3] , \nOut19_31[2] , \nOut19_31[1] , 
        \nOut19_31[0] }), .EastIn({\nOut20_30[7] , \nOut20_30[6] , 
        \nOut20_30[5] , \nOut20_30[4] , \nOut20_30[3] , \nOut20_30[2] , 
        \nOut20_30[1] , \nOut20_30[0] }), .WestIn({\nOut18_30[7] , 
        \nOut18_30[6] , \nOut18_30[5] , \nOut18_30[4] , \nOut18_30[3] , 
        \nOut18_30[2] , \nOut18_30[1] , \nOut18_30[0] }), .Out({\nOut19_30[7] , 
        \nOut19_30[6] , \nOut19_30[5] , \nOut19_30[4] , \nOut19_30[3] , 
        \nOut19_30[2] , \nOut19_30[1] , \nOut19_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_319 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut320[7] , \nScanOut320[6] , 
        \nScanOut320[5] , \nScanOut320[4] , \nScanOut320[3] , \nScanOut320[2] , 
        \nScanOut320[1] , \nScanOut320[0] }), .ScanOut({\nScanOut319[7] , 
        \nScanOut319[6] , \nScanOut319[5] , \nScanOut319[4] , \nScanOut319[3] , 
        \nScanOut319[2] , \nScanOut319[1] , \nScanOut319[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut9_31[7] , \nOut9_31[6] , 
        \nOut9_31[5] , \nOut9_31[4] , \nOut9_31[3] , \nOut9_31[2] , 
        \nOut9_31[1] , \nOut9_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_508 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut509[7] , \nScanOut509[6] , 
        \nScanOut509[5] , \nScanOut509[4] , \nScanOut509[3] , \nScanOut509[2] , 
        \nScanOut509[1] , \nScanOut509[0] }), .ScanOut({\nScanOut508[7] , 
        \nScanOut508[6] , \nScanOut508[5] , \nScanOut508[4] , \nScanOut508[3] , 
        \nScanOut508[2] , \nScanOut508[1] , \nScanOut508[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_27[7] , \nOut15_27[6] , \nOut15_27[5] , \nOut15_27[4] , 
        \nOut15_27[3] , \nOut15_27[2] , \nOut15_27[1] , \nOut15_27[0] }), 
        .SouthIn({\nOut15_29[7] , \nOut15_29[6] , \nOut15_29[5] , 
        \nOut15_29[4] , \nOut15_29[3] , \nOut15_29[2] , \nOut15_29[1] , 
        \nOut15_29[0] }), .EastIn({\nOut16_28[7] , \nOut16_28[6] , 
        \nOut16_28[5] , \nOut16_28[4] , \nOut16_28[3] , \nOut16_28[2] , 
        \nOut16_28[1] , \nOut16_28[0] }), .WestIn({\nOut14_28[7] , 
        \nOut14_28[6] , \nOut14_28[5] , \nOut14_28[4] , \nOut14_28[3] , 
        \nOut14_28[2] , \nOut14_28[1] , \nOut14_28[0] }), .Out({\nOut15_28[7] , 
        \nOut15_28[6] , \nOut15_28[5] , \nOut15_28[4] , \nOut15_28[3] , 
        \nOut15_28[2] , \nOut15_28[1] , \nOut15_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_498 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut499[7] , \nScanOut499[6] , 
        \nScanOut499[5] , \nScanOut499[4] , \nScanOut499[3] , \nScanOut499[2] , 
        \nScanOut499[1] , \nScanOut499[0] }), .ScanOut({\nScanOut498[7] , 
        \nScanOut498[6] , \nScanOut498[5] , \nScanOut498[4] , \nScanOut498[3] , 
        \nScanOut498[2] , \nScanOut498[1] , \nScanOut498[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_17[7] , \nOut15_17[6] , \nOut15_17[5] , \nOut15_17[4] , 
        \nOut15_17[3] , \nOut15_17[2] , \nOut15_17[1] , \nOut15_17[0] }), 
        .SouthIn({\nOut15_19[7] , \nOut15_19[6] , \nOut15_19[5] , 
        \nOut15_19[4] , \nOut15_19[3] , \nOut15_19[2] , \nOut15_19[1] , 
        \nOut15_19[0] }), .EastIn({\nOut16_18[7] , \nOut16_18[6] , 
        \nOut16_18[5] , \nOut16_18[4] , \nOut16_18[3] , \nOut16_18[2] , 
        \nOut16_18[1] , \nOut16_18[0] }), .WestIn({\nOut14_18[7] , 
        \nOut14_18[6] , \nOut14_18[5] , \nOut14_18[4] , \nOut14_18[3] , 
        \nOut14_18[2] , \nOut14_18[1] , \nOut14_18[0] }), .Out({\nOut15_18[7] , 
        \nOut15_18[6] , \nOut15_18[5] , \nOut15_18[4] , \nOut15_18[3] , 
        \nOut15_18[2] , \nOut15_18[1] , \nOut15_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_614 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut615[7] , \nScanOut615[6] , 
        \nScanOut615[5] , \nScanOut615[4] , \nScanOut615[3] , \nScanOut615[2] , 
        \nScanOut615[1] , \nScanOut615[0] }), .ScanOut({\nScanOut614[7] , 
        \nScanOut614[6] , \nScanOut614[5] , \nScanOut614[4] , \nScanOut614[3] , 
        \nScanOut614[2] , \nScanOut614[1] , \nScanOut614[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_5[7] , \nOut19_5[6] , \nOut19_5[5] , \nOut19_5[4] , 
        \nOut19_5[3] , \nOut19_5[2] , \nOut19_5[1] , \nOut19_5[0] }), 
        .SouthIn({\nOut19_7[7] , \nOut19_7[6] , \nOut19_7[5] , \nOut19_7[4] , 
        \nOut19_7[3] , \nOut19_7[2] , \nOut19_7[1] , \nOut19_7[0] }), .EastIn(
        {\nOut20_6[7] , \nOut20_6[6] , \nOut20_6[5] , \nOut20_6[4] , 
        \nOut20_6[3] , \nOut20_6[2] , \nOut20_6[1] , \nOut20_6[0] }), .WestIn(
        {\nOut18_6[7] , \nOut18_6[6] , \nOut18_6[5] , \nOut18_6[4] , 
        \nOut18_6[3] , \nOut18_6[2] , \nOut18_6[1] , \nOut18_6[0] }), .Out({
        \nOut19_6[7] , \nOut19_6[6] , \nOut19_6[5] , \nOut19_6[4] , 
        \nOut19_6[3] , \nOut19_6[2] , \nOut19_6[1] , \nOut19_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_282 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut283[7] , \nScanOut283[6] , 
        \nScanOut283[5] , \nScanOut283[4] , \nScanOut283[3] , \nScanOut283[2] , 
        \nScanOut283[1] , \nScanOut283[0] }), .ScanOut({\nScanOut282[7] , 
        \nScanOut282[6] , \nScanOut282[5] , \nScanOut282[4] , \nScanOut282[3] , 
        \nScanOut282[2] , \nScanOut282[1] , \nScanOut282[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_25[7] , \nOut8_25[6] , \nOut8_25[5] , \nOut8_25[4] , 
        \nOut8_25[3] , \nOut8_25[2] , \nOut8_25[1] , \nOut8_25[0] }), 
        .SouthIn({\nOut8_27[7] , \nOut8_27[6] , \nOut8_27[5] , \nOut8_27[4] , 
        \nOut8_27[3] , \nOut8_27[2] , \nOut8_27[1] , \nOut8_27[0] }), .EastIn(
        {\nOut9_26[7] , \nOut9_26[6] , \nOut9_26[5] , \nOut9_26[4] , 
        \nOut9_26[3] , \nOut9_26[2] , \nOut9_26[1] , \nOut9_26[0] }), .WestIn(
        {\nOut7_26[7] , \nOut7_26[6] , \nOut7_26[5] , \nOut7_26[4] , 
        \nOut7_26[3] , \nOut7_26[2] , \nOut7_26[1] , \nOut7_26[0] }), .Out({
        \nOut8_26[7] , \nOut8_26[6] , \nOut8_26[5] , \nOut8_26[4] , 
        \nOut8_26[3] , \nOut8_26[2] , \nOut8_26[1] , \nOut8_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_312 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut313[7] , \nScanOut313[6] , 
        \nScanOut313[5] , \nScanOut313[4] , \nScanOut313[3] , \nScanOut313[2] , 
        \nScanOut313[1] , \nScanOut313[0] }), .ScanOut({\nScanOut312[7] , 
        \nScanOut312[6] , \nScanOut312[5] , \nScanOut312[4] , \nScanOut312[3] , 
        \nScanOut312[2] , \nScanOut312[1] , \nScanOut312[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_23[7] , \nOut9_23[6] , \nOut9_23[5] , \nOut9_23[4] , 
        \nOut9_23[3] , \nOut9_23[2] , \nOut9_23[1] , \nOut9_23[0] }), 
        .SouthIn({\nOut9_25[7] , \nOut9_25[6] , \nOut9_25[5] , \nOut9_25[4] , 
        \nOut9_25[3] , \nOut9_25[2] , \nOut9_25[1] , \nOut9_25[0] }), .EastIn(
        {\nOut10_24[7] , \nOut10_24[6] , \nOut10_24[5] , \nOut10_24[4] , 
        \nOut10_24[3] , \nOut10_24[2] , \nOut10_24[1] , \nOut10_24[0] }), 
        .WestIn({\nOut8_24[7] , \nOut8_24[6] , \nOut8_24[5] , \nOut8_24[4] , 
        \nOut8_24[3] , \nOut8_24[2] , \nOut8_24[1] , \nOut8_24[0] }), .Out({
        \nOut9_24[7] , \nOut9_24[6] , \nOut9_24[5] , \nOut9_24[4] , 
        \nOut9_24[3] , \nOut9_24[2] , \nOut9_24[1] , \nOut9_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_335 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut336[7] , \nScanOut336[6] , 
        \nScanOut336[5] , \nScanOut336[4] , \nScanOut336[3] , \nScanOut336[2] , 
        \nScanOut336[1] , \nScanOut336[0] }), .ScanOut({\nScanOut335[7] , 
        \nScanOut335[6] , \nScanOut335[5] , \nScanOut335[4] , \nScanOut335[3] , 
        \nScanOut335[2] , \nScanOut335[1] , \nScanOut335[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_14[7] , \nOut10_14[6] , \nOut10_14[5] , \nOut10_14[4] , 
        \nOut10_14[3] , \nOut10_14[2] , \nOut10_14[1] , \nOut10_14[0] }), 
        .SouthIn({\nOut10_16[7] , \nOut10_16[6] , \nOut10_16[5] , 
        \nOut10_16[4] , \nOut10_16[3] , \nOut10_16[2] , \nOut10_16[1] , 
        \nOut10_16[0] }), .EastIn({\nOut11_15[7] , \nOut11_15[6] , 
        \nOut11_15[5] , \nOut11_15[4] , \nOut11_15[3] , \nOut11_15[2] , 
        \nOut11_15[1] , \nOut11_15[0] }), .WestIn({\nOut9_15[7] , 
        \nOut9_15[6] , \nOut9_15[5] , \nOut9_15[4] , \nOut9_15[3] , 
        \nOut9_15[2] , \nOut9_15[1] , \nOut9_15[0] }), .Out({\nOut10_15[7] , 
        \nOut10_15[6] , \nOut10_15[5] , \nOut10_15[4] , \nOut10_15[3] , 
        \nOut10_15[2] , \nOut10_15[1] , \nOut10_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_524 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut525[7] , \nScanOut525[6] , 
        \nScanOut525[5] , \nScanOut525[4] , \nScanOut525[3] , \nScanOut525[2] , 
        \nScanOut525[1] , \nScanOut525[0] }), .ScanOut({\nScanOut524[7] , 
        \nScanOut524[6] , \nScanOut524[5] , \nScanOut524[4] , \nScanOut524[3] , 
        \nScanOut524[2] , \nScanOut524[1] , \nScanOut524[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_11[7] , \nOut16_11[6] , \nOut16_11[5] , \nOut16_11[4] , 
        \nOut16_11[3] , \nOut16_11[2] , \nOut16_11[1] , \nOut16_11[0] }), 
        .SouthIn({\nOut16_13[7] , \nOut16_13[6] , \nOut16_13[5] , 
        \nOut16_13[4] , \nOut16_13[3] , \nOut16_13[2] , \nOut16_13[1] , 
        \nOut16_13[0] }), .EastIn({\nOut17_12[7] , \nOut17_12[6] , 
        \nOut17_12[5] , \nOut17_12[4] , \nOut17_12[3] , \nOut17_12[2] , 
        \nOut17_12[1] , \nOut17_12[0] }), .WestIn({\nOut15_12[7] , 
        \nOut15_12[6] , \nOut15_12[5] , \nOut15_12[4] , \nOut15_12[3] , 
        \nOut15_12[2] , \nOut15_12[1] , \nOut15_12[0] }), .Out({\nOut16_12[7] , 
        \nOut16_12[6] , \nOut16_12[5] , \nOut16_12[4] , \nOut16_12[3] , 
        \nOut16_12[2] , \nOut16_12[1] , \nOut16_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_784 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut785[7] , \nScanOut785[6] , 
        \nScanOut785[5] , \nScanOut785[4] , \nScanOut785[3] , \nScanOut785[2] , 
        \nScanOut785[1] , \nScanOut785[0] }), .ScanOut({\nScanOut784[7] , 
        \nScanOut784[6] , \nScanOut784[5] , \nScanOut784[4] , \nScanOut784[3] , 
        \nScanOut784[2] , \nScanOut784[1] , \nScanOut784[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_15[7] , \nOut24_15[6] , \nOut24_15[5] , \nOut24_15[4] , 
        \nOut24_15[3] , \nOut24_15[2] , \nOut24_15[1] , \nOut24_15[0] }), 
        .SouthIn({\nOut24_17[7] , \nOut24_17[6] , \nOut24_17[5] , 
        \nOut24_17[4] , \nOut24_17[3] , \nOut24_17[2] , \nOut24_17[1] , 
        \nOut24_17[0] }), .EastIn({\nOut25_16[7] , \nOut25_16[6] , 
        \nOut25_16[5] , \nOut25_16[4] , \nOut25_16[3] , \nOut25_16[2] , 
        \nOut25_16[1] , \nOut25_16[0] }), .WestIn({\nOut23_16[7] , 
        \nOut23_16[6] , \nOut23_16[5] , \nOut23_16[4] , \nOut23_16[3] , 
        \nOut23_16[2] , \nOut23_16[1] , \nOut23_16[0] }), .Out({\nOut24_16[7] , 
        \nOut24_16[6] , \nOut24_16[5] , \nOut24_16[4] , \nOut24_16[3] , 
        \nOut24_16[2] , \nOut24_16[1] , \nOut24_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_956 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut957[7] , \nScanOut957[6] , 
        \nScanOut957[5] , \nScanOut957[4] , \nScanOut957[3] , \nScanOut957[2] , 
        \nScanOut957[1] , \nScanOut957[0] }), .ScanOut({\nScanOut956[7] , 
        \nScanOut956[6] , \nScanOut956[5] , \nScanOut956[4] , \nScanOut956[3] , 
        \nScanOut956[2] , \nScanOut956[1] , \nScanOut956[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_27[7] , \nOut29_27[6] , \nOut29_27[5] , \nOut29_27[4] , 
        \nOut29_27[3] , \nOut29_27[2] , \nOut29_27[1] , \nOut29_27[0] }), 
        .SouthIn({\nOut29_29[7] , \nOut29_29[6] , \nOut29_29[5] , 
        \nOut29_29[4] , \nOut29_29[3] , \nOut29_29[2] , \nOut29_29[1] , 
        \nOut29_29[0] }), .EastIn({\nOut30_28[7] , \nOut30_28[6] , 
        \nOut30_28[5] , \nOut30_28[4] , \nOut30_28[3] , \nOut30_28[2] , 
        \nOut30_28[1] , \nOut30_28[0] }), .WestIn({\nOut28_28[7] , 
        \nOut28_28[6] , \nOut28_28[5] , \nOut28_28[4] , \nOut28_28[3] , 
        \nOut28_28[2] , \nOut28_28[1] , \nOut28_28[0] }), .Out({\nOut29_28[7] , 
        \nOut29_28[6] , \nOut29_28[5] , \nOut29_28[4] , \nOut29_28[3] , 
        \nOut29_28[2] , \nOut29_28[1] , \nOut29_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_971 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut972[7] , \nScanOut972[6] , 
        \nScanOut972[5] , \nScanOut972[4] , \nScanOut972[3] , \nScanOut972[2] , 
        \nScanOut972[1] , \nScanOut972[0] }), .ScanOut({\nScanOut971[7] , 
        \nScanOut971[6] , \nScanOut971[5] , \nScanOut971[4] , \nScanOut971[3] , 
        \nScanOut971[2] , \nScanOut971[1] , \nScanOut971[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_10[7] , \nOut30_10[6] , \nOut30_10[5] , \nOut30_10[4] , 
        \nOut30_10[3] , \nOut30_10[2] , \nOut30_10[1] , \nOut30_10[0] }), 
        .SouthIn({\nOut30_12[7] , \nOut30_12[6] , \nOut30_12[5] , 
        \nOut30_12[4] , \nOut30_12[3] , \nOut30_12[2] , \nOut30_12[1] , 
        \nOut30_12[0] }), .EastIn({\nOut31_11[7] , \nOut31_11[6] , 
        \nOut31_11[5] , \nOut31_11[4] , \nOut31_11[3] , \nOut31_11[2] , 
        \nOut31_11[1] , \nOut31_11[0] }), .WestIn({\nOut29_11[7] , 
        \nOut29_11[6] , \nOut29_11[5] , \nOut29_11[4] , \nOut29_11[3] , 
        \nOut29_11[2] , \nOut29_11[1] , \nOut29_11[0] }), .Out({\nOut30_11[7] , 
        \nOut30_11[6] , \nOut30_11[5] , \nOut30_11[4] , \nOut30_11[3] , 
        \nOut30_11[2] , \nOut30_11[1] , \nOut30_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_493 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut494[7] , \nScanOut494[6] , 
        \nScanOut494[5] , \nScanOut494[4] , \nScanOut494[3] , \nScanOut494[2] , 
        \nScanOut494[1] , \nScanOut494[0] }), .ScanOut({\nScanOut493[7] , 
        \nScanOut493[6] , \nScanOut493[5] , \nScanOut493[4] , \nScanOut493[3] , 
        \nScanOut493[2] , \nScanOut493[1] , \nScanOut493[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_12[7] , \nOut15_12[6] , \nOut15_12[5] , \nOut15_12[4] , 
        \nOut15_12[3] , \nOut15_12[2] , \nOut15_12[1] , \nOut15_12[0] }), 
        .SouthIn({\nOut15_14[7] , \nOut15_14[6] , \nOut15_14[5] , 
        \nOut15_14[4] , \nOut15_14[3] , \nOut15_14[2] , \nOut15_14[1] , 
        \nOut15_14[0] }), .EastIn({\nOut16_13[7] , \nOut16_13[6] , 
        \nOut16_13[5] , \nOut16_13[4] , \nOut16_13[3] , \nOut16_13[2] , 
        \nOut16_13[1] , \nOut16_13[0] }), .WestIn({\nOut14_13[7] , 
        \nOut14_13[6] , \nOut14_13[5] , \nOut14_13[4] , \nOut14_13[3] , 
        \nOut14_13[2] , \nOut14_13[1] , \nOut14_13[0] }), .Out({\nOut15_13[7] , 
        \nOut15_13[6] , \nOut15_13[5] , \nOut15_13[4] , \nOut15_13[3] , 
        \nOut15_13[2] , \nOut15_13[1] , \nOut15_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_503 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut504[7] , \nScanOut504[6] , 
        \nScanOut504[5] , \nScanOut504[4] , \nScanOut504[3] , \nScanOut504[2] , 
        \nScanOut504[1] , \nScanOut504[0] }), .ScanOut({\nScanOut503[7] , 
        \nScanOut503[6] , \nScanOut503[5] , \nScanOut503[4] , \nScanOut503[3] , 
        \nScanOut503[2] , \nScanOut503[1] , \nScanOut503[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_22[7] , \nOut15_22[6] , \nOut15_22[5] , \nOut15_22[4] , 
        \nOut15_22[3] , \nOut15_22[2] , \nOut15_22[1] , \nOut15_22[0] }), 
        .SouthIn({\nOut15_24[7] , \nOut15_24[6] , \nOut15_24[5] , 
        \nOut15_24[4] , \nOut15_24[3] , \nOut15_24[2] , \nOut15_24[1] , 
        \nOut15_24[0] }), .EastIn({\nOut16_23[7] , \nOut16_23[6] , 
        \nOut16_23[5] , \nOut16_23[4] , \nOut16_23[3] , \nOut16_23[2] , 
        \nOut16_23[1] , \nOut16_23[0] }), .WestIn({\nOut14_23[7] , 
        \nOut14_23[6] , \nOut14_23[5] , \nOut14_23[4] , \nOut14_23[3] , 
        \nOut14_23[2] , \nOut14_23[1] , \nOut14_23[0] }), .Out({\nOut15_23[7] , 
        \nOut15_23[6] , \nOut15_23[5] , \nOut15_23[4] , \nOut15_23[3] , 
        \nOut15_23[2] , \nOut15_23[1] , \nOut15_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_48 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut49[7] , \nScanOut49[6] , 
        \nScanOut49[5] , \nScanOut49[4] , \nScanOut49[3] , \nScanOut49[2] , 
        \nScanOut49[1] , \nScanOut49[0] }), .ScanOut({\nScanOut48[7] , 
        \nScanOut48[6] , \nScanOut48[5] , \nScanOut48[4] , \nScanOut48[3] , 
        \nScanOut48[2] , \nScanOut48[1] , \nScanOut48[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_15[7] , \nOut1_15[6] , \nOut1_15[5] , \nOut1_15[4] , 
        \nOut1_15[3] , \nOut1_15[2] , \nOut1_15[1] , \nOut1_15[0] }), 
        .SouthIn({\nOut1_17[7] , \nOut1_17[6] , \nOut1_17[5] , \nOut1_17[4] , 
        \nOut1_17[3] , \nOut1_17[2] , \nOut1_17[1] , \nOut1_17[0] }), .EastIn(
        {\nOut2_16[7] , \nOut2_16[6] , \nOut2_16[5] , \nOut2_16[4] , 
        \nOut2_16[3] , \nOut2_16[2] , \nOut2_16[1] , \nOut2_16[0] }), .WestIn(
        {\nOut0_16[7] , \nOut0_16[6] , \nOut0_16[5] , \nOut0_16[4] , 
        \nOut0_16[3] , \nOut0_16[2] , \nOut0_16[1] , \nOut0_16[0] }), .Out({
        \nOut1_16[7] , \nOut1_16[6] , \nOut1_16[5] , \nOut1_16[4] , 
        \nOut1_16[3] , \nOut1_16[2] , \nOut1_16[1] , \nOut1_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_139 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut140[7] , \nScanOut140[6] , 
        \nScanOut140[5] , \nScanOut140[4] , \nScanOut140[3] , \nScanOut140[2] , 
        \nScanOut140[1] , \nScanOut140[0] }), .ScanOut({\nScanOut139[7] , 
        \nScanOut139[6] , \nScanOut139[5] , \nScanOut139[4] , \nScanOut139[3] , 
        \nScanOut139[2] , \nScanOut139[1] , \nScanOut139[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_10[7] , \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , 
        \nOut4_10[3] , \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }), 
        .SouthIn({\nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }), .EastIn(
        {\nOut5_11[7] , \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , 
        \nOut5_11[3] , \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }), .WestIn(
        {\nOut3_11[7] , \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , 
        \nOut3_11[3] , \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }), .Out({
        \nOut4_11[7] , \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , 
        \nOut4_11[3] , \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_209 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut210[7] , \nScanOut210[6] , 
        \nScanOut210[5] , \nScanOut210[4] , \nScanOut210[3] , \nScanOut210[2] , 
        \nScanOut210[1] , \nScanOut210[0] }), .ScanOut({\nScanOut209[7] , 
        \nScanOut209[6] , \nScanOut209[5] , \nScanOut209[4] , \nScanOut209[3] , 
        \nScanOut209[2] , \nScanOut209[1] , \nScanOut209[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_16[7] , \nOut6_16[6] , \nOut6_16[5] , \nOut6_16[4] , 
        \nOut6_16[3] , \nOut6_16[2] , \nOut6_16[1] , \nOut6_16[0] }), 
        .SouthIn({\nOut6_18[7] , \nOut6_18[6] , \nOut6_18[5] , \nOut6_18[4] , 
        \nOut6_18[3] , \nOut6_18[2] , \nOut6_18[1] , \nOut6_18[0] }), .EastIn(
        {\nOut7_17[7] , \nOut7_17[6] , \nOut7_17[5] , \nOut7_17[4] , 
        \nOut7_17[3] , \nOut7_17[2] , \nOut7_17[1] , \nOut7_17[0] }), .WestIn(
        {\nOut5_17[7] , \nOut5_17[6] , \nOut5_17[5] , \nOut5_17[4] , 
        \nOut5_17[3] , \nOut5_17[2] , \nOut5_17[1] , \nOut5_17[0] }), .Out({
        \nOut6_17[7] , \nOut6_17[6] , \nOut6_17[5] , \nOut6_17[4] , 
        \nOut6_17[3] , \nOut6_17[2] , \nOut6_17[1] , \nOut6_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_399 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut400[7] , \nScanOut400[6] , 
        \nScanOut400[5] , \nScanOut400[4] , \nScanOut400[3] , \nScanOut400[2] , 
        \nScanOut400[1] , \nScanOut400[0] }), .ScanOut({\nScanOut399[7] , 
        \nScanOut399[6] , \nScanOut399[5] , \nScanOut399[4] , \nScanOut399[3] , 
        \nScanOut399[2] , \nScanOut399[1] , \nScanOut399[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_14[7] , \nOut12_14[6] , \nOut12_14[5] , \nOut12_14[4] , 
        \nOut12_14[3] , \nOut12_14[2] , \nOut12_14[1] , \nOut12_14[0] }), 
        .SouthIn({\nOut12_16[7] , \nOut12_16[6] , \nOut12_16[5] , 
        \nOut12_16[4] , \nOut12_16[3] , \nOut12_16[2] , \nOut12_16[1] , 
        \nOut12_16[0] }), .EastIn({\nOut13_15[7] , \nOut13_15[6] , 
        \nOut13_15[5] , \nOut13_15[4] , \nOut13_15[3] , \nOut13_15[2] , 
        \nOut13_15[1] , \nOut13_15[0] }), .WestIn({\nOut11_15[7] , 
        \nOut11_15[6] , \nOut11_15[5] , \nOut11_15[4] , \nOut11_15[3] , 
        \nOut11_15[2] , \nOut11_15[1] , \nOut11_15[0] }), .Out({\nOut12_15[7] , 
        \nOut12_15[6] , \nOut12_15[5] , \nOut12_15[4] , \nOut12_15[3] , 
        \nOut12_15[2] , \nOut12_15[1] , \nOut12_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_633 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut634[7] , \nScanOut634[6] , 
        \nScanOut634[5] , \nScanOut634[4] , \nScanOut634[3] , \nScanOut634[2] , 
        \nScanOut634[1] , \nScanOut634[0] }), .ScanOut({\nScanOut633[7] , 
        \nScanOut633[6] , \nScanOut633[5] , \nScanOut633[4] , \nScanOut633[3] , 
        \nScanOut633[2] , \nScanOut633[1] , \nScanOut633[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_24[7] , \nOut19_24[6] , \nOut19_24[5] , \nOut19_24[4] , 
        \nOut19_24[3] , \nOut19_24[2] , \nOut19_24[1] , \nOut19_24[0] }), 
        .SouthIn({\nOut19_26[7] , \nOut19_26[6] , \nOut19_26[5] , 
        \nOut19_26[4] , \nOut19_26[3] , \nOut19_26[2] , \nOut19_26[1] , 
        \nOut19_26[0] }), .EastIn({\nOut20_25[7] , \nOut20_25[6] , 
        \nOut20_25[5] , \nOut20_25[4] , \nOut20_25[3] , \nOut20_25[2] , 
        \nOut20_25[1] , \nOut20_25[0] }), .WestIn({\nOut18_25[7] , 
        \nOut18_25[6] , \nOut18_25[5] , \nOut18_25[4] , \nOut18_25[3] , 
        \nOut18_25[2] , \nOut18_25[1] , \nOut18_25[0] }), .Out({\nOut19_25[7] , 
        \nOut19_25[6] , \nOut19_25[5] , \nOut19_25[4] , \nOut19_25[3] , 
        \nOut19_25[2] , \nOut19_25[1] , \nOut19_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1009 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1010[7] , \nScanOut1010[6] , 
        \nScanOut1010[5] , \nScanOut1010[4] , \nScanOut1010[3] , 
        \nScanOut1010[2] , \nScanOut1010[1] , \nScanOut1010[0] }), .ScanOut({
        \nScanOut1009[7] , \nScanOut1009[6] , \nScanOut1009[5] , 
        \nScanOut1009[4] , \nScanOut1009[3] , \nScanOut1009[2] , 
        \nScanOut1009[1] , \nScanOut1009[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_17[7] , \nOut31_17[6] , \nOut31_17[5] , 
        \nOut31_17[4] , \nOut31_17[3] , \nOut31_17[2] , \nOut31_17[1] , 
        \nOut31_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_418 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut419[7] , \nScanOut419[6] , 
        \nScanOut419[5] , \nScanOut419[4] , \nScanOut419[3] , \nScanOut419[2] , 
        \nScanOut419[1] , \nScanOut419[0] }), .ScanOut({\nScanOut418[7] , 
        \nScanOut418[6] , \nScanOut418[5] , \nScanOut418[4] , \nScanOut418[3] , 
        \nScanOut418[2] , \nScanOut418[1] , \nScanOut418[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_1[7] , \nOut13_1[6] , \nOut13_1[5] , \nOut13_1[4] , 
        \nOut13_1[3] , \nOut13_1[2] , \nOut13_1[1] , \nOut13_1[0] }), 
        .SouthIn({\nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }), .EastIn(
        {\nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }), .WestIn(
        {\nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }), .Out({
        \nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_588 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut589[7] , \nScanOut589[6] , 
        \nScanOut589[5] , \nScanOut589[4] , \nScanOut589[3] , \nScanOut589[2] , 
        \nScanOut589[1] , \nScanOut589[0] }), .ScanOut({\nScanOut588[7] , 
        \nScanOut588[6] , \nScanOut588[5] , \nScanOut588[4] , \nScanOut588[3] , 
        \nScanOut588[2] , \nScanOut588[1] , \nScanOut588[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_11[7] , \nOut18_11[6] , \nOut18_11[5] , \nOut18_11[4] , 
        \nOut18_11[3] , \nOut18_11[2] , \nOut18_11[1] , \nOut18_11[0] }), 
        .SouthIn({\nOut18_13[7] , \nOut18_13[6] , \nOut18_13[5] , 
        \nOut18_13[4] , \nOut18_13[3] , \nOut18_13[2] , \nOut18_13[1] , 
        \nOut18_13[0] }), .EastIn({\nOut19_12[7] , \nOut19_12[6] , 
        \nOut19_12[5] , \nOut19_12[4] , \nOut19_12[3] , \nOut19_12[2] , 
        \nOut19_12[1] , \nOut19_12[0] }), .WestIn({\nOut17_12[7] , 
        \nOut17_12[6] , \nOut17_12[5] , \nOut17_12[4] , \nOut17_12[3] , 
        \nOut17_12[2] , \nOut17_12[1] , \nOut17_12[0] }), .Out({\nOut18_12[7] , 
        \nOut18_12[6] , \nOut18_12[5] , \nOut18_12[4] , \nOut18_12[3] , 
        \nOut18_12[2] , \nOut18_12[1] , \nOut18_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_728 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut729[7] , \nScanOut729[6] , 
        \nScanOut729[5] , \nScanOut729[4] , \nScanOut729[3] , \nScanOut729[2] , 
        \nScanOut729[1] , \nScanOut729[0] }), .ScanOut({\nScanOut728[7] , 
        \nScanOut728[6] , \nScanOut728[5] , \nScanOut728[4] , \nScanOut728[3] , 
        \nScanOut728[2] , \nScanOut728[1] , \nScanOut728[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_23[7] , \nOut22_23[6] , \nOut22_23[5] , \nOut22_23[4] , 
        \nOut22_23[3] , \nOut22_23[2] , \nOut22_23[1] , \nOut22_23[0] }), 
        .SouthIn({\nOut22_25[7] , \nOut22_25[6] , \nOut22_25[5] , 
        \nOut22_25[4] , \nOut22_25[3] , \nOut22_25[2] , \nOut22_25[1] , 
        \nOut22_25[0] }), .EastIn({\nOut23_24[7] , \nOut23_24[6] , 
        \nOut23_24[5] , \nOut23_24[4] , \nOut23_24[3] , \nOut23_24[2] , 
        \nOut23_24[1] , \nOut23_24[0] }), .WestIn({\nOut21_24[7] , 
        \nOut21_24[6] , \nOut21_24[5] , \nOut21_24[4] , \nOut21_24[3] , 
        \nOut21_24[2] , \nOut21_24[1] , \nOut21_24[0] }), .Out({\nOut22_24[7] , 
        \nOut22_24[6] , \nOut22_24[5] , \nOut22_24[4] , \nOut22_24[3] , 
        \nOut22_24[2] , \nOut22_24[1] , \nOut22_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_157 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut158[7] , \nScanOut158[6] , 
        \nScanOut158[5] , \nScanOut158[4] , \nScanOut158[3] , \nScanOut158[2] , 
        \nScanOut158[1] , \nScanOut158[0] }), .ScanOut({\nScanOut157[7] , 
        \nScanOut157[6] , \nScanOut157[5] , \nScanOut157[4] , \nScanOut157[3] , 
        \nScanOut157[2] , \nScanOut157[1] , \nScanOut157[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_28[7] , \nOut4_28[6] , \nOut4_28[5] , \nOut4_28[4] , 
        \nOut4_28[3] , \nOut4_28[2] , \nOut4_28[1] , \nOut4_28[0] }), 
        .SouthIn({\nOut4_30[7] , \nOut4_30[6] , \nOut4_30[5] , \nOut4_30[4] , 
        \nOut4_30[3] , \nOut4_30[2] , \nOut4_30[1] , \nOut4_30[0] }), .EastIn(
        {\nOut5_29[7] , \nOut5_29[6] , \nOut5_29[5] , \nOut5_29[4] , 
        \nOut5_29[3] , \nOut5_29[2] , \nOut5_29[1] , \nOut5_29[0] }), .WestIn(
        {\nOut3_29[7] , \nOut3_29[6] , \nOut3_29[5] , \nOut3_29[4] , 
        \nOut3_29[3] , \nOut3_29[2] , \nOut3_29[1] , \nOut3_29[0] }), .Out({
        \nOut4_29[7] , \nOut4_29[6] , \nOut4_29[5] , \nOut4_29[4] , 
        \nOut4_29[3] , \nOut4_29[2] , \nOut4_29[1] , \nOut4_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_267 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut268[7] , \nScanOut268[6] , 
        \nScanOut268[5] , \nScanOut268[4] , \nScanOut268[3] , \nScanOut268[2] , 
        \nScanOut268[1] , \nScanOut268[0] }), .ScanOut({\nScanOut267[7] , 
        \nScanOut267[6] , \nScanOut267[5] , \nScanOut267[4] , \nScanOut267[3] , 
        \nScanOut267[2] , \nScanOut267[1] , \nScanOut267[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_10[7] , \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , 
        \nOut8_10[3] , \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }), 
        .SouthIn({\nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }), .EastIn(
        {\nOut9_11[7] , \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , 
        \nOut9_11[3] , \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }), .WestIn(
        {\nOut7_11[7] , \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , 
        \nOut7_11[3] , \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }), .Out({
        \nOut8_11[7] , \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , 
        \nOut8_11[3] , \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_804 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut805[7] , \nScanOut805[6] , 
        \nScanOut805[5] , \nScanOut805[4] , \nScanOut805[3] , \nScanOut805[2] , 
        \nScanOut805[1] , \nScanOut805[0] }), .ScanOut({\nScanOut804[7] , 
        \nScanOut804[6] , \nScanOut804[5] , \nScanOut804[4] , \nScanOut804[3] , 
        \nScanOut804[2] , \nScanOut804[1] , \nScanOut804[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_3[7] , \nOut25_3[6] , \nOut25_3[5] , \nOut25_3[4] , 
        \nOut25_3[3] , \nOut25_3[2] , \nOut25_3[1] , \nOut25_3[0] }), 
        .SouthIn({\nOut25_5[7] , \nOut25_5[6] , \nOut25_5[5] , \nOut25_5[4] , 
        \nOut25_5[3] , \nOut25_5[2] , \nOut25_5[1] , \nOut25_5[0] }), .EastIn(
        {\nOut26_4[7] , \nOut26_4[6] , \nOut26_4[5] , \nOut26_4[4] , 
        \nOut26_4[3] , \nOut26_4[2] , \nOut26_4[1] , \nOut26_4[0] }), .WestIn(
        {\nOut24_4[7] , \nOut24_4[6] , \nOut24_4[5] , \nOut24_4[4] , 
        \nOut24_4[3] , \nOut24_4[2] , \nOut24_4[1] , \nOut24_4[0] }), .Out({
        \nOut25_4[7] , \nOut25_4[6] , \nOut25_4[5] , \nOut25_4[4] , 
        \nOut25_4[3] , \nOut25_4[2] , \nOut25_4[1] , \nOut25_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_994 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut995[7] , \nScanOut995[6] , 
        \nScanOut995[5] , \nScanOut995[4] , \nScanOut995[3] , \nScanOut995[2] , 
        \nScanOut995[1] , \nScanOut995[0] }), .ScanOut({\nScanOut994[7] , 
        \nScanOut994[6] , \nScanOut994[5] , \nScanOut994[4] , \nScanOut994[3] , 
        \nScanOut994[2] , \nScanOut994[1] , \nScanOut994[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut31_2[7] , \nOut31_2[6] , 
        \nOut31_2[5] , \nOut31_2[4] , \nOut31_2[3] , \nOut31_2[2] , 
        \nOut31_2[1] , \nOut31_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_476 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut477[7] , \nScanOut477[6] , 
        \nScanOut477[5] , \nScanOut477[4] , \nScanOut477[3] , \nScanOut477[2] , 
        \nScanOut477[1] , \nScanOut477[0] }), .ScanOut({\nScanOut476[7] , 
        \nScanOut476[6] , \nScanOut476[5] , \nScanOut476[4] , \nScanOut476[3] , 
        \nScanOut476[2] , \nScanOut476[1] , \nScanOut476[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_27[7] , \nOut14_27[6] , \nOut14_27[5] , \nOut14_27[4] , 
        \nOut14_27[3] , \nOut14_27[2] , \nOut14_27[1] , \nOut14_27[0] }), 
        .SouthIn({\nOut14_29[7] , \nOut14_29[6] , \nOut14_29[5] , 
        \nOut14_29[4] , \nOut14_29[3] , \nOut14_29[2] , \nOut14_29[1] , 
        \nOut14_29[0] }), .EastIn({\nOut15_28[7] , \nOut15_28[6] , 
        \nOut15_28[5] , \nOut15_28[4] , \nOut15_28[3] , \nOut15_28[2] , 
        \nOut15_28[1] , \nOut15_28[0] }), .WestIn({\nOut13_28[7] , 
        \nOut13_28[6] , \nOut13_28[5] , \nOut13_28[4] , \nOut13_28[3] , 
        \nOut13_28[2] , \nOut13_28[1] , \nOut13_28[0] }), .Out({\nOut14_28[7] , 
        \nOut14_28[6] , \nOut14_28[5] , \nOut14_28[4] , \nOut14_28[3] , 
        \nOut14_28[2] , \nOut14_28[1] , \nOut14_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_170 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut171[7] , \nScanOut171[6] , 
        \nScanOut171[5] , \nScanOut171[4] , \nScanOut171[3] , \nScanOut171[2] , 
        \nScanOut171[1] , \nScanOut171[0] }), .ScanOut({\nScanOut170[7] , 
        \nScanOut170[6] , \nScanOut170[5] , \nScanOut170[4] , \nScanOut170[3] , 
        \nScanOut170[2] , \nScanOut170[1] , \nScanOut170[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_9[7] , \nOut5_9[6] , \nOut5_9[5] , \nOut5_9[4] , \nOut5_9[3] , 
        \nOut5_9[2] , \nOut5_9[1] , \nOut5_9[0] }), .SouthIn({\nOut5_11[7] , 
        \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , \nOut5_11[3] , 
        \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }), .EastIn({\nOut6_10[7] , 
        \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , \nOut6_10[3] , 
        \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }), .WestIn({\nOut4_10[7] , 
        \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , \nOut4_10[3] , 
        \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }), .Out({\nOut5_10[7] , 
        \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , \nOut5_10[3] , 
        \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_746 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut747[7] , \nScanOut747[6] , 
        \nScanOut747[5] , \nScanOut747[4] , \nScanOut747[3] , \nScanOut747[2] , 
        \nScanOut747[1] , \nScanOut747[0] }), .ScanOut({\nScanOut746[7] , 
        \nScanOut746[6] , \nScanOut746[5] , \nScanOut746[4] , \nScanOut746[3] , 
        \nScanOut746[2] , \nScanOut746[1] , \nScanOut746[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_9[7] , \nOut23_9[6] , \nOut23_9[5] , \nOut23_9[4] , 
        \nOut23_9[3] , \nOut23_9[2] , \nOut23_9[1] , \nOut23_9[0] }), 
        .SouthIn({\nOut23_11[7] , \nOut23_11[6] , \nOut23_11[5] , 
        \nOut23_11[4] , \nOut23_11[3] , \nOut23_11[2] , \nOut23_11[1] , 
        \nOut23_11[0] }), .EastIn({\nOut24_10[7] , \nOut24_10[6] , 
        \nOut24_10[5] , \nOut24_10[4] , \nOut24_10[3] , \nOut24_10[2] , 
        \nOut24_10[1] , \nOut24_10[0] }), .WestIn({\nOut22_10[7] , 
        \nOut22_10[6] , \nOut22_10[5] , \nOut22_10[4] , \nOut22_10[3] , 
        \nOut22_10[2] , \nOut22_10[1] , \nOut22_10[0] }), .Out({\nOut23_10[7] , 
        \nOut23_10[6] , \nOut23_10[5] , \nOut23_10[4] , \nOut23_10[3] , 
        \nOut23_10[2] , \nOut23_10[1] , \nOut23_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_761 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut762[7] , \nScanOut762[6] , 
        \nScanOut762[5] , \nScanOut762[4] , \nScanOut762[3] , \nScanOut762[2] , 
        \nScanOut762[1] , \nScanOut762[0] }), .ScanOut({\nScanOut761[7] , 
        \nScanOut761[6] , \nScanOut761[5] , \nScanOut761[4] , \nScanOut761[3] , 
        \nScanOut761[2] , \nScanOut761[1] , \nScanOut761[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_24[7] , \nOut23_24[6] , \nOut23_24[5] , \nOut23_24[4] , 
        \nOut23_24[3] , \nOut23_24[2] , \nOut23_24[1] , \nOut23_24[0] }), 
        .SouthIn({\nOut23_26[7] , \nOut23_26[6] , \nOut23_26[5] , 
        \nOut23_26[4] , \nOut23_26[3] , \nOut23_26[2] , \nOut23_26[1] , 
        \nOut23_26[0] }), .EastIn({\nOut24_25[7] , \nOut24_25[6] , 
        \nOut24_25[5] , \nOut24_25[4] , \nOut24_25[3] , \nOut24_25[2] , 
        \nOut24_25[1] , \nOut24_25[0] }), .WestIn({\nOut22_25[7] , 
        \nOut22_25[6] , \nOut22_25[5] , \nOut22_25[4] , \nOut22_25[3] , 
        \nOut22_25[2] , \nOut22_25[1] , \nOut22_25[0] }), .Out({\nOut23_25[7] , 
        \nOut23_25[6] , \nOut23_25[5] , \nOut23_25[4] , \nOut23_25[3] , 
        \nOut23_25[2] , \nOut23_25[1] , \nOut23_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_240 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut241[7] , \nScanOut241[6] , 
        \nScanOut241[5] , \nScanOut241[4] , \nScanOut241[3] , \nScanOut241[2] , 
        \nScanOut241[1] , \nScanOut241[0] }), .ScanOut({\nScanOut240[7] , 
        \nScanOut240[6] , \nScanOut240[5] , \nScanOut240[4] , \nScanOut240[3] , 
        \nScanOut240[2] , \nScanOut240[1] , \nScanOut240[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_15[7] , \nOut7_15[6] , \nOut7_15[5] , \nOut7_15[4] , 
        \nOut7_15[3] , \nOut7_15[2] , \nOut7_15[1] , \nOut7_15[0] }), 
        .SouthIn({\nOut7_17[7] , \nOut7_17[6] , \nOut7_17[5] , \nOut7_17[4] , 
        \nOut7_17[3] , \nOut7_17[2] , \nOut7_17[1] , \nOut7_17[0] }), .EastIn(
        {\nOut8_16[7] , \nOut8_16[6] , \nOut8_16[5] , \nOut8_16[4] , 
        \nOut8_16[3] , \nOut8_16[2] , \nOut8_16[1] , \nOut8_16[0] }), .WestIn(
        {\nOut6_16[7] , \nOut6_16[6] , \nOut6_16[5] , \nOut6_16[4] , 
        \nOut6_16[3] , \nOut6_16[2] , \nOut6_16[1] , \nOut6_16[0] }), .Out({
        \nOut7_16[7] , \nOut7_16[6] , \nOut7_16[5] , \nOut7_16[4] , 
        \nOut7_16[3] , \nOut7_16[2] , \nOut7_16[1] , \nOut7_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_451 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut452[7] , \nScanOut452[6] , 
        \nScanOut452[5] , \nScanOut452[4] , \nScanOut452[3] , \nScanOut452[2] , 
        \nScanOut452[1] , \nScanOut452[0] }), .ScanOut({\nScanOut451[7] , 
        \nScanOut451[6] , \nScanOut451[5] , \nScanOut451[4] , \nScanOut451[3] , 
        \nScanOut451[2] , \nScanOut451[1] , \nScanOut451[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }), 
        .SouthIn({\nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }), .EastIn(
        {\nOut15_3[7] , \nOut15_3[6] , \nOut15_3[5] , \nOut15_3[4] , 
        \nOut15_3[3] , \nOut15_3[2] , \nOut15_3[1] , \nOut15_3[0] }), .WestIn(
        {\nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }), .Out({
        \nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_823 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut824[7] , \nScanOut824[6] , 
        \nScanOut824[5] , \nScanOut824[4] , \nScanOut824[3] , \nScanOut824[2] , 
        \nScanOut824[1] , \nScanOut824[0] }), .ScanOut({\nScanOut823[7] , 
        \nScanOut823[6] , \nScanOut823[5] , \nScanOut823[4] , \nScanOut823[3] , 
        \nScanOut823[2] , \nScanOut823[1] , \nScanOut823[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_22[7] , \nOut25_22[6] , \nOut25_22[5] , \nOut25_22[4] , 
        \nOut25_22[3] , \nOut25_22[2] , \nOut25_22[1] , \nOut25_22[0] }), 
        .SouthIn({\nOut25_24[7] , \nOut25_24[6] , \nOut25_24[5] , 
        \nOut25_24[4] , \nOut25_24[3] , \nOut25_24[2] , \nOut25_24[1] , 
        \nOut25_24[0] }), .EastIn({\nOut26_23[7] , \nOut26_23[6] , 
        \nOut26_23[5] , \nOut26_23[4] , \nOut26_23[3] , \nOut26_23[2] , 
        \nOut26_23[1] , \nOut26_23[0] }), .WestIn({\nOut24_23[7] , 
        \nOut24_23[6] , \nOut24_23[5] , \nOut24_23[4] , \nOut24_23[3] , 
        \nOut24_23[2] , \nOut24_23[1] , \nOut24_23[0] }), .Out({\nOut25_23[7] , 
        \nOut25_23[6] , \nOut25_23[5] , \nOut25_23[4] , \nOut25_23[3] , 
        \nOut25_23[2] , \nOut25_23[1] , \nOut25_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_53 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut54[7] , \nScanOut54[6] , 
        \nScanOut54[5] , \nScanOut54[4] , \nScanOut54[3] , \nScanOut54[2] , 
        \nScanOut54[1] , \nScanOut54[0] }), .ScanOut({\nScanOut53[7] , 
        \nScanOut53[6] , \nScanOut53[5] , \nScanOut53[4] , \nScanOut53[3] , 
        \nScanOut53[2] , \nScanOut53[1] , \nScanOut53[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_20[7] , \nOut1_20[6] , \nOut1_20[5] , \nOut1_20[4] , 
        \nOut1_20[3] , \nOut1_20[2] , \nOut1_20[1] , \nOut1_20[0] }), 
        .SouthIn({\nOut1_22[7] , \nOut1_22[6] , \nOut1_22[5] , \nOut1_22[4] , 
        \nOut1_22[3] , \nOut1_22[2] , \nOut1_22[1] , \nOut1_22[0] }), .EastIn(
        {\nOut2_21[7] , \nOut2_21[6] , \nOut2_21[5] , \nOut2_21[4] , 
        \nOut2_21[3] , \nOut2_21[2] , \nOut2_21[1] , \nOut2_21[0] }), .WestIn(
        {\nOut0_21[7] , \nOut0_21[6] , \nOut0_21[5] , \nOut0_21[4] , 
        \nOut0_21[3] , \nOut0_21[2] , \nOut0_21[1] , \nOut0_21[0] }), .Out({
        \nOut1_21[7] , \nOut1_21[6] , \nOut1_21[5] , \nOut1_21[4] , 
        \nOut1_21[3] , \nOut1_21[2] , \nOut1_21[1] , \nOut1_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_74 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut75[7] , \nScanOut75[6] , 
        \nScanOut75[5] , \nScanOut75[4] , \nScanOut75[3] , \nScanOut75[2] , 
        \nScanOut75[1] , \nScanOut75[0] }), .ScanOut({\nScanOut74[7] , 
        \nScanOut74[6] , \nScanOut74[5] , \nScanOut74[4] , \nScanOut74[3] , 
        \nScanOut74[2] , \nScanOut74[1] , \nScanOut74[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_9[7] , \nOut2_9[6] , \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , 
        \nOut2_9[2] , \nOut2_9[1] , \nOut2_9[0] }), .SouthIn({\nOut2_11[7] , 
        \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , \nOut2_11[3] , 
        \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), .EastIn({\nOut3_10[7] , 
        \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , \nOut3_10[3] , 
        \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }), .WestIn({\nOut1_10[7] , 
        \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , \nOut1_10[3] , 
        \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), .Out({\nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_340 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut341[7] , \nScanOut341[6] , 
        \nScanOut341[5] , \nScanOut341[4] , \nScanOut341[3] , \nScanOut341[2] , 
        \nScanOut341[1] , \nScanOut341[0] }), .ScanOut({\nScanOut340[7] , 
        \nScanOut340[6] , \nScanOut340[5] , \nScanOut340[4] , \nScanOut340[3] , 
        \nScanOut340[2] , \nScanOut340[1] , \nScanOut340[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_19[7] , \nOut10_19[6] , \nOut10_19[5] , \nOut10_19[4] , 
        \nOut10_19[3] , \nOut10_19[2] , \nOut10_19[1] , \nOut10_19[0] }), 
        .SouthIn({\nOut10_21[7] , \nOut10_21[6] , \nOut10_21[5] , 
        \nOut10_21[4] , \nOut10_21[3] , \nOut10_21[2] , \nOut10_21[1] , 
        \nOut10_21[0] }), .EastIn({\nOut11_20[7] , \nOut11_20[6] , 
        \nOut11_20[5] , \nOut11_20[4] , \nOut11_20[3] , \nOut11_20[2] , 
        \nOut11_20[1] , \nOut11_20[0] }), .WestIn({\nOut9_20[7] , 
        \nOut9_20[6] , \nOut9_20[5] , \nOut9_20[4] , \nOut9_20[3] , 
        \nOut9_20[2] , \nOut9_20[1] , \nOut9_20[0] }), .Out({\nOut10_20[7] , 
        \nOut10_20[6] , \nOut10_20[5] , \nOut10_20[4] , \nOut10_20[3] , 
        \nOut10_20[2] , \nOut10_20[1] , \nOut10_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_923 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut924[7] , \nScanOut924[6] , 
        \nScanOut924[5] , \nScanOut924[4] , \nScanOut924[3] , \nScanOut924[2] , 
        \nScanOut924[1] , \nScanOut924[0] }), .ScanOut({\nScanOut923[7] , 
        \nScanOut923[6] , \nScanOut923[5] , \nScanOut923[4] , \nScanOut923[3] , 
        \nScanOut923[2] , \nScanOut923[1] , \nScanOut923[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_26[7] , \nOut28_26[6] , \nOut28_26[5] , \nOut28_26[4] , 
        \nOut28_26[3] , \nOut28_26[2] , \nOut28_26[1] , \nOut28_26[0] }), 
        .SouthIn({\nOut28_28[7] , \nOut28_28[6] , \nOut28_28[5] , 
        \nOut28_28[4] , \nOut28_28[3] , \nOut28_28[2] , \nOut28_28[1] , 
        \nOut28_28[0] }), .EastIn({\nOut29_27[7] , \nOut29_27[6] , 
        \nOut29_27[5] , \nOut29_27[4] , \nOut29_27[3] , \nOut29_27[2] , 
        \nOut29_27[1] , \nOut29_27[0] }), .WestIn({\nOut27_27[7] , 
        \nOut27_27[6] , \nOut27_27[5] , \nOut27_27[4] , \nOut27_27[3] , 
        \nOut27_27[2] , \nOut27_27[1] , \nOut27_27[0] }), .Out({\nOut28_27[7] , 
        \nOut28_27[6] , \nOut28_27[5] , \nOut28_27[4] , \nOut28_27[3] , 
        \nOut28_27[2] , \nOut28_27[1] , \nOut28_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_938 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut939[7] , \nScanOut939[6] , 
        \nScanOut939[5] , \nScanOut939[4] , \nScanOut939[3] , \nScanOut939[2] , 
        \nScanOut939[1] , \nScanOut939[0] }), .ScanOut({\nScanOut938[7] , 
        \nScanOut938[6] , \nScanOut938[5] , \nScanOut938[4] , \nScanOut938[3] , 
        \nScanOut938[2] , \nScanOut938[1] , \nScanOut938[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_9[7] , \nOut29_9[6] , \nOut29_9[5] , \nOut29_9[4] , 
        \nOut29_9[3] , \nOut29_9[2] , \nOut29_9[1] , \nOut29_9[0] }), 
        .SouthIn({\nOut29_11[7] , \nOut29_11[6] , \nOut29_11[5] , 
        \nOut29_11[4] , \nOut29_11[3] , \nOut29_11[2] , \nOut29_11[1] , 
        \nOut29_11[0] }), .EastIn({\nOut30_10[7] , \nOut30_10[6] , 
        \nOut30_10[5] , \nOut30_10[4] , \nOut30_10[3] , \nOut30_10[2] , 
        \nOut30_10[1] , \nOut30_10[0] }), .WestIn({\nOut28_10[7] , 
        \nOut28_10[6] , \nOut28_10[5] , \nOut28_10[4] , \nOut28_10[3] , 
        \nOut28_10[2] , \nOut28_10[1] , \nOut28_10[0] }), .Out({\nOut29_10[7] , 
        \nOut29_10[6] , \nOut29_10[5] , \nOut29_10[4] , \nOut29_10[3] , 
        \nOut29_10[2] , \nOut29_10[1] , \nOut29_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_551 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut552[7] , \nScanOut552[6] , 
        \nScanOut552[5] , \nScanOut552[4] , \nScanOut552[3] , \nScanOut552[2] , 
        \nScanOut552[1] , \nScanOut552[0] }), .ScanOut({\nScanOut551[7] , 
        \nScanOut551[6] , \nScanOut551[5] , \nScanOut551[4] , \nScanOut551[3] , 
        \nScanOut551[2] , \nScanOut551[1] , \nScanOut551[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_6[7] , \nOut17_6[6] , \nOut17_6[5] , \nOut17_6[4] , 
        \nOut17_6[3] , \nOut17_6[2] , \nOut17_6[1] , \nOut17_6[0] }), 
        .SouthIn({\nOut17_8[7] , \nOut17_8[6] , \nOut17_8[5] , \nOut17_8[4] , 
        \nOut17_8[3] , \nOut17_8[2] , \nOut17_8[1] , \nOut17_8[0] }), .EastIn(
        {\nOut18_7[7] , \nOut18_7[6] , \nOut18_7[5] , \nOut18_7[4] , 
        \nOut18_7[3] , \nOut18_7[2] , \nOut18_7[1] , \nOut18_7[0] }), .WestIn(
        {\nOut16_7[7] , \nOut16_7[6] , \nOut16_7[5] , \nOut16_7[4] , 
        \nOut16_7[3] , \nOut16_7[2] , \nOut16_7[1] , \nOut16_7[0] }), .Out({
        \nOut17_7[7] , \nOut17_7[6] , \nOut17_7[5] , \nOut17_7[4] , 
        \nOut17_7[3] , \nOut17_7[2] , \nOut17_7[1] , \nOut17_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_661 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut662[7] , \nScanOut662[6] , 
        \nScanOut662[5] , \nScanOut662[4] , \nScanOut662[3] , \nScanOut662[2] , 
        \nScanOut662[1] , \nScanOut662[0] }), .ScanOut({\nScanOut661[7] , 
        \nScanOut661[6] , \nScanOut661[5] , \nScanOut661[4] , \nScanOut661[3] , 
        \nScanOut661[2] , \nScanOut661[1] , \nScanOut661[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_20[7] , \nOut20_20[6] , \nOut20_20[5] , \nOut20_20[4] , 
        \nOut20_20[3] , \nOut20_20[2] , \nOut20_20[1] , \nOut20_20[0] }), 
        .SouthIn({\nOut20_22[7] , \nOut20_22[6] , \nOut20_22[5] , 
        \nOut20_22[4] , \nOut20_22[3] , \nOut20_22[2] , \nOut20_22[1] , 
        \nOut20_22[0] }), .EastIn({\nOut21_21[7] , \nOut21_21[6] , 
        \nOut21_21[5] , \nOut21_21[4] , \nOut21_21[3] , \nOut21_21[2] , 
        \nOut21_21[1] , \nOut21_21[0] }), .WestIn({\nOut19_21[7] , 
        \nOut19_21[6] , \nOut19_21[5] , \nOut19_21[4] , \nOut19_21[3] , 
        \nOut19_21[2] , \nOut19_21[1] , \nOut19_21[0] }), .Out({\nOut20_21[7] , 
        \nOut20_21[6] , \nOut20_21[5] , \nOut20_21[4] , \nOut20_21[3] , 
        \nOut20_21[2] , \nOut20_21[1] , \nOut20_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_646 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut647[7] , \nScanOut647[6] , 
        \nScanOut647[5] , \nScanOut647[4] , \nScanOut647[3] , \nScanOut647[2] , 
        \nScanOut647[1] , \nScanOut647[0] }), .ScanOut({\nScanOut646[7] , 
        \nScanOut646[6] , \nScanOut646[5] , \nScanOut646[4] , \nScanOut646[3] , 
        \nScanOut646[2] , \nScanOut646[1] , \nScanOut646[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_5[7] , \nOut20_5[6] , \nOut20_5[5] , \nOut20_5[4] , 
        \nOut20_5[3] , \nOut20_5[2] , \nOut20_5[1] , \nOut20_5[0] }), 
        .SouthIn({\nOut20_7[7] , \nOut20_7[6] , \nOut20_7[5] , \nOut20_7[4] , 
        \nOut20_7[3] , \nOut20_7[2] , \nOut20_7[1] , \nOut20_7[0] }), .EastIn(
        {\nOut21_6[7] , \nOut21_6[6] , \nOut21_6[5] , \nOut21_6[4] , 
        \nOut21_6[3] , \nOut21_6[2] , \nOut21_6[1] , \nOut21_6[0] }), .WestIn(
        {\nOut19_6[7] , \nOut19_6[6] , \nOut19_6[5] , \nOut19_6[4] , 
        \nOut19_6[3] , \nOut19_6[2] , \nOut19_6[1] , \nOut19_6[0] }), .Out({
        \nOut20_6[7] , \nOut20_6[6] , \nOut20_6[5] , \nOut20_6[4] , 
        \nOut20_6[3] , \nOut20_6[2] , \nOut20_6[1] , \nOut20_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_66 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut67[7] , \nScanOut67[6] , 
        \nScanOut67[5] , \nScanOut67[4] , \nScanOut67[3] , \nScanOut67[2] , 
        \nScanOut67[1] , \nScanOut67[0] }), .ScanOut({\nScanOut66[7] , 
        \nScanOut66[6] , \nScanOut66[5] , \nScanOut66[4] , \nScanOut66[3] , 
        \nScanOut66[2] , \nScanOut66[1] , \nScanOut66[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , \nOut2_1[4] , \nOut2_1[3] , 
        \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }), .SouthIn({\nOut2_3[7] , 
        \nOut2_3[6] , \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , 
        \nOut2_3[1] , \nOut2_3[0] }), .EastIn({\nOut3_2[7] , \nOut3_2[6] , 
        \nOut3_2[5] , \nOut3_2[4] , \nOut3_2[3] , \nOut3_2[2] , \nOut3_2[1] , 
        \nOut3_2[0] }), .WestIn({\nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , 
        \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), 
        .Out({\nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , 
        \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_83 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut84[7] , \nScanOut84[6] , 
        \nScanOut84[5] , \nScanOut84[4] , \nScanOut84[3] , \nScanOut84[2] , 
        \nScanOut84[1] , \nScanOut84[0] }), .ScanOut({\nScanOut83[7] , 
        \nScanOut83[6] , \nScanOut83[5] , \nScanOut83[4] , \nScanOut83[3] , 
        \nScanOut83[2] , \nScanOut83[1] , \nScanOut83[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_18[7] , \nOut2_18[6] , \nOut2_18[5] , \nOut2_18[4] , 
        \nOut2_18[3] , \nOut2_18[2] , \nOut2_18[1] , \nOut2_18[0] }), 
        .SouthIn({\nOut2_20[7] , \nOut2_20[6] , \nOut2_20[5] , \nOut2_20[4] , 
        \nOut2_20[3] , \nOut2_20[2] , \nOut2_20[1] , \nOut2_20[0] }), .EastIn(
        {\nOut3_19[7] , \nOut3_19[6] , \nOut3_19[5] , \nOut3_19[4] , 
        \nOut3_19[3] , \nOut3_19[2] , \nOut3_19[1] , \nOut3_19[0] }), .WestIn(
        {\nOut1_19[7] , \nOut1_19[6] , \nOut1_19[5] , \nOut1_19[4] , 
        \nOut1_19[3] , \nOut1_19[2] , \nOut1_19[1] , \nOut1_19[0] }), .Out({
        \nOut2_19[7] , \nOut2_19[6] , \nOut2_19[5] , \nOut2_19[4] , 
        \nOut2_19[3] , \nOut2_19[2] , \nOut2_19[1] , \nOut2_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_91 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut92[7] , \nScanOut92[6] , 
        \nScanOut92[5] , \nScanOut92[4] , \nScanOut92[3] , \nScanOut92[2] , 
        \nScanOut92[1] , \nScanOut92[0] }), .ScanOut({\nScanOut91[7] , 
        \nScanOut91[6] , \nScanOut91[5] , \nScanOut91[4] , \nScanOut91[3] , 
        \nScanOut91[2] , \nScanOut91[1] , \nScanOut91[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_26[7] , \nOut2_26[6] , \nOut2_26[5] , \nOut2_26[4] , 
        \nOut2_26[3] , \nOut2_26[2] , \nOut2_26[1] , \nOut2_26[0] }), 
        .SouthIn({\nOut2_28[7] , \nOut2_28[6] , \nOut2_28[5] , \nOut2_28[4] , 
        \nOut2_28[3] , \nOut2_28[2] , \nOut2_28[1] , \nOut2_28[0] }), .EastIn(
        {\nOut3_27[7] , \nOut3_27[6] , \nOut3_27[5] , \nOut3_27[4] , 
        \nOut3_27[3] , \nOut3_27[2] , \nOut3_27[1] , \nOut3_27[0] }), .WestIn(
        {\nOut1_27[7] , \nOut1_27[6] , \nOut1_27[5] , \nOut1_27[4] , 
        \nOut1_27[3] , \nOut1_27[2] , \nOut1_27[1] , \nOut1_27[0] }), .Out({
        \nOut2_27[7] , \nOut2_27[6] , \nOut2_27[5] , \nOut2_27[4] , 
        \nOut2_27[3] , \nOut2_27[2] , \nOut2_27[1] , \nOut2_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_122 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut123[7] , \nScanOut123[6] , 
        \nScanOut123[5] , \nScanOut123[4] , \nScanOut123[3] , \nScanOut123[2] , 
        \nScanOut123[1] , \nScanOut123[0] }), .ScanOut({\nScanOut122[7] , 
        \nScanOut122[6] , \nScanOut122[5] , \nScanOut122[4] , \nScanOut122[3] , 
        \nScanOut122[2] , \nScanOut122[1] , \nScanOut122[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_25[7] , \nOut3_25[6] , \nOut3_25[5] , \nOut3_25[4] , 
        \nOut3_25[3] , \nOut3_25[2] , \nOut3_25[1] , \nOut3_25[0] }), 
        .SouthIn({\nOut3_27[7] , \nOut3_27[6] , \nOut3_27[5] , \nOut3_27[4] , 
        \nOut3_27[3] , \nOut3_27[2] , \nOut3_27[1] , \nOut3_27[0] }), .EastIn(
        {\nOut4_26[7] , \nOut4_26[6] , \nOut4_26[5] , \nOut4_26[4] , 
        \nOut4_26[3] , \nOut4_26[2] , \nOut4_26[1] , \nOut4_26[0] }), .WestIn(
        {\nOut2_26[7] , \nOut2_26[6] , \nOut2_26[5] , \nOut2_26[4] , 
        \nOut2_26[3] , \nOut2_26[2] , \nOut2_26[1] , \nOut2_26[0] }), .Out({
        \nOut3_26[7] , \nOut3_26[6] , \nOut3_26[5] , \nOut3_26[4] , 
        \nOut3_26[3] , \nOut3_26[2] , \nOut3_26[1] , \nOut3_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_367 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut368[7] , \nScanOut368[6] , 
        \nScanOut368[5] , \nScanOut368[4] , \nScanOut368[3] , \nScanOut368[2] , 
        \nScanOut368[1] , \nScanOut368[0] }), .ScanOut({\nScanOut367[7] , 
        \nScanOut367[6] , \nScanOut367[5] , \nScanOut367[4] , \nScanOut367[3] , 
        \nScanOut367[2] , \nScanOut367[1] , \nScanOut367[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_14[7] , \nOut11_14[6] , \nOut11_14[5] , \nOut11_14[4] , 
        \nOut11_14[3] , \nOut11_14[2] , \nOut11_14[1] , \nOut11_14[0] }), 
        .SouthIn({\nOut11_16[7] , \nOut11_16[6] , \nOut11_16[5] , 
        \nOut11_16[4] , \nOut11_16[3] , \nOut11_16[2] , \nOut11_16[1] , 
        \nOut11_16[0] }), .EastIn({\nOut12_15[7] , \nOut12_15[6] , 
        \nOut12_15[5] , \nOut12_15[4] , \nOut12_15[3] , \nOut12_15[2] , 
        \nOut12_15[1] , \nOut12_15[0] }), .WestIn({\nOut10_15[7] , 
        \nOut10_15[6] , \nOut10_15[5] , \nOut10_15[4] , \nOut10_15[3] , 
        \nOut10_15[2] , \nOut10_15[1] , \nOut10_15[0] }), .Out({\nOut11_15[7] , 
        \nOut11_15[6] , \nOut11_15[5] , \nOut11_15[4] , \nOut11_15[3] , 
        \nOut11_15[2] , \nOut11_15[1] , \nOut11_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_576 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut577[7] , \nScanOut577[6] , 
        \nScanOut577[5] , \nScanOut577[4] , \nScanOut577[3] , \nScanOut577[2] , 
        \nScanOut577[1] , \nScanOut577[0] }), .ScanOut({\nScanOut576[7] , 
        \nScanOut576[6] , \nScanOut576[5] , \nScanOut576[4] , \nScanOut576[3] , 
        \nScanOut576[2] , \nScanOut576[1] , \nScanOut576[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut18_0[7] , \nOut18_0[6] , 
        \nOut18_0[5] , \nOut18_0[4] , \nOut18_0[3] , \nOut18_0[2] , 
        \nOut18_0[1] , \nOut18_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_894 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut895[7] , \nScanOut895[6] , 
        \nScanOut895[5] , \nScanOut895[4] , \nScanOut895[3] , \nScanOut895[2] , 
        \nScanOut895[1] , \nScanOut895[0] }), .ScanOut({\nScanOut894[7] , 
        \nScanOut894[6] , \nScanOut894[5] , \nScanOut894[4] , \nScanOut894[3] , 
        \nScanOut894[2] , \nScanOut894[1] , \nScanOut894[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_29[7] , \nOut27_29[6] , \nOut27_29[5] , \nOut27_29[4] , 
        \nOut27_29[3] , \nOut27_29[2] , \nOut27_29[1] , \nOut27_29[0] }), 
        .SouthIn({\nOut27_31[7] , \nOut27_31[6] , \nOut27_31[5] , 
        \nOut27_31[4] , \nOut27_31[3] , \nOut27_31[2] , \nOut27_31[1] , 
        \nOut27_31[0] }), .EastIn({\nOut28_30[7] , \nOut28_30[6] , 
        \nOut28_30[5] , \nOut28_30[4] , \nOut28_30[3] , \nOut28_30[2] , 
        \nOut28_30[1] , \nOut28_30[0] }), .WestIn({\nOut26_30[7] , 
        \nOut26_30[6] , \nOut26_30[5] , \nOut26_30[4] , \nOut26_30[3] , 
        \nOut26_30[2] , \nOut26_30[1] , \nOut26_30[0] }), .Out({\nOut27_30[7] , 
        \nOut27_30[6] , \nOut27_30[5] , \nOut27_30[4] , \nOut27_30[3] , 
        \nOut27_30[2] , \nOut27_30[1] , \nOut27_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_904 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut905[7] , \nScanOut905[6] , 
        \nScanOut905[5] , \nScanOut905[4] , \nScanOut905[3] , \nScanOut905[2] , 
        \nScanOut905[1] , \nScanOut905[0] }), .ScanOut({\nScanOut904[7] , 
        \nScanOut904[6] , \nScanOut904[5] , \nScanOut904[4] , \nScanOut904[3] , 
        \nScanOut904[2] , \nScanOut904[1] , \nScanOut904[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_7[7] , \nOut28_7[6] , \nOut28_7[5] , \nOut28_7[4] , 
        \nOut28_7[3] , \nOut28_7[2] , \nOut28_7[1] , \nOut28_7[0] }), 
        .SouthIn({\nOut28_9[7] , \nOut28_9[6] , \nOut28_9[5] , \nOut28_9[4] , 
        \nOut28_9[3] , \nOut28_9[2] , \nOut28_9[1] , \nOut28_9[0] }), .EastIn(
        {\nOut29_8[7] , \nOut29_8[6] , \nOut29_8[5] , \nOut29_8[4] , 
        \nOut29_8[3] , \nOut29_8[2] , \nOut29_8[1] , \nOut29_8[0] }), .WestIn(
        {\nOut27_8[7] , \nOut27_8[6] , \nOut27_8[5] , \nOut27_8[4] , 
        \nOut27_8[3] , \nOut27_8[2] , \nOut27_8[1] , \nOut27_8[0] }), .Out({
        \nOut28_8[7] , \nOut28_8[6] , \nOut28_8[5] , \nOut28_8[4] , 
        \nOut28_8[3] , \nOut28_8[2] , \nOut28_8[1] , \nOut28_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_733 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut734[7] , \nScanOut734[6] , 
        \nScanOut734[5] , \nScanOut734[4] , \nScanOut734[3] , \nScanOut734[2] , 
        \nScanOut734[1] , \nScanOut734[0] }), .ScanOut({\nScanOut733[7] , 
        \nScanOut733[6] , \nScanOut733[5] , \nScanOut733[4] , \nScanOut733[3] , 
        \nScanOut733[2] , \nScanOut733[1] , \nScanOut733[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_28[7] , \nOut22_28[6] , \nOut22_28[5] , \nOut22_28[4] , 
        \nOut22_28[3] , \nOut22_28[2] , \nOut22_28[1] , \nOut22_28[0] }), 
        .SouthIn({\nOut22_30[7] , \nOut22_30[6] , \nOut22_30[5] , 
        \nOut22_30[4] , \nOut22_30[3] , \nOut22_30[2] , \nOut22_30[1] , 
        \nOut22_30[0] }), .EastIn({\nOut23_29[7] , \nOut23_29[6] , 
        \nOut23_29[5] , \nOut23_29[4] , \nOut23_29[3] , \nOut23_29[2] , 
        \nOut23_29[1] , \nOut23_29[0] }), .WestIn({\nOut21_29[7] , 
        \nOut21_29[6] , \nOut21_29[5] , \nOut21_29[4] , \nOut21_29[3] , 
        \nOut21_29[2] , \nOut21_29[1] , \nOut21_29[0] }), .Out({\nOut22_29[7] , 
        \nOut22_29[6] , \nOut22_29[5] , \nOut22_29[4] , \nOut22_29[3] , 
        \nOut22_29[2] , \nOut22_29[1] , \nOut22_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_838 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut839[7] , \nScanOut839[6] , 
        \nScanOut839[5] , \nScanOut839[4] , \nScanOut839[3] , \nScanOut839[2] , 
        \nScanOut839[1] , \nScanOut839[0] }), .ScanOut({\nScanOut838[7] , 
        \nScanOut838[6] , \nScanOut838[5] , \nScanOut838[4] , \nScanOut838[3] , 
        \nScanOut838[2] , \nScanOut838[1] , \nScanOut838[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_5[7] , \nOut26_5[6] , \nOut26_5[5] , \nOut26_5[4] , 
        \nOut26_5[3] , \nOut26_5[2] , \nOut26_5[1] , \nOut26_5[0] }), 
        .SouthIn({\nOut26_7[7] , \nOut26_7[6] , \nOut26_7[5] , \nOut26_7[4] , 
        \nOut26_7[3] , \nOut26_7[2] , \nOut26_7[1] , \nOut26_7[0] }), .EastIn(
        {\nOut27_6[7] , \nOut27_6[6] , \nOut27_6[5] , \nOut27_6[4] , 
        \nOut27_6[3] , \nOut27_6[2] , \nOut27_6[1] , \nOut27_6[0] }), .WestIn(
        {\nOut25_6[7] , \nOut25_6[6] , \nOut25_6[5] , \nOut25_6[4] , 
        \nOut25_6[3] , \nOut25_6[2] , \nOut25_6[1] , \nOut25_6[0] }), .Out({
        \nOut26_6[7] , \nOut26_6[6] , \nOut26_6[5] , \nOut26_6[4] , 
        \nOut26_6[3] , \nOut26_6[2] , \nOut26_6[1] , \nOut26_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_212 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut213[7] , \nScanOut213[6] , 
        \nScanOut213[5] , \nScanOut213[4] , \nScanOut213[3] , \nScanOut213[2] , 
        \nScanOut213[1] , \nScanOut213[0] }), .ScanOut({\nScanOut212[7] , 
        \nScanOut212[6] , \nScanOut212[5] , \nScanOut212[4] , \nScanOut212[3] , 
        \nScanOut212[2] , \nScanOut212[1] , \nScanOut212[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_19[7] , \nOut6_19[6] , \nOut6_19[5] , \nOut6_19[4] , 
        \nOut6_19[3] , \nOut6_19[2] , \nOut6_19[1] , \nOut6_19[0] }), 
        .SouthIn({\nOut6_21[7] , \nOut6_21[6] , \nOut6_21[5] , \nOut6_21[4] , 
        \nOut6_21[3] , \nOut6_21[2] , \nOut6_21[1] , \nOut6_21[0] }), .EastIn(
        {\nOut7_20[7] , \nOut7_20[6] , \nOut7_20[5] , \nOut7_20[4] , 
        \nOut7_20[3] , \nOut7_20[2] , \nOut7_20[1] , \nOut7_20[0] }), .WestIn(
        {\nOut5_20[7] , \nOut5_20[6] , \nOut5_20[5] , \nOut5_20[4] , 
        \nOut5_20[3] , \nOut5_20[2] , \nOut5_20[1] , \nOut5_20[0] }), .Out({
        \nOut6_20[7] , \nOut6_20[6] , \nOut6_20[5] , \nOut6_20[4] , 
        \nOut6_20[3] , \nOut6_20[2] , \nOut6_20[1] , \nOut6_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_382 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut383[7] , \nScanOut383[6] , 
        \nScanOut383[5] , \nScanOut383[4] , \nScanOut383[3] , \nScanOut383[2] , 
        \nScanOut383[1] , \nScanOut383[0] }), .ScanOut({\nScanOut382[7] , 
        \nScanOut382[6] , \nScanOut382[5] , \nScanOut382[4] , \nScanOut382[3] , 
        \nScanOut382[2] , \nScanOut382[1] , \nScanOut382[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_29[7] , \nOut11_29[6] , \nOut11_29[5] , \nOut11_29[4] , 
        \nOut11_29[3] , \nOut11_29[2] , \nOut11_29[1] , \nOut11_29[0] }), 
        .SouthIn({\nOut11_31[7] , \nOut11_31[6] , \nOut11_31[5] , 
        \nOut11_31[4] , \nOut11_31[3] , \nOut11_31[2] , \nOut11_31[1] , 
        \nOut11_31[0] }), .EastIn({\nOut12_30[7] , \nOut12_30[6] , 
        \nOut12_30[5] , \nOut12_30[4] , \nOut12_30[3] , \nOut12_30[2] , 
        \nOut12_30[1] , \nOut12_30[0] }), .WestIn({\nOut10_30[7] , 
        \nOut10_30[6] , \nOut10_30[5] , \nOut10_30[4] , \nOut10_30[3] , 
        \nOut10_30[2] , \nOut10_30[1] , \nOut10_30[0] }), .Out({\nOut11_30[7] , 
        \nOut11_30[6] , \nOut11_30[5] , \nOut11_30[4] , \nOut11_30[3] , 
        \nOut11_30[2] , \nOut11_30[1] , \nOut11_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_871 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut872[7] , \nScanOut872[6] , 
        \nScanOut872[5] , \nScanOut872[4] , \nScanOut872[3] , \nScanOut872[2] , 
        \nScanOut872[1] , \nScanOut872[0] }), .ScanOut({\nScanOut871[7] , 
        \nScanOut871[6] , \nScanOut871[5] , \nScanOut871[4] , \nScanOut871[3] , 
        \nScanOut871[2] , \nScanOut871[1] , \nScanOut871[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_6[7] , \nOut27_6[6] , \nOut27_6[5] , \nOut27_6[4] , 
        \nOut27_6[3] , \nOut27_6[2] , \nOut27_6[1] , \nOut27_6[0] }), 
        .SouthIn({\nOut27_8[7] , \nOut27_8[6] , \nOut27_8[5] , \nOut27_8[4] , 
        \nOut27_8[3] , \nOut27_8[2] , \nOut27_8[1] , \nOut27_8[0] }), .EastIn(
        {\nOut28_7[7] , \nOut28_7[6] , \nOut28_7[5] , \nOut28_7[4] , 
        \nOut28_7[3] , \nOut28_7[2] , \nOut28_7[1] , \nOut28_7[0] }), .WestIn(
        {\nOut26_7[7] , \nOut26_7[6] , \nOut26_7[5] , \nOut26_7[4] , 
        \nOut26_7[3] , \nOut26_7[2] , \nOut26_7[1] , \nOut26_7[0] }), .Out({
        \nOut27_7[7] , \nOut27_7[6] , \nOut27_7[5] , \nOut27_7[4] , 
        \nOut27_7[3] , \nOut27_7[2] , \nOut27_7[1] , \nOut27_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_403 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut404[7] , \nScanOut404[6] , 
        \nScanOut404[5] , \nScanOut404[4] , \nScanOut404[3] , \nScanOut404[2] , 
        \nScanOut404[1] , \nScanOut404[0] }), .ScanOut({\nScanOut403[7] , 
        \nScanOut403[6] , \nScanOut403[5] , \nScanOut403[4] , \nScanOut403[3] , 
        \nScanOut403[2] , \nScanOut403[1] , \nScanOut403[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_18[7] , \nOut12_18[6] , \nOut12_18[5] , \nOut12_18[4] , 
        \nOut12_18[3] , \nOut12_18[2] , \nOut12_18[1] , \nOut12_18[0] }), 
        .SouthIn({\nOut12_20[7] , \nOut12_20[6] , \nOut12_20[5] , 
        \nOut12_20[4] , \nOut12_20[3] , \nOut12_20[2] , \nOut12_20[1] , 
        \nOut12_20[0] }), .EastIn({\nOut13_19[7] , \nOut13_19[6] , 
        \nOut13_19[5] , \nOut13_19[4] , \nOut13_19[3] , \nOut13_19[2] , 
        \nOut13_19[1] , \nOut13_19[0] }), .WestIn({\nOut11_19[7] , 
        \nOut11_19[6] , \nOut11_19[5] , \nOut11_19[4] , \nOut11_19[3] , 
        \nOut11_19[2] , \nOut11_19[1] , \nOut11_19[0] }), .Out({\nOut12_19[7] , 
        \nOut12_19[6] , \nOut12_19[5] , \nOut12_19[4] , \nOut12_19[3] , 
        \nOut12_19[2] , \nOut12_19[1] , \nOut12_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_235 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut236[7] , \nScanOut236[6] , 
        \nScanOut236[5] , \nScanOut236[4] , \nScanOut236[3] , \nScanOut236[2] , 
        \nScanOut236[1] , \nScanOut236[0] }), .ScanOut({\nScanOut235[7] , 
        \nScanOut235[6] , \nScanOut235[5] , \nScanOut235[4] , \nScanOut235[3] , 
        \nScanOut235[2] , \nScanOut235[1] , \nScanOut235[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_10[7] , \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , 
        \nOut7_10[3] , \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }), 
        .SouthIn({\nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }), .EastIn(
        {\nOut8_11[7] , \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , 
        \nOut8_11[3] , \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }), .WestIn(
        {\nOut6_11[7] , \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , 
        \nOut6_11[3] , \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }), .Out({
        \nOut7_11[7] , \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , 
        \nOut7_11[3] , \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_593 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut594[7] , \nScanOut594[6] , 
        \nScanOut594[5] , \nScanOut594[4] , \nScanOut594[3] , \nScanOut594[2] , 
        \nScanOut594[1] , \nScanOut594[0] }), .ScanOut({\nScanOut593[7] , 
        \nScanOut593[6] , \nScanOut593[5] , \nScanOut593[4] , \nScanOut593[3] , 
        \nScanOut593[2] , \nScanOut593[1] , \nScanOut593[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_16[7] , \nOut18_16[6] , \nOut18_16[5] , \nOut18_16[4] , 
        \nOut18_16[3] , \nOut18_16[2] , \nOut18_16[1] , \nOut18_16[0] }), 
        .SouthIn({\nOut18_18[7] , \nOut18_18[6] , \nOut18_18[5] , 
        \nOut18_18[4] , \nOut18_18[3] , \nOut18_18[2] , \nOut18_18[1] , 
        \nOut18_18[0] }), .EastIn({\nOut19_17[7] , \nOut19_17[6] , 
        \nOut19_17[5] , \nOut19_17[4] , \nOut19_17[3] , \nOut19_17[2] , 
        \nOut19_17[1] , \nOut19_17[0] }), .WestIn({\nOut17_17[7] , 
        \nOut17_17[6] , \nOut17_17[5] , \nOut17_17[4] , \nOut17_17[3] , 
        \nOut17_17[2] , \nOut17_17[1] , \nOut17_17[0] }), .Out({\nOut18_17[7] , 
        \nOut18_17[6] , \nOut18_17[5] , \nOut18_17[4] , \nOut18_17[3] , 
        \nOut18_17[2] , \nOut18_17[1] , \nOut18_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_856 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut857[7] , \nScanOut857[6] , 
        \nScanOut857[5] , \nScanOut857[4] , \nScanOut857[3] , \nScanOut857[2] , 
        \nScanOut857[1] , \nScanOut857[0] }), .ScanOut({\nScanOut856[7] , 
        \nScanOut856[6] , \nScanOut856[5] , \nScanOut856[4] , \nScanOut856[3] , 
        \nScanOut856[2] , \nScanOut856[1] , \nScanOut856[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_23[7] , \nOut26_23[6] , \nOut26_23[5] , \nOut26_23[4] , 
        \nOut26_23[3] , \nOut26_23[2] , \nOut26_23[1] , \nOut26_23[0] }), 
        .SouthIn({\nOut26_25[7] , \nOut26_25[6] , \nOut26_25[5] , 
        \nOut26_25[4] , \nOut26_25[3] , \nOut26_25[2] , \nOut26_25[1] , 
        \nOut26_25[0] }), .EastIn({\nOut27_24[7] , \nOut27_24[6] , 
        \nOut27_24[5] , \nOut27_24[4] , \nOut27_24[3] , \nOut27_24[2] , 
        \nOut27_24[1] , \nOut27_24[0] }), .WestIn({\nOut25_24[7] , 
        \nOut25_24[6] , \nOut25_24[5] , \nOut25_24[4] , \nOut25_24[3] , 
        \nOut25_24[2] , \nOut25_24[1] , \nOut25_24[0] }), .Out({\nOut26_24[7] , 
        \nOut26_24[6] , \nOut26_24[5] , \nOut26_24[4] , \nOut26_24[3] , 
        \nOut26_24[2] , \nOut26_24[1] , \nOut26_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_424 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut425[7] , \nScanOut425[6] , 
        \nScanOut425[5] , \nScanOut425[4] , \nScanOut425[3] , \nScanOut425[2] , 
        \nScanOut425[1] , \nScanOut425[0] }), .ScanOut({\nScanOut424[7] , 
        \nScanOut424[6] , \nScanOut424[5] , \nScanOut424[4] , \nScanOut424[3] , 
        \nScanOut424[2] , \nScanOut424[1] , \nScanOut424[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }), 
        .SouthIn({\nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , \nOut13_9[4] , 
        \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , \nOut13_9[0] }), .EastIn(
        {\nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }), .WestIn(
        {\nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }), .Out({
        \nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_105 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut106[7] , \nScanOut106[6] , 
        \nScanOut106[5] , \nScanOut106[4] , \nScanOut106[3] , \nScanOut106[2] , 
        \nScanOut106[1] , \nScanOut106[0] }), .ScanOut({\nScanOut105[7] , 
        \nScanOut105[6] , \nScanOut105[5] , \nScanOut105[4] , \nScanOut105[3] , 
        \nScanOut105[2] , \nScanOut105[1] , \nScanOut105[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_8[7] , \nOut3_8[6] , \nOut3_8[5] , \nOut3_8[4] , \nOut3_8[3] , 
        \nOut3_8[2] , \nOut3_8[1] , \nOut3_8[0] }), .SouthIn({\nOut3_10[7] , 
        \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , \nOut3_10[3] , 
        \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }), .EastIn({\nOut4_9[7] , 
        \nOut4_9[6] , \nOut4_9[5] , \nOut4_9[4] , \nOut4_9[3] , \nOut4_9[2] , 
        \nOut4_9[1] , \nOut4_9[0] }), .WestIn({\nOut2_9[7] , \nOut2_9[6] , 
        \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , \nOut2_9[1] , 
        \nOut2_9[0] }), .Out({\nOut3_9[7] , \nOut3_9[6] , \nOut3_9[5] , 
        \nOut3_9[4] , \nOut3_9[3] , \nOut3_9[2] , \nOut3_9[1] , \nOut3_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_684 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut685[7] , \nScanOut685[6] , 
        \nScanOut685[5] , \nScanOut685[4] , \nScanOut685[3] , \nScanOut685[2] , 
        \nScanOut685[1] , \nScanOut685[0] }), .ScanOut({\nScanOut684[7] , 
        \nScanOut684[6] , \nScanOut684[5] , \nScanOut684[4] , \nScanOut684[3] , 
        \nScanOut684[2] , \nScanOut684[1] , \nScanOut684[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_11[7] , \nOut21_11[6] , \nOut21_11[5] , \nOut21_11[4] , 
        \nOut21_11[3] , \nOut21_11[2] , \nOut21_11[1] , \nOut21_11[0] }), 
        .SouthIn({\nOut21_13[7] , \nOut21_13[6] , \nOut21_13[5] , 
        \nOut21_13[4] , \nOut21_13[3] , \nOut21_13[2] , \nOut21_13[1] , 
        \nOut21_13[0] }), .EastIn({\nOut22_12[7] , \nOut22_12[6] , 
        \nOut22_12[5] , \nOut22_12[4] , \nOut22_12[3] , \nOut22_12[2] , 
        \nOut22_12[1] , \nOut22_12[0] }), .WestIn({\nOut20_12[7] , 
        \nOut20_12[6] , \nOut20_12[5] , \nOut20_12[4] , \nOut20_12[3] , 
        \nOut20_12[2] , \nOut20_12[1] , \nOut20_12[0] }), .Out({\nOut21_12[7] , 
        \nOut21_12[6] , \nOut21_12[5] , \nOut21_12[4] , \nOut21_12[3] , 
        \nOut21_12[2] , \nOut21_12[1] , \nOut21_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1012 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1013[7] , \nScanOut1013[6] , 
        \nScanOut1013[5] , \nScanOut1013[4] , \nScanOut1013[3] , 
        \nScanOut1013[2] , \nScanOut1013[1] , \nScanOut1013[0] }), .ScanOut({
        \nScanOut1012[7] , \nScanOut1012[6] , \nScanOut1012[5] , 
        \nScanOut1012[4] , \nScanOut1012[3] , \nScanOut1012[2] , 
        \nScanOut1012[1] , \nScanOut1012[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_20[7] , \nOut31_20[6] , \nOut31_20[5] , 
        \nOut31_20[4] , \nOut31_20[3] , \nOut31_20[2] , \nOut31_20[1] , 
        \nOut31_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_130 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut131[7] , \nScanOut131[6] , 
        \nScanOut131[5] , \nScanOut131[4] , \nScanOut131[3] , \nScanOut131[2] , 
        \nScanOut131[1] , \nScanOut131[0] }), .ScanOut({\nScanOut130[7] , 
        \nScanOut130[6] , \nScanOut130[5] , \nScanOut130[4] , \nScanOut130[3] , 
        \nScanOut130[2] , \nScanOut130[1] , \nScanOut130[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_1[7] , \nOut4_1[6] , \nOut4_1[5] , \nOut4_1[4] , \nOut4_1[3] , 
        \nOut4_1[2] , \nOut4_1[1] , \nOut4_1[0] }), .SouthIn({\nOut4_3[7] , 
        \nOut4_3[6] , \nOut4_3[5] , \nOut4_3[4] , \nOut4_3[3] , \nOut4_3[2] , 
        \nOut4_3[1] , \nOut4_3[0] }), .EastIn({\nOut5_2[7] , \nOut5_2[6] , 
        \nOut5_2[5] , \nOut5_2[4] , \nOut5_2[3] , \nOut5_2[2] , \nOut5_2[1] , 
        \nOut5_2[0] }), .WestIn({\nOut3_2[7] , \nOut3_2[6] , \nOut3_2[5] , 
        \nOut3_2[4] , \nOut3_2[3] , \nOut3_2[2] , \nOut3_2[1] , \nOut3_2[0] }), 
        .Out({\nOut4_2[7] , \nOut4_2[6] , \nOut4_2[5] , \nOut4_2[4] , 
        \nOut4_2[3] , \nOut4_2[2] , \nOut4_2[1] , \nOut4_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_299 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut300[7] , \nScanOut300[6] , 
        \nScanOut300[5] , \nScanOut300[4] , \nScanOut300[3] , \nScanOut300[2] , 
        \nScanOut300[1] , \nScanOut300[0] }), .ScanOut({\nScanOut299[7] , 
        \nScanOut299[6] , \nScanOut299[5] , \nScanOut299[4] , \nScanOut299[3] , 
        \nScanOut299[2] , \nScanOut299[1] , \nScanOut299[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_10[7] , \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , 
        \nOut9_10[3] , \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }), 
        .SouthIn({\nOut9_12[7] , \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , 
        \nOut9_12[3] , \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }), .EastIn(
        {\nOut10_11[7] , \nOut10_11[6] , \nOut10_11[5] , \nOut10_11[4] , 
        \nOut10_11[3] , \nOut10_11[2] , \nOut10_11[1] , \nOut10_11[0] }), 
        .WestIn({\nOut8_11[7] , \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , 
        \nOut8_11[3] , \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }), .Out({
        \nOut9_11[7] , \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , 
        \nOut9_11[3] , \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_309 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut310[7] , \nScanOut310[6] , 
        \nScanOut310[5] , \nScanOut310[4] , \nScanOut310[3] , \nScanOut310[2] , 
        \nScanOut310[1] , \nScanOut310[0] }), .ScanOut({\nScanOut309[7] , 
        \nScanOut309[6] , \nScanOut309[5] , \nScanOut309[4] , \nScanOut309[3] , 
        \nScanOut309[2] , \nScanOut309[1] , \nScanOut309[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_20[7] , \nOut9_20[6] , \nOut9_20[5] , \nOut9_20[4] , 
        \nOut9_20[3] , \nOut9_20[2] , \nOut9_20[1] , \nOut9_20[0] }), 
        .SouthIn({\nOut9_22[7] , \nOut9_22[6] , \nOut9_22[5] , \nOut9_22[4] , 
        \nOut9_22[3] , \nOut9_22[2] , \nOut9_22[1] , \nOut9_22[0] }), .EastIn(
        {\nOut10_21[7] , \nOut10_21[6] , \nOut10_21[5] , \nOut10_21[4] , 
        \nOut10_21[3] , \nOut10_21[2] , \nOut10_21[1] , \nOut10_21[0] }), 
        .WestIn({\nOut8_21[7] , \nOut8_21[6] , \nOut8_21[5] , \nOut8_21[4] , 
        \nOut8_21[3] , \nOut8_21[2] , \nOut8_21[1] , \nOut8_21[0] }), .Out({
        \nOut9_21[7] , \nOut9_21[6] , \nOut9_21[5] , \nOut9_21[4] , 
        \nOut9_21[3] , \nOut9_21[2] , \nOut9_21[1] , \nOut9_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_628 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut629[7] , \nScanOut629[6] , 
        \nScanOut629[5] , \nScanOut629[4] , \nScanOut629[3] , \nScanOut629[2] , 
        \nScanOut629[1] , \nScanOut629[0] }), .ScanOut({\nScanOut628[7] , 
        \nScanOut628[6] , \nScanOut628[5] , \nScanOut628[4] , \nScanOut628[3] , 
        \nScanOut628[2] , \nScanOut628[1] , \nScanOut628[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_19[7] , \nOut19_19[6] , \nOut19_19[5] , \nOut19_19[4] , 
        \nOut19_19[3] , \nOut19_19[2] , \nOut19_19[1] , \nOut19_19[0] }), 
        .SouthIn({\nOut19_21[7] , \nOut19_21[6] , \nOut19_21[5] , 
        \nOut19_21[4] , \nOut19_21[3] , \nOut19_21[2] , \nOut19_21[1] , 
        \nOut19_21[0] }), .EastIn({\nOut20_20[7] , \nOut20_20[6] , 
        \nOut20_20[5] , \nOut20_20[4] , \nOut20_20[3] , \nOut20_20[2] , 
        \nOut20_20[1] , \nOut20_20[0] }), .WestIn({\nOut18_20[7] , 
        \nOut18_20[6] , \nOut18_20[5] , \nOut18_20[4] , \nOut18_20[3] , 
        \nOut18_20[2] , \nOut18_20[1] , \nOut18_20[0] }), .Out({\nOut19_20[7] , 
        \nOut19_20[6] , \nOut19_20[5] , \nOut19_20[4] , \nOut19_20[3] , 
        \nOut19_20[2] , \nOut19_20[1] , \nOut19_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_714 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut715[7] , \nScanOut715[6] , 
        \nScanOut715[5] , \nScanOut715[4] , \nScanOut715[3] , \nScanOut715[2] , 
        \nScanOut715[1] , \nScanOut715[0] }), .ScanOut({\nScanOut714[7] , 
        \nScanOut714[6] , \nScanOut714[5] , \nScanOut714[4] , \nScanOut714[3] , 
        \nScanOut714[2] , \nScanOut714[1] , \nScanOut714[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_9[7] , \nOut22_9[6] , \nOut22_9[5] , \nOut22_9[4] , 
        \nOut22_9[3] , \nOut22_9[2] , \nOut22_9[1] , \nOut22_9[0] }), 
        .SouthIn({\nOut22_11[7] , \nOut22_11[6] , \nOut22_11[5] , 
        \nOut22_11[4] , \nOut22_11[3] , \nOut22_11[2] , \nOut22_11[1] , 
        \nOut22_11[0] }), .EastIn({\nOut23_10[7] , \nOut23_10[6] , 
        \nOut23_10[5] , \nOut23_10[4] , \nOut23_10[3] , \nOut23_10[2] , 
        \nOut23_10[1] , \nOut23_10[0] }), .WestIn({\nOut21_10[7] , 
        \nOut21_10[6] , \nOut21_10[5] , \nOut21_10[4] , \nOut21_10[3] , 
        \nOut21_10[2] , \nOut21_10[1] , \nOut21_10[0] }), .Out({\nOut22_10[7] , 
        \nOut22_10[6] , \nOut22_10[5] , \nOut22_10[4] , \nOut22_10[3] , 
        \nOut22_10[2] , \nOut22_10[1] , \nOut22_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_488 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut489[7] , \nScanOut489[6] , 
        \nScanOut489[5] , \nScanOut489[4] , \nScanOut489[3] , \nScanOut489[2] , 
        \nScanOut489[1] , \nScanOut489[0] }), .ScanOut({\nScanOut488[7] , 
        \nScanOut488[6] , \nScanOut488[5] , \nScanOut488[4] , \nScanOut488[3] , 
        \nScanOut488[2] , \nScanOut488[1] , \nScanOut488[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_7[7] , \nOut15_7[6] , \nOut15_7[5] , \nOut15_7[4] , 
        \nOut15_7[3] , \nOut15_7[2] , \nOut15_7[1] , \nOut15_7[0] }), 
        .SouthIn({\nOut15_9[7] , \nOut15_9[6] , \nOut15_9[5] , \nOut15_9[4] , 
        \nOut15_9[3] , \nOut15_9[2] , \nOut15_9[1] , \nOut15_9[0] }), .EastIn(
        {\nOut16_8[7] , \nOut16_8[6] , \nOut16_8[5] , \nOut16_8[4] , 
        \nOut16_8[3] , \nOut16_8[2] , \nOut16_8[1] , \nOut16_8[0] }), .WestIn(
        {\nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }), .Out({
        \nOut15_8[7] , \nOut15_8[6] , \nOut15_8[5] , \nOut15_8[4] , 
        \nOut15_8[3] , \nOut15_8[2] , \nOut15_8[1] , \nOut15_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_518 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut519[7] , \nScanOut519[6] , 
        \nScanOut519[5] , \nScanOut519[4] , \nScanOut519[3] , \nScanOut519[2] , 
        \nScanOut519[1] , \nScanOut519[0] }), .ScanOut({\nScanOut518[7] , 
        \nScanOut518[6] , \nScanOut518[5] , \nScanOut518[4] , \nScanOut518[3] , 
        \nScanOut518[2] , \nScanOut518[1] , \nScanOut518[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_5[7] , \nOut16_5[6] , \nOut16_5[5] , \nOut16_5[4] , 
        \nOut16_5[3] , \nOut16_5[2] , \nOut16_5[1] , \nOut16_5[0] }), 
        .SouthIn({\nOut16_7[7] , \nOut16_7[6] , \nOut16_7[5] , \nOut16_7[4] , 
        \nOut16_7[3] , \nOut16_7[2] , \nOut16_7[1] , \nOut16_7[0] }), .EastIn(
        {\nOut17_6[7] , \nOut17_6[6] , \nOut17_6[5] , \nOut17_6[4] , 
        \nOut17_6[3] , \nOut17_6[2] , \nOut17_6[1] , \nOut17_6[0] }), .WestIn(
        {\nOut15_6[7] , \nOut15_6[6] , \nOut15_6[5] , \nOut15_6[4] , 
        \nOut15_6[3] , \nOut15_6[2] , \nOut15_6[1] , \nOut15_6[0] }), .Out({
        \nOut16_6[7] , \nOut16_6[6] , \nOut16_6[5] , \nOut16_6[4] , 
        \nOut16_6[3] , \nOut16_6[2] , \nOut16_6[1] , \nOut16_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_978 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut979[7] , \nScanOut979[6] , 
        \nScanOut979[5] , \nScanOut979[4] , \nScanOut979[3] , \nScanOut979[2] , 
        \nScanOut979[1] , \nScanOut979[0] }), .ScanOut({\nScanOut978[7] , 
        \nScanOut978[6] , \nScanOut978[5] , \nScanOut978[4] , \nScanOut978[3] , 
        \nScanOut978[2] , \nScanOut978[1] , \nScanOut978[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_17[7] , \nOut30_17[6] , \nOut30_17[5] , \nOut30_17[4] , 
        \nOut30_17[3] , \nOut30_17[2] , \nOut30_17[1] , \nOut30_17[0] }), 
        .SouthIn({\nOut30_19[7] , \nOut30_19[6] , \nOut30_19[5] , 
        \nOut30_19[4] , \nOut30_19[3] , \nOut30_19[2] , \nOut30_19[1] , 
        \nOut30_19[0] }), .EastIn({\nOut31_18[7] , \nOut31_18[6] , 
        \nOut31_18[5] , \nOut31_18[4] , \nOut31_18[3] , \nOut31_18[2] , 
        \nOut31_18[1] , \nOut31_18[0] }), .WestIn({\nOut29_18[7] , 
        \nOut29_18[6] , \nOut29_18[5] , \nOut29_18[4] , \nOut29_18[3] , 
        \nOut29_18[2] , \nOut29_18[1] , \nOut29_18[0] }), .Out({\nOut30_18[7] , 
        \nOut30_18[6] , \nOut30_18[5] , \nOut30_18[4] , \nOut30_18[3] , 
        \nOut30_18[2] , \nOut30_18[1] , \nOut30_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_200 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut201[7] , \nScanOut201[6] , 
        \nScanOut201[5] , \nScanOut201[4] , \nScanOut201[3] , \nScanOut201[2] , 
        \nScanOut201[1] , \nScanOut201[0] }), .ScanOut({\nScanOut200[7] , 
        \nScanOut200[6] , \nScanOut200[5] , \nScanOut200[4] , \nScanOut200[3] , 
        \nScanOut200[2] , \nScanOut200[1] , \nScanOut200[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_7[7] , \nOut6_7[6] , \nOut6_7[5] , \nOut6_7[4] , \nOut6_7[3] , 
        \nOut6_7[2] , \nOut6_7[1] , \nOut6_7[0] }), .SouthIn({\nOut6_9[7] , 
        \nOut6_9[6] , \nOut6_9[5] , \nOut6_9[4] , \nOut6_9[3] , \nOut6_9[2] , 
        \nOut6_9[1] , \nOut6_9[0] }), .EastIn({\nOut7_8[7] , \nOut7_8[6] , 
        \nOut7_8[5] , \nOut7_8[4] , \nOut7_8[3] , \nOut7_8[2] , \nOut7_8[1] , 
        \nOut7_8[0] }), .WestIn({\nOut5_8[7] , \nOut5_8[6] , \nOut5_8[5] , 
        \nOut5_8[4] , \nOut5_8[3] , \nOut5_8[2] , \nOut5_8[1] , \nOut5_8[0] }), 
        .Out({\nOut6_8[7] , \nOut6_8[6] , \nOut6_8[5] , \nOut6_8[4] , 
        \nOut6_8[3] , \nOut6_8[2] , \nOut6_8[1] , \nOut6_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_721 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut722[7] , \nScanOut722[6] , 
        \nScanOut722[5] , \nScanOut722[4] , \nScanOut722[3] , \nScanOut722[2] , 
        \nScanOut722[1] , \nScanOut722[0] }), .ScanOut({\nScanOut721[7] , 
        \nScanOut721[6] , \nScanOut721[5] , \nScanOut721[4] , \nScanOut721[3] , 
        \nScanOut721[2] , \nScanOut721[1] , \nScanOut721[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_16[7] , \nOut22_16[6] , \nOut22_16[5] , \nOut22_16[4] , 
        \nOut22_16[3] , \nOut22_16[2] , \nOut22_16[1] , \nOut22_16[0] }), 
        .SouthIn({\nOut22_18[7] , \nOut22_18[6] , \nOut22_18[5] , 
        \nOut22_18[4] , \nOut22_18[3] , \nOut22_18[2] , \nOut22_18[1] , 
        \nOut22_18[0] }), .EastIn({\nOut23_17[7] , \nOut23_17[6] , 
        \nOut23_17[5] , \nOut23_17[4] , \nOut23_17[3] , \nOut23_17[2] , 
        \nOut23_17[1] , \nOut23_17[0] }), .WestIn({\nOut21_17[7] , 
        \nOut21_17[6] , \nOut21_17[5] , \nOut21_17[4] , \nOut21_17[3] , 
        \nOut21_17[2] , \nOut21_17[1] , \nOut21_17[0] }), .Out({\nOut22_17[7] , 
        \nOut22_17[6] , \nOut22_17[5] , \nOut22_17[4] , \nOut22_17[3] , 
        \nOut22_17[2] , \nOut22_17[1] , \nOut22_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_227 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut228[7] , \nScanOut228[6] , 
        \nScanOut228[5] , \nScanOut228[4] , \nScanOut228[3] , \nScanOut228[2] , 
        \nScanOut228[1] , \nScanOut228[0] }), .ScanOut({\nScanOut227[7] , 
        \nScanOut227[6] , \nScanOut227[5] , \nScanOut227[4] , \nScanOut227[3] , 
        \nScanOut227[2] , \nScanOut227[1] , \nScanOut227[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_2[7] , \nOut7_2[6] , \nOut7_2[5] , \nOut7_2[4] , \nOut7_2[3] , 
        \nOut7_2[2] , \nOut7_2[1] , \nOut7_2[0] }), .SouthIn({\nOut7_4[7] , 
        \nOut7_4[6] , \nOut7_4[5] , \nOut7_4[4] , \nOut7_4[3] , \nOut7_4[2] , 
        \nOut7_4[1] , \nOut7_4[0] }), .EastIn({\nOut8_3[7] , \nOut8_3[6] , 
        \nOut8_3[5] , \nOut8_3[4] , \nOut8_3[3] , \nOut8_3[2] , \nOut8_3[1] , 
        \nOut8_3[0] }), .WestIn({\nOut6_3[7] , \nOut6_3[6] , \nOut6_3[5] , 
        \nOut6_3[4] , \nOut6_3[3] , \nOut6_3[2] , \nOut6_3[1] , \nOut6_3[0] }), 
        .Out({\nOut7_3[7] , \nOut7_3[6] , \nOut7_3[5] , \nOut7_3[4] , 
        \nOut7_3[3] , \nOut7_3[2] , \nOut7_3[1] , \nOut7_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_390 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut391[7] , \nScanOut391[6] , 
        \nScanOut391[5] , \nScanOut391[4] , \nScanOut391[3] , \nScanOut391[2] , 
        \nScanOut391[1] , \nScanOut391[0] }), .ScanOut({\nScanOut390[7] , 
        \nScanOut390[6] , \nScanOut390[5] , \nScanOut390[4] , \nScanOut390[3] , 
        \nScanOut390[2] , \nScanOut390[1] , \nScanOut390[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }), 
        .SouthIn({\nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }), .EastIn(
        {\nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }), .WestIn(
        {\nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }), .Out({
        \nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_581 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut582[7] , \nScanOut582[6] , 
        \nScanOut582[5] , \nScanOut582[4] , \nScanOut582[3] , \nScanOut582[2] , 
        \nScanOut582[1] , \nScanOut582[0] }), .ScanOut({\nScanOut581[7] , 
        \nScanOut581[6] , \nScanOut581[5] , \nScanOut581[4] , \nScanOut581[3] , 
        \nScanOut581[2] , \nScanOut581[1] , \nScanOut581[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_4[7] , \nOut18_4[6] , \nOut18_4[5] , \nOut18_4[4] , 
        \nOut18_4[3] , \nOut18_4[2] , \nOut18_4[1] , \nOut18_4[0] }), 
        .SouthIn({\nOut18_6[7] , \nOut18_6[6] , \nOut18_6[5] , \nOut18_6[4] , 
        \nOut18_6[3] , \nOut18_6[2] , \nOut18_6[1] , \nOut18_6[0] }), .EastIn(
        {\nOut19_5[7] , \nOut19_5[6] , \nOut19_5[5] , \nOut19_5[4] , 
        \nOut19_5[3] , \nOut19_5[2] , \nOut19_5[1] , \nOut19_5[0] }), .WestIn(
        {\nOut17_5[7] , \nOut17_5[6] , \nOut17_5[5] , \nOut17_5[4] , 
        \nOut17_5[3] , \nOut17_5[2] , \nOut17_5[1] , \nOut17_5[0] }), .Out({
        \nOut18_5[7] , \nOut18_5[6] , \nOut18_5[5] , \nOut18_5[4] , 
        \nOut18_5[3] , \nOut18_5[2] , \nOut18_5[1] , \nOut18_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_411 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut412[7] , \nScanOut412[6] , 
        \nScanOut412[5] , \nScanOut412[4] , \nScanOut412[3] , \nScanOut412[2] , 
        \nScanOut412[1] , \nScanOut412[0] }), .ScanOut({\nScanOut411[7] , 
        \nScanOut411[6] , \nScanOut411[5] , \nScanOut411[4] , \nScanOut411[3] , 
        \nScanOut411[2] , \nScanOut411[1] , \nScanOut411[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_26[7] , \nOut12_26[6] , \nOut12_26[5] , \nOut12_26[4] , 
        \nOut12_26[3] , \nOut12_26[2] , \nOut12_26[1] , \nOut12_26[0] }), 
        .SouthIn({\nOut12_28[7] , \nOut12_28[6] , \nOut12_28[5] , 
        \nOut12_28[4] , \nOut12_28[3] , \nOut12_28[2] , \nOut12_28[1] , 
        \nOut12_28[0] }), .EastIn({\nOut13_27[7] , \nOut13_27[6] , 
        \nOut13_27[5] , \nOut13_27[4] , \nOut13_27[3] , \nOut13_27[2] , 
        \nOut13_27[1] , \nOut13_27[0] }), .WestIn({\nOut11_27[7] , 
        \nOut11_27[6] , \nOut11_27[5] , \nOut11_27[4] , \nOut11_27[3] , 
        \nOut11_27[2] , \nOut11_27[1] , \nOut11_27[0] }), .Out({\nOut12_27[7] , 
        \nOut12_27[6] , \nOut12_27[5] , \nOut12_27[4] , \nOut12_27[3] , 
        \nOut12_27[2] , \nOut12_27[1] , \nOut12_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_436 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut437[7] , \nScanOut437[6] , 
        \nScanOut437[5] , \nScanOut437[4] , \nScanOut437[3] , \nScanOut437[2] , 
        \nScanOut437[1] , \nScanOut437[0] }), .ScanOut({\nScanOut436[7] , 
        \nScanOut436[6] , \nScanOut436[5] , \nScanOut436[4] , \nScanOut436[3] , 
        \nScanOut436[2] , \nScanOut436[1] , \nScanOut436[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_19[7] , \nOut13_19[6] , \nOut13_19[5] , \nOut13_19[4] , 
        \nOut13_19[3] , \nOut13_19[2] , \nOut13_19[1] , \nOut13_19[0] }), 
        .SouthIn({\nOut13_21[7] , \nOut13_21[6] , \nOut13_21[5] , 
        \nOut13_21[4] , \nOut13_21[3] , \nOut13_21[2] , \nOut13_21[1] , 
        \nOut13_21[0] }), .EastIn({\nOut14_20[7] , \nOut14_20[6] , 
        \nOut14_20[5] , \nOut14_20[4] , \nOut14_20[3] , \nOut14_20[2] , 
        \nOut14_20[1] , \nOut14_20[0] }), .WestIn({\nOut12_20[7] , 
        \nOut12_20[6] , \nOut12_20[5] , \nOut12_20[4] , \nOut12_20[3] , 
        \nOut12_20[2] , \nOut12_20[1] , \nOut12_20[0] }), .Out({\nOut13_20[7] , 
        \nOut13_20[6] , \nOut13_20[5] , \nOut13_20[4] , \nOut13_20[3] , 
        \nOut13_20[2] , \nOut13_20[1] , \nOut13_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_863 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut864[7] , \nScanOut864[6] , 
        \nScanOut864[5] , \nScanOut864[4] , \nScanOut864[3] , \nScanOut864[2] , 
        \nScanOut864[1] , \nScanOut864[0] }), .ScanOut({\nScanOut863[7] , 
        \nScanOut863[6] , \nScanOut863[5] , \nScanOut863[4] , \nScanOut863[3] , 
        \nScanOut863[2] , \nScanOut863[1] , \nScanOut863[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut26_31[7] , \nOut26_31[6] , 
        \nOut26_31[5] , \nOut26_31[4] , \nOut26_31[3] , \nOut26_31[2] , 
        \nOut26_31[1] , \nOut26_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_844 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut845[7] , \nScanOut845[6] , 
        \nScanOut845[5] , \nScanOut845[4] , \nScanOut845[3] , \nScanOut845[2] , 
        \nScanOut845[1] , \nScanOut845[0] }), .ScanOut({\nScanOut844[7] , 
        \nScanOut844[6] , \nScanOut844[5] , \nScanOut844[4] , \nScanOut844[3] , 
        \nScanOut844[2] , \nScanOut844[1] , \nScanOut844[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_11[7] , \nOut26_11[6] , \nOut26_11[5] , \nOut26_11[4] , 
        \nOut26_11[3] , \nOut26_11[2] , \nOut26_11[1] , \nOut26_11[0] }), 
        .SouthIn({\nOut26_13[7] , \nOut26_13[6] , \nOut26_13[5] , 
        \nOut26_13[4] , \nOut26_13[3] , \nOut26_13[2] , \nOut26_13[1] , 
        \nOut26_13[0] }), .EastIn({\nOut27_12[7] , \nOut27_12[6] , 
        \nOut27_12[5] , \nOut27_12[4] , \nOut27_12[3] , \nOut27_12[2] , 
        \nOut27_12[1] , \nOut27_12[0] }), .WestIn({\nOut25_12[7] , 
        \nOut25_12[6] , \nOut25_12[5] , \nOut25_12[4] , \nOut25_12[3] , 
        \nOut25_12[2] , \nOut25_12[1] , \nOut25_12[0] }), .Out({\nOut26_12[7] , 
        \nOut26_12[6] , \nOut26_12[5] , \nOut26_12[4] , \nOut26_12[3] , 
        \nOut26_12[2] , \nOut26_12[1] , \nOut26_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_117 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut118[7] , \nScanOut118[6] , 
        \nScanOut118[5] , \nScanOut118[4] , \nScanOut118[3] , \nScanOut118[2] , 
        \nScanOut118[1] , \nScanOut118[0] }), .ScanOut({\nScanOut117[7] , 
        \nScanOut117[6] , \nScanOut117[5] , \nScanOut117[4] , \nScanOut117[3] , 
        \nScanOut117[2] , \nScanOut117[1] , \nScanOut117[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_20[7] , \nOut3_20[6] , \nOut3_20[5] , \nOut3_20[4] , 
        \nOut3_20[3] , \nOut3_20[2] , \nOut3_20[1] , \nOut3_20[0] }), 
        .SouthIn({\nOut3_22[7] , \nOut3_22[6] , \nOut3_22[5] , \nOut3_22[4] , 
        \nOut3_22[3] , \nOut3_22[2] , \nOut3_22[1] , \nOut3_22[0] }), .EastIn(
        {\nOut4_21[7] , \nOut4_21[6] , \nOut4_21[5] , \nOut4_21[4] , 
        \nOut4_21[3] , \nOut4_21[2] , \nOut4_21[1] , \nOut4_21[0] }), .WestIn(
        {\nOut2_21[7] , \nOut2_21[6] , \nOut2_21[5] , \nOut2_21[4] , 
        \nOut2_21[3] , \nOut2_21[2] , \nOut2_21[1] , \nOut2_21[0] }), .Out({
        \nOut3_21[7] , \nOut3_21[6] , \nOut3_21[5] , \nOut3_21[4] , 
        \nOut3_21[3] , \nOut3_21[2] , \nOut3_21[1] , \nOut3_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_696 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut697[7] , \nScanOut697[6] , 
        \nScanOut697[5] , \nScanOut697[4] , \nScanOut697[3] , \nScanOut697[2] , 
        \nScanOut697[1] , \nScanOut697[0] }), .ScanOut({\nScanOut696[7] , 
        \nScanOut696[6] , \nScanOut696[5] , \nScanOut696[4] , \nScanOut696[3] , 
        \nScanOut696[2] , \nScanOut696[1] , \nScanOut696[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_23[7] , \nOut21_23[6] , \nOut21_23[5] , \nOut21_23[4] , 
        \nOut21_23[3] , \nOut21_23[2] , \nOut21_23[1] , \nOut21_23[0] }), 
        .SouthIn({\nOut21_25[7] , \nOut21_25[6] , \nOut21_25[5] , 
        \nOut21_25[4] , \nOut21_25[3] , \nOut21_25[2] , \nOut21_25[1] , 
        \nOut21_25[0] }), .EastIn({\nOut22_24[7] , \nOut22_24[6] , 
        \nOut22_24[5] , \nOut22_24[4] , \nOut22_24[3] , \nOut22_24[2] , 
        \nOut22_24[1] , \nOut22_24[0] }), .WestIn({\nOut20_24[7] , 
        \nOut20_24[6] , \nOut20_24[5] , \nOut20_24[4] , \nOut20_24[3] , 
        \nOut20_24[2] , \nOut20_24[1] , \nOut20_24[0] }), .Out({\nOut21_24[7] , 
        \nOut21_24[6] , \nOut21_24[5] , \nOut21_24[4] , \nOut21_24[3] , 
        \nOut21_24[2] , \nOut21_24[1] , \nOut21_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_706 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut707[7] , \nScanOut707[6] , 
        \nScanOut707[5] , \nScanOut707[4] , \nScanOut707[3] , \nScanOut707[2] , 
        \nScanOut707[1] , \nScanOut707[0] }), .ScanOut({\nScanOut706[7] , 
        \nScanOut706[6] , \nScanOut706[5] , \nScanOut706[4] , \nScanOut706[3] , 
        \nScanOut706[2] , \nScanOut706[1] , \nScanOut706[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_1[7] , \nOut22_1[6] , \nOut22_1[5] , \nOut22_1[4] , 
        \nOut22_1[3] , \nOut22_1[2] , \nOut22_1[1] , \nOut22_1[0] }), 
        .SouthIn({\nOut22_3[7] , \nOut22_3[6] , \nOut22_3[5] , \nOut22_3[4] , 
        \nOut22_3[3] , \nOut22_3[2] , \nOut22_3[1] , \nOut22_3[0] }), .EastIn(
        {\nOut23_2[7] , \nOut23_2[6] , \nOut23_2[5] , \nOut23_2[4] , 
        \nOut23_2[3] , \nOut23_2[2] , \nOut23_2[1] , \nOut23_2[0] }), .WestIn(
        {\nOut21_2[7] , \nOut21_2[6] , \nOut21_2[5] , \nOut21_2[4] , 
        \nOut21_2[3] , \nOut21_2[2] , \nOut21_2[1] , \nOut21_2[0] }), .Out({
        \nOut22_2[7] , \nOut22_2[6] , \nOut22_2[5] , \nOut22_2[4] , 
        \nOut22_2[3] , \nOut22_2[2] , \nOut22_2[1] , \nOut22_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1000 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1001[7] , \nScanOut1001[6] , 
        \nScanOut1001[5] , \nScanOut1001[4] , \nScanOut1001[3] , 
        \nScanOut1001[2] , \nScanOut1001[1] , \nScanOut1001[0] }), .ScanOut({
        \nScanOut1000[7] , \nScanOut1000[6] , \nScanOut1000[5] , 
        \nScanOut1000[4] , \nScanOut1000[3] , \nScanOut1000[2] , 
        \nScanOut1000[1] , \nScanOut1000[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_8[7] , \nOut31_8[6] , \nOut31_8[5] , 
        \nOut31_8[4] , \nOut31_8[3] , \nOut31_8[2] , \nOut31_8[1] , 
        \nOut31_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_179 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut180[7] , \nScanOut180[6] , 
        \nScanOut180[5] , \nScanOut180[4] , \nScanOut180[3] , \nScanOut180[2] , 
        \nScanOut180[1] , \nScanOut180[0] }), .ScanOut({\nScanOut179[7] , 
        \nScanOut179[6] , \nScanOut179[5] , \nScanOut179[4] , \nScanOut179[3] , 
        \nScanOut179[2] , \nScanOut179[1] , \nScanOut179[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_18[7] , \nOut5_18[6] , \nOut5_18[5] , \nOut5_18[4] , 
        \nOut5_18[3] , \nOut5_18[2] , \nOut5_18[1] , \nOut5_18[0] }), 
        .SouthIn({\nOut5_20[7] , \nOut5_20[6] , \nOut5_20[5] , \nOut5_20[4] , 
        \nOut5_20[3] , \nOut5_20[2] , \nOut5_20[1] , \nOut5_20[0] }), .EastIn(
        {\nOut6_19[7] , \nOut6_19[6] , \nOut6_19[5] , \nOut6_19[4] , 
        \nOut6_19[3] , \nOut6_19[2] , \nOut6_19[1] , \nOut6_19[0] }), .WestIn(
        {\nOut4_19[7] , \nOut4_19[6] , \nOut4_19[5] , \nOut4_19[4] , 
        \nOut4_19[3] , \nOut4_19[2] , \nOut4_19[1] , \nOut4_19[0] }), .Out({
        \nOut5_19[7] , \nOut5_19[6] , \nOut5_19[5] , \nOut5_19[4] , 
        \nOut5_19[3] , \nOut5_19[2] , \nOut5_19[1] , \nOut5_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_249 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut250[7] , \nScanOut250[6] , 
        \nScanOut250[5] , \nScanOut250[4] , \nScanOut250[3] , \nScanOut250[2] , 
        \nScanOut250[1] , \nScanOut250[0] }), .ScanOut({\nScanOut249[7] , 
        \nScanOut249[6] , \nScanOut249[5] , \nScanOut249[4] , \nScanOut249[3] , 
        \nScanOut249[2] , \nScanOut249[1] , \nScanOut249[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_24[7] , \nOut7_24[6] , \nOut7_24[5] , \nOut7_24[4] , 
        \nOut7_24[3] , \nOut7_24[2] , \nOut7_24[1] , \nOut7_24[0] }), 
        .SouthIn({\nOut7_26[7] , \nOut7_26[6] , \nOut7_26[5] , \nOut7_26[4] , 
        \nOut7_26[3] , \nOut7_26[2] , \nOut7_26[1] , \nOut7_26[0] }), .EastIn(
        {\nOut8_25[7] , \nOut8_25[6] , \nOut8_25[5] , \nOut8_25[4] , 
        \nOut8_25[3] , \nOut8_25[2] , \nOut8_25[1] , \nOut8_25[0] }), .WestIn(
        {\nOut6_25[7] , \nOut6_25[6] , \nOut6_25[5] , \nOut6_25[4] , 
        \nOut6_25[3] , \nOut6_25[2] , \nOut6_25[1] , \nOut6_25[0] }), .Out({
        \nOut7_25[7] , \nOut7_25[6] , \nOut7_25[5] , \nOut7_25[4] , 
        \nOut7_25[3] , \nOut7_25[2] , \nOut7_25[1] , \nOut7_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_458 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut459[7] , \nScanOut459[6] , 
        \nScanOut459[5] , \nScanOut459[4] , \nScanOut459[3] , \nScanOut459[2] , 
        \nScanOut459[1] , \nScanOut459[0] }), .ScanOut({\nScanOut458[7] , 
        \nScanOut458[6] , \nScanOut458[5] , \nScanOut458[4] , \nScanOut458[3] , 
        \nScanOut458[2] , \nScanOut458[1] , \nScanOut458[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , \nOut14_9[4] , 
        \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , \nOut14_9[0] }), 
        .SouthIn({\nOut14_11[7] , \nOut14_11[6] , \nOut14_11[5] , 
        \nOut14_11[4] , \nOut14_11[3] , \nOut14_11[2] , \nOut14_11[1] , 
        \nOut14_11[0] }), .EastIn({\nOut15_10[7] , \nOut15_10[6] , 
        \nOut15_10[5] , \nOut15_10[4] , \nOut15_10[3] , \nOut15_10[2] , 
        \nOut15_10[1] , \nOut15_10[0] }), .WestIn({\nOut13_10[7] , 
        \nOut13_10[6] , \nOut13_10[5] , \nOut13_10[4] , \nOut13_10[3] , 
        \nOut13_10[2] , \nOut13_10[1] , \nOut13_10[0] }), .Out({\nOut14_10[7] , 
        \nOut14_10[6] , \nOut14_10[5] , \nOut14_10[4] , \nOut14_10[3] , 
        \nOut14_10[2] , \nOut14_10[1] , \nOut14_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_352 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut353[7] , \nScanOut353[6] , 
        \nScanOut353[5] , \nScanOut353[4] , \nScanOut353[3] , \nScanOut353[2] , 
        \nScanOut353[1] , \nScanOut353[0] }), .ScanOut({\nScanOut352[7] , 
        \nScanOut352[6] , \nScanOut352[5] , \nScanOut352[4] , \nScanOut352[3] , 
        \nScanOut352[2] , \nScanOut352[1] , \nScanOut352[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut11_0[7] , \nOut11_0[6] , 
        \nOut11_0[5] , \nOut11_0[4] , \nOut11_0[3] , \nOut11_0[2] , 
        \nOut11_0[1] , \nOut11_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_543 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut544[7] , \nScanOut544[6] , 
        \nScanOut544[5] , \nScanOut544[4] , \nScanOut544[3] , \nScanOut544[2] , 
        \nScanOut544[1] , \nScanOut544[0] }), .ScanOut({\nScanOut543[7] , 
        \nScanOut543[6] , \nScanOut543[5] , \nScanOut543[4] , \nScanOut543[3] , 
        \nScanOut543[2] , \nScanOut543[1] , \nScanOut543[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut16_31[7] , \nOut16_31[6] , 
        \nOut16_31[5] , \nOut16_31[4] , \nOut16_31[3] , \nOut16_31[2] , 
        \nOut16_31[1] , \nOut16_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_768 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut769[7] , \nScanOut769[6] , 
        \nScanOut769[5] , \nScanOut769[4] , \nScanOut769[3] , \nScanOut769[2] , 
        \nScanOut769[1] , \nScanOut769[0] }), .ScanOut({\nScanOut768[7] , 
        \nScanOut768[6] , \nScanOut768[5] , \nScanOut768[4] , \nScanOut768[3] , 
        \nScanOut768[2] , \nScanOut768[1] , \nScanOut768[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut24_0[7] , \nOut24_0[6] , 
        \nOut24_0[5] , \nOut24_0[4] , \nOut24_0[3] , \nOut24_0[2] , 
        \nOut24_0[1] , \nOut24_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_673 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut674[7] , \nScanOut674[6] , 
        \nScanOut674[5] , \nScanOut674[4] , \nScanOut674[3] , \nScanOut674[2] , 
        \nScanOut674[1] , \nScanOut674[0] }), .ScanOut({\nScanOut673[7] , 
        \nScanOut673[6] , \nScanOut673[5] , \nScanOut673[4] , \nScanOut673[3] , 
        \nScanOut673[2] , \nScanOut673[1] , \nScanOut673[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_0[7] , \nOut21_0[6] , \nOut21_0[5] , \nOut21_0[4] , 
        \nOut21_0[3] , \nOut21_0[2] , \nOut21_0[1] , \nOut21_0[0] }), 
        .SouthIn({\nOut21_2[7] , \nOut21_2[6] , \nOut21_2[5] , \nOut21_2[4] , 
        \nOut21_2[3] , \nOut21_2[2] , \nOut21_2[1] , \nOut21_2[0] }), .EastIn(
        {\nOut22_1[7] , \nOut22_1[6] , \nOut22_1[5] , \nOut22_1[4] , 
        \nOut22_1[3] , \nOut22_1[2] , \nOut22_1[1] , \nOut22_1[0] }), .WestIn(
        {\nOut20_1[7] , \nOut20_1[6] , \nOut20_1[5] , \nOut20_1[4] , 
        \nOut20_1[3] , \nOut20_1[2] , \nOut20_1[1] , \nOut20_1[0] }), .Out({
        \nOut21_1[7] , \nOut21_1[6] , \nOut21_1[5] , \nOut21_1[4] , 
        \nOut21_1[3] , \nOut21_1[2] , \nOut21_1[1] , \nOut21_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_931 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut932[7] , \nScanOut932[6] , 
        \nScanOut932[5] , \nScanOut932[4] , \nScanOut932[3] , \nScanOut932[2] , 
        \nScanOut932[1] , \nScanOut932[0] }), .ScanOut({\nScanOut931[7] , 
        \nScanOut931[6] , \nScanOut931[5] , \nScanOut931[4] , \nScanOut931[3] , 
        \nScanOut931[2] , \nScanOut931[1] , \nScanOut931[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_2[7] , \nOut29_2[6] , \nOut29_2[5] , \nOut29_2[4] , 
        \nOut29_2[3] , \nOut29_2[2] , \nOut29_2[1] , \nOut29_2[0] }), 
        .SouthIn({\nOut29_4[7] , \nOut29_4[6] , \nOut29_4[5] , \nOut29_4[4] , 
        \nOut29_4[3] , \nOut29_4[2] , \nOut29_4[1] , \nOut29_4[0] }), .EastIn(
        {\nOut30_3[7] , \nOut30_3[6] , \nOut30_3[5] , \nOut30_3[4] , 
        \nOut30_3[3] , \nOut30_3[2] , \nOut30_3[1] , \nOut30_3[0] }), .WestIn(
        {\nOut28_3[7] , \nOut28_3[6] , \nOut28_3[5] , \nOut28_3[4] , 
        \nOut28_3[3] , \nOut28_3[2] , \nOut28_3[1] , \nOut28_3[0] }), .Out({
        \nOut29_3[7] , \nOut29_3[6] , \nOut29_3[5] , \nOut29_3[4] , 
        \nOut29_3[3] , \nOut29_3[2] , \nOut29_3[1] , \nOut29_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_654 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut655[7] , \nScanOut655[6] , 
        \nScanOut655[5] , \nScanOut655[4] , \nScanOut655[3] , \nScanOut655[2] , 
        \nScanOut655[1] , \nScanOut655[0] }), .ScanOut({\nScanOut654[7] , 
        \nScanOut654[6] , \nScanOut654[5] , \nScanOut654[4] , \nScanOut654[3] , 
        \nScanOut654[2] , \nScanOut654[1] , \nScanOut654[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_13[7] , \nOut20_13[6] , \nOut20_13[5] , \nOut20_13[4] , 
        \nOut20_13[3] , \nOut20_13[2] , \nOut20_13[1] , \nOut20_13[0] }), 
        .SouthIn({\nOut20_15[7] , \nOut20_15[6] , \nOut20_15[5] , 
        \nOut20_15[4] , \nOut20_15[3] , \nOut20_15[2] , \nOut20_15[1] , 
        \nOut20_15[0] }), .EastIn({\nOut21_14[7] , \nOut21_14[6] , 
        \nOut21_14[5] , \nOut21_14[4] , \nOut21_14[3] , \nOut21_14[2] , 
        \nOut21_14[1] , \nOut21_14[0] }), .WestIn({\nOut19_14[7] , 
        \nOut19_14[6] , \nOut19_14[5] , \nOut19_14[4] , \nOut19_14[3] , 
        \nOut19_14[2] , \nOut19_14[1] , \nOut19_14[0] }), .Out({\nOut20_14[7] , 
        \nOut20_14[6] , \nOut20_14[5] , \nOut20_14[4] , \nOut20_14[3] , 
        \nOut20_14[2] , \nOut20_14[1] , \nOut20_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_13 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut14[7] , \nScanOut14[6] , 
        \nScanOut14[5] , \nScanOut14[4] , \nScanOut14[3] , \nScanOut14[2] , 
        \nScanOut14[1] , \nScanOut14[0] }), .ScanOut({\nScanOut13[7] , 
        \nScanOut13[6] , \nScanOut13[5] , \nScanOut13[4] , \nScanOut13[3] , 
        \nScanOut13[2] , \nScanOut13[1] , \nScanOut13[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_13[7] , \nOut0_13[6] , 
        \nOut0_13[5] , \nOut0_13[4] , \nOut0_13[3] , \nOut0_13[2] , 
        \nOut0_13[1] , \nOut0_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_41 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut42[7] , \nScanOut42[6] , 
        \nScanOut42[5] , \nScanOut42[4] , \nScanOut42[3] , \nScanOut42[2] , 
        \nScanOut42[1] , \nScanOut42[0] }), .ScanOut({\nScanOut41[7] , 
        \nScanOut41[6] , \nScanOut41[5] , \nScanOut41[4] , \nScanOut41[3] , 
        \nScanOut41[2] , \nScanOut41[1] , \nScanOut41[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , \nOut1_8[4] , \nOut1_8[3] , 
        \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }), .SouthIn({\nOut1_10[7] , 
        \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , \nOut1_10[3] , 
        \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), .EastIn({\nOut2_9[7] , 
        \nOut2_9[6] , \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , 
        \nOut2_9[1] , \nOut2_9[0] }), .WestIn({\nOut0_9[7] , \nOut0_9[6] , 
        \nOut0_9[5] , \nOut0_9[4] , \nOut0_9[3] , \nOut0_9[2] , \nOut0_9[1] , 
        \nOut0_9[0] }), .Out({\nOut1_9[7] , \nOut1_9[6] , \nOut1_9[5] , 
        \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , \nOut1_9[1] , \nOut1_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_98 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut99[7] , \nScanOut99[6] , 
        \nScanOut99[5] , \nScanOut99[4] , \nScanOut99[3] , \nScanOut99[2] , 
        \nScanOut99[1] , \nScanOut99[0] }), .ScanOut({\nScanOut98[7] , 
        \nScanOut98[6] , \nScanOut98[5] , \nScanOut98[4] , \nScanOut98[3] , 
        \nScanOut98[2] , \nScanOut98[1] , \nScanOut98[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_1[7] , \nOut3_1[6] , \nOut3_1[5] , \nOut3_1[4] , \nOut3_1[3] , 
        \nOut3_1[2] , \nOut3_1[1] , \nOut3_1[0] }), .SouthIn({\nOut3_3[7] , 
        \nOut3_3[6] , \nOut3_3[5] , \nOut3_3[4] , \nOut3_3[3] , \nOut3_3[2] , 
        \nOut3_3[1] , \nOut3_3[0] }), .EastIn({\nOut4_2[7] , \nOut4_2[6] , 
        \nOut4_2[5] , \nOut4_2[4] , \nOut4_2[3] , \nOut4_2[2] , \nOut4_2[1] , 
        \nOut4_2[0] }), .WestIn({\nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , 
        \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }), 
        .Out({\nOut3_2[7] , \nOut3_2[6] , \nOut3_2[5] , \nOut3_2[4] , 
        \nOut3_2[3] , \nOut3_2[2] , \nOut3_2[1] , \nOut3_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_145 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut146[7] , \nScanOut146[6] , 
        \nScanOut146[5] , \nScanOut146[4] , \nScanOut146[3] , \nScanOut146[2] , 
        \nScanOut146[1] , \nScanOut146[0] }), .ScanOut({\nScanOut145[7] , 
        \nScanOut145[6] , \nScanOut145[5] , \nScanOut145[4] , \nScanOut145[3] , 
        \nScanOut145[2] , \nScanOut145[1] , \nScanOut145[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_16[7] , \nOut4_16[6] , \nOut4_16[5] , \nOut4_16[4] , 
        \nOut4_16[3] , \nOut4_16[2] , \nOut4_16[1] , \nOut4_16[0] }), 
        .SouthIn({\nOut4_18[7] , \nOut4_18[6] , \nOut4_18[5] , \nOut4_18[4] , 
        \nOut4_18[3] , \nOut4_18[2] , \nOut4_18[1] , \nOut4_18[0] }), .EastIn(
        {\nOut5_17[7] , \nOut5_17[6] , \nOut5_17[5] , \nOut5_17[4] , 
        \nOut5_17[3] , \nOut5_17[2] , \nOut5_17[1] , \nOut5_17[0] }), .WestIn(
        {\nOut3_17[7] , \nOut3_17[6] , \nOut3_17[5] , \nOut3_17[4] , 
        \nOut3_17[3] , \nOut3_17[2] , \nOut3_17[1] , \nOut3_17[0] }), .Out({
        \nOut4_17[7] , \nOut4_17[6] , \nOut4_17[5] , \nOut4_17[4] , 
        \nOut4_17[3] , \nOut4_17[2] , \nOut4_17[1] , \nOut4_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_275 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut276[7] , \nScanOut276[6] , 
        \nScanOut276[5] , \nScanOut276[4] , \nScanOut276[3] , \nScanOut276[2] , 
        \nScanOut276[1] , \nScanOut276[0] }), .ScanOut({\nScanOut275[7] , 
        \nScanOut275[6] , \nScanOut275[5] , \nScanOut275[4] , \nScanOut275[3] , 
        \nScanOut275[2] , \nScanOut275[1] , \nScanOut275[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_18[7] , \nOut8_18[6] , \nOut8_18[5] , \nOut8_18[4] , 
        \nOut8_18[3] , \nOut8_18[2] , \nOut8_18[1] , \nOut8_18[0] }), 
        .SouthIn({\nOut8_20[7] , \nOut8_20[6] , \nOut8_20[5] , \nOut8_20[4] , 
        \nOut8_20[3] , \nOut8_20[2] , \nOut8_20[1] , \nOut8_20[0] }), .EastIn(
        {\nOut9_19[7] , \nOut9_19[6] , \nOut9_19[5] , \nOut9_19[4] , 
        \nOut9_19[3] , \nOut9_19[2] , \nOut9_19[1] , \nOut9_19[0] }), .WestIn(
        {\nOut7_19[7] , \nOut7_19[6] , \nOut7_19[5] , \nOut7_19[4] , 
        \nOut7_19[3] , \nOut7_19[2] , \nOut7_19[1] , \nOut7_19[0] }), .Out({
        \nOut8_19[7] , \nOut8_19[6] , \nOut8_19[5] , \nOut8_19[4] , 
        \nOut8_19[3] , \nOut8_19[2] , \nOut8_19[1] , \nOut8_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_349 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut350[7] , \nScanOut350[6] , 
        \nScanOut350[5] , \nScanOut350[4] , \nScanOut350[3] , \nScanOut350[2] , 
        \nScanOut350[1] , \nScanOut350[0] }), .ScanOut({\nScanOut349[7] , 
        \nScanOut349[6] , \nScanOut349[5] , \nScanOut349[4] , \nScanOut349[3] , 
        \nScanOut349[2] , \nScanOut349[1] , \nScanOut349[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_28[7] , \nOut10_28[6] , \nOut10_28[5] , \nOut10_28[4] , 
        \nOut10_28[3] , \nOut10_28[2] , \nOut10_28[1] , \nOut10_28[0] }), 
        .SouthIn({\nOut10_30[7] , \nOut10_30[6] , \nOut10_30[5] , 
        \nOut10_30[4] , \nOut10_30[3] , \nOut10_30[2] , \nOut10_30[1] , 
        \nOut10_30[0] }), .EastIn({\nOut11_29[7] , \nOut11_29[6] , 
        \nOut11_29[5] , \nOut11_29[4] , \nOut11_29[3] , \nOut11_29[2] , 
        \nOut11_29[1] , \nOut11_29[0] }), .WestIn({\nOut9_29[7] , 
        \nOut9_29[6] , \nOut9_29[5] , \nOut9_29[4] , \nOut9_29[3] , 
        \nOut9_29[2] , \nOut9_29[1] , \nOut9_29[0] }), .Out({\nOut10_29[7] , 
        \nOut10_29[6] , \nOut10_29[5] , \nOut10_29[4] , \nOut10_29[3] , 
        \nOut10_29[2] , \nOut10_29[1] , \nOut10_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_375 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut376[7] , \nScanOut376[6] , 
        \nScanOut376[5] , \nScanOut376[4] , \nScanOut376[3] , \nScanOut376[2] , 
        \nScanOut376[1] , \nScanOut376[0] }), .ScanOut({\nScanOut375[7] , 
        \nScanOut375[6] , \nScanOut375[5] , \nScanOut375[4] , \nScanOut375[3] , 
        \nScanOut375[2] , \nScanOut375[1] , \nScanOut375[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_22[7] , \nOut11_22[6] , \nOut11_22[5] , \nOut11_22[4] , 
        \nOut11_22[3] , \nOut11_22[2] , \nOut11_22[1] , \nOut11_22[0] }), 
        .SouthIn({\nOut11_24[7] , \nOut11_24[6] , \nOut11_24[5] , 
        \nOut11_24[4] , \nOut11_24[3] , \nOut11_24[2] , \nOut11_24[1] , 
        \nOut11_24[0] }), .EastIn({\nOut12_23[7] , \nOut12_23[6] , 
        \nOut12_23[5] , \nOut12_23[4] , \nOut12_23[3] , \nOut12_23[2] , 
        \nOut12_23[1] , \nOut12_23[0] }), .WestIn({\nOut10_23[7] , 
        \nOut10_23[6] , \nOut10_23[5] , \nOut10_23[4] , \nOut10_23[3] , 
        \nOut10_23[2] , \nOut10_23[1] , \nOut10_23[0] }), .Out({\nOut11_23[7] , 
        \nOut11_23[6] , \nOut11_23[5] , \nOut11_23[4] , \nOut11_23[3] , 
        \nOut11_23[2] , \nOut11_23[1] , \nOut11_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_558 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut559[7] , \nScanOut559[6] , 
        \nScanOut559[5] , \nScanOut559[4] , \nScanOut559[3] , \nScanOut559[2] , 
        \nScanOut559[1] , \nScanOut559[0] }), .ScanOut({\nScanOut558[7] , 
        \nScanOut558[6] , \nScanOut558[5] , \nScanOut558[4] , \nScanOut558[3] , 
        \nScanOut558[2] , \nScanOut558[1] , \nScanOut558[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_13[7] , \nOut17_13[6] , \nOut17_13[5] , \nOut17_13[4] , 
        \nOut17_13[3] , \nOut17_13[2] , \nOut17_13[1] , \nOut17_13[0] }), 
        .SouthIn({\nOut17_15[7] , \nOut17_15[6] , \nOut17_15[5] , 
        \nOut17_15[4] , \nOut17_15[3] , \nOut17_15[2] , \nOut17_15[1] , 
        \nOut17_15[0] }), .EastIn({\nOut18_14[7] , \nOut18_14[6] , 
        \nOut18_14[5] , \nOut18_14[4] , \nOut18_14[3] , \nOut18_14[2] , 
        \nOut18_14[1] , \nOut18_14[0] }), .WestIn({\nOut16_14[7] , 
        \nOut16_14[6] , \nOut16_14[5] , \nOut16_14[4] , \nOut16_14[3] , 
        \nOut16_14[2] , \nOut16_14[1] , \nOut16_14[0] }), .Out({\nOut17_14[7] , 
        \nOut17_14[6] , \nOut17_14[5] , \nOut17_14[4] , \nOut17_14[3] , 
        \nOut17_14[2] , \nOut17_14[1] , \nOut17_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_564 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut565[7] , \nScanOut565[6] , 
        \nScanOut565[5] , \nScanOut565[4] , \nScanOut565[3] , \nScanOut565[2] , 
        \nScanOut565[1] , \nScanOut565[0] }), .ScanOut({\nScanOut564[7] , 
        \nScanOut564[6] , \nScanOut564[5] , \nScanOut564[4] , \nScanOut564[3] , 
        \nScanOut564[2] , \nScanOut564[1] , \nScanOut564[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_19[7] , \nOut17_19[6] , \nOut17_19[5] , \nOut17_19[4] , 
        \nOut17_19[3] , \nOut17_19[2] , \nOut17_19[1] , \nOut17_19[0] }), 
        .SouthIn({\nOut17_21[7] , \nOut17_21[6] , \nOut17_21[5] , 
        \nOut17_21[4] , \nOut17_21[3] , \nOut17_21[2] , \nOut17_21[1] , 
        \nOut17_21[0] }), .EastIn({\nOut18_20[7] , \nOut18_20[6] , 
        \nOut18_20[5] , \nOut18_20[4] , \nOut18_20[3] , \nOut18_20[2] , 
        \nOut18_20[1] , \nOut18_20[0] }), .WestIn({\nOut16_20[7] , 
        \nOut16_20[6] , \nOut16_20[5] , \nOut16_20[4] , \nOut16_20[3] , 
        \nOut16_20[2] , \nOut16_20[1] , \nOut16_20[0] }), .Out({\nOut17_20[7] , 
        \nOut17_20[6] , \nOut17_20[5] , \nOut17_20[4] , \nOut17_20[3] , 
        \nOut17_20[2] , \nOut17_20[1] , \nOut17_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_668 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut669[7] , \nScanOut669[6] , 
        \nScanOut669[5] , \nScanOut669[4] , \nScanOut669[3] , \nScanOut669[2] , 
        \nScanOut669[1] , \nScanOut669[0] }), .ScanOut({\nScanOut668[7] , 
        \nScanOut668[6] , \nScanOut668[5] , \nScanOut668[4] , \nScanOut668[3] , 
        \nScanOut668[2] , \nScanOut668[1] , \nScanOut668[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_27[7] , \nOut20_27[6] , \nOut20_27[5] , \nOut20_27[4] , 
        \nOut20_27[3] , \nOut20_27[2] , \nOut20_27[1] , \nOut20_27[0] }), 
        .SouthIn({\nOut20_29[7] , \nOut20_29[6] , \nOut20_29[5] , 
        \nOut20_29[4] , \nOut20_29[3] , \nOut20_29[2] , \nOut20_29[1] , 
        \nOut20_29[0] }), .EastIn({\nOut21_28[7] , \nOut21_28[6] , 
        \nOut21_28[5] , \nOut21_28[4] , \nOut21_28[3] , \nOut21_28[2] , 
        \nOut21_28[1] , \nOut21_28[0] }), .WestIn({\nOut19_28[7] , 
        \nOut19_28[6] , \nOut19_28[5] , \nOut19_28[4] , \nOut19_28[3] , 
        \nOut19_28[2] , \nOut19_28[1] , \nOut19_28[0] }), .Out({\nOut20_28[7] , 
        \nOut20_28[6] , \nOut20_28[5] , \nOut20_28[4] , \nOut20_28[3] , 
        \nOut20_28[2] , \nOut20_28[1] , \nOut20_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_886 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut887[7] , \nScanOut887[6] , 
        \nScanOut887[5] , \nScanOut887[4] , \nScanOut887[3] , \nScanOut887[2] , 
        \nScanOut887[1] , \nScanOut887[0] }), .ScanOut({\nScanOut886[7] , 
        \nScanOut886[6] , \nScanOut886[5] , \nScanOut886[4] , \nScanOut886[3] , 
        \nScanOut886[2] , \nScanOut886[1] , \nScanOut886[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_21[7] , \nOut27_21[6] , \nOut27_21[5] , \nOut27_21[4] , 
        \nOut27_21[3] , \nOut27_21[2] , \nOut27_21[1] , \nOut27_21[0] }), 
        .SouthIn({\nOut27_23[7] , \nOut27_23[6] , \nOut27_23[5] , 
        \nOut27_23[4] , \nOut27_23[3] , \nOut27_23[2] , \nOut27_23[1] , 
        \nOut27_23[0] }), .EastIn({\nOut28_22[7] , \nOut28_22[6] , 
        \nOut28_22[5] , \nOut28_22[4] , \nOut28_22[3] , \nOut28_22[2] , 
        \nOut28_22[1] , \nOut28_22[0] }), .WestIn({\nOut26_22[7] , 
        \nOut26_22[6] , \nOut26_22[5] , \nOut26_22[4] , \nOut26_22[3] , 
        \nOut26_22[2] , \nOut26_22[1] , \nOut26_22[0] }), .Out({\nOut27_22[7] , 
        \nOut27_22[6] , \nOut27_22[5] , \nOut27_22[4] , \nOut27_22[3] , 
        \nOut27_22[2] , \nOut27_22[1] , \nOut27_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_916 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut917[7] , \nScanOut917[6] , 
        \nScanOut917[5] , \nScanOut917[4] , \nScanOut917[3] , \nScanOut917[2] , 
        \nScanOut917[1] , \nScanOut917[0] }), .ScanOut({\nScanOut916[7] , 
        \nScanOut916[6] , \nScanOut916[5] , \nScanOut916[4] , \nScanOut916[3] , 
        \nScanOut916[2] , \nScanOut916[1] , \nScanOut916[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_19[7] , \nOut28_19[6] , \nOut28_19[5] , \nOut28_19[4] , 
        \nOut28_19[3] , \nOut28_19[2] , \nOut28_19[1] , \nOut28_19[0] }), 
        .SouthIn({\nOut28_21[7] , \nOut28_21[6] , \nOut28_21[5] , 
        \nOut28_21[4] , \nOut28_21[3] , \nOut28_21[2] , \nOut28_21[1] , 
        \nOut28_21[0] }), .EastIn({\nOut29_20[7] , \nOut29_20[6] , 
        \nOut29_20[5] , \nOut29_20[4] , \nOut29_20[3] , \nOut29_20[2] , 
        \nOut29_20[1] , \nOut29_20[0] }), .WestIn({\nOut27_20[7] , 
        \nOut27_20[6] , \nOut27_20[5] , \nOut27_20[4] , \nOut27_20[3] , 
        \nOut27_20[2] , \nOut27_20[1] , \nOut27_20[0] }), .Out({\nOut28_20[7] , 
        \nOut28_20[6] , \nOut28_20[5] , \nOut28_20[4] , \nOut28_20[3] , 
        \nOut28_20[2] , \nOut28_20[1] , \nOut28_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_464 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut465[7] , \nScanOut465[6] , 
        \nScanOut465[5] , \nScanOut465[4] , \nScanOut465[3] , \nScanOut465[2] , 
        \nScanOut465[1] , \nScanOut465[0] }), .ScanOut({\nScanOut464[7] , 
        \nScanOut464[6] , \nScanOut464[5] , \nScanOut464[4] , \nScanOut464[3] , 
        \nScanOut464[2] , \nScanOut464[1] , \nScanOut464[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_15[7] , \nOut14_15[6] , \nOut14_15[5] , \nOut14_15[4] , 
        \nOut14_15[3] , \nOut14_15[2] , \nOut14_15[1] , \nOut14_15[0] }), 
        .SouthIn({\nOut14_17[7] , \nOut14_17[6] , \nOut14_17[5] , 
        \nOut14_17[4] , \nOut14_17[3] , \nOut14_17[2] , \nOut14_17[1] , 
        \nOut14_17[0] }), .EastIn({\nOut15_16[7] , \nOut15_16[6] , 
        \nOut15_16[5] , \nOut15_16[4] , \nOut15_16[3] , \nOut15_16[2] , 
        \nOut15_16[1] , \nOut15_16[0] }), .WestIn({\nOut13_16[7] , 
        \nOut13_16[6] , \nOut13_16[5] , \nOut13_16[4] , \nOut13_16[3] , 
        \nOut13_16[2] , \nOut13_16[1] , \nOut13_16[0] }), .Out({\nOut14_16[7] , 
        \nOut14_16[6] , \nOut14_16[5] , \nOut14_16[4] , \nOut14_16[3] , 
        \nOut14_16[2] , \nOut14_16[1] , \nOut14_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_754 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut755[7] , \nScanOut755[6] , 
        \nScanOut755[5] , \nScanOut755[4] , \nScanOut755[3] , \nScanOut755[2] , 
        \nScanOut755[1] , \nScanOut755[0] }), .ScanOut({\nScanOut754[7] , 
        \nScanOut754[6] , \nScanOut754[5] , \nScanOut754[4] , \nScanOut754[3] , 
        \nScanOut754[2] , \nScanOut754[1] , \nScanOut754[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_17[7] , \nOut23_17[6] , \nOut23_17[5] , \nOut23_17[4] , 
        \nOut23_17[3] , \nOut23_17[2] , \nOut23_17[1] , \nOut23_17[0] }), 
        .SouthIn({\nOut23_19[7] , \nOut23_19[6] , \nOut23_19[5] , 
        \nOut23_19[4] , \nOut23_19[3] , \nOut23_19[2] , \nOut23_19[1] , 
        \nOut23_19[0] }), .EastIn({\nOut24_18[7] , \nOut24_18[6] , 
        \nOut24_18[5] , \nOut24_18[4] , \nOut24_18[3] , \nOut24_18[2] , 
        \nOut24_18[1] , \nOut24_18[0] }), .WestIn({\nOut22_18[7] , 
        \nOut22_18[6] , \nOut22_18[5] , \nOut22_18[4] , \nOut22_18[3] , 
        \nOut22_18[2] , \nOut22_18[1] , \nOut22_18[0] }), .Out({\nOut23_18[7] , 
        \nOut23_18[6] , \nOut23_18[5] , \nOut23_18[4] , \nOut23_18[3] , 
        \nOut23_18[2] , \nOut23_18[1] , \nOut23_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_816 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut817[7] , \nScanOut817[6] , 
        \nScanOut817[5] , \nScanOut817[4] , \nScanOut817[3] , \nScanOut817[2] , 
        \nScanOut817[1] , \nScanOut817[0] }), .ScanOut({\nScanOut816[7] , 
        \nScanOut816[6] , \nScanOut816[5] , \nScanOut816[4] , \nScanOut816[3] , 
        \nScanOut816[2] , \nScanOut816[1] , \nScanOut816[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_15[7] , \nOut25_15[6] , \nOut25_15[5] , \nOut25_15[4] , 
        \nOut25_15[3] , \nOut25_15[2] , \nOut25_15[1] , \nOut25_15[0] }), 
        .SouthIn({\nOut25_17[7] , \nOut25_17[6] , \nOut25_17[5] , 
        \nOut25_17[4] , \nOut25_17[3] , \nOut25_17[2] , \nOut25_17[1] , 
        \nOut25_17[0] }), .EastIn({\nOut26_16[7] , \nOut26_16[6] , 
        \nOut26_16[5] , \nOut26_16[4] , \nOut26_16[3] , \nOut26_16[2] , 
        \nOut26_16[1] , \nOut26_16[0] }), .WestIn({\nOut24_16[7] , 
        \nOut24_16[6] , \nOut24_16[5] , \nOut24_16[4] , \nOut24_16[3] , 
        \nOut24_16[2] , \nOut24_16[1] , \nOut24_16[0] }), .Out({\nOut25_16[7] , 
        \nOut25_16[6] , \nOut25_16[5] , \nOut25_16[4] , \nOut25_16[3] , 
        \nOut25_16[2] , \nOut25_16[1] , \nOut25_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_986 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut987[7] , \nScanOut987[6] , 
        \nScanOut987[5] , \nScanOut987[4] , \nScanOut987[3] , \nScanOut987[2] , 
        \nScanOut987[1] , \nScanOut987[0] }), .ScanOut({\nScanOut986[7] , 
        \nScanOut986[6] , \nScanOut986[5] , \nScanOut986[4] , \nScanOut986[3] , 
        \nScanOut986[2] , \nScanOut986[1] , \nScanOut986[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_25[7] , \nOut30_25[6] , \nOut30_25[5] , \nOut30_25[4] , 
        \nOut30_25[3] , \nOut30_25[2] , \nOut30_25[1] , \nOut30_25[0] }), 
        .SouthIn({\nOut30_27[7] , \nOut30_27[6] , \nOut30_27[5] , 
        \nOut30_27[4] , \nOut30_27[3] , \nOut30_27[2] , \nOut30_27[1] , 
        \nOut30_27[0] }), .EastIn({\nOut31_26[7] , \nOut31_26[6] , 
        \nOut31_26[5] , \nOut31_26[4] , \nOut31_26[3] , \nOut31_26[2] , 
        \nOut31_26[1] , \nOut31_26[0] }), .WestIn({\nOut29_26[7] , 
        \nOut29_26[6] , \nOut29_26[5] , \nOut29_26[4] , \nOut29_26[3] , 
        \nOut29_26[2] , \nOut29_26[1] , \nOut29_26[0] }), .Out({\nOut30_26[7] , 
        \nOut30_26[6] , \nOut30_26[5] , \nOut30_26[4] , \nOut30_26[3] , 
        \nOut30_26[2] , \nOut30_26[1] , \nOut30_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_162 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut163[7] , \nScanOut163[6] , 
        \nScanOut163[5] , \nScanOut163[4] , \nScanOut163[3] , \nScanOut163[2] , 
        \nScanOut163[1] , \nScanOut163[0] }), .ScanOut({\nScanOut162[7] , 
        \nScanOut162[6] , \nScanOut162[5] , \nScanOut162[4] , \nScanOut162[3] , 
        \nScanOut162[2] , \nScanOut162[1] , \nScanOut162[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_1[7] , \nOut5_1[6] , \nOut5_1[5] , \nOut5_1[4] , \nOut5_1[3] , 
        \nOut5_1[2] , \nOut5_1[1] , \nOut5_1[0] }), .SouthIn({\nOut5_3[7] , 
        \nOut5_3[6] , \nOut5_3[5] , \nOut5_3[4] , \nOut5_3[3] , \nOut5_3[2] , 
        \nOut5_3[1] , \nOut5_3[0] }), .EastIn({\nOut6_2[7] , \nOut6_2[6] , 
        \nOut6_2[5] , \nOut6_2[4] , \nOut6_2[3] , \nOut6_2[2] , \nOut6_2[1] , 
        \nOut6_2[0] }), .WestIn({\nOut4_2[7] , \nOut4_2[6] , \nOut4_2[5] , 
        \nOut4_2[4] , \nOut4_2[3] , \nOut4_2[2] , \nOut4_2[1] , \nOut4_2[0] }), 
        .Out({\nOut5_2[7] , \nOut5_2[6] , \nOut5_2[5] , \nOut5_2[4] , 
        \nOut5_2[3] , \nOut5_2[2] , \nOut5_2[1] , \nOut5_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_252 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut253[7] , \nScanOut253[6] , 
        \nScanOut253[5] , \nScanOut253[4] , \nScanOut253[3] , \nScanOut253[2] , 
        \nScanOut253[1] , \nScanOut253[0] }), .ScanOut({\nScanOut252[7] , 
        \nScanOut252[6] , \nScanOut252[5] , \nScanOut252[4] , \nScanOut252[3] , 
        \nScanOut252[2] , \nScanOut252[1] , \nScanOut252[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_27[7] , \nOut7_27[6] , \nOut7_27[5] , \nOut7_27[4] , 
        \nOut7_27[3] , \nOut7_27[2] , \nOut7_27[1] , \nOut7_27[0] }), 
        .SouthIn({\nOut7_29[7] , \nOut7_29[6] , \nOut7_29[5] , \nOut7_29[4] , 
        \nOut7_29[3] , \nOut7_29[2] , \nOut7_29[1] , \nOut7_29[0] }), .EastIn(
        {\nOut8_28[7] , \nOut8_28[6] , \nOut8_28[5] , \nOut8_28[4] , 
        \nOut8_28[3] , \nOut8_28[2] , \nOut8_28[1] , \nOut8_28[0] }), .WestIn(
        {\nOut6_28[7] , \nOut6_28[6] , \nOut6_28[5] , \nOut6_28[4] , 
        \nOut6_28[3] , \nOut6_28[2] , \nOut6_28[1] , \nOut6_28[0] }), .Out({
        \nOut7_28[7] , \nOut7_28[6] , \nOut7_28[5] , \nOut7_28[4] , 
        \nOut7_28[3] , \nOut7_28[2] , \nOut7_28[1] , \nOut7_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_773 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut774[7] , \nScanOut774[6] , 
        \nScanOut774[5] , \nScanOut774[4] , \nScanOut774[3] , \nScanOut774[2] , 
        \nScanOut774[1] , \nScanOut774[0] }), .ScanOut({\nScanOut773[7] , 
        \nScanOut773[6] , \nScanOut773[5] , \nScanOut773[4] , \nScanOut773[3] , 
        \nScanOut773[2] , \nScanOut773[1] , \nScanOut773[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_4[7] , \nOut24_4[6] , \nOut24_4[5] , \nOut24_4[4] , 
        \nOut24_4[3] , \nOut24_4[2] , \nOut24_4[1] , \nOut24_4[0] }), 
        .SouthIn({\nOut24_6[7] , \nOut24_6[6] , \nOut24_6[5] , \nOut24_6[4] , 
        \nOut24_6[3] , \nOut24_6[2] , \nOut24_6[1] , \nOut24_6[0] }), .EastIn(
        {\nOut25_5[7] , \nOut25_5[6] , \nOut25_5[5] , \nOut25_5[4] , 
        \nOut25_5[3] , \nOut25_5[2] , \nOut25_5[1] , \nOut25_5[0] }), .WestIn(
        {\nOut23_5[7] , \nOut23_5[6] , \nOut23_5[5] , \nOut23_5[4] , 
        \nOut23_5[3] , \nOut23_5[2] , \nOut23_5[1] , \nOut23_5[0] }), .Out({
        \nOut24_5[7] , \nOut24_5[6] , \nOut24_5[5] , \nOut24_5[4] , 
        \nOut24_5[3] , \nOut24_5[2] , \nOut24_5[1] , \nOut24_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_443 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut444[7] , \nScanOut444[6] , 
        \nScanOut444[5] , \nScanOut444[4] , \nScanOut444[3] , \nScanOut444[2] , 
        \nScanOut444[1] , \nScanOut444[0] }), .ScanOut({\nScanOut443[7] , 
        \nScanOut443[6] , \nScanOut443[5] , \nScanOut443[4] , \nScanOut443[3] , 
        \nScanOut443[2] , \nScanOut443[1] , \nScanOut443[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_26[7] , \nOut13_26[6] , \nOut13_26[5] , \nOut13_26[4] , 
        \nOut13_26[3] , \nOut13_26[2] , \nOut13_26[1] , \nOut13_26[0] }), 
        .SouthIn({\nOut13_28[7] , \nOut13_28[6] , \nOut13_28[5] , 
        \nOut13_28[4] , \nOut13_28[3] , \nOut13_28[2] , \nOut13_28[1] , 
        \nOut13_28[0] }), .EastIn({\nOut14_27[7] , \nOut14_27[6] , 
        \nOut14_27[5] , \nOut14_27[4] , \nOut14_27[3] , \nOut14_27[2] , 
        \nOut14_27[1] , \nOut14_27[0] }), .WestIn({\nOut12_27[7] , 
        \nOut12_27[6] , \nOut12_27[5] , \nOut12_27[4] , \nOut12_27[3] , 
        \nOut12_27[2] , \nOut12_27[1] , \nOut12_27[0] }), .Out({\nOut13_27[7] , 
        \nOut13_27[6] , \nOut13_27[5] , \nOut13_27[4] , \nOut13_27[3] , 
        \nOut13_27[2] , \nOut13_27[1] , \nOut13_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_831 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut832[7] , \nScanOut832[6] , 
        \nScanOut832[5] , \nScanOut832[4] , \nScanOut832[3] , \nScanOut832[2] , 
        \nScanOut832[1] , \nScanOut832[0] }), .ScanOut({\nScanOut831[7] , 
        \nScanOut831[6] , \nScanOut831[5] , \nScanOut831[4] , \nScanOut831[3] , 
        \nScanOut831[2] , \nScanOut831[1] , \nScanOut831[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut25_31[7] , \nOut25_31[6] , 
        \nOut25_31[5] , \nOut25_31[4] , \nOut25_31[3] , \nOut25_31[2] , 
        \nOut25_31[1] , \nOut25_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_878 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut879[7] , \nScanOut879[6] , 
        \nScanOut879[5] , \nScanOut879[4] , \nScanOut879[3] , \nScanOut879[2] , 
        \nScanOut879[1] , \nScanOut879[0] }), .ScanOut({\nScanOut878[7] , 
        \nScanOut878[6] , \nScanOut878[5] , \nScanOut878[4] , \nScanOut878[3] , 
        \nScanOut878[2] , \nScanOut878[1] , \nScanOut878[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_13[7] , \nOut27_13[6] , \nOut27_13[5] , \nOut27_13[4] , 
        \nOut27_13[3] , \nOut27_13[2] , \nOut27_13[1] , \nOut27_13[0] }), 
        .SouthIn({\nOut27_15[7] , \nOut27_15[6] , \nOut27_15[5] , 
        \nOut27_15[4] , \nOut27_15[3] , \nOut27_15[2] , \nOut27_15[1] , 
        \nOut27_15[0] }), .EastIn({\nOut28_14[7] , \nOut28_14[6] , 
        \nOut28_14[5] , \nOut28_14[4] , \nOut28_14[3] , \nOut28_14[2] , 
        \nOut28_14[1] , \nOut28_14[0] }), .WestIn({\nOut26_14[7] , 
        \nOut26_14[6] , \nOut26_14[5] , \nOut26_14[4] , \nOut26_14[3] , 
        \nOut26_14[2] , \nOut26_14[1] , \nOut26_14[0] }), .Out({\nOut27_14[7] , 
        \nOut27_14[6] , \nOut27_14[5] , \nOut27_14[4] , \nOut27_14[3] , 
        \nOut27_14[2] , \nOut27_14[1] , \nOut27_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_14 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut15[7] , \nScanOut15[6] , 
        \nScanOut15[5] , \nScanOut15[4] , \nScanOut15[3] , \nScanOut15[2] , 
        \nScanOut15[1] , \nScanOut15[0] }), .ScanOut({\nScanOut14[7] , 
        \nScanOut14[6] , \nScanOut14[5] , \nScanOut14[4] , \nScanOut14[3] , 
        \nScanOut14[2] , \nScanOut14[1] , \nScanOut14[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_14[7] , \nOut0_14[6] , 
        \nOut0_14[5] , \nOut0_14[4] , \nOut0_14[3] , \nOut0_14[2] , 
        \nOut0_14[1] , \nOut0_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_33 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut34[7] , \nScanOut34[6] , 
        \nScanOut34[5] , \nScanOut34[4] , \nScanOut34[3] , \nScanOut34[2] , 
        \nScanOut34[1] , \nScanOut34[0] }), .ScanOut({\nScanOut33[7] , 
        \nScanOut33[6] , \nScanOut33[5] , \nScanOut33[4] , \nScanOut33[3] , 
        \nScanOut33[2] , \nScanOut33[1] , \nScanOut33[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_0[7] , \nOut1_0[6] , \nOut1_0[5] , \nOut1_0[4] , \nOut1_0[3] , 
        \nOut1_0[2] , \nOut1_0[1] , \nOut1_0[0] }), .SouthIn({\nOut1_2[7] , 
        \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , 
        \nOut1_2[1] , \nOut1_2[0] }), .EastIn({\nOut2_1[7] , \nOut2_1[6] , 
        \nOut2_1[5] , \nOut2_1[4] , \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , 
        \nOut2_1[0] }), .WestIn({\nOut0_1[7] , \nOut0_1[6] , \nOut0_1[5] , 
        \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , \nOut0_1[0] }), 
        .Out({\nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , \nOut1_1[4] , 
        \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_34 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut35[7] , \nScanOut35[6] , 
        \nScanOut35[5] , \nScanOut35[4] , \nScanOut35[3] , \nScanOut35[2] , 
        \nScanOut35[1] , \nScanOut35[0] }), .ScanOut({\nScanOut34[7] , 
        \nScanOut34[6] , \nScanOut34[5] , \nScanOut34[4] , \nScanOut34[3] , 
        \nScanOut34[2] , \nScanOut34[1] , \nScanOut34[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , \nOut1_1[4] , \nOut1_1[3] , 
        \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), .SouthIn({\nOut1_3[7] , 
        \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , 
        \nOut1_3[1] , \nOut1_3[0] }), .EastIn({\nOut2_2[7] , \nOut2_2[6] , 
        \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , 
        \nOut2_2[0] }), .WestIn({\nOut0_2[7] , \nOut0_2[6] , \nOut0_2[5] , 
        \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , \nOut0_2[0] }), 
        .Out({\nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , 
        \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_187 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut188[7] , \nScanOut188[6] , 
        \nScanOut188[5] , \nScanOut188[4] , \nScanOut188[3] , \nScanOut188[2] , 
        \nScanOut188[1] , \nScanOut188[0] }), .ScanOut({\nScanOut187[7] , 
        \nScanOut187[6] , \nScanOut187[5] , \nScanOut187[4] , \nScanOut187[3] , 
        \nScanOut187[2] , \nScanOut187[1] , \nScanOut187[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_26[7] , \nOut5_26[6] , \nOut5_26[5] , \nOut5_26[4] , 
        \nOut5_26[3] , \nOut5_26[2] , \nOut5_26[1] , \nOut5_26[0] }), 
        .SouthIn({\nOut5_28[7] , \nOut5_28[6] , \nOut5_28[5] , \nOut5_28[4] , 
        \nOut5_28[3] , \nOut5_28[2] , \nOut5_28[1] , \nOut5_28[0] }), .EastIn(
        {\nOut6_27[7] , \nOut6_27[6] , \nOut6_27[5] , \nOut6_27[4] , 
        \nOut6_27[3] , \nOut6_27[2] , \nOut6_27[1] , \nOut6_27[0] }), .WestIn(
        {\nOut4_27[7] , \nOut4_27[6] , \nOut4_27[5] , \nOut4_27[4] , 
        \nOut4_27[3] , \nOut4_27[2] , \nOut4_27[1] , \nOut4_27[0] }), .Out({
        \nOut5_27[7] , \nOut5_27[6] , \nOut5_27[5] , \nOut5_27[4] , 
        \nOut5_27[3] , \nOut5_27[2] , \nOut5_27[1] , \nOut5_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_606 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut607[7] , \nScanOut607[6] , 
        \nScanOut607[5] , \nScanOut607[4] , \nScanOut607[3] , \nScanOut607[2] , 
        \nScanOut607[1] , \nScanOut607[0] }), .ScanOut({\nScanOut606[7] , 
        \nScanOut606[6] , \nScanOut606[5] , \nScanOut606[4] , \nScanOut606[3] , 
        \nScanOut606[2] , \nScanOut606[1] , \nScanOut606[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_29[7] , \nOut18_29[6] , \nOut18_29[5] , \nOut18_29[4] , 
        \nOut18_29[3] , \nOut18_29[2] , \nOut18_29[1] , \nOut18_29[0] }), 
        .SouthIn({\nOut18_31[7] , \nOut18_31[6] , \nOut18_31[5] , 
        \nOut18_31[4] , \nOut18_31[3] , \nOut18_31[2] , \nOut18_31[1] , 
        \nOut18_31[0] }), .EastIn({\nOut19_30[7] , \nOut19_30[6] , 
        \nOut19_30[5] , \nOut19_30[4] , \nOut19_30[3] , \nOut19_30[2] , 
        \nOut19_30[1] , \nOut19_30[0] }), .WestIn({\nOut17_30[7] , 
        \nOut17_30[6] , \nOut17_30[5] , \nOut17_30[4] , \nOut17_30[3] , 
        \nOut17_30[2] , \nOut17_30[1] , \nOut17_30[0] }), .Out({\nOut18_30[7] , 
        \nOut18_30[6] , \nOut18_30[5] , \nOut18_30[4] , \nOut18_30[3] , 
        \nOut18_30[2] , \nOut18_30[1] , \nOut18_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_796 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut797[7] , \nScanOut797[6] , 
        \nScanOut797[5] , \nScanOut797[4] , \nScanOut797[3] , \nScanOut797[2] , 
        \nScanOut797[1] , \nScanOut797[0] }), .ScanOut({\nScanOut796[7] , 
        \nScanOut796[6] , \nScanOut796[5] , \nScanOut796[4] , \nScanOut796[3] , 
        \nScanOut796[2] , \nScanOut796[1] , \nScanOut796[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_27[7] , \nOut24_27[6] , \nOut24_27[5] , \nOut24_27[4] , 
        \nOut24_27[3] , \nOut24_27[2] , \nOut24_27[1] , \nOut24_27[0] }), 
        .SouthIn({\nOut24_29[7] , \nOut24_29[6] , \nOut24_29[5] , 
        \nOut24_29[4] , \nOut24_29[3] , \nOut24_29[2] , \nOut24_29[1] , 
        \nOut24_29[0] }), .EastIn({\nOut25_28[7] , \nOut25_28[6] , 
        \nOut25_28[5] , \nOut25_28[4] , \nOut25_28[3] , \nOut25_28[2] , 
        \nOut25_28[1] , \nOut25_28[0] }), .WestIn({\nOut23_28[7] , 
        \nOut23_28[6] , \nOut23_28[5] , \nOut23_28[4] , \nOut23_28[3] , 
        \nOut23_28[2] , \nOut23_28[1] , \nOut23_28[0] }), .Out({\nOut24_28[7] , 
        \nOut24_28[6] , \nOut24_28[5] , \nOut24_28[4] , \nOut24_28[3] , 
        \nOut24_28[2] , \nOut24_28[1] , \nOut24_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_290 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut291[7] , \nScanOut291[6] , 
        \nScanOut291[5] , \nScanOut291[4] , \nScanOut291[3] , \nScanOut291[2] , 
        \nScanOut291[1] , \nScanOut291[0] }), .ScanOut({\nScanOut290[7] , 
        \nScanOut290[6] , \nScanOut290[5] , \nScanOut290[4] , \nScanOut290[3] , 
        \nScanOut290[2] , \nScanOut290[1] , \nScanOut290[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_1[7] , \nOut9_1[6] , \nOut9_1[5] , \nOut9_1[4] , \nOut9_1[3] , 
        \nOut9_1[2] , \nOut9_1[1] , \nOut9_1[0] }), .SouthIn({\nOut9_3[7] , 
        \nOut9_3[6] , \nOut9_3[5] , \nOut9_3[4] , \nOut9_3[3] , \nOut9_3[2] , 
        \nOut9_3[1] , \nOut9_3[0] }), .EastIn({\nOut10_2[7] , \nOut10_2[6] , 
        \nOut10_2[5] , \nOut10_2[4] , \nOut10_2[3] , \nOut10_2[2] , 
        \nOut10_2[1] , \nOut10_2[0] }), .WestIn({\nOut8_2[7] , \nOut8_2[6] , 
        \nOut8_2[5] , \nOut8_2[4] , \nOut8_2[3] , \nOut8_2[2] , \nOut8_2[1] , 
        \nOut8_2[0] }), .Out({\nOut9_2[7] , \nOut9_2[6] , \nOut9_2[5] , 
        \nOut9_2[4] , \nOut9_2[3] , \nOut9_2[2] , \nOut9_2[1] , \nOut9_2[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_327 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut328[7] , \nScanOut328[6] , 
        \nScanOut328[5] , \nScanOut328[4] , \nScanOut328[3] , \nScanOut328[2] , 
        \nScanOut328[1] , \nScanOut328[0] }), .ScanOut({\nScanOut327[7] , 
        \nScanOut327[6] , \nScanOut327[5] , \nScanOut327[4] , \nScanOut327[3] , 
        \nScanOut327[2] , \nScanOut327[1] , \nScanOut327[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_6[7] , \nOut10_6[6] , \nOut10_6[5] , \nOut10_6[4] , 
        \nOut10_6[3] , \nOut10_6[2] , \nOut10_6[1] , \nOut10_6[0] }), 
        .SouthIn({\nOut10_8[7] , \nOut10_8[6] , \nOut10_8[5] , \nOut10_8[4] , 
        \nOut10_8[3] , \nOut10_8[2] , \nOut10_8[1] , \nOut10_8[0] }), .EastIn(
        {\nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }), .WestIn(
        {\nOut9_7[7] , \nOut9_7[6] , \nOut9_7[5] , \nOut9_7[4] , \nOut9_7[3] , 
        \nOut9_7[2] , \nOut9_7[1] , \nOut9_7[0] }), .Out({\nOut10_7[7] , 
        \nOut10_7[6] , \nOut10_7[5] , \nOut10_7[4] , \nOut10_7[3] , 
        \nOut10_7[2] , \nOut10_7[1] , \nOut10_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_536 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut537[7] , \nScanOut537[6] , 
        \nScanOut537[5] , \nScanOut537[4] , \nScanOut537[3] , \nScanOut537[2] , 
        \nScanOut537[1] , \nScanOut537[0] }), .ScanOut({\nScanOut536[7] , 
        \nScanOut536[6] , \nScanOut536[5] , \nScanOut536[4] , \nScanOut536[3] , 
        \nScanOut536[2] , \nScanOut536[1] , \nScanOut536[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_23[7] , \nOut16_23[6] , \nOut16_23[5] , \nOut16_23[4] , 
        \nOut16_23[3] , \nOut16_23[2] , \nOut16_23[1] , \nOut16_23[0] }), 
        .SouthIn({\nOut16_25[7] , \nOut16_25[6] , \nOut16_25[5] , 
        \nOut16_25[4] , \nOut16_25[3] , \nOut16_25[2] , \nOut16_25[1] , 
        \nOut16_25[0] }), .EastIn({\nOut17_24[7] , \nOut17_24[6] , 
        \nOut17_24[5] , \nOut17_24[4] , \nOut17_24[3] , \nOut17_24[2] , 
        \nOut17_24[1] , \nOut17_24[0] }), .WestIn({\nOut15_24[7] , 
        \nOut15_24[6] , \nOut15_24[5] , \nOut15_24[4] , \nOut15_24[3] , 
        \nOut15_24[2] , \nOut15_24[1] , \nOut15_24[0] }), .Out({\nOut16_24[7] , 
        \nOut16_24[6] , \nOut16_24[5] , \nOut16_24[4] , \nOut16_24[3] , 
        \nOut16_24[2] , \nOut16_24[1] , \nOut16_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_944 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut945[7] , \nScanOut945[6] , 
        \nScanOut945[5] , \nScanOut945[4] , \nScanOut945[3] , \nScanOut945[2] , 
        \nScanOut945[1] , \nScanOut945[0] }), .ScanOut({\nScanOut944[7] , 
        \nScanOut944[6] , \nScanOut944[5] , \nScanOut944[4] , \nScanOut944[3] , 
        \nScanOut944[2] , \nScanOut944[1] , \nScanOut944[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_15[7] , \nOut29_15[6] , \nOut29_15[5] , \nOut29_15[4] , 
        \nOut29_15[3] , \nOut29_15[2] , \nOut29_15[1] , \nOut29_15[0] }), 
        .SouthIn({\nOut29_17[7] , \nOut29_17[6] , \nOut29_17[5] , 
        \nOut29_17[4] , \nOut29_17[3] , \nOut29_17[2] , \nOut29_17[1] , 
        \nOut29_17[0] }), .EastIn({\nOut30_16[7] , \nOut30_16[6] , 
        \nOut30_16[5] , \nOut30_16[4] , \nOut30_16[3] , \nOut30_16[2] , 
        \nOut30_16[1] , \nOut30_16[0] }), .WestIn({\nOut28_16[7] , 
        \nOut28_16[6] , \nOut28_16[5] , \nOut28_16[4] , \nOut28_16[3] , 
        \nOut28_16[2] , \nOut28_16[1] , \nOut28_16[0] }), .Out({\nOut29_16[7] , 
        \nOut29_16[6] , \nOut29_16[5] , \nOut29_16[4] , \nOut29_16[3] , 
        \nOut29_16[2] , \nOut29_16[1] , \nOut29_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_300 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut301[7] , \nScanOut301[6] , 
        \nScanOut301[5] , \nScanOut301[4] , \nScanOut301[3] , \nScanOut301[2] , 
        \nScanOut301[1] , \nScanOut301[0] }), .ScanOut({\nScanOut300[7] , 
        \nScanOut300[6] , \nScanOut300[5] , \nScanOut300[4] , \nScanOut300[3] , 
        \nScanOut300[2] , \nScanOut300[1] , \nScanOut300[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_11[7] , \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , 
        \nOut9_11[3] , \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }), 
        .SouthIn({\nOut9_13[7] , \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , 
        \nOut9_13[3] , \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }), .EastIn(
        {\nOut10_12[7] , \nOut10_12[6] , \nOut10_12[5] , \nOut10_12[4] , 
        \nOut10_12[3] , \nOut10_12[2] , \nOut10_12[1] , \nOut10_12[0] }), 
        .WestIn({\nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }), .Out({
        \nOut9_12[7] , \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , 
        \nOut9_12[3] , \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_511 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut512[7] , \nScanOut512[6] , 
        \nScanOut512[5] , \nScanOut512[4] , \nScanOut512[3] , \nScanOut512[2] , 
        \nScanOut512[1] , \nScanOut512[0] }), .ScanOut({\nScanOut511[7] , 
        \nScanOut511[6] , \nScanOut511[5] , \nScanOut511[4] , \nScanOut511[3] , 
        \nScanOut511[2] , \nScanOut511[1] , \nScanOut511[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_31[7] , \nOut15_31[6] , 
        \nOut15_31[5] , \nOut15_31[4] , \nOut15_31[3] , \nOut15_31[2] , 
        \nOut15_31[1] , \nOut15_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_481 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut482[7] , \nScanOut482[6] , 
        \nScanOut482[5] , \nScanOut482[4] , \nScanOut482[3] , \nScanOut482[2] , 
        \nScanOut482[1] , \nScanOut482[0] }), .ScanOut({\nScanOut481[7] , 
        \nScanOut481[6] , \nScanOut481[5] , \nScanOut481[4] , \nScanOut481[3] , 
        \nScanOut481[2] , \nScanOut481[1] , \nScanOut481[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_0[7] , \nOut15_0[6] , \nOut15_0[5] , \nOut15_0[4] , 
        \nOut15_0[3] , \nOut15_0[2] , \nOut15_0[1] , \nOut15_0[0] }), 
        .SouthIn({\nOut15_2[7] , \nOut15_2[6] , \nOut15_2[5] , \nOut15_2[4] , 
        \nOut15_2[3] , \nOut15_2[2] , \nOut15_2[1] , \nOut15_2[0] }), .EastIn(
        {\nOut16_1[7] , \nOut16_1[6] , \nOut16_1[5] , \nOut16_1[4] , 
        \nOut16_1[3] , \nOut16_1[2] , \nOut16_1[1] , \nOut16_1[0] }), .WestIn(
        {\nOut14_1[7] , \nOut14_1[6] , \nOut14_1[5] , \nOut14_1[4] , 
        \nOut14_1[3] , \nOut14_1[2] , \nOut14_1[1] , \nOut14_1[0] }), .Out({
        \nOut15_1[7] , \nOut15_1[6] , \nOut15_1[5] , \nOut15_1[4] , 
        \nOut15_1[3] , \nOut15_1[2] , \nOut15_1[1] , \nOut15_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_963 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut964[7] , \nScanOut964[6] , 
        \nScanOut964[5] , \nScanOut964[4] , \nScanOut964[3] , \nScanOut964[2] , 
        \nScanOut964[1] , \nScanOut964[0] }), .ScanOut({\nScanOut963[7] , 
        \nScanOut963[6] , \nScanOut963[5] , \nScanOut963[4] , \nScanOut963[3] , 
        \nScanOut963[2] , \nScanOut963[1] , \nScanOut963[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_2[7] , \nOut30_2[6] , \nOut30_2[5] , \nOut30_2[4] , 
        \nOut30_2[3] , \nOut30_2[2] , \nOut30_2[1] , \nOut30_2[0] }), 
        .SouthIn({\nOut30_4[7] , \nOut30_4[6] , \nOut30_4[5] , \nOut30_4[4] , 
        \nOut30_4[3] , \nOut30_4[2] , \nOut30_4[1] , \nOut30_4[0] }), .EastIn(
        {\nOut31_3[7] , \nOut31_3[6] , \nOut31_3[5] , \nOut31_3[4] , 
        \nOut31_3[3] , \nOut31_3[2] , \nOut31_3[1] , \nOut31_3[0] }), .WestIn(
        {\nOut29_3[7] , \nOut29_3[6] , \nOut29_3[5] , \nOut29_3[4] , 
        \nOut29_3[3] , \nOut29_3[2] , \nOut29_3[1] , \nOut29_3[0] }), .Out({
        \nOut30_3[7] , \nOut30_3[6] , \nOut30_3[5] , \nOut30_3[4] , 
        \nOut30_3[3] , \nOut30_3[2] , \nOut30_3[1] , \nOut30_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_621 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut622[7] , \nScanOut622[6] , 
        \nScanOut622[5] , \nScanOut622[4] , \nScanOut622[3] , \nScanOut622[2] , 
        \nScanOut622[1] , \nScanOut622[0] }), .ScanOut({\nScanOut621[7] , 
        \nScanOut621[6] , \nScanOut621[5] , \nScanOut621[4] , \nScanOut621[3] , 
        \nScanOut621[2] , \nScanOut621[1] , \nScanOut621[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_12[7] , \nOut19_12[6] , \nOut19_12[5] , \nOut19_12[4] , 
        \nOut19_12[3] , \nOut19_12[2] , \nOut19_12[1] , \nOut19_12[0] }), 
        .SouthIn({\nOut19_14[7] , \nOut19_14[6] , \nOut19_14[5] , 
        \nOut19_14[4] , \nOut19_14[3] , \nOut19_14[2] , \nOut19_14[1] , 
        \nOut19_14[0] }), .EastIn({\nOut20_13[7] , \nOut20_13[6] , 
        \nOut20_13[5] , \nOut20_13[4] , \nOut20_13[3] , \nOut20_13[2] , 
        \nOut20_13[1] , \nOut20_13[0] }), .WestIn({\nOut18_13[7] , 
        \nOut18_13[6] , \nOut18_13[5] , \nOut18_13[4] , \nOut18_13[3] , 
        \nOut18_13[2] , \nOut18_13[1] , \nOut18_13[0] }), .Out({\nOut19_13[7] , 
        \nOut19_13[6] , \nOut19_13[5] , \nOut19_13[4] , \nOut19_13[3] , 
        \nOut19_13[2] , \nOut19_13[1] , \nOut19_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_626 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut627[7] , \nScanOut627[6] , 
        \nScanOut627[5] , \nScanOut627[4] , \nScanOut627[3] , \nScanOut627[2] , 
        \nScanOut627[1] , \nScanOut627[0] }), .ScanOut({\nScanOut626[7] , 
        \nScanOut626[6] , \nScanOut626[5] , \nScanOut626[4] , \nScanOut626[3] , 
        \nScanOut626[2] , \nScanOut626[1] , \nScanOut626[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_17[7] , \nOut19_17[6] , \nOut19_17[5] , \nOut19_17[4] , 
        \nOut19_17[3] , \nOut19_17[2] , \nOut19_17[1] , \nOut19_17[0] }), 
        .SouthIn({\nOut19_19[7] , \nOut19_19[6] , \nOut19_19[5] , 
        \nOut19_19[4] , \nOut19_19[3] , \nOut19_19[2] , \nOut19_19[1] , 
        \nOut19_19[0] }), .EastIn({\nOut20_18[7] , \nOut20_18[6] , 
        \nOut20_18[5] , \nOut20_18[4] , \nOut20_18[3] , \nOut20_18[2] , 
        \nOut20_18[1] , \nOut20_18[0] }), .WestIn({\nOut18_18[7] , 
        \nOut18_18[6] , \nOut18_18[5] , \nOut18_18[4] , \nOut18_18[3] , 
        \nOut18_18[2] , \nOut18_18[1] , \nOut18_18[0] }), .Out({\nOut19_18[7] , 
        \nOut19_18[6] , \nOut19_18[5] , \nOut19_18[4] , \nOut19_18[3] , 
        \nOut19_18[2] , \nOut19_18[1] , \nOut19_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_858 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut859[7] , \nScanOut859[6] , 
        \nScanOut859[5] , \nScanOut859[4] , \nScanOut859[3] , \nScanOut859[2] , 
        \nScanOut859[1] , \nScanOut859[0] }), .ScanOut({\nScanOut858[7] , 
        \nScanOut858[6] , \nScanOut858[5] , \nScanOut858[4] , \nScanOut858[3] , 
        \nScanOut858[2] , \nScanOut858[1] , \nScanOut858[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_25[7] , \nOut26_25[6] , \nOut26_25[5] , \nOut26_25[4] , 
        \nOut26_25[3] , \nOut26_25[2] , \nOut26_25[1] , \nOut26_25[0] }), 
        .SouthIn({\nOut26_27[7] , \nOut26_27[6] , \nOut26_27[5] , 
        \nOut26_27[4] , \nOut26_27[3] , \nOut26_27[2] , \nOut26_27[1] , 
        \nOut26_27[0] }), .EastIn({\nOut27_26[7] , \nOut27_26[6] , 
        \nOut27_26[5] , \nOut27_26[4] , \nOut27_26[3] , \nOut27_26[2] , 
        \nOut27_26[1] , \nOut27_26[0] }), .WestIn({\nOut25_26[7] , 
        \nOut25_26[6] , \nOut25_26[5] , \nOut25_26[4] , \nOut25_26[3] , 
        \nOut25_26[2] , \nOut25_26[1] , \nOut25_26[0] }), .Out({\nOut26_26[7] , 
        \nOut26_26[6] , \nOut26_26[5] , \nOut26_26[4] , \nOut26_26[3] , 
        \nOut26_26[2] , \nOut26_26[1] , \nOut26_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_180 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut181[7] , \nScanOut181[6] , 
        \nScanOut181[5] , \nScanOut181[4] , \nScanOut181[3] , \nScanOut181[2] , 
        \nScanOut181[1] , \nScanOut181[0] }), .ScanOut({\nScanOut180[7] , 
        \nScanOut180[6] , \nScanOut180[5] , \nScanOut180[4] , \nScanOut180[3] , 
        \nScanOut180[2] , \nScanOut180[1] , \nScanOut180[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_19[7] , \nOut5_19[6] , \nOut5_19[5] , \nOut5_19[4] , 
        \nOut5_19[3] , \nOut5_19[2] , \nOut5_19[1] , \nOut5_19[0] }), 
        .SouthIn({\nOut5_21[7] , \nOut5_21[6] , \nOut5_21[5] , \nOut5_21[4] , 
        \nOut5_21[3] , \nOut5_21[2] , \nOut5_21[1] , \nOut5_21[0] }), .EastIn(
        {\nOut6_20[7] , \nOut6_20[6] , \nOut6_20[5] , \nOut6_20[4] , 
        \nOut6_20[3] , \nOut6_20[2] , \nOut6_20[1] , \nOut6_20[0] }), .WestIn(
        {\nOut4_20[7] , \nOut4_20[6] , \nOut4_20[5] , \nOut4_20[4] , 
        \nOut4_20[3] , \nOut4_20[2] , \nOut4_20[1] , \nOut4_20[0] }), .Out({
        \nOut5_20[7] , \nOut5_20[6] , \nOut5_20[5] , \nOut5_20[4] , 
        \nOut5_20[3] , \nOut5_20[2] , \nOut5_20[1] , \nOut5_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_297 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut298[7] , \nScanOut298[6] , 
        \nScanOut298[5] , \nScanOut298[4] , \nScanOut298[3] , \nScanOut298[2] , 
        \nScanOut298[1] , \nScanOut298[0] }), .ScanOut({\nScanOut297[7] , 
        \nScanOut297[6] , \nScanOut297[5] , \nScanOut297[4] , \nScanOut297[3] , 
        \nScanOut297[2] , \nScanOut297[1] , \nScanOut297[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_8[7] , \nOut9_8[6] , \nOut9_8[5] , \nOut9_8[4] , \nOut9_8[3] , 
        \nOut9_8[2] , \nOut9_8[1] , \nOut9_8[0] }), .SouthIn({\nOut9_10[7] , 
        \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , \nOut9_10[3] , 
        \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }), .EastIn({\nOut10_9[7] , 
        \nOut10_9[6] , \nOut10_9[5] , \nOut10_9[4] , \nOut10_9[3] , 
        \nOut10_9[2] , \nOut10_9[1] , \nOut10_9[0] }), .WestIn({\nOut8_9[7] , 
        \nOut8_9[6] , \nOut8_9[5] , \nOut8_9[4] , \nOut8_9[3] , \nOut8_9[2] , 
        \nOut8_9[1] , \nOut8_9[0] }), .Out({\nOut9_9[7] , \nOut9_9[6] , 
        \nOut9_9[5] , \nOut9_9[4] , \nOut9_9[3] , \nOut9_9[2] , \nOut9_9[1] , 
        \nOut9_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_307 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut308[7] , \nScanOut308[6] , 
        \nScanOut308[5] , \nScanOut308[4] , \nScanOut308[3] , \nScanOut308[2] , 
        \nScanOut308[1] , \nScanOut308[0] }), .ScanOut({\nScanOut307[7] , 
        \nScanOut307[6] , \nScanOut307[5] , \nScanOut307[4] , \nScanOut307[3] , 
        \nScanOut307[2] , \nScanOut307[1] , \nScanOut307[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_18[7] , \nOut9_18[6] , \nOut9_18[5] , \nOut9_18[4] , 
        \nOut9_18[3] , \nOut9_18[2] , \nOut9_18[1] , \nOut9_18[0] }), 
        .SouthIn({\nOut9_20[7] , \nOut9_20[6] , \nOut9_20[5] , \nOut9_20[4] , 
        \nOut9_20[3] , \nOut9_20[2] , \nOut9_20[1] , \nOut9_20[0] }), .EastIn(
        {\nOut10_19[7] , \nOut10_19[6] , \nOut10_19[5] , \nOut10_19[4] , 
        \nOut10_19[3] , \nOut10_19[2] , \nOut10_19[1] , \nOut10_19[0] }), 
        .WestIn({\nOut8_19[7] , \nOut8_19[6] , \nOut8_19[5] , \nOut8_19[4] , 
        \nOut8_19[3] , \nOut8_19[2] , \nOut8_19[1] , \nOut8_19[0] }), .Out({
        \nOut9_19[7] , \nOut9_19[6] , \nOut9_19[5] , \nOut9_19[4] , 
        \nOut9_19[3] , \nOut9_19[2] , \nOut9_19[1] , \nOut9_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_486 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut487[7] , \nScanOut487[6] , 
        \nScanOut487[5] , \nScanOut487[4] , \nScanOut487[3] , \nScanOut487[2] , 
        \nScanOut487[1] , \nScanOut487[0] }), .ScanOut({\nScanOut486[7] , 
        \nScanOut486[6] , \nScanOut486[5] , \nScanOut486[4] , \nScanOut486[3] , 
        \nScanOut486[2] , \nScanOut486[1] , \nScanOut486[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_5[7] , \nOut15_5[6] , \nOut15_5[5] , \nOut15_5[4] , 
        \nOut15_5[3] , \nOut15_5[2] , \nOut15_5[1] , \nOut15_5[0] }), 
        .SouthIn({\nOut15_7[7] , \nOut15_7[6] , \nOut15_7[5] , \nOut15_7[4] , 
        \nOut15_7[3] , \nOut15_7[2] , \nOut15_7[1] , \nOut15_7[0] }), .EastIn(
        {\nOut16_6[7] , \nOut16_6[6] , \nOut16_6[5] , \nOut16_6[4] , 
        \nOut16_6[3] , \nOut16_6[2] , \nOut16_6[1] , \nOut16_6[0] }), .WestIn(
        {\nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }), .Out({
        \nOut15_6[7] , \nOut15_6[6] , \nOut15_6[5] , \nOut15_6[4] , 
        \nOut15_6[3] , \nOut15_6[2] , \nOut15_6[1] , \nOut15_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_964 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut965[7] , \nScanOut965[6] , 
        \nScanOut965[5] , \nScanOut965[4] , \nScanOut965[3] , \nScanOut965[2] , 
        \nScanOut965[1] , \nScanOut965[0] }), .ScanOut({\nScanOut964[7] , 
        \nScanOut964[6] , \nScanOut964[5] , \nScanOut964[4] , \nScanOut964[3] , 
        \nScanOut964[2] , \nScanOut964[1] , \nScanOut964[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_3[7] , \nOut30_3[6] , \nOut30_3[5] , \nOut30_3[4] , 
        \nOut30_3[3] , \nOut30_3[2] , \nOut30_3[1] , \nOut30_3[0] }), 
        .SouthIn({\nOut30_5[7] , \nOut30_5[6] , \nOut30_5[5] , \nOut30_5[4] , 
        \nOut30_5[3] , \nOut30_5[2] , \nOut30_5[1] , \nOut30_5[0] }), .EastIn(
        {\nOut31_4[7] , \nOut31_4[6] , \nOut31_4[5] , \nOut31_4[4] , 
        \nOut31_4[3] , \nOut31_4[2] , \nOut31_4[1] , \nOut31_4[0] }), .WestIn(
        {\nOut29_4[7] , \nOut29_4[6] , \nOut29_4[5] , \nOut29_4[4] , 
        \nOut29_4[3] , \nOut29_4[2] , \nOut29_4[1] , \nOut29_4[0] }), .Out({
        \nOut30_4[7] , \nOut30_4[6] , \nOut30_4[5] , \nOut30_4[4] , 
        \nOut30_4[3] , \nOut30_4[2] , \nOut30_4[1] , \nOut30_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_516 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut517[7] , \nScanOut517[6] , 
        \nScanOut517[5] , \nScanOut517[4] , \nScanOut517[3] , \nScanOut517[2] , 
        \nScanOut517[1] , \nScanOut517[0] }), .ScanOut({\nScanOut516[7] , 
        \nScanOut516[6] , \nScanOut516[5] , \nScanOut516[4] , \nScanOut516[3] , 
        \nScanOut516[2] , \nScanOut516[1] , \nScanOut516[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_3[7] , \nOut16_3[6] , \nOut16_3[5] , \nOut16_3[4] , 
        \nOut16_3[3] , \nOut16_3[2] , \nOut16_3[1] , \nOut16_3[0] }), 
        .SouthIn({\nOut16_5[7] , \nOut16_5[6] , \nOut16_5[5] , \nOut16_5[4] , 
        \nOut16_5[3] , \nOut16_5[2] , \nOut16_5[1] , \nOut16_5[0] }), .EastIn(
        {\nOut17_4[7] , \nOut17_4[6] , \nOut17_4[5] , \nOut17_4[4] , 
        \nOut17_4[3] , \nOut17_4[2] , \nOut17_4[1] , \nOut17_4[0] }), .WestIn(
        {\nOut15_4[7] , \nOut15_4[6] , \nOut15_4[5] , \nOut15_4[4] , 
        \nOut15_4[3] , \nOut15_4[2] , \nOut15_4[1] , \nOut15_4[0] }), .Out({
        \nOut16_4[7] , \nOut16_4[6] , \nOut16_4[5] , \nOut16_4[4] , 
        \nOut16_4[3] , \nOut16_4[2] , \nOut16_4[1] , \nOut16_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_320 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut321[7] , \nScanOut321[6] , 
        \nScanOut321[5] , \nScanOut321[4] , \nScanOut321[3] , \nScanOut321[2] , 
        \nScanOut321[1] , \nScanOut321[0] }), .ScanOut({\nScanOut320[7] , 
        \nScanOut320[6] , \nScanOut320[5] , \nScanOut320[4] , \nScanOut320[3] , 
        \nScanOut320[2] , \nScanOut320[1] , \nScanOut320[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut10_0[7] , \nOut10_0[6] , 
        \nOut10_0[5] , \nOut10_0[4] , \nOut10_0[3] , \nOut10_0[2] , 
        \nOut10_0[1] , \nOut10_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_531 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut532[7] , \nScanOut532[6] , 
        \nScanOut532[5] , \nScanOut532[4] , \nScanOut532[3] , \nScanOut532[2] , 
        \nScanOut532[1] , \nScanOut532[0] }), .ScanOut({\nScanOut531[7] , 
        \nScanOut531[6] , \nScanOut531[5] , \nScanOut531[4] , \nScanOut531[3] , 
        \nScanOut531[2] , \nScanOut531[1] , \nScanOut531[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_18[7] , \nOut16_18[6] , \nOut16_18[5] , \nOut16_18[4] , 
        \nOut16_18[3] , \nOut16_18[2] , \nOut16_18[1] , \nOut16_18[0] }), 
        .SouthIn({\nOut16_20[7] , \nOut16_20[6] , \nOut16_20[5] , 
        \nOut16_20[4] , \nOut16_20[3] , \nOut16_20[2] , \nOut16_20[1] , 
        \nOut16_20[0] }), .EastIn({\nOut17_19[7] , \nOut17_19[6] , 
        \nOut17_19[5] , \nOut17_19[4] , \nOut17_19[3] , \nOut17_19[2] , 
        \nOut17_19[1] , \nOut17_19[0] }), .WestIn({\nOut15_19[7] , 
        \nOut15_19[6] , \nOut15_19[5] , \nOut15_19[4] , \nOut15_19[3] , 
        \nOut15_19[2] , \nOut15_19[1] , \nOut15_19[0] }), .Out({\nOut16_19[7] , 
        \nOut16_19[6] , \nOut16_19[5] , \nOut16_19[4] , \nOut16_19[3] , 
        \nOut16_19[2] , \nOut16_19[1] , \nOut16_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_943 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut944[7] , \nScanOut944[6] , 
        \nScanOut944[5] , \nScanOut944[4] , \nScanOut944[3] , \nScanOut944[2] , 
        \nScanOut944[1] , \nScanOut944[0] }), .ScanOut({\nScanOut943[7] , 
        \nScanOut943[6] , \nScanOut943[5] , \nScanOut943[4] , \nScanOut943[3] , 
        \nScanOut943[2] , \nScanOut943[1] , \nScanOut943[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_14[7] , \nOut29_14[6] , \nOut29_14[5] , \nOut29_14[4] , 
        \nOut29_14[3] , \nOut29_14[2] , \nOut29_14[1] , \nOut29_14[0] }), 
        .SouthIn({\nOut29_16[7] , \nOut29_16[6] , \nOut29_16[5] , 
        \nOut29_16[4] , \nOut29_16[3] , \nOut29_16[2] , \nOut29_16[1] , 
        \nOut29_16[0] }), .EastIn({\nOut30_15[7] , \nOut30_15[6] , 
        \nOut30_15[5] , \nOut30_15[4] , \nOut30_15[3] , \nOut30_15[2] , 
        \nOut30_15[1] , \nOut30_15[0] }), .WestIn({\nOut28_15[7] , 
        \nOut28_15[6] , \nOut28_15[5] , \nOut28_15[4] , \nOut28_15[3] , 
        \nOut28_15[2] , \nOut28_15[1] , \nOut28_15[0] }), .Out({\nOut29_15[7] , 
        \nOut29_15[6] , \nOut29_15[5] , \nOut29_15[4] , \nOut29_15[3] , 
        \nOut29_15[2] , \nOut29_15[1] , \nOut29_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_601 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut602[7] , \nScanOut602[6] , 
        \nScanOut602[5] , \nScanOut602[4] , \nScanOut602[3] , \nScanOut602[2] , 
        \nScanOut602[1] , \nScanOut602[0] }), .ScanOut({\nScanOut601[7] , 
        \nScanOut601[6] , \nScanOut601[5] , \nScanOut601[4] , \nScanOut601[3] , 
        \nScanOut601[2] , \nScanOut601[1] , \nScanOut601[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_24[7] , \nOut18_24[6] , \nOut18_24[5] , \nOut18_24[4] , 
        \nOut18_24[3] , \nOut18_24[2] , \nOut18_24[1] , \nOut18_24[0] }), 
        .SouthIn({\nOut18_26[7] , \nOut18_26[6] , \nOut18_26[5] , 
        \nOut18_26[4] , \nOut18_26[3] , \nOut18_26[2] , \nOut18_26[1] , 
        \nOut18_26[0] }), .EastIn({\nOut19_25[7] , \nOut19_25[6] , 
        \nOut19_25[5] , \nOut19_25[4] , \nOut19_25[3] , \nOut19_25[2] , 
        \nOut19_25[1] , \nOut19_25[0] }), .WestIn({\nOut17_25[7] , 
        \nOut17_25[6] , \nOut17_25[5] , \nOut17_25[4] , \nOut17_25[3] , 
        \nOut17_25[2] , \nOut17_25[1] , \nOut17_25[0] }), .Out({\nOut18_25[7] , 
        \nOut18_25[6] , \nOut18_25[5] , \nOut18_25[4] , \nOut18_25[3] , 
        \nOut18_25[2] , \nOut18_25[1] , \nOut18_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_791 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut792[7] , \nScanOut792[6] , 
        \nScanOut792[5] , \nScanOut792[4] , \nScanOut792[3] , \nScanOut792[2] , 
        \nScanOut792[1] , \nScanOut792[0] }), .ScanOut({\nScanOut791[7] , 
        \nScanOut791[6] , \nScanOut791[5] , \nScanOut791[4] , \nScanOut791[3] , 
        \nScanOut791[2] , \nScanOut791[1] , \nScanOut791[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_22[7] , \nOut24_22[6] , \nOut24_22[5] , \nOut24_22[4] , 
        \nOut24_22[3] , \nOut24_22[2] , \nOut24_22[1] , \nOut24_22[0] }), 
        .SouthIn({\nOut24_24[7] , \nOut24_24[6] , \nOut24_24[5] , 
        \nOut24_24[4] , \nOut24_24[3] , \nOut24_24[2] , \nOut24_24[1] , 
        \nOut24_24[0] }), .EastIn({\nOut25_23[7] , \nOut25_23[6] , 
        \nOut25_23[5] , \nOut25_23[4] , \nOut25_23[3] , \nOut25_23[2] , 
        \nOut25_23[1] , \nOut25_23[0] }), .WestIn({\nOut23_23[7] , 
        \nOut23_23[6] , \nOut23_23[5] , \nOut23_23[4] , \nOut23_23[3] , 
        \nOut23_23[2] , \nOut23_23[1] , \nOut23_23[0] }), .Out({\nOut24_23[7] , 
        \nOut24_23[6] , \nOut24_23[5] , \nOut24_23[4] , \nOut24_23[3] , 
        \nOut24_23[2] , \nOut24_23[1] , \nOut24_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_46 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut47[7] , \nScanOut47[6] , 
        \nScanOut47[5] , \nScanOut47[4] , \nScanOut47[3] , \nScanOut47[2] , 
        \nScanOut47[1] , \nScanOut47[0] }), .ScanOut({\nScanOut46[7] , 
        \nScanOut46[6] , \nScanOut46[5] , \nScanOut46[4] , \nScanOut46[3] , 
        \nScanOut46[2] , \nScanOut46[1] , \nScanOut46[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), 
        .SouthIn({\nOut1_15[7] , \nOut1_15[6] , \nOut1_15[5] , \nOut1_15[4] , 
        \nOut1_15[3] , \nOut1_15[2] , \nOut1_15[1] , \nOut1_15[0] }), .EastIn(
        {\nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), .WestIn(
        {\nOut0_14[7] , \nOut0_14[6] , \nOut0_14[5] , \nOut0_14[4] , 
        \nOut0_14[3] , \nOut0_14[2] , \nOut0_14[1] , \nOut0_14[0] }), .Out({
        \nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_142 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut143[7] , \nScanOut143[6] , 
        \nScanOut143[5] , \nScanOut143[4] , \nScanOut143[3] , \nScanOut143[2] , 
        \nScanOut143[1] , \nScanOut143[0] }), .ScanOut({\nScanOut142[7] , 
        \nScanOut142[6] , \nScanOut142[5] , \nScanOut142[4] , \nScanOut142[3] , 
        \nScanOut142[2] , \nScanOut142[1] , \nScanOut142[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }), 
        .SouthIn({\nOut4_15[7] , \nOut4_15[6] , \nOut4_15[5] , \nOut4_15[4] , 
        \nOut4_15[3] , \nOut4_15[2] , \nOut4_15[1] , \nOut4_15[0] }), .EastIn(
        {\nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }), .WestIn(
        {\nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }), .Out({
        \nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_165 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut166[7] , \nScanOut166[6] , 
        \nScanOut166[5] , \nScanOut166[4] , \nScanOut166[3] , \nScanOut166[2] , 
        \nScanOut166[1] , \nScanOut166[0] }), .ScanOut({\nScanOut165[7] , 
        \nScanOut165[6] , \nScanOut165[5] , \nScanOut165[4] , \nScanOut165[3] , 
        \nScanOut165[2] , \nScanOut165[1] , \nScanOut165[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_4[7] , \nOut5_4[6] , \nOut5_4[5] , \nOut5_4[4] , \nOut5_4[3] , 
        \nOut5_4[2] , \nOut5_4[1] , \nOut5_4[0] }), .SouthIn({\nOut5_6[7] , 
        \nOut5_6[6] , \nOut5_6[5] , \nOut5_6[4] , \nOut5_6[3] , \nOut5_6[2] , 
        \nOut5_6[1] , \nOut5_6[0] }), .EastIn({\nOut6_5[7] , \nOut6_5[6] , 
        \nOut6_5[5] , \nOut6_5[4] , \nOut6_5[3] , \nOut6_5[2] , \nOut6_5[1] , 
        \nOut6_5[0] }), .WestIn({\nOut4_5[7] , \nOut4_5[6] , \nOut4_5[5] , 
        \nOut4_5[4] , \nOut4_5[3] , \nOut4_5[2] , \nOut4_5[1] , \nOut4_5[0] }), 
        .Out({\nOut5_5[7] , \nOut5_5[6] , \nOut5_5[5] , \nOut5_5[4] , 
        \nOut5_5[3] , \nOut5_5[2] , \nOut5_5[1] , \nOut5_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_255 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut256[7] , \nScanOut256[6] , 
        \nScanOut256[5] , \nScanOut256[4] , \nScanOut256[3] , \nScanOut256[2] , 
        \nScanOut256[1] , \nScanOut256[0] }), .ScanOut({\nScanOut255[7] , 
        \nScanOut255[6] , \nScanOut255[5] , \nScanOut255[4] , \nScanOut255[3] , 
        \nScanOut255[2] , \nScanOut255[1] , \nScanOut255[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut7_31[7] , \nOut7_31[6] , 
        \nOut7_31[5] , \nOut7_31[4] , \nOut7_31[3] , \nOut7_31[2] , 
        \nOut7_31[1] , \nOut7_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_369 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut370[7] , \nScanOut370[6] , 
        \nScanOut370[5] , \nScanOut370[4] , \nScanOut370[3] , \nScanOut370[2] , 
        \nScanOut370[1] , \nScanOut370[0] }), .ScanOut({\nScanOut369[7] , 
        \nScanOut369[6] , \nScanOut369[5] , \nScanOut369[4] , \nScanOut369[3] , 
        \nScanOut369[2] , \nScanOut369[1] , \nScanOut369[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_16[7] , \nOut11_16[6] , \nOut11_16[5] , \nOut11_16[4] , 
        \nOut11_16[3] , \nOut11_16[2] , \nOut11_16[1] , \nOut11_16[0] }), 
        .SouthIn({\nOut11_18[7] , \nOut11_18[6] , \nOut11_18[5] , 
        \nOut11_18[4] , \nOut11_18[3] , \nOut11_18[2] , \nOut11_18[1] , 
        \nOut11_18[0] }), .EastIn({\nOut12_17[7] , \nOut12_17[6] , 
        \nOut12_17[5] , \nOut12_17[4] , \nOut12_17[3] , \nOut12_17[2] , 
        \nOut12_17[1] , \nOut12_17[0] }), .WestIn({\nOut10_17[7] , 
        \nOut10_17[6] , \nOut10_17[5] , \nOut10_17[4] , \nOut10_17[3] , 
        \nOut10_17[2] , \nOut10_17[1] , \nOut10_17[0] }), .Out({\nOut11_17[7] , 
        \nOut11_17[6] , \nOut11_17[5] , \nOut11_17[4] , \nOut11_17[3] , 
        \nOut11_17[2] , \nOut11_17[1] , \nOut11_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_578 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut579[7] , \nScanOut579[6] , 
        \nScanOut579[5] , \nScanOut579[4] , \nScanOut579[3] , \nScanOut579[2] , 
        \nScanOut579[1] , \nScanOut579[0] }), .ScanOut({\nScanOut578[7] , 
        \nScanOut578[6] , \nScanOut578[5] , \nScanOut578[4] , \nScanOut578[3] , 
        \nScanOut578[2] , \nScanOut578[1] , \nScanOut578[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_1[7] , \nOut18_1[6] , \nOut18_1[5] , \nOut18_1[4] , 
        \nOut18_1[3] , \nOut18_1[2] , \nOut18_1[1] , \nOut18_1[0] }), 
        .SouthIn({\nOut18_3[7] , \nOut18_3[6] , \nOut18_3[5] , \nOut18_3[4] , 
        \nOut18_3[3] , \nOut18_3[2] , \nOut18_3[1] , \nOut18_3[0] }), .EastIn(
        {\nOut19_2[7] , \nOut19_2[6] , \nOut19_2[5] , \nOut19_2[4] , 
        \nOut19_2[3] , \nOut19_2[2] , \nOut19_2[1] , \nOut19_2[0] }), .WestIn(
        {\nOut17_2[7] , \nOut17_2[6] , \nOut17_2[5] , \nOut17_2[4] , 
        \nOut17_2[3] , \nOut17_2[2] , \nOut17_2[1] , \nOut17_2[0] }), .Out({
        \nOut18_2[7] , \nOut18_2[6] , \nOut18_2[5] , \nOut18_2[4] , 
        \nOut18_2[3] , \nOut18_2[2] , \nOut18_2[1] , \nOut18_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_648 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut649[7] , \nScanOut649[6] , 
        \nScanOut649[5] , \nScanOut649[4] , \nScanOut649[3] , \nScanOut649[2] , 
        \nScanOut649[1] , \nScanOut649[0] }), .ScanOut({\nScanOut648[7] , 
        \nScanOut648[6] , \nScanOut648[5] , \nScanOut648[4] , \nScanOut648[3] , 
        \nScanOut648[2] , \nScanOut648[1] , \nScanOut648[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_7[7] , \nOut20_7[6] , \nOut20_7[5] , \nOut20_7[4] , 
        \nOut20_7[3] , \nOut20_7[2] , \nOut20_7[1] , \nOut20_7[0] }), 
        .SouthIn({\nOut20_9[7] , \nOut20_9[6] , \nOut20_9[5] , \nOut20_9[4] , 
        \nOut20_9[3] , \nOut20_9[2] , \nOut20_9[1] , \nOut20_9[0] }), .EastIn(
        {\nOut21_8[7] , \nOut21_8[6] , \nOut21_8[5] , \nOut21_8[4] , 
        \nOut21_8[3] , \nOut21_8[2] , \nOut21_8[1] , \nOut21_8[0] }), .WestIn(
        {\nOut19_8[7] , \nOut19_8[6] , \nOut19_8[5] , \nOut19_8[4] , 
        \nOut19_8[3] , \nOut19_8[2] , \nOut19_8[1] , \nOut19_8[0] }), .Out({
        \nOut20_8[7] , \nOut20_8[6] , \nOut20_8[5] , \nOut20_8[4] , 
        \nOut20_8[3] , \nOut20_8[2] , \nOut20_8[1] , \nOut20_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_444 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut445[7] , \nScanOut445[6] , 
        \nScanOut445[5] , \nScanOut445[4] , \nScanOut445[3] , \nScanOut445[2] , 
        \nScanOut445[1] , \nScanOut445[0] }), .ScanOut({\nScanOut444[7] , 
        \nScanOut444[6] , \nScanOut444[5] , \nScanOut444[4] , \nScanOut444[3] , 
        \nScanOut444[2] , \nScanOut444[1] , \nScanOut444[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_27[7] , \nOut13_27[6] , \nOut13_27[5] , \nOut13_27[4] , 
        \nOut13_27[3] , \nOut13_27[2] , \nOut13_27[1] , \nOut13_27[0] }), 
        .SouthIn({\nOut13_29[7] , \nOut13_29[6] , \nOut13_29[5] , 
        \nOut13_29[4] , \nOut13_29[3] , \nOut13_29[2] , \nOut13_29[1] , 
        \nOut13_29[0] }), .EastIn({\nOut14_28[7] , \nOut14_28[6] , 
        \nOut14_28[5] , \nOut14_28[4] , \nOut14_28[3] , \nOut14_28[2] , 
        \nOut14_28[1] , \nOut14_28[0] }), .WestIn({\nOut12_28[7] , 
        \nOut12_28[6] , \nOut12_28[5] , \nOut12_28[4] , \nOut12_28[3] , 
        \nOut12_28[2] , \nOut12_28[1] , \nOut12_28[0] }), .Out({\nOut13_28[7] , 
        \nOut13_28[6] , \nOut13_28[5] , \nOut13_28[4] , \nOut13_28[3] , 
        \nOut13_28[2] , \nOut13_28[1] , \nOut13_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_836 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut837[7] , \nScanOut837[6] , 
        \nScanOut837[5] , \nScanOut837[4] , \nScanOut837[3] , \nScanOut837[2] , 
        \nScanOut837[1] , \nScanOut837[0] }), .ScanOut({\nScanOut836[7] , 
        \nScanOut836[6] , \nScanOut836[5] , \nScanOut836[4] , \nScanOut836[3] , 
        \nScanOut836[2] , \nScanOut836[1] , \nScanOut836[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_3[7] , \nOut26_3[6] , \nOut26_3[5] , \nOut26_3[4] , 
        \nOut26_3[3] , \nOut26_3[2] , \nOut26_3[1] , \nOut26_3[0] }), 
        .SouthIn({\nOut26_5[7] , \nOut26_5[6] , \nOut26_5[5] , \nOut26_5[4] , 
        \nOut26_5[3] , \nOut26_5[2] , \nOut26_5[1] , \nOut26_5[0] }), .EastIn(
        {\nOut27_4[7] , \nOut27_4[6] , \nOut27_4[5] , \nOut27_4[4] , 
        \nOut27_4[3] , \nOut27_4[2] , \nOut27_4[1] , \nOut27_4[0] }), .WestIn(
        {\nOut25_4[7] , \nOut25_4[6] , \nOut25_4[5] , \nOut25_4[4] , 
        \nOut25_4[3] , \nOut25_4[2] , \nOut25_4[1] , \nOut25_4[0] }), .Out({
        \nOut26_4[7] , \nOut26_4[6] , \nOut26_4[5] , \nOut26_4[4] , 
        \nOut26_4[3] , \nOut26_4[2] , \nOut26_4[1] , \nOut26_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_774 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut775[7] , \nScanOut775[6] , 
        \nScanOut775[5] , \nScanOut775[4] , \nScanOut775[3] , \nScanOut775[2] , 
        \nScanOut775[1] , \nScanOut775[0] }), .ScanOut({\nScanOut774[7] , 
        \nScanOut774[6] , \nScanOut774[5] , \nScanOut774[4] , \nScanOut774[3] , 
        \nScanOut774[2] , \nScanOut774[1] , \nScanOut774[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_5[7] , \nOut24_5[6] , \nOut24_5[5] , \nOut24_5[4] , 
        \nOut24_5[3] , \nOut24_5[2] , \nOut24_5[1] , \nOut24_5[0] }), 
        .SouthIn({\nOut24_7[7] , \nOut24_7[6] , \nOut24_7[5] , \nOut24_7[4] , 
        \nOut24_7[3] , \nOut24_7[2] , \nOut24_7[1] , \nOut24_7[0] }), .EastIn(
        {\nOut25_6[7] , \nOut25_6[6] , \nOut25_6[5] , \nOut25_6[4] , 
        \nOut25_6[3] , \nOut25_6[2] , \nOut25_6[1] , \nOut25_6[0] }), .WestIn(
        {\nOut23_6[7] , \nOut23_6[6] , \nOut23_6[5] , \nOut23_6[4] , 
        \nOut23_6[3] , \nOut23_6[2] , \nOut23_6[1] , \nOut23_6[0] }), .Out({
        \nOut24_6[7] , \nOut24_6[6] , \nOut24_6[5] , \nOut24_6[4] , 
        \nOut24_6[3] , \nOut24_6[2] , \nOut24_6[1] , \nOut24_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_159 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut160[7] , \nScanOut160[6] , 
        \nScanOut160[5] , \nScanOut160[4] , \nScanOut160[3] , \nScanOut160[2] , 
        \nScanOut160[1] , \nScanOut160[0] }), .ScanOut({\nScanOut159[7] , 
        \nScanOut159[6] , \nScanOut159[5] , \nScanOut159[4] , \nScanOut159[3] , 
        \nScanOut159[2] , \nScanOut159[1] , \nScanOut159[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut4_31[7] , \nOut4_31[6] , 
        \nOut4_31[5] , \nOut4_31[4] , \nOut4_31[3] , \nOut4_31[2] , 
        \nOut4_31[1] , \nOut4_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_269 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut270[7] , \nScanOut270[6] , 
        \nScanOut270[5] , \nScanOut270[4] , \nScanOut270[3] , \nScanOut270[2] , 
        \nScanOut270[1] , \nScanOut270[0] }), .ScanOut({\nScanOut269[7] , 
        \nScanOut269[6] , \nScanOut269[5] , \nScanOut269[4] , \nScanOut269[3] , 
        \nScanOut269[2] , \nScanOut269[1] , \nScanOut269[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }), 
        .SouthIn({\nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }), .EastIn(
        {\nOut9_13[7] , \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , 
        \nOut9_13[3] , \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }), .WestIn(
        {\nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }), .Out({
        \nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_272 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut273[7] , \nScanOut273[6] , 
        \nScanOut273[5] , \nScanOut273[4] , \nScanOut273[3] , \nScanOut273[2] , 
        \nScanOut273[1] , \nScanOut273[0] }), .ScanOut({\nScanOut272[7] , 
        \nScanOut272[6] , \nScanOut272[5] , \nScanOut272[4] , \nScanOut272[3] , 
        \nScanOut272[2] , \nScanOut272[1] , \nScanOut272[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_15[7] , \nOut8_15[6] , \nOut8_15[5] , \nOut8_15[4] , 
        \nOut8_15[3] , \nOut8_15[2] , \nOut8_15[1] , \nOut8_15[0] }), 
        .SouthIn({\nOut8_17[7] , \nOut8_17[6] , \nOut8_17[5] , \nOut8_17[4] , 
        \nOut8_17[3] , \nOut8_17[2] , \nOut8_17[1] , \nOut8_17[0] }), .EastIn(
        {\nOut9_16[7] , \nOut9_16[6] , \nOut9_16[5] , \nOut9_16[4] , 
        \nOut9_16[3] , \nOut9_16[2] , \nOut9_16[1] , \nOut9_16[0] }), .WestIn(
        {\nOut7_16[7] , \nOut7_16[6] , \nOut7_16[5] , \nOut7_16[4] , 
        \nOut7_16[3] , \nOut7_16[2] , \nOut7_16[1] , \nOut7_16[0] }), .Out({
        \nOut8_16[7] , \nOut8_16[6] , \nOut8_16[5] , \nOut8_16[4] , 
        \nOut8_16[3] , \nOut8_16[2] , \nOut8_16[1] , \nOut8_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_753 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut754[7] , \nScanOut754[6] , 
        \nScanOut754[5] , \nScanOut754[4] , \nScanOut754[3] , \nScanOut754[2] , 
        \nScanOut754[1] , \nScanOut754[0] }), .ScanOut({\nScanOut753[7] , 
        \nScanOut753[6] , \nScanOut753[5] , \nScanOut753[4] , \nScanOut753[3] , 
        \nScanOut753[2] , \nScanOut753[1] , \nScanOut753[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_16[7] , \nOut23_16[6] , \nOut23_16[5] , \nOut23_16[4] , 
        \nOut23_16[3] , \nOut23_16[2] , \nOut23_16[1] , \nOut23_16[0] }), 
        .SouthIn({\nOut23_18[7] , \nOut23_18[6] , \nOut23_18[5] , 
        \nOut23_18[4] , \nOut23_18[3] , \nOut23_18[2] , \nOut23_18[1] , 
        \nOut23_18[0] }), .EastIn({\nOut24_17[7] , \nOut24_17[6] , 
        \nOut24_17[5] , \nOut24_17[4] , \nOut24_17[3] , \nOut24_17[2] , 
        \nOut24_17[1] , \nOut24_17[0] }), .WestIn({\nOut22_17[7] , 
        \nOut22_17[6] , \nOut22_17[5] , \nOut22_17[4] , \nOut22_17[3] , 
        \nOut22_17[2] , \nOut22_17[1] , \nOut22_17[0] }), .Out({\nOut23_17[7] , 
        \nOut23_17[6] , \nOut23_17[5] , \nOut23_17[4] , \nOut23_17[3] , 
        \nOut23_17[2] , \nOut23_17[1] , \nOut23_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_811 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut812[7] , \nScanOut812[6] , 
        \nScanOut812[5] , \nScanOut812[4] , \nScanOut812[3] , \nScanOut812[2] , 
        \nScanOut812[1] , \nScanOut812[0] }), .ScanOut({\nScanOut811[7] , 
        \nScanOut811[6] , \nScanOut811[5] , \nScanOut811[4] , \nScanOut811[3] , 
        \nScanOut811[2] , \nScanOut811[1] , \nScanOut811[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_10[7] , \nOut25_10[6] , \nOut25_10[5] , \nOut25_10[4] , 
        \nOut25_10[3] , \nOut25_10[2] , \nOut25_10[1] , \nOut25_10[0] }), 
        .SouthIn({\nOut25_12[7] , \nOut25_12[6] , \nOut25_12[5] , 
        \nOut25_12[4] , \nOut25_12[3] , \nOut25_12[2] , \nOut25_12[1] , 
        \nOut25_12[0] }), .EastIn({\nOut26_11[7] , \nOut26_11[6] , 
        \nOut26_11[5] , \nOut26_11[4] , \nOut26_11[3] , \nOut26_11[2] , 
        \nOut26_11[1] , \nOut26_11[0] }), .WestIn({\nOut24_11[7] , 
        \nOut24_11[6] , \nOut24_11[5] , \nOut24_11[4] , \nOut24_11[3] , 
        \nOut24_11[2] , \nOut24_11[1] , \nOut24_11[0] }), .Out({\nOut25_11[7] , 
        \nOut25_11[6] , \nOut25_11[5] , \nOut25_11[4] , \nOut25_11[3] , 
        \nOut25_11[2] , \nOut25_11[1] , \nOut25_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_981 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut982[7] , \nScanOut982[6] , 
        \nScanOut982[5] , \nScanOut982[4] , \nScanOut982[3] , \nScanOut982[2] , 
        \nScanOut982[1] , \nScanOut982[0] }), .ScanOut({\nScanOut981[7] , 
        \nScanOut981[6] , \nScanOut981[5] , \nScanOut981[4] , \nScanOut981[3] , 
        \nScanOut981[2] , \nScanOut981[1] , \nScanOut981[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_20[7] , \nOut30_20[6] , \nOut30_20[5] , \nOut30_20[4] , 
        \nOut30_20[3] , \nOut30_20[2] , \nOut30_20[1] , \nOut30_20[0] }), 
        .SouthIn({\nOut30_22[7] , \nOut30_22[6] , \nOut30_22[5] , 
        \nOut30_22[4] , \nOut30_22[3] , \nOut30_22[2] , \nOut30_22[1] , 
        \nOut30_22[0] }), .EastIn({\nOut31_21[7] , \nOut31_21[6] , 
        \nOut31_21[5] , \nOut31_21[4] , \nOut31_21[3] , \nOut31_21[2] , 
        \nOut31_21[1] , \nOut31_21[0] }), .WestIn({\nOut29_21[7] , 
        \nOut29_21[6] , \nOut29_21[5] , \nOut29_21[4] , \nOut29_21[3] , 
        \nOut29_21[2] , \nOut29_21[1] , \nOut29_21[0] }), .Out({\nOut30_21[7] , 
        \nOut30_21[6] , \nOut30_21[5] , \nOut30_21[4] , \nOut30_21[3] , 
        \nOut30_21[2] , \nOut30_21[1] , \nOut30_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_463 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut464[7] , \nScanOut464[6] , 
        \nScanOut464[5] , \nScanOut464[4] , \nScanOut464[3] , \nScanOut464[2] , 
        \nScanOut464[1] , \nScanOut464[0] }), .ScanOut({\nScanOut463[7] , 
        \nScanOut463[6] , \nScanOut463[5] , \nScanOut463[4] , \nScanOut463[3] , 
        \nScanOut463[2] , \nScanOut463[1] , \nScanOut463[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_14[7] , \nOut14_14[6] , \nOut14_14[5] , \nOut14_14[4] , 
        \nOut14_14[3] , \nOut14_14[2] , \nOut14_14[1] , \nOut14_14[0] }), 
        .SouthIn({\nOut14_16[7] , \nOut14_16[6] , \nOut14_16[5] , 
        \nOut14_16[4] , \nOut14_16[3] , \nOut14_16[2] , \nOut14_16[1] , 
        \nOut14_16[0] }), .EastIn({\nOut15_15[7] , \nOut15_15[6] , 
        \nOut15_15[5] , \nOut15_15[4] , \nOut15_15[3] , \nOut15_15[2] , 
        \nOut15_15[1] , \nOut15_15[0] }), .WestIn({\nOut13_15[7] , 
        \nOut13_15[6] , \nOut13_15[5] , \nOut13_15[4] , \nOut13_15[3] , 
        \nOut13_15[2] , \nOut13_15[1] , \nOut13_15[0] }), .Out({\nOut14_15[7] , 
        \nOut14_15[6] , \nOut14_15[5] , \nOut14_15[4] , \nOut14_15[3] , 
        \nOut14_15[2] , \nOut14_15[1] , \nOut14_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_478 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut479[7] , \nScanOut479[6] , 
        \nScanOut479[5] , \nScanOut479[4] , \nScanOut479[3] , \nScanOut479[2] , 
        \nScanOut479[1] , \nScanOut479[0] }), .ScanOut({\nScanOut478[7] , 
        \nScanOut478[6] , \nScanOut478[5] , \nScanOut478[4] , \nScanOut478[3] , 
        \nScanOut478[2] , \nScanOut478[1] , \nScanOut478[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_29[7] , \nOut14_29[6] , \nOut14_29[5] , \nOut14_29[4] , 
        \nOut14_29[3] , \nOut14_29[2] , \nOut14_29[1] , \nOut14_29[0] }), 
        .SouthIn({\nOut14_31[7] , \nOut14_31[6] , \nOut14_31[5] , 
        \nOut14_31[4] , \nOut14_31[3] , \nOut14_31[2] , \nOut14_31[1] , 
        \nOut14_31[0] }), .EastIn({\nOut15_30[7] , \nOut15_30[6] , 
        \nOut15_30[5] , \nOut15_30[4] , \nOut15_30[3] , \nOut15_30[2] , 
        \nOut15_30[1] , \nOut15_30[0] }), .WestIn({\nOut13_30[7] , 
        \nOut13_30[6] , \nOut13_30[5] , \nOut13_30[4] , \nOut13_30[3] , 
        \nOut13_30[2] , \nOut13_30[1] , \nOut13_30[0] }), .Out({\nOut14_30[7] , 
        \nOut14_30[6] , \nOut14_30[5] , \nOut14_30[4] , \nOut14_30[3] , 
        \nOut14_30[2] , \nOut14_30[1] , \nOut14_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_372 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut373[7] , \nScanOut373[6] , 
        \nScanOut373[5] , \nScanOut373[4] , \nScanOut373[3] , \nScanOut373[2] , 
        \nScanOut373[1] , \nScanOut373[0] }), .ScanOut({\nScanOut372[7] , 
        \nScanOut372[6] , \nScanOut372[5] , \nScanOut372[4] , \nScanOut372[3] , 
        \nScanOut372[2] , \nScanOut372[1] , \nScanOut372[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_19[7] , \nOut11_19[6] , \nOut11_19[5] , \nOut11_19[4] , 
        \nOut11_19[3] , \nOut11_19[2] , \nOut11_19[1] , \nOut11_19[0] }), 
        .SouthIn({\nOut11_21[7] , \nOut11_21[6] , \nOut11_21[5] , 
        \nOut11_21[4] , \nOut11_21[3] , \nOut11_21[2] , \nOut11_21[1] , 
        \nOut11_21[0] }), .EastIn({\nOut12_20[7] , \nOut12_20[6] , 
        \nOut12_20[5] , \nOut12_20[4] , \nOut12_20[3] , \nOut12_20[2] , 
        \nOut12_20[1] , \nOut12_20[0] }), .WestIn({\nOut10_20[7] , 
        \nOut10_20[6] , \nOut10_20[5] , \nOut10_20[4] , \nOut10_20[3] , 
        \nOut10_20[2] , \nOut10_20[1] , \nOut10_20[0] }), .Out({\nOut11_20[7] , 
        \nOut11_20[6] , \nOut11_20[5] , \nOut11_20[4] , \nOut11_20[3] , 
        \nOut11_20[2] , \nOut11_20[1] , \nOut11_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_563 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut564[7] , \nScanOut564[6] , 
        \nScanOut564[5] , \nScanOut564[4] , \nScanOut564[3] , \nScanOut564[2] , 
        \nScanOut564[1] , \nScanOut564[0] }), .ScanOut({\nScanOut563[7] , 
        \nScanOut563[6] , \nScanOut563[5] , \nScanOut563[4] , \nScanOut563[3] , 
        \nScanOut563[2] , \nScanOut563[1] , \nScanOut563[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_18[7] , \nOut17_18[6] , \nOut17_18[5] , \nOut17_18[4] , 
        \nOut17_18[3] , \nOut17_18[2] , \nOut17_18[1] , \nOut17_18[0] }), 
        .SouthIn({\nOut17_20[7] , \nOut17_20[6] , \nOut17_20[5] , 
        \nOut17_20[4] , \nOut17_20[3] , \nOut17_20[2] , \nOut17_20[1] , 
        \nOut17_20[0] }), .EastIn({\nOut18_19[7] , \nOut18_19[6] , 
        \nOut18_19[5] , \nOut18_19[4] , \nOut18_19[3] , \nOut18_19[2] , 
        \nOut18_19[1] , \nOut18_19[0] }), .WestIn({\nOut16_19[7] , 
        \nOut16_19[6] , \nOut16_19[5] , \nOut16_19[4] , \nOut16_19[3] , 
        \nOut16_19[2] , \nOut16_19[1] , \nOut16_19[0] }), .Out({\nOut17_19[7] , 
        \nOut17_19[6] , \nOut17_19[5] , \nOut17_19[4] , \nOut17_19[3] , 
        \nOut17_19[2] , \nOut17_19[1] , \nOut17_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_748 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut749[7] , \nScanOut749[6] , 
        \nScanOut749[5] , \nScanOut749[4] , \nScanOut749[3] , \nScanOut749[2] , 
        \nScanOut749[1] , \nScanOut749[0] }), .ScanOut({\nScanOut748[7] , 
        \nScanOut748[6] , \nScanOut748[5] , \nScanOut748[4] , \nScanOut748[3] , 
        \nScanOut748[2] , \nScanOut748[1] , \nScanOut748[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_11[7] , \nOut23_11[6] , \nOut23_11[5] , \nOut23_11[4] , 
        \nOut23_11[3] , \nOut23_11[2] , \nOut23_11[1] , \nOut23_11[0] }), 
        .SouthIn({\nOut23_13[7] , \nOut23_13[6] , \nOut23_13[5] , 
        \nOut23_13[4] , \nOut23_13[3] , \nOut23_13[2] , \nOut23_13[1] , 
        \nOut23_13[0] }), .EastIn({\nOut24_12[7] , \nOut24_12[6] , 
        \nOut24_12[5] , \nOut24_12[4] , \nOut24_12[3] , \nOut24_12[2] , 
        \nOut24_12[1] , \nOut24_12[0] }), .WestIn({\nOut22_12[7] , 
        \nOut22_12[6] , \nOut22_12[5] , \nOut22_12[4] , \nOut22_12[3] , 
        \nOut22_12[2] , \nOut22_12[1] , \nOut22_12[0] }), .Out({\nOut23_12[7] , 
        \nOut23_12[6] , \nOut23_12[5] , \nOut23_12[4] , \nOut23_12[3] , 
        \nOut23_12[2] , \nOut23_12[1] , \nOut23_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_881 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut882[7] , \nScanOut882[6] , 
        \nScanOut882[5] , \nScanOut882[4] , \nScanOut882[3] , \nScanOut882[2] , 
        \nScanOut882[1] , \nScanOut882[0] }), .ScanOut({\nScanOut881[7] , 
        \nScanOut881[6] , \nScanOut881[5] , \nScanOut881[4] , \nScanOut881[3] , 
        \nScanOut881[2] , \nScanOut881[1] , \nScanOut881[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_16[7] , \nOut27_16[6] , \nOut27_16[5] , \nOut27_16[4] , 
        \nOut27_16[3] , \nOut27_16[2] , \nOut27_16[1] , \nOut27_16[0] }), 
        .SouthIn({\nOut27_18[7] , \nOut27_18[6] , \nOut27_18[5] , 
        \nOut27_18[4] , \nOut27_18[3] , \nOut27_18[2] , \nOut27_18[1] , 
        \nOut27_18[0] }), .EastIn({\nOut28_17[7] , \nOut28_17[6] , 
        \nOut28_17[5] , \nOut28_17[4] , \nOut28_17[3] , \nOut28_17[2] , 
        \nOut28_17[1] , \nOut28_17[0] }), .WestIn({\nOut26_17[7] , 
        \nOut26_17[6] , \nOut26_17[5] , \nOut26_17[4] , \nOut26_17[3] , 
        \nOut26_17[2] , \nOut26_17[1] , \nOut26_17[0] }), .Out({\nOut27_17[7] , 
        \nOut27_17[6] , \nOut27_17[5] , \nOut27_17[4] , \nOut27_17[3] , 
        \nOut27_17[2] , \nOut27_17[1] , \nOut27_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_911 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut912[7] , \nScanOut912[6] , 
        \nScanOut912[5] , \nScanOut912[4] , \nScanOut912[3] , \nScanOut912[2] , 
        \nScanOut912[1] , \nScanOut912[0] }), .ScanOut({\nScanOut911[7] , 
        \nScanOut911[6] , \nScanOut911[5] , \nScanOut911[4] , \nScanOut911[3] , 
        \nScanOut911[2] , \nScanOut911[1] , \nScanOut911[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_14[7] , \nOut28_14[6] , \nOut28_14[5] , \nOut28_14[4] , 
        \nOut28_14[3] , \nOut28_14[2] , \nOut28_14[1] , \nOut28_14[0] }), 
        .SouthIn({\nOut28_16[7] , \nOut28_16[6] , \nOut28_16[5] , 
        \nOut28_16[4] , \nOut28_16[3] , \nOut28_16[2] , \nOut28_16[1] , 
        \nOut28_16[0] }), .EastIn({\nOut29_15[7] , \nOut29_15[6] , 
        \nOut29_15[5] , \nOut29_15[4] , \nOut29_15[3] , \nOut29_15[2] , 
        \nOut29_15[1] , \nOut29_15[0] }), .WestIn({\nOut27_15[7] , 
        \nOut27_15[6] , \nOut27_15[5] , \nOut27_15[4] , \nOut27_15[3] , 
        \nOut27_15[2] , \nOut27_15[1] , \nOut27_15[0] }), .Out({\nOut28_15[7] , 
        \nOut28_15[6] , \nOut28_15[5] , \nOut28_15[4] , \nOut28_15[3] , 
        \nOut28_15[2] , \nOut28_15[1] , \nOut28_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut2[7] , \nScanOut2[6] , 
        \nScanOut2[5] , \nScanOut2[4] , \nScanOut2[3] , \nScanOut2[2] , 
        \nScanOut2[1] , \nScanOut2[0] }), .ScanOut({\nScanOut1[7] , 
        \nScanOut1[6] , \nScanOut1[5] , \nScanOut1[4] , \nScanOut1[3] , 
        \nScanOut1[2] , \nScanOut1[1] , \nScanOut1[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_1[7] , \nOut0_1[6] , 
        \nOut0_1[5] , \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , 
        \nOut0_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_9 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut10[7] , \nScanOut10[6] , 
        \nScanOut10[5] , \nScanOut10[4] , \nScanOut10[3] , \nScanOut10[2] , 
        \nScanOut10[1] , \nScanOut10[0] }), .ScanOut({\nScanOut9[7] , 
        \nScanOut9[6] , \nScanOut9[5] , \nScanOut9[4] , \nScanOut9[3] , 
        \nScanOut9[2] , \nScanOut9[1] , \nScanOut9[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_9[7] , \nOut0_9[6] , 
        \nOut0_9[5] , \nOut0_9[4] , \nOut0_9[3] , \nOut0_9[2] , \nOut0_9[1] , 
        \nOut0_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_28 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut29[7] , \nScanOut29[6] , 
        \nScanOut29[5] , \nScanOut29[4] , \nScanOut29[3] , \nScanOut29[2] , 
        \nScanOut29[1] , \nScanOut29[0] }), .ScanOut({\nScanOut28[7] , 
        \nScanOut28[6] , \nScanOut28[5] , \nScanOut28[4] , \nScanOut28[3] , 
        \nScanOut28[2] , \nScanOut28[1] , \nScanOut28[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_28[7] , \nOut0_28[6] , 
        \nOut0_28[5] , \nOut0_28[4] , \nOut0_28[3] , \nOut0_28[2] , 
        \nOut0_28[1] , \nOut0_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_61 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut62[7] , \nScanOut62[6] , 
        \nScanOut62[5] , \nScanOut62[4] , \nScanOut62[3] , \nScanOut62[2] , 
        \nScanOut62[1] , \nScanOut62[0] }), .ScanOut({\nScanOut61[7] , 
        \nScanOut61[6] , \nScanOut61[5] , \nScanOut61[4] , \nScanOut61[3] , 
        \nScanOut61[2] , \nScanOut61[1] , \nScanOut61[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_28[7] , \nOut1_28[6] , \nOut1_28[5] , \nOut1_28[4] , 
        \nOut1_28[3] , \nOut1_28[2] , \nOut1_28[1] , \nOut1_28[0] }), 
        .SouthIn({\nOut1_30[7] , \nOut1_30[6] , \nOut1_30[5] , \nOut1_30[4] , 
        \nOut1_30[3] , \nOut1_30[2] , \nOut1_30[1] , \nOut1_30[0] }), .EastIn(
        {\nOut2_29[7] , \nOut2_29[6] , \nOut2_29[5] , \nOut2_29[4] , 
        \nOut2_29[3] , \nOut2_29[2] , \nOut2_29[1] , \nOut2_29[0] }), .WestIn(
        {\nOut0_29[7] , \nOut0_29[6] , \nOut0_29[5] , \nOut0_29[4] , 
        \nOut0_29[3] , \nOut0_29[2] , \nOut0_29[1] , \nOut0_29[0] }), .Out({
        \nOut1_29[7] , \nOut1_29[6] , \nOut1_29[5] , \nOut1_29[4] , 
        \nOut1_29[3] , \nOut1_29[2] , \nOut1_29[1] , \nOut1_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_653 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut654[7] , \nScanOut654[6] , 
        \nScanOut654[5] , \nScanOut654[4] , \nScanOut654[3] , \nScanOut654[2] , 
        \nScanOut654[1] , \nScanOut654[0] }), .ScanOut({\nScanOut653[7] , 
        \nScanOut653[6] , \nScanOut653[5] , \nScanOut653[4] , \nScanOut653[3] , 
        \nScanOut653[2] , \nScanOut653[1] , \nScanOut653[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_12[7] , \nOut20_12[6] , \nOut20_12[5] , \nOut20_12[4] , 
        \nOut20_12[3] , \nOut20_12[2] , \nOut20_12[1] , \nOut20_12[0] }), 
        .SouthIn({\nOut20_14[7] , \nOut20_14[6] , \nOut20_14[5] , 
        \nOut20_14[4] , \nOut20_14[3] , \nOut20_14[2] , \nOut20_14[1] , 
        \nOut20_14[0] }), .EastIn({\nOut21_13[7] , \nOut21_13[6] , 
        \nOut21_13[5] , \nOut21_13[4] , \nOut21_13[3] , \nOut21_13[2] , 
        \nOut21_13[1] , \nOut21_13[0] }), .WestIn({\nOut19_13[7] , 
        \nOut19_13[6] , \nOut19_13[5] , \nOut19_13[4] , \nOut19_13[3] , 
        \nOut19_13[2] , \nOut19_13[1] , \nOut19_13[0] }), .Out({\nOut20_13[7] , 
        \nOut20_13[6] , \nOut20_13[5] , \nOut20_13[4] , \nOut20_13[3] , 
        \nOut20_13[2] , \nOut20_13[1] , \nOut20_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_355 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut356[7] , \nScanOut356[6] , 
        \nScanOut356[5] , \nScanOut356[4] , \nScanOut356[3] , \nScanOut356[2] , 
        \nScanOut356[1] , \nScanOut356[0] }), .ScanOut({\nScanOut355[7] , 
        \nScanOut355[6] , \nScanOut355[5] , \nScanOut355[4] , \nScanOut355[3] , 
        \nScanOut355[2] , \nScanOut355[1] , \nScanOut355[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }), 
        .SouthIn({\nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }), .EastIn(
        {\nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }), .WestIn(
        {\nOut10_3[7] , \nOut10_3[6] , \nOut10_3[5] , \nOut10_3[4] , 
        \nOut10_3[3] , \nOut10_3[2] , \nOut10_3[1] , \nOut10_3[0] }), .Out({
        \nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_674 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut675[7] , \nScanOut675[6] , 
        \nScanOut675[5] , \nScanOut675[4] , \nScanOut675[3] , \nScanOut675[2] , 
        \nScanOut675[1] , \nScanOut675[0] }), .ScanOut({\nScanOut674[7] , 
        \nScanOut674[6] , \nScanOut674[5] , \nScanOut674[4] , \nScanOut674[3] , 
        \nScanOut674[2] , \nScanOut674[1] , \nScanOut674[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_1[7] , \nOut21_1[6] , \nOut21_1[5] , \nOut21_1[4] , 
        \nOut21_1[3] , \nOut21_1[2] , \nOut21_1[1] , \nOut21_1[0] }), 
        .SouthIn({\nOut21_3[7] , \nOut21_3[6] , \nOut21_3[5] , \nOut21_3[4] , 
        \nOut21_3[3] , \nOut21_3[2] , \nOut21_3[1] , \nOut21_3[0] }), .EastIn(
        {\nOut22_2[7] , \nOut22_2[6] , \nOut22_2[5] , \nOut22_2[4] , 
        \nOut22_2[3] , \nOut22_2[2] , \nOut22_2[1] , \nOut22_2[0] }), .WestIn(
        {\nOut20_2[7] , \nOut20_2[6] , \nOut20_2[5] , \nOut20_2[4] , 
        \nOut20_2[3] , \nOut20_2[2] , \nOut20_2[1] , \nOut20_2[0] }), .Out({
        \nOut21_2[7] , \nOut21_2[6] , \nOut21_2[5] , \nOut21_2[4] , 
        \nOut21_2[3] , \nOut21_2[2] , \nOut21_2[1] , \nOut21_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_936 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut937[7] , \nScanOut937[6] , 
        \nScanOut937[5] , \nScanOut937[4] , \nScanOut937[3] , \nScanOut937[2] , 
        \nScanOut937[1] , \nScanOut937[0] }), .ScanOut({\nScanOut936[7] , 
        \nScanOut936[6] , \nScanOut936[5] , \nScanOut936[4] , \nScanOut936[3] , 
        \nScanOut936[2] , \nScanOut936[1] , \nScanOut936[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_7[7] , \nOut29_7[6] , \nOut29_7[5] , \nOut29_7[4] , 
        \nOut29_7[3] , \nOut29_7[2] , \nOut29_7[1] , \nOut29_7[0] }), 
        .SouthIn({\nOut29_9[7] , \nOut29_9[6] , \nOut29_9[5] , \nOut29_9[4] , 
        \nOut29_9[3] , \nOut29_9[2] , \nOut29_9[1] , \nOut29_9[0] }), .EastIn(
        {\nOut30_8[7] , \nOut30_8[6] , \nOut30_8[5] , \nOut30_8[4] , 
        \nOut30_8[3] , \nOut30_8[2] , \nOut30_8[1] , \nOut30_8[0] }), .WestIn(
        {\nOut28_8[7] , \nOut28_8[6] , \nOut28_8[5] , \nOut28_8[4] , 
        \nOut28_8[3] , \nOut28_8[2] , \nOut28_8[1] , \nOut28_8[0] }), .Out({
        \nOut29_8[7] , \nOut29_8[6] , \nOut29_8[5] , \nOut29_8[4] , 
        \nOut29_8[3] , \nOut29_8[2] , \nOut29_8[1] , \nOut29_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_544 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut545[7] , \nScanOut545[6] , 
        \nScanOut545[5] , \nScanOut545[4] , \nScanOut545[3] , \nScanOut545[2] , 
        \nScanOut545[1] , \nScanOut545[0] }), .ScanOut({\nScanOut544[7] , 
        \nScanOut544[6] , \nScanOut544[5] , \nScanOut544[4] , \nScanOut544[3] , 
        \nScanOut544[2] , \nScanOut544[1] , \nScanOut544[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut17_0[7] , \nOut17_0[6] , 
        \nOut17_0[5] , \nOut17_0[4] , \nOut17_0[3] , \nOut17_0[2] , 
        \nOut17_0[1] , \nOut17_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_958 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut959[7] , \nScanOut959[6] , 
        \nScanOut959[5] , \nScanOut959[4] , \nScanOut959[3] , \nScanOut959[2] , 
        \nScanOut959[1] , \nScanOut959[0] }), .ScanOut({\nScanOut958[7] , 
        \nScanOut958[6] , \nScanOut958[5] , \nScanOut958[4] , \nScanOut958[3] , 
        \nScanOut958[2] , \nScanOut958[1] , \nScanOut958[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_29[7] , \nOut29_29[6] , \nOut29_29[5] , \nOut29_29[4] , 
        \nOut29_29[3] , \nOut29_29[2] , \nOut29_29[1] , \nOut29_29[0] }), 
        .SouthIn({\nOut29_31[7] , \nOut29_31[6] , \nOut29_31[5] , 
        \nOut29_31[4] , \nOut29_31[3] , \nOut29_31[2] , \nOut29_31[1] , 
        \nOut29_31[0] }), .EastIn({\nOut30_30[7] , \nOut30_30[6] , 
        \nOut30_30[5] , \nOut30_30[4] , \nOut30_30[3] , \nOut30_30[2] , 
        \nOut30_30[1] , \nOut30_30[0] }), .WestIn({\nOut28_30[7] , 
        \nOut28_30[6] , \nOut28_30[5] , \nOut28_30[4] , \nOut28_30[3] , 
        \nOut28_30[2] , \nOut28_30[1] , \nOut28_30[0] }), .Out({\nOut29_30[7] , 
        \nOut29_30[6] , \nOut29_30[5] , \nOut29_30[4] , \nOut29_30[3] , 
        \nOut29_30[2] , \nOut29_30[1] , \nOut29_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_54 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut55[7] , \nScanOut55[6] , 
        \nScanOut55[5] , \nScanOut55[4] , \nScanOut55[3] , \nScanOut55[2] , 
        \nScanOut55[1] , \nScanOut55[0] }), .ScanOut({\nScanOut54[7] , 
        \nScanOut54[6] , \nScanOut54[5] , \nScanOut54[4] , \nScanOut54[3] , 
        \nScanOut54[2] , \nScanOut54[1] , \nScanOut54[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_21[7] , \nOut1_21[6] , \nOut1_21[5] , \nOut1_21[4] , 
        \nOut1_21[3] , \nOut1_21[2] , \nOut1_21[1] , \nOut1_21[0] }), 
        .SouthIn({\nOut1_23[7] , \nOut1_23[6] , \nOut1_23[5] , \nOut1_23[4] , 
        \nOut1_23[3] , \nOut1_23[2] , \nOut1_23[1] , \nOut1_23[0] }), .EastIn(
        {\nOut2_22[7] , \nOut2_22[6] , \nOut2_22[5] , \nOut2_22[4] , 
        \nOut2_22[3] , \nOut2_22[2] , \nOut2_22[1] , \nOut2_22[0] }), .WestIn(
        {\nOut0_22[7] , \nOut0_22[6] , \nOut0_22[5] , \nOut0_22[4] , 
        \nOut0_22[3] , \nOut0_22[2] , \nOut0_22[1] , \nOut0_22[0] }), .Out({
        \nOut1_22[7] , \nOut1_22[6] , \nOut1_22[5] , \nOut1_22[4] , 
        \nOut1_22[3] , \nOut1_22[2] , \nOut1_22[1] , \nOut1_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_84 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut85[7] , \nScanOut85[6] , 
        \nScanOut85[5] , \nScanOut85[4] , \nScanOut85[3] , \nScanOut85[2] , 
        \nScanOut85[1] , \nScanOut85[0] }), .ScanOut({\nScanOut84[7] , 
        \nScanOut84[6] , \nScanOut84[5] , \nScanOut84[4] , \nScanOut84[3] , 
        \nScanOut84[2] , \nScanOut84[1] , \nScanOut84[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_19[7] , \nOut2_19[6] , \nOut2_19[5] , \nOut2_19[4] , 
        \nOut2_19[3] , \nOut2_19[2] , \nOut2_19[1] , \nOut2_19[0] }), 
        .SouthIn({\nOut2_21[7] , \nOut2_21[6] , \nOut2_21[5] , \nOut2_21[4] , 
        \nOut2_21[3] , \nOut2_21[2] , \nOut2_21[1] , \nOut2_21[0] }), .EastIn(
        {\nOut3_20[7] , \nOut3_20[6] , \nOut3_20[5] , \nOut3_20[4] , 
        \nOut3_20[3] , \nOut3_20[2] , \nOut3_20[1] , \nOut3_20[0] }), .WestIn(
        {\nOut1_20[7] , \nOut1_20[6] , \nOut1_20[5] , \nOut1_20[4] , 
        \nOut1_20[3] , \nOut1_20[2] , \nOut1_20[1] , \nOut1_20[0] }), .Out({
        \nOut2_20[7] , \nOut2_20[6] , \nOut2_20[5] , \nOut2_20[4] , 
        \nOut2_20[3] , \nOut2_20[2] , \nOut2_20[1] , \nOut2_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_110 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut111[7] , \nScanOut111[6] , 
        \nScanOut111[5] , \nScanOut111[4] , \nScanOut111[3] , \nScanOut111[2] , 
        \nScanOut111[1] , \nScanOut111[0] }), .ScanOut({\nScanOut110[7] , 
        \nScanOut110[6] , \nScanOut110[5] , \nScanOut110[4] , \nScanOut110[3] , 
        \nScanOut110[2] , \nScanOut110[1] , \nScanOut110[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }), 
        .SouthIn({\nOut3_15[7] , \nOut3_15[6] , \nOut3_15[5] , \nOut3_15[4] , 
        \nOut3_15[3] , \nOut3_15[2] , \nOut3_15[1] , \nOut3_15[0] }), .EastIn(
        {\nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }), .WestIn(
        {\nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), .Out({
        \nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_691 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut692[7] , \nScanOut692[6] , 
        \nScanOut692[5] , \nScanOut692[4] , \nScanOut692[3] , \nScanOut692[2] , 
        \nScanOut692[1] , \nScanOut692[0] }), .ScanOut({\nScanOut691[7] , 
        \nScanOut691[6] , \nScanOut691[5] , \nScanOut691[4] , \nScanOut691[3] , 
        \nScanOut691[2] , \nScanOut691[1] , \nScanOut691[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_18[7] , \nOut21_18[6] , \nOut21_18[5] , \nOut21_18[4] , 
        \nOut21_18[3] , \nOut21_18[2] , \nOut21_18[1] , \nOut21_18[0] }), 
        .SouthIn({\nOut21_20[7] , \nOut21_20[6] , \nOut21_20[5] , 
        \nOut21_20[4] , \nOut21_20[3] , \nOut21_20[2] , \nOut21_20[1] , 
        \nOut21_20[0] }), .EastIn({\nOut22_19[7] , \nOut22_19[6] , 
        \nOut22_19[5] , \nOut22_19[4] , \nOut22_19[3] , \nOut22_19[2] , 
        \nOut22_19[1] , \nOut22_19[0] }), .WestIn({\nOut20_19[7] , 
        \nOut20_19[6] , \nOut20_19[5] , \nOut20_19[4] , \nOut20_19[3] , 
        \nOut20_19[2] , \nOut20_19[1] , \nOut20_19[0] }), .Out({\nOut21_19[7] , 
        \nOut21_19[6] , \nOut21_19[5] , \nOut21_19[4] , \nOut21_19[3] , 
        \nOut21_19[2] , \nOut21_19[1] , \nOut21_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_701 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut702[7] , \nScanOut702[6] , 
        \nScanOut702[5] , \nScanOut702[4] , \nScanOut702[3] , \nScanOut702[2] , 
        \nScanOut702[1] , \nScanOut702[0] }), .ScanOut({\nScanOut701[7] , 
        \nScanOut701[6] , \nScanOut701[5] , \nScanOut701[4] , \nScanOut701[3] , 
        \nScanOut701[2] , \nScanOut701[1] , \nScanOut701[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_28[7] , \nOut21_28[6] , \nOut21_28[5] , \nOut21_28[4] , 
        \nOut21_28[3] , \nOut21_28[2] , \nOut21_28[1] , \nOut21_28[0] }), 
        .SouthIn({\nOut21_30[7] , \nOut21_30[6] , \nOut21_30[5] , 
        \nOut21_30[4] , \nOut21_30[3] , \nOut21_30[2] , \nOut21_30[1] , 
        \nOut21_30[0] }), .EastIn({\nOut22_29[7] , \nOut22_29[6] , 
        \nOut22_29[5] , \nOut22_29[4] , \nOut22_29[3] , \nOut22_29[2] , 
        \nOut22_29[1] , \nOut22_29[0] }), .WestIn({\nOut20_29[7] , 
        \nOut20_29[6] , \nOut20_29[5] , \nOut20_29[4] , \nOut20_29[3] , 
        \nOut20_29[2] , \nOut20_29[1] , \nOut20_29[0] }), .Out({\nOut21_29[7] , 
        \nOut21_29[6] , \nOut21_29[5] , \nOut21_29[4] , \nOut21_29[3] , 
        \nOut21_29[2] , \nOut21_29[1] , \nOut21_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1007 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1008[7] , \nScanOut1008[6] , 
        \nScanOut1008[5] , \nScanOut1008[4] , \nScanOut1008[3] , 
        \nScanOut1008[2] , \nScanOut1008[1] , \nScanOut1008[0] }), .ScanOut({
        \nScanOut1007[7] , \nScanOut1007[6] , \nScanOut1007[5] , 
        \nScanOut1007[4] , \nScanOut1007[3] , \nScanOut1007[2] , 
        \nScanOut1007[1] , \nScanOut1007[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_15[7] , \nOut31_15[6] , \nOut31_15[5] , 
        \nOut31_15[4] , \nOut31_15[3] , \nOut31_15[2] , \nOut31_15[1] , 
        \nOut31_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_96 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut97[7] , \nScanOut97[6] , 
        \nScanOut97[5] , \nScanOut97[4] , \nScanOut97[3] , \nScanOut97[2] , 
        \nScanOut97[1] , \nScanOut97[0] }), .ScanOut({\nScanOut96[7] , 
        \nScanOut96[6] , \nScanOut96[5] , \nScanOut96[4] , \nScanOut96[3] , 
        \nScanOut96[2] , \nScanOut96[1] , \nScanOut96[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut3_0[7] , \nOut3_0[6] , 
        \nOut3_0[5] , \nOut3_0[4] , \nOut3_0[3] , \nOut3_0[2] , \nOut3_0[1] , 
        \nOut3_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_102 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut103[7] , \nScanOut103[6] , 
        \nScanOut103[5] , \nScanOut103[4] , \nScanOut103[3] , \nScanOut103[2] , 
        \nScanOut103[1] , \nScanOut103[0] }), .ScanOut({\nScanOut102[7] , 
        \nScanOut102[6] , \nScanOut102[5] , \nScanOut102[4] , \nScanOut102[3] , 
        \nScanOut102[2] , \nScanOut102[1] , \nScanOut102[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_5[7] , \nOut3_5[6] , \nOut3_5[5] , \nOut3_5[4] , \nOut3_5[3] , 
        \nOut3_5[2] , \nOut3_5[1] , \nOut3_5[0] }), .SouthIn({\nOut3_7[7] , 
        \nOut3_7[6] , \nOut3_7[5] , \nOut3_7[4] , \nOut3_7[3] , \nOut3_7[2] , 
        \nOut3_7[1] , \nOut3_7[0] }), .EastIn({\nOut4_6[7] , \nOut4_6[6] , 
        \nOut4_6[5] , \nOut4_6[4] , \nOut4_6[3] , \nOut4_6[2] , \nOut4_6[1] , 
        \nOut4_6[0] }), .WestIn({\nOut2_6[7] , \nOut2_6[6] , \nOut2_6[5] , 
        \nOut2_6[4] , \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , \nOut2_6[0] }), 
        .Out({\nOut3_6[7] , \nOut3_6[6] , \nOut3_6[5] , \nOut3_6[4] , 
        \nOut3_6[3] , \nOut3_6[2] , \nOut3_6[1] , \nOut3_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_137 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut138[7] , \nScanOut138[6] , 
        \nScanOut138[5] , \nScanOut138[4] , \nScanOut138[3] , \nScanOut138[2] , 
        \nScanOut138[1] , \nScanOut138[0] }), .ScanOut({\nScanOut137[7] , 
        \nScanOut137[6] , \nScanOut137[5] , \nScanOut137[4] , \nScanOut137[3] , 
        \nScanOut137[2] , \nScanOut137[1] , \nScanOut137[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_8[7] , \nOut4_8[6] , \nOut4_8[5] , \nOut4_8[4] , \nOut4_8[3] , 
        \nOut4_8[2] , \nOut4_8[1] , \nOut4_8[0] }), .SouthIn({\nOut4_10[7] , 
        \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , \nOut4_10[3] , 
        \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }), .EastIn({\nOut5_9[7] , 
        \nOut5_9[6] , \nOut5_9[5] , \nOut5_9[4] , \nOut5_9[3] , \nOut5_9[2] , 
        \nOut5_9[1] , \nOut5_9[0] }), .WestIn({\nOut3_9[7] , \nOut3_9[6] , 
        \nOut3_9[5] , \nOut3_9[4] , \nOut3_9[3] , \nOut3_9[2] , \nOut3_9[1] , 
        \nOut3_9[0] }), .Out({\nOut4_9[7] , \nOut4_9[6] , \nOut4_9[5] , 
        \nOut4_9[4] , \nOut4_9[3] , \nOut4_9[2] , \nOut4_9[1] , \nOut4_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_207 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut208[7] , \nScanOut208[6] , 
        \nScanOut208[5] , \nScanOut208[4] , \nScanOut208[3] , \nScanOut208[2] , 
        \nScanOut208[1] , \nScanOut208[0] }), .ScanOut({\nScanOut207[7] , 
        \nScanOut207[6] , \nScanOut207[5] , \nScanOut207[4] , \nScanOut207[3] , 
        \nScanOut207[2] , \nScanOut207[1] , \nScanOut207[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }), 
        .SouthIn({\nOut6_16[7] , \nOut6_16[6] , \nOut6_16[5] , \nOut6_16[4] , 
        \nOut6_16[3] , \nOut6_16[2] , \nOut6_16[1] , \nOut6_16[0] }), .EastIn(
        {\nOut7_15[7] , \nOut7_15[6] , \nOut7_15[5] , \nOut7_15[4] , 
        \nOut7_15[3] , \nOut7_15[2] , \nOut7_15[1] , \nOut7_15[0] }), .WestIn(
        {\nOut5_15[7] , \nOut5_15[6] , \nOut5_15[5] , \nOut5_15[4] , 
        \nOut5_15[3] , \nOut5_15[2] , \nOut5_15[1] , \nOut5_15[0] }), .Out({
        \nOut6_15[7] , \nOut6_15[6] , \nOut6_15[5] , \nOut6_15[4] , 
        \nOut6_15[3] , \nOut6_15[2] , \nOut6_15[1] , \nOut6_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_220 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut221[7] , \nScanOut221[6] , 
        \nScanOut221[5] , \nScanOut221[4] , \nScanOut221[3] , \nScanOut221[2] , 
        \nScanOut221[1] , \nScanOut221[0] }), .ScanOut({\nScanOut220[7] , 
        \nScanOut220[6] , \nScanOut220[5] , \nScanOut220[4] , \nScanOut220[3] , 
        \nScanOut220[2] , \nScanOut220[1] , \nScanOut220[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_27[7] , \nOut6_27[6] , \nOut6_27[5] , \nOut6_27[4] , 
        \nOut6_27[3] , \nOut6_27[2] , \nOut6_27[1] , \nOut6_27[0] }), 
        .SouthIn({\nOut6_29[7] , \nOut6_29[6] , \nOut6_29[5] , \nOut6_29[4] , 
        \nOut6_29[3] , \nOut6_29[2] , \nOut6_29[1] , \nOut6_29[0] }), .EastIn(
        {\nOut7_28[7] , \nOut7_28[6] , \nOut7_28[5] , \nOut7_28[4] , 
        \nOut7_28[3] , \nOut7_28[2] , \nOut7_28[1] , \nOut7_28[0] }), .WestIn(
        {\nOut5_28[7] , \nOut5_28[6] , \nOut5_28[5] , \nOut5_28[4] , 
        \nOut5_28[3] , \nOut5_28[2] , \nOut5_28[1] , \nOut5_28[0] }), .Out({
        \nOut6_28[7] , \nOut6_28[6] , \nOut6_28[5] , \nOut6_28[4] , 
        \nOut6_28[3] , \nOut6_28[2] , \nOut6_28[1] , \nOut6_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_843 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut844[7] , \nScanOut844[6] , 
        \nScanOut844[5] , \nScanOut844[4] , \nScanOut844[3] , \nScanOut844[2] , 
        \nScanOut844[1] , \nScanOut844[0] }), .ScanOut({\nScanOut843[7] , 
        \nScanOut843[6] , \nScanOut843[5] , \nScanOut843[4] , \nScanOut843[3] , 
        \nScanOut843[2] , \nScanOut843[1] , \nScanOut843[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_10[7] , \nOut26_10[6] , \nOut26_10[5] , \nOut26_10[4] , 
        \nOut26_10[3] , \nOut26_10[2] , \nOut26_10[1] , \nOut26_10[0] }), 
        .SouthIn({\nOut26_12[7] , \nOut26_12[6] , \nOut26_12[5] , 
        \nOut26_12[4] , \nOut26_12[3] , \nOut26_12[2] , \nOut26_12[1] , 
        \nOut26_12[0] }), .EastIn({\nOut27_11[7] , \nOut27_11[6] , 
        \nOut27_11[5] , \nOut27_11[4] , \nOut27_11[3] , \nOut27_11[2] , 
        \nOut27_11[1] , \nOut27_11[0] }), .WestIn({\nOut25_11[7] , 
        \nOut25_11[6] , \nOut25_11[5] , \nOut25_11[4] , \nOut25_11[3] , 
        \nOut25_11[2] , \nOut25_11[1] , \nOut25_11[0] }), .Out({\nOut26_11[7] , 
        \nOut26_11[6] , \nOut26_11[5] , \nOut26_11[4] , \nOut26_11[3] , 
        \nOut26_11[2] , \nOut26_11[1] , \nOut26_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_397 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut398[7] , \nScanOut398[6] , 
        \nScanOut398[5] , \nScanOut398[4] , \nScanOut398[3] , \nScanOut398[2] , 
        \nScanOut398[1] , \nScanOut398[0] }), .ScanOut({\nScanOut397[7] , 
        \nScanOut397[6] , \nScanOut397[5] , \nScanOut397[4] , \nScanOut397[3] , 
        \nScanOut397[2] , \nScanOut397[1] , \nScanOut397[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_12[7] , \nOut12_12[6] , \nOut12_12[5] , \nOut12_12[4] , 
        \nOut12_12[3] , \nOut12_12[2] , \nOut12_12[1] , \nOut12_12[0] }), 
        .SouthIn({\nOut12_14[7] , \nOut12_14[6] , \nOut12_14[5] , 
        \nOut12_14[4] , \nOut12_14[3] , \nOut12_14[2] , \nOut12_14[1] , 
        \nOut12_14[0] }), .EastIn({\nOut13_13[7] , \nOut13_13[6] , 
        \nOut13_13[5] , \nOut13_13[4] , \nOut13_13[3] , \nOut13_13[2] , 
        \nOut13_13[1] , \nOut13_13[0] }), .WestIn({\nOut11_13[7] , 
        \nOut11_13[6] , \nOut11_13[5] , \nOut11_13[4] , \nOut11_13[3] , 
        \nOut11_13[2] , \nOut11_13[1] , \nOut11_13[0] }), .Out({\nOut12_13[7] , 
        \nOut12_13[6] , \nOut12_13[5] , \nOut12_13[4] , \nOut12_13[3] , 
        \nOut12_13[2] , \nOut12_13[1] , \nOut12_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_416 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut417[7] , \nScanOut417[6] , 
        \nScanOut417[5] , \nScanOut417[4] , \nScanOut417[3] , \nScanOut417[2] , 
        \nScanOut417[1] , \nScanOut417[0] }), .ScanOut({\nScanOut416[7] , 
        \nScanOut416[6] , \nScanOut416[5] , \nScanOut416[4] , \nScanOut416[3] , 
        \nScanOut416[2] , \nScanOut416[1] , \nScanOut416[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut13_0[7] , \nOut13_0[6] , 
        \nOut13_0[5] , \nOut13_0[4] , \nOut13_0[3] , \nOut13_0[2] , 
        \nOut13_0[1] , \nOut13_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_431 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut432[7] , \nScanOut432[6] , 
        \nScanOut432[5] , \nScanOut432[4] , \nScanOut432[3] , \nScanOut432[2] , 
        \nScanOut432[1] , \nScanOut432[0] }), .ScanOut({\nScanOut431[7] , 
        \nScanOut431[6] , \nScanOut431[5] , \nScanOut431[4] , \nScanOut431[3] , 
        \nScanOut431[2] , \nScanOut431[1] , \nScanOut431[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_14[7] , \nOut13_14[6] , \nOut13_14[5] , \nOut13_14[4] , 
        \nOut13_14[3] , \nOut13_14[2] , \nOut13_14[1] , \nOut13_14[0] }), 
        .SouthIn({\nOut13_16[7] , \nOut13_16[6] , \nOut13_16[5] , 
        \nOut13_16[4] , \nOut13_16[3] , \nOut13_16[2] , \nOut13_16[1] , 
        \nOut13_16[0] }), .EastIn({\nOut14_15[7] , \nOut14_15[6] , 
        \nOut14_15[5] , \nOut14_15[4] , \nOut14_15[3] , \nOut14_15[2] , 
        \nOut14_15[1] , \nOut14_15[0] }), .WestIn({\nOut12_15[7] , 
        \nOut12_15[6] , \nOut12_15[5] , \nOut12_15[4] , \nOut12_15[3] , 
        \nOut12_15[2] , \nOut12_15[1] , \nOut12_15[0] }), .Out({\nOut13_15[7] , 
        \nOut13_15[6] , \nOut13_15[5] , \nOut13_15[4] , \nOut13_15[3] , 
        \nOut13_15[2] , \nOut13_15[1] , \nOut13_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_864 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut865[7] , \nScanOut865[6] , 
        \nScanOut865[5] , \nScanOut865[4] , \nScanOut865[3] , \nScanOut865[2] , 
        \nScanOut865[1] , \nScanOut865[0] }), .ScanOut({\nScanOut864[7] , 
        \nScanOut864[6] , \nScanOut864[5] , \nScanOut864[4] , \nScanOut864[3] , 
        \nScanOut864[2] , \nScanOut864[1] , \nScanOut864[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut27_0[7] , \nOut27_0[6] , 
        \nOut27_0[5] , \nOut27_0[4] , \nOut27_0[3] , \nOut27_0[2] , 
        \nOut27_0[1] , \nOut27_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_586 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut587[7] , \nScanOut587[6] , 
        \nScanOut587[5] , \nScanOut587[4] , \nScanOut587[3] , \nScanOut587[2] , 
        \nScanOut587[1] , \nScanOut587[0] }), .ScanOut({\nScanOut586[7] , 
        \nScanOut586[6] , \nScanOut586[5] , \nScanOut586[4] , \nScanOut586[3] , 
        \nScanOut586[2] , \nScanOut586[1] , \nScanOut586[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_9[7] , \nOut18_9[6] , \nOut18_9[5] , \nOut18_9[4] , 
        \nOut18_9[3] , \nOut18_9[2] , \nOut18_9[1] , \nOut18_9[0] }), 
        .SouthIn({\nOut18_11[7] , \nOut18_11[6] , \nOut18_11[5] , 
        \nOut18_11[4] , \nOut18_11[3] , \nOut18_11[2] , \nOut18_11[1] , 
        \nOut18_11[0] }), .EastIn({\nOut19_10[7] , \nOut19_10[6] , 
        \nOut19_10[5] , \nOut19_10[4] , \nOut19_10[3] , \nOut19_10[2] , 
        \nOut19_10[1] , \nOut19_10[0] }), .WestIn({\nOut17_10[7] , 
        \nOut17_10[6] , \nOut17_10[5] , \nOut17_10[4] , \nOut17_10[3] , 
        \nOut17_10[2] , \nOut17_10[1] , \nOut17_10[0] }), .Out({\nOut18_10[7] , 
        \nOut18_10[6] , \nOut18_10[5] , \nOut18_10[4] , \nOut18_10[3] , 
        \nOut18_10[2] , \nOut18_10[1] , \nOut18_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_726 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut727[7] , \nScanOut727[6] , 
        \nScanOut727[5] , \nScanOut727[4] , \nScanOut727[3] , \nScanOut727[2] , 
        \nScanOut727[1] , \nScanOut727[0] }), .ScanOut({\nScanOut726[7] , 
        \nScanOut726[6] , \nScanOut726[5] , \nScanOut726[4] , \nScanOut726[3] , 
        \nScanOut726[2] , \nScanOut726[1] , \nScanOut726[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_21[7] , \nOut22_21[6] , \nOut22_21[5] , \nOut22_21[4] , 
        \nOut22_21[3] , \nOut22_21[2] , \nOut22_21[1] , \nOut22_21[0] }), 
        .SouthIn({\nOut22_23[7] , \nOut22_23[6] , \nOut22_23[5] , 
        \nOut22_23[4] , \nOut22_23[3] , \nOut22_23[2] , \nOut22_23[1] , 
        \nOut22_23[0] }), .EastIn({\nOut23_22[7] , \nOut23_22[6] , 
        \nOut23_22[5] , \nOut23_22[4] , \nOut23_22[3] , \nOut23_22[2] , 
        \nOut23_22[1] , \nOut23_22[0] }), .WestIn({\nOut21_22[7] , 
        \nOut21_22[6] , \nOut21_22[5] , \nOut21_22[4] , \nOut21_22[3] , 
        \nOut21_22[2] , \nOut21_22[1] , \nOut21_22[0] }), .Out({\nOut22_22[7] , 
        \nOut22_22[6] , \nOut22_22[5] , \nOut22_22[4] , \nOut22_22[3] , 
        \nOut22_22[2] , \nOut22_22[1] , \nOut22_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_713 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut714[7] , \nScanOut714[6] , 
        \nScanOut714[5] , \nScanOut714[4] , \nScanOut714[3] , \nScanOut714[2] , 
        \nScanOut714[1] , \nScanOut714[0] }), .ScanOut({\nScanOut713[7] , 
        \nScanOut713[6] , \nScanOut713[5] , \nScanOut713[4] , \nScanOut713[3] , 
        \nScanOut713[2] , \nScanOut713[1] , \nScanOut713[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_8[7] , \nOut22_8[6] , \nOut22_8[5] , \nOut22_8[4] , 
        \nOut22_8[3] , \nOut22_8[2] , \nOut22_8[1] , \nOut22_8[0] }), 
        .SouthIn({\nOut22_10[7] , \nOut22_10[6] , \nOut22_10[5] , 
        \nOut22_10[4] , \nOut22_10[3] , \nOut22_10[2] , \nOut22_10[1] , 
        \nOut22_10[0] }), .EastIn({\nOut23_9[7] , \nOut23_9[6] , \nOut23_9[5] , 
        \nOut23_9[4] , \nOut23_9[3] , \nOut23_9[2] , \nOut23_9[1] , 
        \nOut23_9[0] }), .WestIn({\nOut21_9[7] , \nOut21_9[6] , \nOut21_9[5] , 
        \nOut21_9[4] , \nOut21_9[3] , \nOut21_9[2] , \nOut21_9[1] , 
        \nOut21_9[0] }), .Out({\nOut22_9[7] , \nOut22_9[6] , \nOut22_9[5] , 
        \nOut22_9[4] , \nOut22_9[3] , \nOut22_9[2] , \nOut22_9[1] , 
        \nOut22_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1020 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1021[7] , \nScanOut1021[6] , 
        \nScanOut1021[5] , \nScanOut1021[4] , \nScanOut1021[3] , 
        \nScanOut1021[2] , \nScanOut1021[1] , \nScanOut1021[0] }), .ScanOut({
        \nScanOut1020[7] , \nScanOut1020[6] , \nScanOut1020[5] , 
        \nScanOut1020[4] , \nScanOut1020[3] , \nScanOut1020[2] , 
        \nScanOut1020[1] , \nScanOut1020[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_28[7] , \nOut31_28[6] , \nOut31_28[5] , 
        \nOut31_28[4] , \nOut31_28[3] , \nOut31_28[2] , \nOut31_28[1] , 
        \nOut31_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_683 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut684[7] , \nScanOut684[6] , 
        \nScanOut684[5] , \nScanOut684[4] , \nScanOut684[3] , \nScanOut684[2] , 
        \nScanOut684[1] , \nScanOut684[0] }), .ScanOut({\nScanOut683[7] , 
        \nScanOut683[6] , \nScanOut683[5] , \nScanOut683[4] , \nScanOut683[3] , 
        \nScanOut683[2] , \nScanOut683[1] , \nScanOut683[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_10[7] , \nOut21_10[6] , \nOut21_10[5] , \nOut21_10[4] , 
        \nOut21_10[3] , \nOut21_10[2] , \nOut21_10[1] , \nOut21_10[0] }), 
        .SouthIn({\nOut21_12[7] , \nOut21_12[6] , \nOut21_12[5] , 
        \nOut21_12[4] , \nOut21_12[3] , \nOut21_12[2] , \nOut21_12[1] , 
        \nOut21_12[0] }), .EastIn({\nOut22_11[7] , \nOut22_11[6] , 
        \nOut22_11[5] , \nOut22_11[4] , \nOut22_11[3] , \nOut22_11[2] , 
        \nOut22_11[1] , \nOut22_11[0] }), .WestIn({\nOut20_11[7] , 
        \nOut20_11[6] , \nOut20_11[5] , \nOut20_11[4] , \nOut20_11[3] , 
        \nOut20_11[2] , \nOut20_11[1] , \nOut20_11[0] }), .Out({\nOut21_11[7] , 
        \nOut21_11[6] , \nOut21_11[5] , \nOut21_11[4] , \nOut21_11[3] , 
        \nOut21_11[2] , \nOut21_11[1] , \nOut21_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1015 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1016[7] , \nScanOut1016[6] , 
        \nScanOut1016[5] , \nScanOut1016[4] , \nScanOut1016[3] , 
        \nScanOut1016[2] , \nScanOut1016[1] , \nScanOut1016[0] }), .ScanOut({
        \nScanOut1015[7] , \nScanOut1015[6] , \nScanOut1015[5] , 
        \nScanOut1015[4] , \nScanOut1015[3] , \nScanOut1015[2] , 
        \nScanOut1015[1] , \nScanOut1015[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_23[7] , \nOut31_23[6] , \nOut31_23[5] , 
        \nOut31_23[4] , \nOut31_23[3] , \nOut31_23[2] , \nOut31_23[1] , 
        \nOut31_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_125 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut126[7] , \nScanOut126[6] , 
        \nScanOut126[5] , \nScanOut126[4] , \nScanOut126[3] , \nScanOut126[2] , 
        \nScanOut126[1] , \nScanOut126[0] }), .ScanOut({\nScanOut125[7] , 
        \nScanOut125[6] , \nScanOut125[5] , \nScanOut125[4] , \nScanOut125[3] , 
        \nScanOut125[2] , \nScanOut125[1] , \nScanOut125[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_28[7] , \nOut3_28[6] , \nOut3_28[5] , \nOut3_28[4] , 
        \nOut3_28[3] , \nOut3_28[2] , \nOut3_28[1] , \nOut3_28[0] }), 
        .SouthIn({\nOut3_30[7] , \nOut3_30[6] , \nOut3_30[5] , \nOut3_30[4] , 
        \nOut3_30[3] , \nOut3_30[2] , \nOut3_30[1] , \nOut3_30[0] }), .EastIn(
        {\nOut4_29[7] , \nOut4_29[6] , \nOut4_29[5] , \nOut4_29[4] , 
        \nOut4_29[3] , \nOut4_29[2] , \nOut4_29[1] , \nOut4_29[0] }), .WestIn(
        {\nOut2_29[7] , \nOut2_29[6] , \nOut2_29[5] , \nOut2_29[4] , 
        \nOut2_29[3] , \nOut2_29[2] , \nOut2_29[1] , \nOut2_29[0] }), .Out({
        \nOut3_29[7] , \nOut3_29[6] , \nOut3_29[5] , \nOut3_29[4] , 
        \nOut3_29[3] , \nOut3_29[2] , \nOut3_29[1] , \nOut3_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_215 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut216[7] , \nScanOut216[6] , 
        \nScanOut216[5] , \nScanOut216[4] , \nScanOut216[3] , \nScanOut216[2] , 
        \nScanOut216[1] , \nScanOut216[0] }), .ScanOut({\nScanOut215[7] , 
        \nScanOut215[6] , \nScanOut215[5] , \nScanOut215[4] , \nScanOut215[3] , 
        \nScanOut215[2] , \nScanOut215[1] , \nScanOut215[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_22[7] , \nOut6_22[6] , \nOut6_22[5] , \nOut6_22[4] , 
        \nOut6_22[3] , \nOut6_22[2] , \nOut6_22[1] , \nOut6_22[0] }), 
        .SouthIn({\nOut6_24[7] , \nOut6_24[6] , \nOut6_24[5] , \nOut6_24[4] , 
        \nOut6_24[3] , \nOut6_24[2] , \nOut6_24[1] , \nOut6_24[0] }), .EastIn(
        {\nOut7_23[7] , \nOut7_23[6] , \nOut7_23[5] , \nOut7_23[4] , 
        \nOut7_23[3] , \nOut7_23[2] , \nOut7_23[1] , \nOut7_23[0] }), .WestIn(
        {\nOut5_23[7] , \nOut5_23[6] , \nOut5_23[5] , \nOut5_23[4] , 
        \nOut5_23[3] , \nOut5_23[2] , \nOut5_23[1] , \nOut5_23[0] }), .Out({
        \nOut6_23[7] , \nOut6_23[6] , \nOut6_23[5] , \nOut6_23[4] , 
        \nOut6_23[3] , \nOut6_23[2] , \nOut6_23[1] , \nOut6_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_232 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut233[7] , \nScanOut233[6] , 
        \nScanOut233[5] , \nScanOut233[4] , \nScanOut233[3] , \nScanOut233[2] , 
        \nScanOut233[1] , \nScanOut233[0] }), .ScanOut({\nScanOut232[7] , 
        \nScanOut232[6] , \nScanOut232[5] , \nScanOut232[4] , \nScanOut232[3] , 
        \nScanOut232[2] , \nScanOut232[1] , \nScanOut232[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_7[7] , \nOut7_7[6] , \nOut7_7[5] , \nOut7_7[4] , \nOut7_7[3] , 
        \nOut7_7[2] , \nOut7_7[1] , \nOut7_7[0] }), .SouthIn({\nOut7_9[7] , 
        \nOut7_9[6] , \nOut7_9[5] , \nOut7_9[4] , \nOut7_9[3] , \nOut7_9[2] , 
        \nOut7_9[1] , \nOut7_9[0] }), .EastIn({\nOut8_8[7] , \nOut8_8[6] , 
        \nOut8_8[5] , \nOut8_8[4] , \nOut8_8[3] , \nOut8_8[2] , \nOut8_8[1] , 
        \nOut8_8[0] }), .WestIn({\nOut6_8[7] , \nOut6_8[6] , \nOut6_8[5] , 
        \nOut6_8[4] , \nOut6_8[3] , \nOut6_8[2] , \nOut6_8[1] , \nOut6_8[0] }), 
        .Out({\nOut7_8[7] , \nOut7_8[6] , \nOut7_8[5] , \nOut7_8[4] , 
        \nOut7_8[3] , \nOut7_8[2] , \nOut7_8[1] , \nOut7_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_423 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut424[7] , \nScanOut424[6] , 
        \nScanOut424[5] , \nScanOut424[4] , \nScanOut424[3] , \nScanOut424[2] , 
        \nScanOut424[1] , \nScanOut424[0] }), .ScanOut({\nScanOut423[7] , 
        \nScanOut423[6] , \nScanOut423[5] , \nScanOut423[4] , \nScanOut423[3] , 
        \nScanOut423[2] , \nScanOut423[1] , \nScanOut423[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }), 
        .SouthIn({\nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }), .EastIn(
        {\nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }), .WestIn(
        {\nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }), .Out({
        \nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_594 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut595[7] , \nScanOut595[6] , 
        \nScanOut595[5] , \nScanOut595[4] , \nScanOut595[3] , \nScanOut595[2] , 
        \nScanOut595[1] , \nScanOut595[0] }), .ScanOut({\nScanOut594[7] , 
        \nScanOut594[6] , \nScanOut594[5] , \nScanOut594[4] , \nScanOut594[3] , 
        \nScanOut594[2] , \nScanOut594[1] , \nScanOut594[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_17[7] , \nOut18_17[6] , \nOut18_17[5] , \nOut18_17[4] , 
        \nOut18_17[3] , \nOut18_17[2] , \nOut18_17[1] , \nOut18_17[0] }), 
        .SouthIn({\nOut18_19[7] , \nOut18_19[6] , \nOut18_19[5] , 
        \nOut18_19[4] , \nOut18_19[3] , \nOut18_19[2] , \nOut18_19[1] , 
        \nOut18_19[0] }), .EastIn({\nOut19_18[7] , \nOut19_18[6] , 
        \nOut19_18[5] , \nOut19_18[4] , \nOut19_18[3] , \nOut19_18[2] , 
        \nOut19_18[1] , \nOut19_18[0] }), .WestIn({\nOut17_18[7] , 
        \nOut17_18[6] , \nOut17_18[5] , \nOut17_18[4] , \nOut17_18[3] , 
        \nOut17_18[2] , \nOut17_18[1] , \nOut17_18[0] }), .Out({\nOut18_18[7] , 
        \nOut18_18[6] , \nOut18_18[5] , \nOut18_18[4] , \nOut18_18[3] , 
        \nOut18_18[2] , \nOut18_18[1] , \nOut18_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_851 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut852[7] , \nScanOut852[6] , 
        \nScanOut852[5] , \nScanOut852[4] , \nScanOut852[3] , \nScanOut852[2] , 
        \nScanOut852[1] , \nScanOut852[0] }), .ScanOut({\nScanOut851[7] , 
        \nScanOut851[6] , \nScanOut851[5] , \nScanOut851[4] , \nScanOut851[3] , 
        \nScanOut851[2] , \nScanOut851[1] , \nScanOut851[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_18[7] , \nOut26_18[6] , \nOut26_18[5] , \nOut26_18[4] , 
        \nOut26_18[3] , \nOut26_18[2] , \nOut26_18[1] , \nOut26_18[0] }), 
        .SouthIn({\nOut26_20[7] , \nOut26_20[6] , \nOut26_20[5] , 
        \nOut26_20[4] , \nOut26_20[3] , \nOut26_20[2] , \nOut26_20[1] , 
        \nOut26_20[0] }), .EastIn({\nOut27_19[7] , \nOut27_19[6] , 
        \nOut27_19[5] , \nOut27_19[4] , \nOut27_19[3] , \nOut27_19[2] , 
        \nOut27_19[1] , \nOut27_19[0] }), .WestIn({\nOut25_19[7] , 
        \nOut25_19[6] , \nOut25_19[5] , \nOut25_19[4] , \nOut25_19[3] , 
        \nOut25_19[2] , \nOut25_19[1] , \nOut25_19[0] }), .Out({\nOut26_19[7] , 
        \nOut26_19[6] , \nOut26_19[5] , \nOut26_19[4] , \nOut26_19[3] , 
        \nOut26_19[2] , \nOut26_19[1] , \nOut26_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_385 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut386[7] , \nScanOut386[6] , 
        \nScanOut386[5] , \nScanOut386[4] , \nScanOut386[3] , \nScanOut386[2] , 
        \nScanOut386[1] , \nScanOut386[0] }), .ScanOut({\nScanOut385[7] , 
        \nScanOut385[6] , \nScanOut385[5] , \nScanOut385[4] , \nScanOut385[3] , 
        \nScanOut385[2] , \nScanOut385[1] , \nScanOut385[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_0[7] , \nOut12_0[6] , \nOut12_0[5] , \nOut12_0[4] , 
        \nOut12_0[3] , \nOut12_0[2] , \nOut12_0[1] , \nOut12_0[0] }), 
        .SouthIn({\nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }), .EastIn(
        {\nOut13_1[7] , \nOut13_1[6] , \nOut13_1[5] , \nOut13_1[4] , 
        \nOut13_1[3] , \nOut13_1[2] , \nOut13_1[1] , \nOut13_1[0] }), .WestIn(
        {\nOut11_1[7] , \nOut11_1[6] , \nOut11_1[5] , \nOut11_1[4] , 
        \nOut11_1[3] , \nOut11_1[2] , \nOut11_1[1] , \nOut11_1[0] }), .Out({
        \nOut12_1[7] , \nOut12_1[6] , \nOut12_1[5] , \nOut12_1[4] , 
        \nOut12_1[3] , \nOut12_1[2] , \nOut12_1[1] , \nOut12_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_404 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut405[7] , \nScanOut405[6] , 
        \nScanOut405[5] , \nScanOut405[4] , \nScanOut405[3] , \nScanOut405[2] , 
        \nScanOut405[1] , \nScanOut405[0] }), .ScanOut({\nScanOut404[7] , 
        \nScanOut404[6] , \nScanOut404[5] , \nScanOut404[4] , \nScanOut404[3] , 
        \nScanOut404[2] , \nScanOut404[1] , \nScanOut404[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_19[7] , \nOut12_19[6] , \nOut12_19[5] , \nOut12_19[4] , 
        \nOut12_19[3] , \nOut12_19[2] , \nOut12_19[1] , \nOut12_19[0] }), 
        .SouthIn({\nOut12_21[7] , \nOut12_21[6] , \nOut12_21[5] , 
        \nOut12_21[4] , \nOut12_21[3] , \nOut12_21[2] , \nOut12_21[1] , 
        \nOut12_21[0] }), .EastIn({\nOut13_20[7] , \nOut13_20[6] , 
        \nOut13_20[5] , \nOut13_20[4] , \nOut13_20[3] , \nOut13_20[2] , 
        \nOut13_20[1] , \nOut13_20[0] }), .WestIn({\nOut11_20[7] , 
        \nOut11_20[6] , \nOut11_20[5] , \nOut11_20[4] , \nOut11_20[3] , 
        \nOut11_20[2] , \nOut11_20[1] , \nOut11_20[0] }), .Out({\nOut12_20[7] , 
        \nOut12_20[6] , \nOut12_20[5] , \nOut12_20[4] , \nOut12_20[3] , 
        \nOut12_20[2] , \nOut12_20[1] , \nOut12_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_876 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut877[7] , \nScanOut877[6] , 
        \nScanOut877[5] , \nScanOut877[4] , \nScanOut877[3] , \nScanOut877[2] , 
        \nScanOut877[1] , \nScanOut877[0] }), .ScanOut({\nScanOut876[7] , 
        \nScanOut876[6] , \nScanOut876[5] , \nScanOut876[4] , \nScanOut876[3] , 
        \nScanOut876[2] , \nScanOut876[1] , \nScanOut876[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_11[7] , \nOut27_11[6] , \nOut27_11[5] , \nOut27_11[4] , 
        \nOut27_11[3] , \nOut27_11[2] , \nOut27_11[1] , \nOut27_11[0] }), 
        .SouthIn({\nOut27_13[7] , \nOut27_13[6] , \nOut27_13[5] , 
        \nOut27_13[4] , \nOut27_13[3] , \nOut27_13[2] , \nOut27_13[1] , 
        \nOut27_13[0] }), .EastIn({\nOut28_12[7] , \nOut28_12[6] , 
        \nOut28_12[5] , \nOut28_12[4] , \nOut28_12[3] , \nOut28_12[2] , 
        \nOut28_12[1] , \nOut28_12[0] }), .WestIn({\nOut26_12[7] , 
        \nOut26_12[6] , \nOut26_12[5] , \nOut26_12[4] , \nOut26_12[3] , 
        \nOut26_12[2] , \nOut26_12[1] , \nOut26_12[0] }), .Out({\nOut27_12[7] , 
        \nOut27_12[6] , \nOut27_12[5] , \nOut27_12[4] , \nOut27_12[3] , 
        \nOut27_12[2] , \nOut27_12[1] , \nOut27_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_189 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut190[7] , \nScanOut190[6] , 
        \nScanOut190[5] , \nScanOut190[4] , \nScanOut190[3] , \nScanOut190[2] , 
        \nScanOut190[1] , \nScanOut190[0] }), .ScanOut({\nScanOut189[7] , 
        \nScanOut189[6] , \nScanOut189[5] , \nScanOut189[4] , \nScanOut189[3] , 
        \nScanOut189[2] , \nScanOut189[1] , \nScanOut189[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_28[7] , \nOut5_28[6] , \nOut5_28[5] , \nOut5_28[4] , 
        \nOut5_28[3] , \nOut5_28[2] , \nOut5_28[1] , \nOut5_28[0] }), 
        .SouthIn({\nOut5_30[7] , \nOut5_30[6] , \nOut5_30[5] , \nOut5_30[4] , 
        \nOut5_30[3] , \nOut5_30[2] , \nOut5_30[1] , \nOut5_30[0] }), .EastIn(
        {\nOut6_29[7] , \nOut6_29[6] , \nOut6_29[5] , \nOut6_29[4] , 
        \nOut6_29[3] , \nOut6_29[2] , \nOut6_29[1] , \nOut6_29[0] }), .WestIn(
        {\nOut4_29[7] , \nOut4_29[6] , \nOut4_29[5] , \nOut4_29[4] , 
        \nOut4_29[3] , \nOut4_29[2] , \nOut4_29[1] , \nOut4_29[0] }), .Out({
        \nOut5_29[7] , \nOut5_29[6] , \nOut5_29[5] , \nOut5_29[4] , 
        \nOut5_29[3] , \nOut5_29[2] , \nOut5_29[1] , \nOut5_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_734 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut735[7] , \nScanOut735[6] , 
        \nScanOut735[5] , \nScanOut735[4] , \nScanOut735[3] , \nScanOut735[2] , 
        \nScanOut735[1] , \nScanOut735[0] }), .ScanOut({\nScanOut734[7] , 
        \nScanOut734[6] , \nScanOut734[5] , \nScanOut734[4] , \nScanOut734[3] , 
        \nScanOut734[2] , \nScanOut734[1] , \nScanOut734[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_29[7] , \nOut22_29[6] , \nOut22_29[5] , \nOut22_29[4] , 
        \nOut22_29[3] , \nOut22_29[2] , \nOut22_29[1] , \nOut22_29[0] }), 
        .SouthIn({\nOut22_31[7] , \nOut22_31[6] , \nOut22_31[5] , 
        \nOut22_31[4] , \nOut22_31[3] , \nOut22_31[2] , \nOut22_31[1] , 
        \nOut22_31[0] }), .EastIn({\nOut23_30[7] , \nOut23_30[6] , 
        \nOut23_30[5] , \nOut23_30[4] , \nOut23_30[3] , \nOut23_30[2] , 
        \nOut23_30[1] , \nOut23_30[0] }), .WestIn({\nOut21_30[7] , 
        \nOut21_30[6] , \nOut21_30[5] , \nOut21_30[4] , \nOut21_30[3] , 
        \nOut21_30[2] , \nOut21_30[1] , \nOut21_30[0] }), .Out({\nOut22_30[7] , 
        \nOut22_30[6] , \nOut22_30[5] , \nOut22_30[4] , \nOut22_30[3] , 
        \nOut22_30[2] , \nOut22_30[1] , \nOut22_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_798 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut799[7] , \nScanOut799[6] , 
        \nScanOut799[5] , \nScanOut799[4] , \nScanOut799[3] , \nScanOut799[2] , 
        \nScanOut799[1] , \nScanOut799[0] }), .ScanOut({\nScanOut798[7] , 
        \nScanOut798[6] , \nScanOut798[5] , \nScanOut798[4] , \nScanOut798[3] , 
        \nScanOut798[2] , \nScanOut798[1] , \nScanOut798[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_29[7] , \nOut24_29[6] , \nOut24_29[5] , \nOut24_29[4] , 
        \nOut24_29[3] , \nOut24_29[2] , \nOut24_29[1] , \nOut24_29[0] }), 
        .SouthIn({\nOut24_31[7] , \nOut24_31[6] , \nOut24_31[5] , 
        \nOut24_31[4] , \nOut24_31[3] , \nOut24_31[2] , \nOut24_31[1] , 
        \nOut24_31[0] }), .EastIn({\nOut25_30[7] , \nOut25_30[6] , 
        \nOut25_30[5] , \nOut25_30[4] , \nOut25_30[3] , \nOut25_30[2] , 
        \nOut25_30[1] , \nOut25_30[0] }), .WestIn({\nOut23_30[7] , 
        \nOut23_30[6] , \nOut23_30[5] , \nOut23_30[4] , \nOut23_30[3] , 
        \nOut23_30[2] , \nOut23_30[1] , \nOut23_30[0] }), .Out({\nOut24_30[7] , 
        \nOut24_30[6] , \nOut24_30[5] , \nOut24_30[4] , \nOut24_30[3] , 
        \nOut24_30[2] , \nOut24_30[1] , \nOut24_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_329 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut330[7] , \nScanOut330[6] , 
        \nScanOut330[5] , \nScanOut330[4] , \nScanOut330[3] , \nScanOut330[2] , 
        \nScanOut330[1] , \nScanOut330[0] }), .ScanOut({\nScanOut329[7] , 
        \nScanOut329[6] , \nScanOut329[5] , \nScanOut329[4] , \nScanOut329[3] , 
        \nScanOut329[2] , \nScanOut329[1] , \nScanOut329[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_8[7] , \nOut10_8[6] , \nOut10_8[5] , \nOut10_8[4] , 
        \nOut10_8[3] , \nOut10_8[2] , \nOut10_8[1] , \nOut10_8[0] }), 
        .SouthIn({\nOut10_10[7] , \nOut10_10[6] , \nOut10_10[5] , 
        \nOut10_10[4] , \nOut10_10[3] , \nOut10_10[2] , \nOut10_10[1] , 
        \nOut10_10[0] }), .EastIn({\nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , 
        \nOut11_9[4] , \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , 
        \nOut11_9[0] }), .WestIn({\nOut9_9[7] , \nOut9_9[6] , \nOut9_9[5] , 
        \nOut9_9[4] , \nOut9_9[3] , \nOut9_9[2] , \nOut9_9[1] , \nOut9_9[0] }), 
        .Out({\nOut10_9[7] , \nOut10_9[6] , \nOut10_9[5] , \nOut10_9[4] , 
        \nOut10_9[3] , \nOut10_9[2] , \nOut10_9[1] , \nOut10_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_608 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut609[7] , \nScanOut609[6] , 
        \nScanOut609[5] , \nScanOut609[4] , \nScanOut609[3] , \nScanOut609[2] , 
        \nScanOut609[1] , \nScanOut609[0] }), .ScanOut({\nScanOut608[7] , 
        \nScanOut608[6] , \nScanOut608[5] , \nScanOut608[4] , \nScanOut608[3] , 
        \nScanOut608[2] , \nScanOut608[1] , \nScanOut608[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut19_0[7] , \nOut19_0[6] , 
        \nOut19_0[5] , \nOut19_0[4] , \nOut19_0[3] , \nOut19_0[2] , 
        \nOut19_0[1] , \nOut19_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_360 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut361[7] , \nScanOut361[6] , 
        \nScanOut361[5] , \nScanOut361[4] , \nScanOut361[3] , \nScanOut361[2] , 
        \nScanOut361[1] , \nScanOut361[0] }), .ScanOut({\nScanOut360[7] , 
        \nScanOut360[6] , \nScanOut360[5] , \nScanOut360[4] , \nScanOut360[3] , 
        \nScanOut360[2] , \nScanOut360[1] , \nScanOut360[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }), 
        .SouthIn({\nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , \nOut11_9[4] , 
        \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , \nOut11_9[0] }), .EastIn(
        {\nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }), .WestIn(
        {\nOut10_8[7] , \nOut10_8[6] , \nOut10_8[5] , \nOut10_8[4] , 
        \nOut10_8[3] , \nOut10_8[2] , \nOut10_8[1] , \nOut10_8[0] }), .Out({
        \nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_538 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut539[7] , \nScanOut539[6] , 
        \nScanOut539[5] , \nScanOut539[4] , \nScanOut539[3] , \nScanOut539[2] , 
        \nScanOut539[1] , \nScanOut539[0] }), .ScanOut({\nScanOut538[7] , 
        \nScanOut538[6] , \nScanOut538[5] , \nScanOut538[4] , \nScanOut538[3] , 
        \nScanOut538[2] , \nScanOut538[1] , \nScanOut538[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_25[7] , \nOut16_25[6] , \nOut16_25[5] , \nOut16_25[4] , 
        \nOut16_25[3] , \nOut16_25[2] , \nOut16_25[1] , \nOut16_25[0] }), 
        .SouthIn({\nOut16_27[7] , \nOut16_27[6] , \nOut16_27[5] , 
        \nOut16_27[4] , \nOut16_27[3] , \nOut16_27[2] , \nOut16_27[1] , 
        \nOut16_27[0] }), .EastIn({\nOut17_26[7] , \nOut17_26[6] , 
        \nOut17_26[5] , \nOut17_26[4] , \nOut17_26[3] , \nOut17_26[2] , 
        \nOut17_26[1] , \nOut17_26[0] }), .WestIn({\nOut15_26[7] , 
        \nOut15_26[6] , \nOut15_26[5] , \nOut15_26[4] , \nOut15_26[3] , 
        \nOut15_26[2] , \nOut15_26[1] , \nOut15_26[0] }), .Out({\nOut16_26[7] , 
        \nOut16_26[6] , \nOut16_26[5] , \nOut16_26[4] , \nOut16_26[3] , 
        \nOut16_26[2] , \nOut16_26[1] , \nOut16_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_571 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut572[7] , \nScanOut572[6] , 
        \nScanOut572[5] , \nScanOut572[4] , \nScanOut572[3] , \nScanOut572[2] , 
        \nScanOut572[1] , \nScanOut572[0] }), .ScanOut({\nScanOut571[7] , 
        \nScanOut571[6] , \nScanOut571[5] , \nScanOut571[4] , \nScanOut571[3] , 
        \nScanOut571[2] , \nScanOut571[1] , \nScanOut571[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_26[7] , \nOut17_26[6] , \nOut17_26[5] , \nOut17_26[4] , 
        \nOut17_26[3] , \nOut17_26[2] , \nOut17_26[1] , \nOut17_26[0] }), 
        .SouthIn({\nOut17_28[7] , \nOut17_28[6] , \nOut17_28[5] , 
        \nOut17_28[4] , \nOut17_28[3] , \nOut17_28[2] , \nOut17_28[1] , 
        \nOut17_28[0] }), .EastIn({\nOut18_27[7] , \nOut18_27[6] , 
        \nOut18_27[5] , \nOut18_27[4] , \nOut18_27[3] , \nOut18_27[2] , 
        \nOut18_27[1] , \nOut18_27[0] }), .WestIn({\nOut16_27[7] , 
        \nOut16_27[6] , \nOut16_27[5] , \nOut16_27[4] , \nOut16_27[3] , 
        \nOut16_27[2] , \nOut16_27[1] , \nOut16_27[0] }), .Out({\nOut17_27[7] , 
        \nOut17_27[6] , \nOut17_27[5] , \nOut17_27[4] , \nOut17_27[3] , 
        \nOut17_27[2] , \nOut17_27[1] , \nOut17_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_893 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut894[7] , \nScanOut894[6] , 
        \nScanOut894[5] , \nScanOut894[4] , \nScanOut894[3] , \nScanOut894[2] , 
        \nScanOut894[1] , \nScanOut894[0] }), .ScanOut({\nScanOut893[7] , 
        \nScanOut893[6] , \nScanOut893[5] , \nScanOut893[4] , \nScanOut893[3] , 
        \nScanOut893[2] , \nScanOut893[1] , \nScanOut893[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_28[7] , \nOut27_28[6] , \nOut27_28[5] , \nOut27_28[4] , 
        \nOut27_28[3] , \nOut27_28[2] , \nOut27_28[1] , \nOut27_28[0] }), 
        .SouthIn({\nOut27_30[7] , \nOut27_30[6] , \nOut27_30[5] , 
        \nOut27_30[4] , \nOut27_30[3] , \nOut27_30[2] , \nOut27_30[1] , 
        \nOut27_30[0] }), .EastIn({\nOut28_29[7] , \nOut28_29[6] , 
        \nOut28_29[5] , \nOut28_29[4] , \nOut28_29[3] , \nOut28_29[2] , 
        \nOut28_29[1] , \nOut28_29[0] }), .WestIn({\nOut26_29[7] , 
        \nOut26_29[6] , \nOut26_29[5] , \nOut26_29[4] , \nOut26_29[3] , 
        \nOut26_29[2] , \nOut26_29[1] , \nOut26_29[0] }), .Out({\nOut27_29[7] , 
        \nOut27_29[6] , \nOut27_29[5] , \nOut27_29[4] , \nOut27_29[3] , 
        \nOut27_29[2] , \nOut27_29[1] , \nOut27_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_903 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut904[7] , \nScanOut904[6] , 
        \nScanOut904[5] , \nScanOut904[4] , \nScanOut904[3] , \nScanOut904[2] , 
        \nScanOut904[1] , \nScanOut904[0] }), .ScanOut({\nScanOut903[7] , 
        \nScanOut903[6] , \nScanOut903[5] , \nScanOut903[4] , \nScanOut903[3] , 
        \nScanOut903[2] , \nScanOut903[1] , \nScanOut903[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_6[7] , \nOut28_6[6] , \nOut28_6[5] , \nOut28_6[4] , 
        \nOut28_6[3] , \nOut28_6[2] , \nOut28_6[1] , \nOut28_6[0] }), 
        .SouthIn({\nOut28_8[7] , \nOut28_8[6] , \nOut28_8[5] , \nOut28_8[4] , 
        \nOut28_8[3] , \nOut28_8[2] , \nOut28_8[1] , \nOut28_8[0] }), .EastIn(
        {\nOut29_7[7] , \nOut29_7[6] , \nOut29_7[5] , \nOut29_7[4] , 
        \nOut29_7[3] , \nOut29_7[2] , \nOut29_7[1] , \nOut29_7[0] }), .WestIn(
        {\nOut27_7[7] , \nOut27_7[6] , \nOut27_7[5] , \nOut27_7[4] , 
        \nOut27_7[3] , \nOut27_7[2] , \nOut27_7[1] , \nOut27_7[0] }), .Out({
        \nOut28_7[7] , \nOut28_7[6] , \nOut28_7[5] , \nOut28_7[4] , 
        \nOut28_7[3] , \nOut28_7[2] , \nOut28_7[1] , \nOut28_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_68 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut69[7] , \nScanOut69[6] , 
        \nScanOut69[5] , \nScanOut69[4] , \nScanOut69[3] , \nScanOut69[2] , 
        \nScanOut69[1] , \nScanOut69[0] }), .ScanOut({\nScanOut68[7] , 
        \nScanOut68[6] , \nScanOut68[5] , \nScanOut68[4] , \nScanOut68[3] , 
        \nScanOut68[2] , \nScanOut68[1] , \nScanOut68[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_3[7] , \nOut2_3[6] , \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , 
        \nOut2_3[2] , \nOut2_3[1] , \nOut2_3[0] }), .SouthIn({\nOut2_5[7] , 
        \nOut2_5[6] , \nOut2_5[5] , \nOut2_5[4] , \nOut2_5[3] , \nOut2_5[2] , 
        \nOut2_5[1] , \nOut2_5[0] }), .EastIn({\nOut3_4[7] , \nOut3_4[6] , 
        \nOut3_4[5] , \nOut3_4[4] , \nOut3_4[3] , \nOut3_4[2] , \nOut3_4[1] , 
        \nOut3_4[0] }), .WestIn({\nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , 
        \nOut1_4[4] , \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }), 
        .Out({\nOut2_4[7] , \nOut2_4[6] , \nOut2_4[5] , \nOut2_4[4] , 
        \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , \nOut2_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_73 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut74[7] , \nScanOut74[6] , 
        \nScanOut74[5] , \nScanOut74[4] , \nScanOut74[3] , \nScanOut74[2] , 
        \nScanOut74[1] , \nScanOut74[0] }), .ScanOut({\nScanOut73[7] , 
        \nScanOut73[6] , \nScanOut73[5] , \nScanOut73[4] , \nScanOut73[3] , 
        \nScanOut73[2] , \nScanOut73[1] , \nScanOut73[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_8[7] , \nOut2_8[6] , \nOut2_8[5] , \nOut2_8[4] , \nOut2_8[3] , 
        \nOut2_8[2] , \nOut2_8[1] , \nOut2_8[0] }), .SouthIn({\nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), .EastIn({\nOut3_9[7] , 
        \nOut3_9[6] , \nOut3_9[5] , \nOut3_9[4] , \nOut3_9[3] , \nOut3_9[2] , 
        \nOut3_9[1] , \nOut3_9[0] }), .WestIn({\nOut1_9[7] , \nOut1_9[6] , 
        \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , \nOut1_9[1] , 
        \nOut1_9[0] }), .Out({\nOut2_9[7] , \nOut2_9[6] , \nOut2_9[5] , 
        \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , \nOut2_9[1] , \nOut2_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_641 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut642[7] , \nScanOut642[6] , 
        \nScanOut642[5] , \nScanOut642[4] , \nScanOut642[3] , \nScanOut642[2] , 
        \nScanOut642[1] , \nScanOut642[0] }), .ScanOut({\nScanOut641[7] , 
        \nScanOut641[6] , \nScanOut641[5] , \nScanOut641[4] , \nScanOut641[3] , 
        \nScanOut641[2] , \nScanOut641[1] , \nScanOut641[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_0[7] , \nOut20_0[6] , \nOut20_0[5] , \nOut20_0[4] , 
        \nOut20_0[3] , \nOut20_0[2] , \nOut20_0[1] , \nOut20_0[0] }), 
        .SouthIn({\nOut20_2[7] , \nOut20_2[6] , \nOut20_2[5] , \nOut20_2[4] , 
        \nOut20_2[3] , \nOut20_2[2] , \nOut20_2[1] , \nOut20_2[0] }), .EastIn(
        {\nOut21_1[7] , \nOut21_1[6] , \nOut21_1[5] , \nOut21_1[4] , 
        \nOut21_1[3] , \nOut21_1[2] , \nOut21_1[1] , \nOut21_1[0] }), .WestIn(
        {\nOut19_1[7] , \nOut19_1[6] , \nOut19_1[5] , \nOut19_1[4] , 
        \nOut19_1[3] , \nOut19_1[2] , \nOut19_1[1] , \nOut19_1[0] }), .Out({
        \nOut20_1[7] , \nOut20_1[6] , \nOut20_1[5] , \nOut20_1[4] , 
        \nOut20_1[3] , \nOut20_1[2] , \nOut20_1[1] , \nOut20_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_150 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut151[7] , \nScanOut151[6] , 
        \nScanOut151[5] , \nScanOut151[4] , \nScanOut151[3] , \nScanOut151[2] , 
        \nScanOut151[1] , \nScanOut151[0] }), .ScanOut({\nScanOut150[7] , 
        \nScanOut150[6] , \nScanOut150[5] , \nScanOut150[4] , \nScanOut150[3] , 
        \nScanOut150[2] , \nScanOut150[1] , \nScanOut150[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_21[7] , \nOut4_21[6] , \nOut4_21[5] , \nOut4_21[4] , 
        \nOut4_21[3] , \nOut4_21[2] , \nOut4_21[1] , \nOut4_21[0] }), 
        .SouthIn({\nOut4_23[7] , \nOut4_23[6] , \nOut4_23[5] , \nOut4_23[4] , 
        \nOut4_23[3] , \nOut4_23[2] , \nOut4_23[1] , \nOut4_23[0] }), .EastIn(
        {\nOut5_22[7] , \nOut5_22[6] , \nOut5_22[5] , \nOut5_22[4] , 
        \nOut5_22[3] , \nOut5_22[2] , \nOut5_22[1] , \nOut5_22[0] }), .WestIn(
        {\nOut3_22[7] , \nOut3_22[6] , \nOut3_22[5] , \nOut3_22[4] , 
        \nOut3_22[3] , \nOut3_22[2] , \nOut3_22[1] , \nOut3_22[0] }), .Out({
        \nOut4_22[7] , \nOut4_22[6] , \nOut4_22[5] , \nOut4_22[4] , 
        \nOut4_22[3] , \nOut4_22[2] , \nOut4_22[1] , \nOut4_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_177 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut178[7] , \nScanOut178[6] , 
        \nScanOut178[5] , \nScanOut178[4] , \nScanOut178[3] , \nScanOut178[2] , 
        \nScanOut178[1] , \nScanOut178[0] }), .ScanOut({\nScanOut177[7] , 
        \nScanOut177[6] , \nScanOut177[5] , \nScanOut177[4] , \nScanOut177[3] , 
        \nScanOut177[2] , \nScanOut177[1] , \nScanOut177[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_16[7] , \nOut5_16[6] , \nOut5_16[5] , \nOut5_16[4] , 
        \nOut5_16[3] , \nOut5_16[2] , \nOut5_16[1] , \nOut5_16[0] }), 
        .SouthIn({\nOut5_18[7] , \nOut5_18[6] , \nOut5_18[5] , \nOut5_18[4] , 
        \nOut5_18[3] , \nOut5_18[2] , \nOut5_18[1] , \nOut5_18[0] }), .EastIn(
        {\nOut6_17[7] , \nOut6_17[6] , \nOut6_17[5] , \nOut6_17[4] , 
        \nOut6_17[3] , \nOut6_17[2] , \nOut6_17[1] , \nOut6_17[0] }), .WestIn(
        {\nOut4_17[7] , \nOut4_17[6] , \nOut4_17[5] , \nOut4_17[4] , 
        \nOut4_17[3] , \nOut4_17[2] , \nOut4_17[1] , \nOut4_17[0] }), .Out({
        \nOut5_17[7] , \nOut5_17[6] , \nOut5_17[5] , \nOut5_17[4] , 
        \nOut5_17[3] , \nOut5_17[2] , \nOut5_17[1] , \nOut5_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_247 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut248[7] , \nScanOut248[6] , 
        \nScanOut248[5] , \nScanOut248[4] , \nScanOut248[3] , \nScanOut248[2] , 
        \nScanOut248[1] , \nScanOut248[0] }), .ScanOut({\nScanOut247[7] , 
        \nScanOut247[6] , \nScanOut247[5] , \nScanOut247[4] , \nScanOut247[3] , 
        \nScanOut247[2] , \nScanOut247[1] , \nScanOut247[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_22[7] , \nOut7_22[6] , \nOut7_22[5] , \nOut7_22[4] , 
        \nOut7_22[3] , \nOut7_22[2] , \nOut7_22[1] , \nOut7_22[0] }), 
        .SouthIn({\nOut7_24[7] , \nOut7_24[6] , \nOut7_24[5] , \nOut7_24[4] , 
        \nOut7_24[3] , \nOut7_24[2] , \nOut7_24[1] , \nOut7_24[0] }), .EastIn(
        {\nOut8_23[7] , \nOut8_23[6] , \nOut8_23[5] , \nOut8_23[4] , 
        \nOut8_23[3] , \nOut8_23[2] , \nOut8_23[1] , \nOut8_23[0] }), .WestIn(
        {\nOut6_23[7] , \nOut6_23[6] , \nOut6_23[5] , \nOut6_23[4] , 
        \nOut6_23[3] , \nOut6_23[2] , \nOut6_23[1] , \nOut6_23[0] }), .Out({
        \nOut7_23[7] , \nOut7_23[6] , \nOut7_23[5] , \nOut7_23[4] , 
        \nOut7_23[3] , \nOut7_23[2] , \nOut7_23[1] , \nOut7_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_347 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut348[7] , \nScanOut348[6] , 
        \nScanOut348[5] , \nScanOut348[4] , \nScanOut348[3] , \nScanOut348[2] , 
        \nScanOut348[1] , \nScanOut348[0] }), .ScanOut({\nScanOut347[7] , 
        \nScanOut347[6] , \nScanOut347[5] , \nScanOut347[4] , \nScanOut347[3] , 
        \nScanOut347[2] , \nScanOut347[1] , \nScanOut347[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_26[7] , \nOut10_26[6] , \nOut10_26[5] , \nOut10_26[4] , 
        \nOut10_26[3] , \nOut10_26[2] , \nOut10_26[1] , \nOut10_26[0] }), 
        .SouthIn({\nOut10_28[7] , \nOut10_28[6] , \nOut10_28[5] , 
        \nOut10_28[4] , \nOut10_28[3] , \nOut10_28[2] , \nOut10_28[1] , 
        \nOut10_28[0] }), .EastIn({\nOut11_27[7] , \nOut11_27[6] , 
        \nOut11_27[5] , \nOut11_27[4] , \nOut11_27[3] , \nOut11_27[2] , 
        \nOut11_27[1] , \nOut11_27[0] }), .WestIn({\nOut9_27[7] , 
        \nOut9_27[6] , \nOut9_27[5] , \nOut9_27[4] , \nOut9_27[3] , 
        \nOut9_27[2] , \nOut9_27[1] , \nOut9_27[0] }), .Out({\nOut10_27[7] , 
        \nOut10_27[6] , \nOut10_27[5] , \nOut10_27[4] , \nOut10_27[3] , 
        \nOut10_27[2] , \nOut10_27[1] , \nOut10_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_556 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut557[7] , \nScanOut557[6] , 
        \nScanOut557[5] , \nScanOut557[4] , \nScanOut557[3] , \nScanOut557[2] , 
        \nScanOut557[1] , \nScanOut557[0] }), .ScanOut({\nScanOut556[7] , 
        \nScanOut556[6] , \nScanOut556[5] , \nScanOut556[4] , \nScanOut556[3] , 
        \nScanOut556[2] , \nScanOut556[1] , \nScanOut556[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_11[7] , \nOut17_11[6] , \nOut17_11[5] , \nOut17_11[4] , 
        \nOut17_11[3] , \nOut17_11[2] , \nOut17_11[1] , \nOut17_11[0] }), 
        .SouthIn({\nOut17_13[7] , \nOut17_13[6] , \nOut17_13[5] , 
        \nOut17_13[4] , \nOut17_13[3] , \nOut17_13[2] , \nOut17_13[1] , 
        \nOut17_13[0] }), .EastIn({\nOut18_12[7] , \nOut18_12[6] , 
        \nOut18_12[5] , \nOut18_12[4] , \nOut18_12[3] , \nOut18_12[2] , 
        \nOut18_12[1] , \nOut18_12[0] }), .WestIn({\nOut16_12[7] , 
        \nOut16_12[6] , \nOut16_12[5] , \nOut16_12[4] , \nOut16_12[3] , 
        \nOut16_12[2] , \nOut16_12[1] , \nOut16_12[0] }), .Out({\nOut17_12[7] , 
        \nOut17_12[6] , \nOut17_12[5] , \nOut17_12[4] , \nOut17_12[3] , 
        \nOut17_12[2] , \nOut17_12[1] , \nOut17_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_666 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut667[7] , \nScanOut667[6] , 
        \nScanOut667[5] , \nScanOut667[4] , \nScanOut667[3] , \nScanOut667[2] , 
        \nScanOut667[1] , \nScanOut667[0] }), .ScanOut({\nScanOut666[7] , 
        \nScanOut666[6] , \nScanOut666[5] , \nScanOut666[4] , \nScanOut666[3] , 
        \nScanOut666[2] , \nScanOut666[1] , \nScanOut666[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_25[7] , \nOut20_25[6] , \nOut20_25[5] , \nOut20_25[4] , 
        \nOut20_25[3] , \nOut20_25[2] , \nOut20_25[1] , \nOut20_25[0] }), 
        .SouthIn({\nOut20_27[7] , \nOut20_27[6] , \nOut20_27[5] , 
        \nOut20_27[4] , \nOut20_27[3] , \nOut20_27[2] , \nOut20_27[1] , 
        \nOut20_27[0] }), .EastIn({\nOut21_26[7] , \nOut21_26[6] , 
        \nOut21_26[5] , \nOut21_26[4] , \nOut21_26[3] , \nOut21_26[2] , 
        \nOut21_26[1] , \nOut21_26[0] }), .WestIn({\nOut19_26[7] , 
        \nOut19_26[6] , \nOut19_26[5] , \nOut19_26[4] , \nOut19_26[3] , 
        \nOut19_26[2] , \nOut19_26[1] , \nOut19_26[0] }), .Out({\nOut20_26[7] , 
        \nOut20_26[6] , \nOut20_26[5] , \nOut20_26[4] , \nOut20_26[3] , 
        \nOut20_26[2] , \nOut20_26[1] , \nOut20_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_818 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut819[7] , \nScanOut819[6] , 
        \nScanOut819[5] , \nScanOut819[4] , \nScanOut819[3] , \nScanOut819[2] , 
        \nScanOut819[1] , \nScanOut819[0] }), .ScanOut({\nScanOut818[7] , 
        \nScanOut818[6] , \nScanOut818[5] , \nScanOut818[4] , \nScanOut818[3] , 
        \nScanOut818[2] , \nScanOut818[1] , \nScanOut818[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_17[7] , \nOut25_17[6] , \nOut25_17[5] , \nOut25_17[4] , 
        \nOut25_17[3] , \nOut25_17[2] , \nOut25_17[1] , \nOut25_17[0] }), 
        .SouthIn({\nOut25_19[7] , \nOut25_19[6] , \nOut25_19[5] , 
        \nOut25_19[4] , \nOut25_19[3] , \nOut25_19[2] , \nOut25_19[1] , 
        \nOut25_19[0] }), .EastIn({\nOut26_18[7] , \nOut26_18[6] , 
        \nOut26_18[5] , \nOut26_18[4] , \nOut26_18[3] , \nOut26_18[2] , 
        \nOut26_18[1] , \nOut26_18[0] }), .WestIn({\nOut24_18[7] , 
        \nOut24_18[6] , \nOut24_18[5] , \nOut24_18[4] , \nOut24_18[3] , 
        \nOut24_18[2] , \nOut24_18[1] , \nOut24_18[0] }), .Out({\nOut25_18[7] , 
        \nOut25_18[6] , \nOut25_18[5] , \nOut25_18[4] , \nOut25_18[3] , 
        \nOut25_18[2] , \nOut25_18[1] , \nOut25_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_924 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut925[7] , \nScanOut925[6] , 
        \nScanOut925[5] , \nScanOut925[4] , \nScanOut925[3] , \nScanOut925[2] , 
        \nScanOut925[1] , \nScanOut925[0] }), .ScanOut({\nScanOut924[7] , 
        \nScanOut924[6] , \nScanOut924[5] , \nScanOut924[4] , \nScanOut924[3] , 
        \nScanOut924[2] , \nScanOut924[1] , \nScanOut924[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_27[7] , \nOut28_27[6] , \nOut28_27[5] , \nOut28_27[4] , 
        \nOut28_27[3] , \nOut28_27[2] , \nOut28_27[1] , \nOut28_27[0] }), 
        .SouthIn({\nOut28_29[7] , \nOut28_29[6] , \nOut28_29[5] , 
        \nOut28_29[4] , \nOut28_29[3] , \nOut28_29[2] , \nOut28_29[1] , 
        \nOut28_29[0] }), .EastIn({\nOut29_28[7] , \nOut29_28[6] , 
        \nOut29_28[5] , \nOut29_28[4] , \nOut29_28[3] , \nOut29_28[2] , 
        \nOut29_28[1] , \nOut29_28[0] }), .WestIn({\nOut27_28[7] , 
        \nOut27_28[6] , \nOut27_28[5] , \nOut27_28[4] , \nOut27_28[3] , 
        \nOut27_28[2] , \nOut27_28[1] , \nOut27_28[0] }), .Out({\nOut28_28[7] , 
        \nOut28_28[6] , \nOut28_28[5] , \nOut28_28[4] , \nOut28_28[3] , 
        \nOut28_28[2] , \nOut28_28[1] , \nOut28_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_988 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut989[7] , \nScanOut989[6] , 
        \nScanOut989[5] , \nScanOut989[4] , \nScanOut989[3] , \nScanOut989[2] , 
        \nScanOut989[1] , \nScanOut989[0] }), .ScanOut({\nScanOut988[7] , 
        \nScanOut988[6] , \nScanOut988[5] , \nScanOut988[4] , \nScanOut988[3] , 
        \nScanOut988[2] , \nScanOut988[1] , \nScanOut988[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_27[7] , \nOut30_27[6] , \nOut30_27[5] , \nOut30_27[4] , 
        \nOut30_27[3] , \nOut30_27[2] , \nOut30_27[1] , \nOut30_27[0] }), 
        .SouthIn({\nOut30_29[7] , \nOut30_29[6] , \nOut30_29[5] , 
        \nOut30_29[4] , \nOut30_29[3] , \nOut30_29[2] , \nOut30_29[1] , 
        \nOut30_29[0] }), .EastIn({\nOut31_28[7] , \nOut31_28[6] , 
        \nOut31_28[5] , \nOut31_28[4] , \nOut31_28[3] , \nOut31_28[2] , 
        \nOut31_28[1] , \nOut31_28[0] }), .WestIn({\nOut29_28[7] , 
        \nOut29_28[6] , \nOut29_28[5] , \nOut29_28[4] , \nOut29_28[3] , 
        \nOut29_28[2] , \nOut29_28[1] , \nOut29_28[0] }), .Out({\nOut30_28[7] , 
        \nOut30_28[6] , \nOut30_28[5] , \nOut30_28[4] , \nOut30_28[3] , 
        \nOut30_28[2] , \nOut30_28[1] , \nOut30_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_456 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut457[7] , \nScanOut457[6] , 
        \nScanOut457[5] , \nScanOut457[4] , \nScanOut457[3] , \nScanOut457[2] , 
        \nScanOut457[1] , \nScanOut457[0] }), .ScanOut({\nScanOut456[7] , 
        \nScanOut456[6] , \nScanOut456[5] , \nScanOut456[4] , \nScanOut456[3] , 
        \nScanOut456[2] , \nScanOut456[1] , \nScanOut456[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }), 
        .SouthIn({\nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , \nOut14_9[4] , 
        \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , \nOut14_9[0] }), .EastIn(
        {\nOut15_8[7] , \nOut15_8[6] , \nOut15_8[5] , \nOut15_8[4] , 
        \nOut15_8[3] , \nOut15_8[2] , \nOut15_8[1] , \nOut15_8[0] }), .WestIn(
        {\nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }), .Out({
        \nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_824 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut825[7] , \nScanOut825[6] , 
        \nScanOut825[5] , \nScanOut825[4] , \nScanOut825[3] , \nScanOut825[2] , 
        \nScanOut825[1] , \nScanOut825[0] }), .ScanOut({\nScanOut824[7] , 
        \nScanOut824[6] , \nScanOut824[5] , \nScanOut824[4] , \nScanOut824[3] , 
        \nScanOut824[2] , \nScanOut824[1] , \nScanOut824[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_23[7] , \nOut25_23[6] , \nOut25_23[5] , \nOut25_23[4] , 
        \nOut25_23[3] , \nOut25_23[2] , \nOut25_23[1] , \nOut25_23[0] }), 
        .SouthIn({\nOut25_25[7] , \nOut25_25[6] , \nOut25_25[5] , 
        \nOut25_25[4] , \nOut25_25[3] , \nOut25_25[2] , \nOut25_25[1] , 
        \nOut25_25[0] }), .EastIn({\nOut26_24[7] , \nOut26_24[6] , 
        \nOut26_24[5] , \nOut26_24[4] , \nOut26_24[3] , \nOut26_24[2] , 
        \nOut26_24[1] , \nOut26_24[0] }), .WestIn({\nOut24_24[7] , 
        \nOut24_24[6] , \nOut24_24[5] , \nOut24_24[4] , \nOut24_24[3] , 
        \nOut24_24[2] , \nOut24_24[1] , \nOut24_24[0] }), .Out({\nOut25_24[7] , 
        \nOut25_24[6] , \nOut25_24[5] , \nOut25_24[4] , \nOut25_24[3] , 
        \nOut25_24[2] , \nOut25_24[1] , \nOut25_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_741 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut742[7] , \nScanOut742[6] , 
        \nScanOut742[5] , \nScanOut742[4] , \nScanOut742[3] , \nScanOut742[2] , 
        \nScanOut742[1] , \nScanOut742[0] }), .ScanOut({\nScanOut741[7] , 
        \nScanOut741[6] , \nScanOut741[5] , \nScanOut741[4] , \nScanOut741[3] , 
        \nScanOut741[2] , \nScanOut741[1] , \nScanOut741[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_4[7] , \nOut23_4[6] , \nOut23_4[5] , \nOut23_4[4] , 
        \nOut23_4[3] , \nOut23_4[2] , \nOut23_4[1] , \nOut23_4[0] }), 
        .SouthIn({\nOut23_6[7] , \nOut23_6[6] , \nOut23_6[5] , \nOut23_6[4] , 
        \nOut23_6[3] , \nOut23_6[2] , \nOut23_6[1] , \nOut23_6[0] }), .EastIn(
        {\nOut24_5[7] , \nOut24_5[6] , \nOut24_5[5] , \nOut24_5[4] , 
        \nOut24_5[3] , \nOut24_5[2] , \nOut24_5[1] , \nOut24_5[0] }), .WestIn(
        {\nOut22_5[7] , \nOut22_5[6] , \nOut22_5[5] , \nOut22_5[4] , 
        \nOut22_5[3] , \nOut22_5[2] , \nOut22_5[1] , \nOut22_5[0] }), .Out({
        \nOut23_5[7] , \nOut23_5[6] , \nOut23_5[5] , \nOut23_5[4] , 
        \nOut23_5[3] , \nOut23_5[2] , \nOut23_5[1] , \nOut23_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_766 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut767[7] , \nScanOut767[6] , 
        \nScanOut767[5] , \nScanOut767[4] , \nScanOut767[3] , \nScanOut767[2] , 
        \nScanOut767[1] , \nScanOut767[0] }), .ScanOut({\nScanOut766[7] , 
        \nScanOut766[6] , \nScanOut766[5] , \nScanOut766[4] , \nScanOut766[3] , 
        \nScanOut766[2] , \nScanOut766[1] , \nScanOut766[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_29[7] , \nOut23_29[6] , \nOut23_29[5] , \nOut23_29[4] , 
        \nOut23_29[3] , \nOut23_29[2] , \nOut23_29[1] , \nOut23_29[0] }), 
        .SouthIn({\nOut23_31[7] , \nOut23_31[6] , \nOut23_31[5] , 
        \nOut23_31[4] , \nOut23_31[3] , \nOut23_31[2] , \nOut23_31[1] , 
        \nOut23_31[0] }), .EastIn({\nOut24_30[7] , \nOut24_30[6] , 
        \nOut24_30[5] , \nOut24_30[4] , \nOut24_30[3] , \nOut24_30[2] , 
        \nOut24_30[1] , \nOut24_30[0] }), .WestIn({\nOut22_30[7] , 
        \nOut22_30[6] , \nOut22_30[5] , \nOut22_30[4] , \nOut22_30[3] , 
        \nOut22_30[2] , \nOut22_30[1] , \nOut22_30[0] }), .Out({\nOut23_30[7] , 
        \nOut23_30[6] , \nOut23_30[5] , \nOut23_30[4] , \nOut23_30[3] , 
        \nOut23_30[2] , \nOut23_30[1] , \nOut23_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_260 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut261[7] , \nScanOut261[6] , 
        \nScanOut261[5] , \nScanOut261[4] , \nScanOut261[3] , \nScanOut261[2] , 
        \nScanOut261[1] , \nScanOut261[0] }), .ScanOut({\nScanOut260[7] , 
        \nScanOut260[6] , \nScanOut260[5] , \nScanOut260[4] , \nScanOut260[3] , 
        \nScanOut260[2] , \nScanOut260[1] , \nScanOut260[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_3[7] , \nOut8_3[6] , \nOut8_3[5] , \nOut8_3[4] , \nOut8_3[3] , 
        \nOut8_3[2] , \nOut8_3[1] , \nOut8_3[0] }), .SouthIn({\nOut8_5[7] , 
        \nOut8_5[6] , \nOut8_5[5] , \nOut8_5[4] , \nOut8_5[3] , \nOut8_5[2] , 
        \nOut8_5[1] , \nOut8_5[0] }), .EastIn({\nOut9_4[7] , \nOut9_4[6] , 
        \nOut9_4[5] , \nOut9_4[4] , \nOut9_4[3] , \nOut9_4[2] , \nOut9_4[1] , 
        \nOut9_4[0] }), .WestIn({\nOut7_4[7] , \nOut7_4[6] , \nOut7_4[5] , 
        \nOut7_4[4] , \nOut7_4[3] , \nOut7_4[2] , \nOut7_4[1] , \nOut7_4[0] }), 
        .Out({\nOut8_4[7] , \nOut8_4[6] , \nOut8_4[5] , \nOut8_4[4] , 
        \nOut8_4[3] , \nOut8_4[2] , \nOut8_4[1] , \nOut8_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_471 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut472[7] , \nScanOut472[6] , 
        \nScanOut472[5] , \nScanOut472[4] , \nScanOut472[3] , \nScanOut472[2] , 
        \nScanOut472[1] , \nScanOut472[0] }), .ScanOut({\nScanOut471[7] , 
        \nScanOut471[6] , \nScanOut471[5] , \nScanOut471[4] , \nScanOut471[3] , 
        \nScanOut471[2] , \nScanOut471[1] , \nScanOut471[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_22[7] , \nOut14_22[6] , \nOut14_22[5] , \nOut14_22[4] , 
        \nOut14_22[3] , \nOut14_22[2] , \nOut14_22[1] , \nOut14_22[0] }), 
        .SouthIn({\nOut14_24[7] , \nOut14_24[6] , \nOut14_24[5] , 
        \nOut14_24[4] , \nOut14_24[3] , \nOut14_24[2] , \nOut14_24[1] , 
        \nOut14_24[0] }), .EastIn({\nOut15_23[7] , \nOut15_23[6] , 
        \nOut15_23[5] , \nOut15_23[4] , \nOut15_23[3] , \nOut15_23[2] , 
        \nOut15_23[1] , \nOut15_23[0] }), .WestIn({\nOut13_23[7] , 
        \nOut13_23[6] , \nOut13_23[5] , \nOut13_23[4] , \nOut13_23[3] , 
        \nOut13_23[2] , \nOut13_23[1] , \nOut13_23[0] }), .Out({\nOut14_23[7] , 
        \nOut14_23[6] , \nOut14_23[5] , \nOut14_23[4] , \nOut14_23[3] , 
        \nOut14_23[2] , \nOut14_23[1] , \nOut14_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_803 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut804[7] , \nScanOut804[6] , 
        \nScanOut804[5] , \nScanOut804[4] , \nScanOut804[3] , \nScanOut804[2] , 
        \nScanOut804[1] , \nScanOut804[0] }), .ScanOut({\nScanOut803[7] , 
        \nScanOut803[6] , \nScanOut803[5] , \nScanOut803[4] , \nScanOut803[3] , 
        \nScanOut803[2] , \nScanOut803[1] , \nScanOut803[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_2[7] , \nOut25_2[6] , \nOut25_2[5] , \nOut25_2[4] , 
        \nOut25_2[3] , \nOut25_2[2] , \nOut25_2[1] , \nOut25_2[0] }), 
        .SouthIn({\nOut25_4[7] , \nOut25_4[6] , \nOut25_4[5] , \nOut25_4[4] , 
        \nOut25_4[3] , \nOut25_4[2] , \nOut25_4[1] , \nOut25_4[0] }), .EastIn(
        {\nOut26_3[7] , \nOut26_3[6] , \nOut26_3[5] , \nOut26_3[4] , 
        \nOut26_3[3] , \nOut26_3[2] , \nOut26_3[1] , \nOut26_3[0] }), .WestIn(
        {\nOut24_3[7] , \nOut24_3[6] , \nOut24_3[5] , \nOut24_3[4] , 
        \nOut24_3[3] , \nOut24_3[2] , \nOut24_3[1] , \nOut24_3[0] }), .Out({
        \nOut25_3[7] , \nOut25_3[6] , \nOut25_3[5] , \nOut25_3[4] , 
        \nOut25_3[3] , \nOut25_3[2] , \nOut25_3[1] , \nOut25_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_993 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut994[7] , \nScanOut994[6] , 
        \nScanOut994[5] , \nScanOut994[4] , \nScanOut994[3] , \nScanOut994[2] , 
        \nScanOut994[1] , \nScanOut994[0] }), .ScanOut({\nScanOut993[7] , 
        \nScanOut993[6] , \nScanOut993[5] , \nScanOut993[4] , \nScanOut993[3] , 
        \nScanOut993[2] , \nScanOut993[1] , \nScanOut993[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut31_1[7] , \nOut31_1[6] , 
        \nOut31_1[5] , \nOut31_1[4] , \nOut31_1[3] , \nOut31_1[2] , 
        \nOut31_1[1] , \nOut31_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_21 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut22[7] , \nScanOut22[6] , 
        \nScanOut22[5] , \nScanOut22[4] , \nScanOut22[3] , \nScanOut22[2] , 
        \nScanOut22[1] , \nScanOut22[0] }), .ScanOut({\nScanOut21[7] , 
        \nScanOut21[6] , \nScanOut21[5] , \nScanOut21[4] , \nScanOut21[3] , 
        \nScanOut21[2] , \nScanOut21[1] , \nScanOut21[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_21[7] , \nOut0_21[6] , 
        \nOut0_21[5] , \nOut0_21[4] , \nOut0_21[3] , \nOut0_21[2] , 
        \nOut0_21[1] , \nOut0_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_634 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut635[7] , \nScanOut635[6] , 
        \nScanOut635[5] , \nScanOut635[4] , \nScanOut635[3] , \nScanOut635[2] , 
        \nScanOut635[1] , \nScanOut635[0] }), .ScanOut({\nScanOut634[7] , 
        \nScanOut634[6] , \nScanOut634[5] , \nScanOut634[4] , \nScanOut634[3] , 
        \nScanOut634[2] , \nScanOut634[1] , \nScanOut634[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_25[7] , \nOut19_25[6] , \nOut19_25[5] , \nOut19_25[4] , 
        \nOut19_25[3] , \nOut19_25[2] , \nOut19_25[1] , \nOut19_25[0] }), 
        .SouthIn({\nOut19_27[7] , \nOut19_27[6] , \nOut19_27[5] , 
        \nOut19_27[4] , \nOut19_27[3] , \nOut19_27[2] , \nOut19_27[1] , 
        \nOut19_27[0] }), .EastIn({\nOut20_26[7] , \nOut20_26[6] , 
        \nOut20_26[5] , \nOut20_26[4] , \nOut20_26[3] , \nOut20_26[2] , 
        \nOut20_26[1] , \nOut20_26[0] }), .WestIn({\nOut18_26[7] , 
        \nOut18_26[6] , \nOut18_26[5] , \nOut18_26[4] , \nOut18_26[3] , 
        \nOut18_26[2] , \nOut18_26[1] , \nOut18_26[0] }), .Out({\nOut19_26[7] , 
        \nOut19_26[6] , \nOut19_26[5] , \nOut19_26[4] , \nOut19_26[3] , 
        \nOut19_26[2] , \nOut19_26[1] , \nOut19_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_888 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut889[7] , \nScanOut889[6] , 
        \nScanOut889[5] , \nScanOut889[4] , \nScanOut889[3] , \nScanOut889[2] , 
        \nScanOut889[1] , \nScanOut889[0] }), .ScanOut({\nScanOut888[7] , 
        \nScanOut888[6] , \nScanOut888[5] , \nScanOut888[4] , \nScanOut888[3] , 
        \nScanOut888[2] , \nScanOut888[1] , \nScanOut888[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_23[7] , \nOut27_23[6] , \nOut27_23[5] , \nOut27_23[4] , 
        \nOut27_23[3] , \nOut27_23[2] , \nOut27_23[1] , \nOut27_23[0] }), 
        .SouthIn({\nOut27_25[7] , \nOut27_25[6] , \nOut27_25[5] , 
        \nOut27_25[4] , \nOut27_25[3] , \nOut27_25[2] , \nOut27_25[1] , 
        \nOut27_25[0] }), .EastIn({\nOut28_24[7] , \nOut28_24[6] , 
        \nOut28_24[5] , \nOut28_24[4] , \nOut28_24[3] , \nOut28_24[2] , 
        \nOut28_24[1] , \nOut28_24[0] }), .WestIn({\nOut26_24[7] , 
        \nOut26_24[6] , \nOut26_24[5] , \nOut26_24[4] , \nOut26_24[3] , 
        \nOut26_24[2] , \nOut26_24[1] , \nOut26_24[0] }), .Out({\nOut27_24[7] , 
        \nOut27_24[6] , \nOut27_24[5] , \nOut27_24[4] , \nOut27_24[3] , 
        \nOut27_24[2] , \nOut27_24[1] , \nOut27_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_918 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut919[7] , \nScanOut919[6] , 
        \nScanOut919[5] , \nScanOut919[4] , \nScanOut919[3] , \nScanOut919[2] , 
        \nScanOut919[1] , \nScanOut919[0] }), .ScanOut({\nScanOut918[7] , 
        \nScanOut918[6] , \nScanOut918[5] , \nScanOut918[4] , \nScanOut918[3] , 
        \nScanOut918[2] , \nScanOut918[1] , \nScanOut918[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_21[7] , \nOut28_21[6] , \nOut28_21[5] , \nOut28_21[4] , 
        \nOut28_21[3] , \nOut28_21[2] , \nOut28_21[1] , \nOut28_21[0] }), 
        .SouthIn({\nOut28_23[7] , \nOut28_23[6] , \nOut28_23[5] , 
        \nOut28_23[4] , \nOut28_23[3] , \nOut28_23[2] , \nOut28_23[1] , 
        \nOut28_23[0] }), .EastIn({\nOut29_22[7] , \nOut29_22[6] , 
        \nOut29_22[5] , \nOut29_22[4] , \nOut29_22[3] , \nOut29_22[2] , 
        \nOut29_22[1] , \nOut29_22[0] }), .WestIn({\nOut27_22[7] , 
        \nOut27_22[6] , \nOut27_22[5] , \nOut27_22[4] , \nOut27_22[3] , 
        \nOut27_22[2] , \nOut27_22[1] , \nOut27_22[0] }), .Out({\nOut28_22[7] , 
        \nOut28_22[6] , \nOut28_22[5] , \nOut28_22[4] , \nOut28_22[3] , 
        \nOut28_22[2] , \nOut28_22[1] , \nOut28_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_29 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut30[7] , \nScanOut30[6] , 
        \nScanOut30[5] , \nScanOut30[4] , \nScanOut30[3] , \nScanOut30[2] , 
        \nScanOut30[1] , \nScanOut30[0] }), .ScanOut({\nScanOut29[7] , 
        \nScanOut29[6] , \nScanOut29[5] , \nScanOut29[4] , \nScanOut29[3] , 
        \nScanOut29[2] , \nScanOut29[1] , \nScanOut29[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_29[7] , \nOut0_29[6] , 
        \nOut0_29[5] , \nOut0_29[4] , \nOut0_29[3] , \nOut0_29[2] , 
        \nOut0_29[1] , \nOut0_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_119 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut120[7] , \nScanOut120[6] , 
        \nScanOut120[5] , \nScanOut120[4] , \nScanOut120[3] , \nScanOut120[2] , 
        \nScanOut120[1] , \nScanOut120[0] }), .ScanOut({\nScanOut119[7] , 
        \nScanOut119[6] , \nScanOut119[5] , \nScanOut119[4] , \nScanOut119[3] , 
        \nScanOut119[2] , \nScanOut119[1] , \nScanOut119[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_22[7] , \nOut3_22[6] , \nOut3_22[5] , \nOut3_22[4] , 
        \nOut3_22[3] , \nOut3_22[2] , \nOut3_22[1] , \nOut3_22[0] }), 
        .SouthIn({\nOut3_24[7] , \nOut3_24[6] , \nOut3_24[5] , \nOut3_24[4] , 
        \nOut3_24[3] , \nOut3_24[2] , \nOut3_24[1] , \nOut3_24[0] }), .EastIn(
        {\nOut4_23[7] , \nOut4_23[6] , \nOut4_23[5] , \nOut4_23[4] , 
        \nOut4_23[3] , \nOut4_23[2] , \nOut4_23[1] , \nOut4_23[0] }), .WestIn(
        {\nOut2_23[7] , \nOut2_23[6] , \nOut2_23[5] , \nOut2_23[4] , 
        \nOut2_23[3] , \nOut2_23[2] , \nOut2_23[1] , \nOut2_23[0] }), .Out({
        \nOut3_23[7] , \nOut3_23[6] , \nOut3_23[5] , \nOut3_23[4] , 
        \nOut3_23[3] , \nOut3_23[2] , \nOut3_23[1] , \nOut3_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_192 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut193[7] , \nScanOut193[6] , 
        \nScanOut193[5] , \nScanOut193[4] , \nScanOut193[3] , \nScanOut193[2] , 
        \nScanOut193[1] , \nScanOut193[0] }), .ScanOut({\nScanOut192[7] , 
        \nScanOut192[6] , \nScanOut192[5] , \nScanOut192[4] , \nScanOut192[3] , 
        \nScanOut192[2] , \nScanOut192[1] , \nScanOut192[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut6_0[7] , \nOut6_0[6] , 
        \nOut6_0[5] , \nOut6_0[4] , \nOut6_0[3] , \nOut6_0[2] , \nOut6_0[1] , 
        \nOut6_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_285 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut286[7] , \nScanOut286[6] , 
        \nScanOut286[5] , \nScanOut286[4] , \nScanOut286[3] , \nScanOut286[2] , 
        \nScanOut286[1] , \nScanOut286[0] }), .ScanOut({\nScanOut285[7] , 
        \nScanOut285[6] , \nScanOut285[5] , \nScanOut285[4] , \nScanOut285[3] , 
        \nScanOut285[2] , \nScanOut285[1] , \nScanOut285[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_28[7] , \nOut8_28[6] , \nOut8_28[5] , \nOut8_28[4] , 
        \nOut8_28[3] , \nOut8_28[2] , \nOut8_28[1] , \nOut8_28[0] }), 
        .SouthIn({\nOut8_30[7] , \nOut8_30[6] , \nOut8_30[5] , \nOut8_30[4] , 
        \nOut8_30[3] , \nOut8_30[2] , \nOut8_30[1] , \nOut8_30[0] }), .EastIn(
        {\nOut9_29[7] , \nOut9_29[6] , \nOut9_29[5] , \nOut9_29[4] , 
        \nOut9_29[3] , \nOut9_29[2] , \nOut9_29[1] , \nOut9_29[0] }), .WestIn(
        {\nOut7_29[7] , \nOut7_29[6] , \nOut7_29[5] , \nOut7_29[4] , 
        \nOut7_29[3] , \nOut7_29[2] , \nOut7_29[1] , \nOut7_29[0] }), .Out({
        \nOut8_29[7] , \nOut8_29[6] , \nOut8_29[5] , \nOut8_29[4] , 
        \nOut8_29[3] , \nOut8_29[2] , \nOut8_29[1] , \nOut8_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_504 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut505[7] , \nScanOut505[6] , 
        \nScanOut505[5] , \nScanOut505[4] , \nScanOut505[3] , \nScanOut505[2] , 
        \nScanOut505[1] , \nScanOut505[0] }), .ScanOut({\nScanOut504[7] , 
        \nScanOut504[6] , \nScanOut504[5] , \nScanOut504[4] , \nScanOut504[3] , 
        \nScanOut504[2] , \nScanOut504[1] , \nScanOut504[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_23[7] , \nOut15_23[6] , \nOut15_23[5] , \nOut15_23[4] , 
        \nOut15_23[3] , \nOut15_23[2] , \nOut15_23[1] , \nOut15_23[0] }), 
        .SouthIn({\nOut15_25[7] , \nOut15_25[6] , \nOut15_25[5] , 
        \nOut15_25[4] , \nOut15_25[3] , \nOut15_25[2] , \nOut15_25[1] , 
        \nOut15_25[0] }), .EastIn({\nOut16_24[7] , \nOut16_24[6] , 
        \nOut16_24[5] , \nOut16_24[4] , \nOut16_24[3] , \nOut16_24[2] , 
        \nOut16_24[1] , \nOut16_24[0] }), .WestIn({\nOut14_24[7] , 
        \nOut14_24[6] , \nOut14_24[5] , \nOut14_24[4] , \nOut14_24[3] , 
        \nOut14_24[2] , \nOut14_24[1] , \nOut14_24[0] }), .Out({\nOut15_24[7] , 
        \nOut15_24[6] , \nOut15_24[5] , \nOut15_24[4] , \nOut15_24[3] , 
        \nOut15_24[2] , \nOut15_24[1] , \nOut15_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_315 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut316[7] , \nScanOut316[6] , 
        \nScanOut316[5] , \nScanOut316[4] , \nScanOut316[3] , \nScanOut316[2] , 
        \nScanOut316[1] , \nScanOut316[0] }), .ScanOut({\nScanOut315[7] , 
        \nScanOut315[6] , \nScanOut315[5] , \nScanOut315[4] , \nScanOut315[3] , 
        \nScanOut315[2] , \nScanOut315[1] , \nScanOut315[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_26[7] , \nOut9_26[6] , \nOut9_26[5] , \nOut9_26[4] , 
        \nOut9_26[3] , \nOut9_26[2] , \nOut9_26[1] , \nOut9_26[0] }), 
        .SouthIn({\nOut9_28[7] , \nOut9_28[6] , \nOut9_28[5] , \nOut9_28[4] , 
        \nOut9_28[3] , \nOut9_28[2] , \nOut9_28[1] , \nOut9_28[0] }), .EastIn(
        {\nOut10_27[7] , \nOut10_27[6] , \nOut10_27[5] , \nOut10_27[4] , 
        \nOut10_27[3] , \nOut10_27[2] , \nOut10_27[1] , \nOut10_27[0] }), 
        .WestIn({\nOut8_27[7] , \nOut8_27[6] , \nOut8_27[5] , \nOut8_27[4] , 
        \nOut8_27[3] , \nOut8_27[2] , \nOut8_27[1] , \nOut8_27[0] }), .Out({
        \nOut9_27[7] , \nOut9_27[6] , \nOut9_27[5] , \nOut9_27[4] , 
        \nOut9_27[3] , \nOut9_27[2] , \nOut9_27[1] , \nOut9_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_494 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut495[7] , \nScanOut495[6] , 
        \nScanOut495[5] , \nScanOut495[4] , \nScanOut495[3] , \nScanOut495[2] , 
        \nScanOut495[1] , \nScanOut495[0] }), .ScanOut({\nScanOut494[7] , 
        \nScanOut494[6] , \nScanOut494[5] , \nScanOut494[4] , \nScanOut494[3] , 
        \nScanOut494[2] , \nScanOut494[1] , \nScanOut494[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_13[7] , \nOut15_13[6] , \nOut15_13[5] , \nOut15_13[4] , 
        \nOut15_13[3] , \nOut15_13[2] , \nOut15_13[1] , \nOut15_13[0] }), 
        .SouthIn({\nOut15_15[7] , \nOut15_15[6] , \nOut15_15[5] , 
        \nOut15_15[4] , \nOut15_15[3] , \nOut15_15[2] , \nOut15_15[1] , 
        \nOut15_15[0] }), .EastIn({\nOut16_14[7] , \nOut16_14[6] , 
        \nOut16_14[5] , \nOut16_14[4] , \nOut16_14[3] , \nOut16_14[2] , 
        \nOut16_14[1] , \nOut16_14[0] }), .WestIn({\nOut14_14[7] , 
        \nOut14_14[6] , \nOut14_14[5] , \nOut14_14[4] , \nOut14_14[3] , 
        \nOut14_14[2] , \nOut14_14[1] , \nOut14_14[0] }), .Out({\nOut15_14[7] , 
        \nOut15_14[6] , \nOut15_14[5] , \nOut15_14[4] , \nOut15_14[3] , 
        \nOut15_14[2] , \nOut15_14[1] , \nOut15_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_332 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut333[7] , \nScanOut333[6] , 
        \nScanOut333[5] , \nScanOut333[4] , \nScanOut333[3] , \nScanOut333[2] , 
        \nScanOut333[1] , \nScanOut333[0] }), .ScanOut({\nScanOut332[7] , 
        \nScanOut332[6] , \nScanOut332[5] , \nScanOut332[4] , \nScanOut332[3] , 
        \nScanOut332[2] , \nScanOut332[1] , \nScanOut332[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_11[7] , \nOut10_11[6] , \nOut10_11[5] , \nOut10_11[4] , 
        \nOut10_11[3] , \nOut10_11[2] , \nOut10_11[1] , \nOut10_11[0] }), 
        .SouthIn({\nOut10_13[7] , \nOut10_13[6] , \nOut10_13[5] , 
        \nOut10_13[4] , \nOut10_13[3] , \nOut10_13[2] , \nOut10_13[1] , 
        \nOut10_13[0] }), .EastIn({\nOut11_12[7] , \nOut11_12[6] , 
        \nOut11_12[5] , \nOut11_12[4] , \nOut11_12[3] , \nOut11_12[2] , 
        \nOut11_12[1] , \nOut11_12[0] }), .WestIn({\nOut9_12[7] , 
        \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , \nOut9_12[3] , 
        \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }), .Out({\nOut10_12[7] , 
        \nOut10_12[6] , \nOut10_12[5] , \nOut10_12[4] , \nOut10_12[3] , 
        \nOut10_12[2] , \nOut10_12[1] , \nOut10_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_976 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut977[7] , \nScanOut977[6] , 
        \nScanOut977[5] , \nScanOut977[4] , \nScanOut977[3] , \nScanOut977[2] , 
        \nScanOut977[1] , \nScanOut977[0] }), .ScanOut({\nScanOut976[7] , 
        \nScanOut976[6] , \nScanOut976[5] , \nScanOut976[4] , \nScanOut976[3] , 
        \nScanOut976[2] , \nScanOut976[1] , \nScanOut976[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_15[7] , \nOut30_15[6] , \nOut30_15[5] , \nOut30_15[4] , 
        \nOut30_15[3] , \nOut30_15[2] , \nOut30_15[1] , \nOut30_15[0] }), 
        .SouthIn({\nOut30_17[7] , \nOut30_17[6] , \nOut30_17[5] , 
        \nOut30_17[4] , \nOut30_17[3] , \nOut30_17[2] , \nOut30_17[1] , 
        \nOut30_17[0] }), .EastIn({\nOut31_16[7] , \nOut31_16[6] , 
        \nOut31_16[5] , \nOut31_16[4] , \nOut31_16[3] , \nOut31_16[2] , 
        \nOut31_16[1] , \nOut31_16[0] }), .WestIn({\nOut29_16[7] , 
        \nOut29_16[6] , \nOut29_16[5] , \nOut29_16[4] , \nOut29_16[3] , 
        \nOut29_16[2] , \nOut29_16[1] , \nOut29_16[0] }), .Out({\nOut30_16[7] , 
        \nOut30_16[6] , \nOut30_16[5] , \nOut30_16[4] , \nOut30_16[3] , 
        \nOut30_16[2] , \nOut30_16[1] , \nOut30_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_523 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut524[7] , \nScanOut524[6] , 
        \nScanOut524[5] , \nScanOut524[4] , \nScanOut524[3] , \nScanOut524[2] , 
        \nScanOut524[1] , \nScanOut524[0] }), .ScanOut({\nScanOut523[7] , 
        \nScanOut523[6] , \nScanOut523[5] , \nScanOut523[4] , \nScanOut523[3] , 
        \nScanOut523[2] , \nScanOut523[1] , \nScanOut523[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_10[7] , \nOut16_10[6] , \nOut16_10[5] , \nOut16_10[4] , 
        \nOut16_10[3] , \nOut16_10[2] , \nOut16_10[1] , \nOut16_10[0] }), 
        .SouthIn({\nOut16_12[7] , \nOut16_12[6] , \nOut16_12[5] , 
        \nOut16_12[4] , \nOut16_12[3] , \nOut16_12[2] , \nOut16_12[1] , 
        \nOut16_12[0] }), .EastIn({\nOut17_11[7] , \nOut17_11[6] , 
        \nOut17_11[5] , \nOut17_11[4] , \nOut17_11[3] , \nOut17_11[2] , 
        \nOut17_11[1] , \nOut17_11[0] }), .WestIn({\nOut15_11[7] , 
        \nOut15_11[6] , \nOut15_11[5] , \nOut15_11[4] , \nOut15_11[3] , 
        \nOut15_11[2] , \nOut15_11[1] , \nOut15_11[0] }), .Out({\nOut16_11[7] , 
        \nOut16_11[6] , \nOut16_11[5] , \nOut16_11[4] , \nOut16_11[3] , 
        \nOut16_11[2] , \nOut16_11[1] , \nOut16_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_783 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut784[7] , \nScanOut784[6] , 
        \nScanOut784[5] , \nScanOut784[4] , \nScanOut784[3] , \nScanOut784[2] , 
        \nScanOut784[1] , \nScanOut784[0] }), .ScanOut({\nScanOut783[7] , 
        \nScanOut783[6] , \nScanOut783[5] , \nScanOut783[4] , \nScanOut783[3] , 
        \nScanOut783[2] , \nScanOut783[1] , \nScanOut783[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_14[7] , \nOut24_14[6] , \nOut24_14[5] , \nOut24_14[4] , 
        \nOut24_14[3] , \nOut24_14[2] , \nOut24_14[1] , \nOut24_14[0] }), 
        .SouthIn({\nOut24_16[7] , \nOut24_16[6] , \nOut24_16[5] , 
        \nOut24_16[4] , \nOut24_16[3] , \nOut24_16[2] , \nOut24_16[1] , 
        \nOut24_16[0] }), .EastIn({\nOut25_15[7] , \nOut25_15[6] , 
        \nOut25_15[5] , \nOut25_15[4] , \nOut25_15[3] , \nOut25_15[2] , 
        \nOut25_15[1] , \nOut25_15[0] }), .WestIn({\nOut23_15[7] , 
        \nOut23_15[6] , \nOut23_15[5] , \nOut23_15[4] , \nOut23_15[3] , 
        \nOut23_15[2] , \nOut23_15[1] , \nOut23_15[0] }), .Out({\nOut24_15[7] , 
        \nOut24_15[6] , \nOut24_15[5] , \nOut24_15[4] , \nOut24_15[3] , 
        \nOut24_15[2] , \nOut24_15[1] , \nOut24_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_951 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut952[7] , \nScanOut952[6] , 
        \nScanOut952[5] , \nScanOut952[4] , \nScanOut952[3] , \nScanOut952[2] , 
        \nScanOut952[1] , \nScanOut952[0] }), .ScanOut({\nScanOut951[7] , 
        \nScanOut951[6] , \nScanOut951[5] , \nScanOut951[4] , \nScanOut951[3] , 
        \nScanOut951[2] , \nScanOut951[1] , \nScanOut951[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_22[7] , \nOut29_22[6] , \nOut29_22[5] , \nOut29_22[4] , 
        \nOut29_22[3] , \nOut29_22[2] , \nOut29_22[1] , \nOut29_22[0] }), 
        .SouthIn({\nOut29_24[7] , \nOut29_24[6] , \nOut29_24[5] , 
        \nOut29_24[4] , \nOut29_24[3] , \nOut29_24[2] , \nOut29_24[1] , 
        \nOut29_24[0] }), .EastIn({\nOut30_23[7] , \nOut30_23[6] , 
        \nOut30_23[5] , \nOut30_23[4] , \nOut30_23[3] , \nOut30_23[2] , 
        \nOut30_23[1] , \nOut30_23[0] }), .WestIn({\nOut28_23[7] , 
        \nOut28_23[6] , \nOut28_23[5] , \nOut28_23[4] , \nOut28_23[3] , 
        \nOut28_23[2] , \nOut28_23[1] , \nOut28_23[0] }), .Out({\nOut29_23[7] , 
        \nOut29_23[6] , \nOut29_23[5] , \nOut29_23[4] , \nOut29_23[3] , 
        \nOut29_23[2] , \nOut29_23[1] , \nOut29_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_229 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut230[7] , \nScanOut230[6] , 
        \nScanOut230[5] , \nScanOut230[4] , \nScanOut230[3] , \nScanOut230[2] , 
        \nScanOut230[1] , \nScanOut230[0] }), .ScanOut({\nScanOut229[7] , 
        \nScanOut229[6] , \nScanOut229[5] , \nScanOut229[4] , \nScanOut229[3] , 
        \nScanOut229[2] , \nScanOut229[1] , \nScanOut229[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_4[7] , \nOut7_4[6] , \nOut7_4[5] , \nOut7_4[4] , \nOut7_4[3] , 
        \nOut7_4[2] , \nOut7_4[1] , \nOut7_4[0] }), .SouthIn({\nOut7_6[7] , 
        \nOut7_6[6] , \nOut7_6[5] , \nOut7_6[4] , \nOut7_6[3] , \nOut7_6[2] , 
        \nOut7_6[1] , \nOut7_6[0] }), .EastIn({\nOut8_5[7] , \nOut8_5[6] , 
        \nOut8_5[5] , \nOut8_5[4] , \nOut8_5[3] , \nOut8_5[2] , \nOut8_5[1] , 
        \nOut8_5[0] }), .WestIn({\nOut6_5[7] , \nOut6_5[6] , \nOut6_5[5] , 
        \nOut6_5[4] , \nOut6_5[3] , \nOut6_5[2] , \nOut6_5[1] , \nOut6_5[0] }), 
        .Out({\nOut7_5[7] , \nOut7_5[6] , \nOut7_5[5] , \nOut7_5[4] , 
        \nOut7_5[3] , \nOut7_5[2] , \nOut7_5[1] , \nOut7_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_438 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut439[7] , \nScanOut439[6] , 
        \nScanOut439[5] , \nScanOut439[4] , \nScanOut439[3] , \nScanOut439[2] , 
        \nScanOut439[1] , \nScanOut439[0] }), .ScanOut({\nScanOut438[7] , 
        \nScanOut438[6] , \nScanOut438[5] , \nScanOut438[4] , \nScanOut438[3] , 
        \nScanOut438[2] , \nScanOut438[1] , \nScanOut438[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_21[7] , \nOut13_21[6] , \nOut13_21[5] , \nOut13_21[4] , 
        \nOut13_21[3] , \nOut13_21[2] , \nOut13_21[1] , \nOut13_21[0] }), 
        .SouthIn({\nOut13_23[7] , \nOut13_23[6] , \nOut13_23[5] , 
        \nOut13_23[4] , \nOut13_23[3] , \nOut13_23[2] , \nOut13_23[1] , 
        \nOut13_23[0] }), .EastIn({\nOut14_22[7] , \nOut14_22[6] , 
        \nOut14_22[5] , \nOut14_22[4] , \nOut14_22[3] , \nOut14_22[2] , 
        \nOut14_22[1] , \nOut14_22[0] }), .WestIn({\nOut12_22[7] , 
        \nOut12_22[6] , \nOut12_22[5] , \nOut12_22[4] , \nOut12_22[3] , 
        \nOut12_22[2] , \nOut12_22[1] , \nOut12_22[0] }), .Out({\nOut13_22[7] , 
        \nOut13_22[6] , \nOut13_22[5] , \nOut13_22[4] , \nOut13_22[3] , 
        \nOut13_22[2] , \nOut13_22[1] , \nOut13_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_613 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut614[7] , \nScanOut614[6] , 
        \nScanOut614[5] , \nScanOut614[4] , \nScanOut614[3] , \nScanOut614[2] , 
        \nScanOut614[1] , \nScanOut614[0] }), .ScanOut({\nScanOut613[7] , 
        \nScanOut613[6] , \nScanOut613[5] , \nScanOut613[4] , \nScanOut613[3] , 
        \nScanOut613[2] , \nScanOut613[1] , \nScanOut613[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_4[7] , \nOut19_4[6] , \nOut19_4[5] , \nOut19_4[4] , 
        \nOut19_4[3] , \nOut19_4[2] , \nOut19_4[1] , \nOut19_4[0] }), 
        .SouthIn({\nOut19_6[7] , \nOut19_6[6] , \nOut19_6[5] , \nOut19_6[4] , 
        \nOut19_6[3] , \nOut19_6[2] , \nOut19_6[1] , \nOut19_6[0] }), .EastIn(
        {\nOut20_5[7] , \nOut20_5[6] , \nOut20_5[5] , \nOut20_5[4] , 
        \nOut20_5[3] , \nOut20_5[2] , \nOut20_5[1] , \nOut20_5[0] }), .WestIn(
        {\nOut18_5[7] , \nOut18_5[6] , \nOut18_5[5] , \nOut18_5[4] , 
        \nOut18_5[3] , \nOut18_5[2] , \nOut18_5[1] , \nOut18_5[0] }), .Out({
        \nOut19_5[7] , \nOut19_5[6] , \nOut19_5[5] , \nOut19_5[4] , 
        \nOut19_5[3] , \nOut19_5[2] , \nOut19_5[1] , \nOut19_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_708 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut709[7] , \nScanOut709[6] , 
        \nScanOut709[5] , \nScanOut709[4] , \nScanOut709[3] , \nScanOut709[2] , 
        \nScanOut709[1] , \nScanOut709[0] }), .ScanOut({\nScanOut708[7] , 
        \nScanOut708[6] , \nScanOut708[5] , \nScanOut708[4] , \nScanOut708[3] , 
        \nScanOut708[2] , \nScanOut708[1] , \nScanOut708[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_3[7] , \nOut22_3[6] , \nOut22_3[5] , \nOut22_3[4] , 
        \nOut22_3[3] , \nOut22_3[2] , \nOut22_3[1] , \nOut22_3[0] }), 
        .SouthIn({\nOut22_5[7] , \nOut22_5[6] , \nOut22_5[5] , \nOut22_5[4] , 
        \nOut22_5[3] , \nOut22_5[2] , \nOut22_5[1] , \nOut22_5[0] }), .EastIn(
        {\nOut23_4[7] , \nOut23_4[6] , \nOut23_4[5] , \nOut23_4[4] , 
        \nOut23_4[3] , \nOut23_4[2] , \nOut23_4[1] , \nOut23_4[0] }), .WestIn(
        {\nOut21_4[7] , \nOut21_4[6] , \nOut21_4[5] , \nOut21_4[4] , 
        \nOut21_4[3] , \nOut21_4[2] , \nOut21_4[1] , \nOut21_4[0] }), .Out({
        \nOut22_4[7] , \nOut22_4[6] , \nOut22_4[5] , \nOut22_4[4] , 
        \nOut22_4[3] , \nOut22_4[2] , \nOut22_4[1] , \nOut22_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_698 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut699[7] , \nScanOut699[6] , 
        \nScanOut699[5] , \nScanOut699[4] , \nScanOut699[3] , \nScanOut699[2] , 
        \nScanOut699[1] , \nScanOut699[0] }), .ScanOut({\nScanOut698[7] , 
        \nScanOut698[6] , \nScanOut698[5] , \nScanOut698[4] , \nScanOut698[3] , 
        \nScanOut698[2] , \nScanOut698[1] , \nScanOut698[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_25[7] , \nOut21_25[6] , \nOut21_25[5] , \nOut21_25[4] , 
        \nOut21_25[3] , \nOut21_25[2] , \nOut21_25[1] , \nOut21_25[0] }), 
        .SouthIn({\nOut21_27[7] , \nOut21_27[6] , \nOut21_27[5] , 
        \nOut21_27[4] , \nOut21_27[3] , \nOut21_27[2] , \nOut21_27[1] , 
        \nOut21_27[0] }), .EastIn({\nOut22_26[7] , \nOut22_26[6] , 
        \nOut22_26[5] , \nOut22_26[4] , \nOut22_26[3] , \nOut22_26[2] , 
        \nOut22_26[1] , \nOut22_26[0] }), .WestIn({\nOut20_26[7] , 
        \nOut20_26[6] , \nOut20_26[5] , \nOut20_26[4] , \nOut20_26[3] , 
        \nOut20_26[2] , \nOut20_26[1] , \nOut20_26[0] }), .Out({\nOut21_26[7] , 
        \nOut21_26[6] , \nOut21_26[5] , \nOut21_26[4] , \nOut21_26[3] , 
        \nOut21_26[2] , \nOut21_26[1] , \nOut21_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_959 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut960[7] , \nScanOut960[6] , 
        \nScanOut960[5] , \nScanOut960[4] , \nScanOut960[3] , \nScanOut960[2] , 
        \nScanOut960[1] , \nScanOut960[0] }), .ScanOut({\nScanOut959[7] , 
        \nScanOut959[6] , \nScanOut959[5] , \nScanOut959[4] , \nScanOut959[3] , 
        \nScanOut959[2] , \nScanOut959[1] , \nScanOut959[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut29_31[7] , \nOut29_31[6] , 
        \nOut29_31[5] , \nOut29_31[4] , \nOut29_31[3] , \nOut29_31[2] , 
        \nOut29_31[1] , \nOut29_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_85 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut86[7] , \nScanOut86[6] , 
        \nScanOut86[5] , \nScanOut86[4] , \nScanOut86[3] , \nScanOut86[2] , 
        \nScanOut86[1] , \nScanOut86[0] }), .ScanOut({\nScanOut85[7] , 
        \nScanOut85[6] , \nScanOut85[5] , \nScanOut85[4] , \nScanOut85[3] , 
        \nScanOut85[2] , \nScanOut85[1] , \nScanOut85[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_20[7] , \nOut2_20[6] , \nOut2_20[5] , \nOut2_20[4] , 
        \nOut2_20[3] , \nOut2_20[2] , \nOut2_20[1] , \nOut2_20[0] }), 
        .SouthIn({\nOut2_22[7] , \nOut2_22[6] , \nOut2_22[5] , \nOut2_22[4] , 
        \nOut2_22[3] , \nOut2_22[2] , \nOut2_22[1] , \nOut2_22[0] }), .EastIn(
        {\nOut3_21[7] , \nOut3_21[6] , \nOut3_21[5] , \nOut3_21[4] , 
        \nOut3_21[3] , \nOut3_21[2] , \nOut3_21[1] , \nOut3_21[0] }), .WestIn(
        {\nOut1_21[7] , \nOut1_21[6] , \nOut1_21[5] , \nOut1_21[4] , 
        \nOut1_21[3] , \nOut1_21[2] , \nOut1_21[1] , \nOut1_21[0] }), .Out({
        \nOut2_21[7] , \nOut2_21[6] , \nOut2_21[5] , \nOut2_21[4] , 
        \nOut2_21[3] , \nOut2_21[2] , \nOut2_21[1] , \nOut2_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_111 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut112[7] , \nScanOut112[6] , 
        \nScanOut112[5] , \nScanOut112[4] , \nScanOut112[3] , \nScanOut112[2] , 
        \nScanOut112[1] , \nScanOut112[0] }), .ScanOut({\nScanOut111[7] , 
        \nScanOut111[6] , \nScanOut111[5] , \nScanOut111[4] , \nScanOut111[3] , 
        \nScanOut111[2] , \nScanOut111[1] , \nScanOut111[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }), 
        .SouthIn({\nOut3_16[7] , \nOut3_16[6] , \nOut3_16[5] , \nOut3_16[4] , 
        \nOut3_16[3] , \nOut3_16[2] , \nOut3_16[1] , \nOut3_16[0] }), .EastIn(
        {\nOut4_15[7] , \nOut4_15[6] , \nOut4_15[5] , \nOut4_15[4] , 
        \nOut4_15[3] , \nOut4_15[2] , \nOut4_15[1] , \nOut4_15[0] }), .WestIn(
        {\nOut2_15[7] , \nOut2_15[6] , \nOut2_15[5] , \nOut2_15[4] , 
        \nOut2_15[3] , \nOut2_15[2] , \nOut2_15[1] , \nOut2_15[0] }), .Out({
        \nOut3_15[7] , \nOut3_15[6] , \nOut3_15[5] , \nOut3_15[4] , 
        \nOut3_15[3] , \nOut3_15[2] , \nOut3_15[1] , \nOut3_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_690 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut691[7] , \nScanOut691[6] , 
        \nScanOut691[5] , \nScanOut691[4] , \nScanOut691[3] , \nScanOut691[2] , 
        \nScanOut691[1] , \nScanOut691[0] }), .ScanOut({\nScanOut690[7] , 
        \nScanOut690[6] , \nScanOut690[5] , \nScanOut690[4] , \nScanOut690[3] , 
        \nScanOut690[2] , \nScanOut690[1] , \nScanOut690[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_17[7] , \nOut21_17[6] , \nOut21_17[5] , \nOut21_17[4] , 
        \nOut21_17[3] , \nOut21_17[2] , \nOut21_17[1] , \nOut21_17[0] }), 
        .SouthIn({\nOut21_19[7] , \nOut21_19[6] , \nOut21_19[5] , 
        \nOut21_19[4] , \nOut21_19[3] , \nOut21_19[2] , \nOut21_19[1] , 
        \nOut21_19[0] }), .EastIn({\nOut22_18[7] , \nOut22_18[6] , 
        \nOut22_18[5] , \nOut22_18[4] , \nOut22_18[3] , \nOut22_18[2] , 
        \nOut22_18[1] , \nOut22_18[0] }), .WestIn({\nOut20_18[7] , 
        \nOut20_18[6] , \nOut20_18[5] , \nOut20_18[4] , \nOut20_18[3] , 
        \nOut20_18[2] , \nOut20_18[1] , \nOut20_18[0] }), .Out({\nOut21_18[7] , 
        \nOut21_18[6] , \nOut21_18[5] , \nOut21_18[4] , \nOut21_18[3] , 
        \nOut21_18[2] , \nOut21_18[1] , \nOut21_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_700 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut701[7] , \nScanOut701[6] , 
        \nScanOut701[5] , \nScanOut701[4] , \nScanOut701[3] , \nScanOut701[2] , 
        \nScanOut701[1] , \nScanOut701[0] }), .ScanOut({\nScanOut700[7] , 
        \nScanOut700[6] , \nScanOut700[5] , \nScanOut700[4] , \nScanOut700[3] , 
        \nScanOut700[2] , \nScanOut700[1] , \nScanOut700[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_27[7] , \nOut21_27[6] , \nOut21_27[5] , \nOut21_27[4] , 
        \nOut21_27[3] , \nOut21_27[2] , \nOut21_27[1] , \nOut21_27[0] }), 
        .SouthIn({\nOut21_29[7] , \nOut21_29[6] , \nOut21_29[5] , 
        \nOut21_29[4] , \nOut21_29[3] , \nOut21_29[2] , \nOut21_29[1] , 
        \nOut21_29[0] }), .EastIn({\nOut22_28[7] , \nOut22_28[6] , 
        \nOut22_28[5] , \nOut22_28[4] , \nOut22_28[3] , \nOut22_28[2] , 
        \nOut22_28[1] , \nOut22_28[0] }), .WestIn({\nOut20_28[7] , 
        \nOut20_28[6] , \nOut20_28[5] , \nOut20_28[4] , \nOut20_28[3] , 
        \nOut20_28[2] , \nOut20_28[1] , \nOut20_28[0] }), .Out({\nOut21_28[7] , 
        \nOut21_28[6] , \nOut21_28[5] , \nOut21_28[4] , \nOut21_28[3] , 
        \nOut21_28[2] , \nOut21_28[1] , \nOut21_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1006 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1007[7] , \nScanOut1007[6] , 
        \nScanOut1007[5] , \nScanOut1007[4] , \nScanOut1007[3] , 
        \nScanOut1007[2] , \nScanOut1007[1] , \nScanOut1007[0] }), .ScanOut({
        \nScanOut1006[7] , \nScanOut1006[6] , \nScanOut1006[5] , 
        \nScanOut1006[4] , \nScanOut1006[3] , \nScanOut1006[2] , 
        \nScanOut1006[1] , \nScanOut1006[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_14[7] , \nOut31_14[6] , \nOut31_14[5] , 
        \nOut31_14[4] , \nOut31_14[3] , \nOut31_14[2] , \nOut31_14[1] , 
        \nOut31_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_136 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut137[7] , \nScanOut137[6] , 
        \nScanOut137[5] , \nScanOut137[4] , \nScanOut137[3] , \nScanOut137[2] , 
        \nScanOut137[1] , \nScanOut137[0] }), .ScanOut({\nScanOut136[7] , 
        \nScanOut136[6] , \nScanOut136[5] , \nScanOut136[4] , \nScanOut136[3] , 
        \nScanOut136[2] , \nScanOut136[1] , \nScanOut136[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_7[7] , \nOut4_7[6] , \nOut4_7[5] , \nOut4_7[4] , \nOut4_7[3] , 
        \nOut4_7[2] , \nOut4_7[1] , \nOut4_7[0] }), .SouthIn({\nOut4_9[7] , 
        \nOut4_9[6] , \nOut4_9[5] , \nOut4_9[4] , \nOut4_9[3] , \nOut4_9[2] , 
        \nOut4_9[1] , \nOut4_9[0] }), .EastIn({\nOut5_8[7] , \nOut5_8[6] , 
        \nOut5_8[5] , \nOut5_8[4] , \nOut5_8[3] , \nOut5_8[2] , \nOut5_8[1] , 
        \nOut5_8[0] }), .WestIn({\nOut3_8[7] , \nOut3_8[6] , \nOut3_8[5] , 
        \nOut3_8[4] , \nOut3_8[3] , \nOut3_8[2] , \nOut3_8[1] , \nOut3_8[0] }), 
        .Out({\nOut4_8[7] , \nOut4_8[6] , \nOut4_8[5] , \nOut4_8[4] , 
        \nOut4_8[3] , \nOut4_8[2] , \nOut4_8[1] , \nOut4_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_206 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut207[7] , \nScanOut207[6] , 
        \nScanOut207[5] , \nScanOut207[4] , \nScanOut207[3] , \nScanOut207[2] , 
        \nScanOut207[1] , \nScanOut207[0] }), .ScanOut({\nScanOut206[7] , 
        \nScanOut206[6] , \nScanOut206[5] , \nScanOut206[4] , \nScanOut206[3] , 
        \nScanOut206[2] , \nScanOut206[1] , \nScanOut206[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }), 
        .SouthIn({\nOut6_15[7] , \nOut6_15[6] , \nOut6_15[5] , \nOut6_15[4] , 
        \nOut6_15[3] , \nOut6_15[2] , \nOut6_15[1] , \nOut6_15[0] }), .EastIn(
        {\nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }), .WestIn(
        {\nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }), .Out({
        \nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_221 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut222[7] , \nScanOut222[6] , 
        \nScanOut222[5] , \nScanOut222[4] , \nScanOut222[3] , \nScanOut222[2] , 
        \nScanOut222[1] , \nScanOut222[0] }), .ScanOut({\nScanOut221[7] , 
        \nScanOut221[6] , \nScanOut221[5] , \nScanOut221[4] , \nScanOut221[3] , 
        \nScanOut221[2] , \nScanOut221[1] , \nScanOut221[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_28[7] , \nOut6_28[6] , \nOut6_28[5] , \nOut6_28[4] , 
        \nOut6_28[3] , \nOut6_28[2] , \nOut6_28[1] , \nOut6_28[0] }), 
        .SouthIn({\nOut6_30[7] , \nOut6_30[6] , \nOut6_30[5] , \nOut6_30[4] , 
        \nOut6_30[3] , \nOut6_30[2] , \nOut6_30[1] , \nOut6_30[0] }), .EastIn(
        {\nOut7_29[7] , \nOut7_29[6] , \nOut7_29[5] , \nOut7_29[4] , 
        \nOut7_29[3] , \nOut7_29[2] , \nOut7_29[1] , \nOut7_29[0] }), .WestIn(
        {\nOut5_29[7] , \nOut5_29[6] , \nOut5_29[5] , \nOut5_29[4] , 
        \nOut5_29[3] , \nOut5_29[2] , \nOut5_29[1] , \nOut5_29[0] }), .Out({
        \nOut6_29[7] , \nOut6_29[6] , \nOut6_29[5] , \nOut6_29[4] , 
        \nOut6_29[3] , \nOut6_29[2] , \nOut6_29[1] , \nOut6_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_430 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut431[7] , \nScanOut431[6] , 
        \nScanOut431[5] , \nScanOut431[4] , \nScanOut431[3] , \nScanOut431[2] , 
        \nScanOut431[1] , \nScanOut431[0] }), .ScanOut({\nScanOut430[7] , 
        \nScanOut430[6] , \nScanOut430[5] , \nScanOut430[4] , \nScanOut430[3] , 
        \nScanOut430[2] , \nScanOut430[1] , \nScanOut430[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_13[7] , \nOut13_13[6] , \nOut13_13[5] , \nOut13_13[4] , 
        \nOut13_13[3] , \nOut13_13[2] , \nOut13_13[1] , \nOut13_13[0] }), 
        .SouthIn({\nOut13_15[7] , \nOut13_15[6] , \nOut13_15[5] , 
        \nOut13_15[4] , \nOut13_15[3] , \nOut13_15[2] , \nOut13_15[1] , 
        \nOut13_15[0] }), .EastIn({\nOut14_14[7] , \nOut14_14[6] , 
        \nOut14_14[5] , \nOut14_14[4] , \nOut14_14[3] , \nOut14_14[2] , 
        \nOut14_14[1] , \nOut14_14[0] }), .WestIn({\nOut12_14[7] , 
        \nOut12_14[6] , \nOut12_14[5] , \nOut12_14[4] , \nOut12_14[3] , 
        \nOut12_14[2] , \nOut12_14[1] , \nOut12_14[0] }), .Out({\nOut13_14[7] , 
        \nOut13_14[6] , \nOut13_14[5] , \nOut13_14[4] , \nOut13_14[3] , 
        \nOut13_14[2] , \nOut13_14[1] , \nOut13_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_842 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut843[7] , \nScanOut843[6] , 
        \nScanOut843[5] , \nScanOut843[4] , \nScanOut843[3] , \nScanOut843[2] , 
        \nScanOut843[1] , \nScanOut843[0] }), .ScanOut({\nScanOut842[7] , 
        \nScanOut842[6] , \nScanOut842[5] , \nScanOut842[4] , \nScanOut842[3] , 
        \nScanOut842[2] , \nScanOut842[1] , \nScanOut842[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_9[7] , \nOut26_9[6] , \nOut26_9[5] , \nOut26_9[4] , 
        \nOut26_9[3] , \nOut26_9[2] , \nOut26_9[1] , \nOut26_9[0] }), 
        .SouthIn({\nOut26_11[7] , \nOut26_11[6] , \nOut26_11[5] , 
        \nOut26_11[4] , \nOut26_11[3] , \nOut26_11[2] , \nOut26_11[1] , 
        \nOut26_11[0] }), .EastIn({\nOut27_10[7] , \nOut27_10[6] , 
        \nOut27_10[5] , \nOut27_10[4] , \nOut27_10[3] , \nOut27_10[2] , 
        \nOut27_10[1] , \nOut27_10[0] }), .WestIn({\nOut25_10[7] , 
        \nOut25_10[6] , \nOut25_10[5] , \nOut25_10[4] , \nOut25_10[3] , 
        \nOut25_10[2] , \nOut25_10[1] , \nOut25_10[0] }), .Out({\nOut26_10[7] , 
        \nOut26_10[6] , \nOut26_10[5] , \nOut26_10[4] , \nOut26_10[3] , 
        \nOut26_10[2] , \nOut26_10[1] , \nOut26_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_865 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut866[7] , \nScanOut866[6] , 
        \nScanOut866[5] , \nScanOut866[4] , \nScanOut866[3] , \nScanOut866[2] , 
        \nScanOut866[1] , \nScanOut866[0] }), .ScanOut({\nScanOut865[7] , 
        \nScanOut865[6] , \nScanOut865[5] , \nScanOut865[4] , \nScanOut865[3] , 
        \nScanOut865[2] , \nScanOut865[1] , \nScanOut865[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_0[7] , \nOut27_0[6] , \nOut27_0[5] , \nOut27_0[4] , 
        \nOut27_0[3] , \nOut27_0[2] , \nOut27_0[1] , \nOut27_0[0] }), 
        .SouthIn({\nOut27_2[7] , \nOut27_2[6] , \nOut27_2[5] , \nOut27_2[4] , 
        \nOut27_2[3] , \nOut27_2[2] , \nOut27_2[1] , \nOut27_2[0] }), .EastIn(
        {\nOut28_1[7] , \nOut28_1[6] , \nOut28_1[5] , \nOut28_1[4] , 
        \nOut28_1[3] , \nOut28_1[2] , \nOut28_1[1] , \nOut28_1[0] }), .WestIn(
        {\nOut26_1[7] , \nOut26_1[6] , \nOut26_1[5] , \nOut26_1[4] , 
        \nOut26_1[3] , \nOut26_1[2] , \nOut26_1[1] , \nOut26_1[0] }), .Out({
        \nOut27_1[7] , \nOut27_1[6] , \nOut27_1[5] , \nOut27_1[4] , 
        \nOut27_1[3] , \nOut27_1[2] , \nOut27_1[1] , \nOut27_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_396 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut397[7] , \nScanOut397[6] , 
        \nScanOut397[5] , \nScanOut397[4] , \nScanOut397[3] , \nScanOut397[2] , 
        \nScanOut397[1] , \nScanOut397[0] }), .ScanOut({\nScanOut396[7] , 
        \nScanOut396[6] , \nScanOut396[5] , \nScanOut396[4] , \nScanOut396[3] , 
        \nScanOut396[2] , \nScanOut396[1] , \nScanOut396[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_11[7] , \nOut12_11[6] , \nOut12_11[5] , \nOut12_11[4] , 
        \nOut12_11[3] , \nOut12_11[2] , \nOut12_11[1] , \nOut12_11[0] }), 
        .SouthIn({\nOut12_13[7] , \nOut12_13[6] , \nOut12_13[5] , 
        \nOut12_13[4] , \nOut12_13[3] , \nOut12_13[2] , \nOut12_13[1] , 
        \nOut12_13[0] }), .EastIn({\nOut13_12[7] , \nOut13_12[6] , 
        \nOut13_12[5] , \nOut13_12[4] , \nOut13_12[3] , \nOut13_12[2] , 
        \nOut13_12[1] , \nOut13_12[0] }), .WestIn({\nOut11_12[7] , 
        \nOut11_12[6] , \nOut11_12[5] , \nOut11_12[4] , \nOut11_12[3] , 
        \nOut11_12[2] , \nOut11_12[1] , \nOut11_12[0] }), .Out({\nOut12_12[7] , 
        \nOut12_12[6] , \nOut12_12[5] , \nOut12_12[4] , \nOut12_12[3] , 
        \nOut12_12[2] , \nOut12_12[1] , \nOut12_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_587 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut588[7] , \nScanOut588[6] , 
        \nScanOut588[5] , \nScanOut588[4] , \nScanOut588[3] , \nScanOut588[2] , 
        \nScanOut588[1] , \nScanOut588[0] }), .ScanOut({\nScanOut587[7] , 
        \nScanOut587[6] , \nScanOut587[5] , \nScanOut587[4] , \nScanOut587[3] , 
        \nScanOut587[2] , \nScanOut587[1] , \nScanOut587[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_10[7] , \nOut18_10[6] , \nOut18_10[5] , \nOut18_10[4] , 
        \nOut18_10[3] , \nOut18_10[2] , \nOut18_10[1] , \nOut18_10[0] }), 
        .SouthIn({\nOut18_12[7] , \nOut18_12[6] , \nOut18_12[5] , 
        \nOut18_12[4] , \nOut18_12[3] , \nOut18_12[2] , \nOut18_12[1] , 
        \nOut18_12[0] }), .EastIn({\nOut19_11[7] , \nOut19_11[6] , 
        \nOut19_11[5] , \nOut19_11[4] , \nOut19_11[3] , \nOut19_11[2] , 
        \nOut19_11[1] , \nOut19_11[0] }), .WestIn({\nOut17_11[7] , 
        \nOut17_11[6] , \nOut17_11[5] , \nOut17_11[4] , \nOut17_11[3] , 
        \nOut17_11[2] , \nOut17_11[1] , \nOut17_11[0] }), .Out({\nOut18_11[7] , 
        \nOut18_11[6] , \nOut18_11[5] , \nOut18_11[4] , \nOut18_11[3] , 
        \nOut18_11[2] , \nOut18_11[1] , \nOut18_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_417 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut418[7] , \nScanOut418[6] , 
        \nScanOut418[5] , \nScanOut418[4] , \nScanOut418[3] , \nScanOut418[2] , 
        \nScanOut418[1] , \nScanOut418[0] }), .ScanOut({\nScanOut417[7] , 
        \nScanOut417[6] , \nScanOut417[5] , \nScanOut417[4] , \nScanOut417[3] , 
        \nScanOut417[2] , \nScanOut417[1] , \nScanOut417[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_0[7] , \nOut13_0[6] , \nOut13_0[5] , \nOut13_0[4] , 
        \nOut13_0[3] , \nOut13_0[2] , \nOut13_0[1] , \nOut13_0[0] }), 
        .SouthIn({\nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }), .EastIn(
        {\nOut14_1[7] , \nOut14_1[6] , \nOut14_1[5] , \nOut14_1[4] , 
        \nOut14_1[3] , \nOut14_1[2] , \nOut14_1[1] , \nOut14_1[0] }), .WestIn(
        {\nOut12_1[7] , \nOut12_1[6] , \nOut12_1[5] , \nOut12_1[4] , 
        \nOut12_1[3] , \nOut12_1[2] , \nOut12_1[1] , \nOut12_1[0] }), .Out({
        \nOut13_1[7] , \nOut13_1[6] , \nOut13_1[5] , \nOut13_1[4] , 
        \nOut13_1[3] , \nOut13_1[2] , \nOut13_1[1] , \nOut13_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1021 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1022[7] , \nScanOut1022[6] , 
        \nScanOut1022[5] , \nScanOut1022[4] , \nScanOut1022[3] , 
        \nScanOut1022[2] , \nScanOut1022[1] , \nScanOut1022[0] }), .ScanOut({
        \nScanOut1021[7] , \nScanOut1021[6] , \nScanOut1021[5] , 
        \nScanOut1021[4] , \nScanOut1021[3] , \nScanOut1021[2] , 
        \nScanOut1021[1] , \nScanOut1021[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_29[7] , \nOut31_29[6] , \nOut31_29[5] , 
        \nOut31_29[4] , \nOut31_29[3] , \nOut31_29[2] , \nOut31_29[1] , 
        \nOut31_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_158 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut159[7] , \nScanOut159[6] , 
        \nScanOut159[5] , \nScanOut159[4] , \nScanOut159[3] , \nScanOut159[2] , 
        \nScanOut159[1] , \nScanOut159[0] }), .ScanOut({\nScanOut158[7] , 
        \nScanOut158[6] , \nScanOut158[5] , \nScanOut158[4] , \nScanOut158[3] , 
        \nScanOut158[2] , \nScanOut158[1] , \nScanOut158[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_29[7] , \nOut4_29[6] , \nOut4_29[5] , \nOut4_29[4] , 
        \nOut4_29[3] , \nOut4_29[2] , \nOut4_29[1] , \nOut4_29[0] }), 
        .SouthIn({\nOut4_31[7] , \nOut4_31[6] , \nOut4_31[5] , \nOut4_31[4] , 
        \nOut4_31[3] , \nOut4_31[2] , \nOut4_31[1] , \nOut4_31[0] }), .EastIn(
        {\nOut5_30[7] , \nOut5_30[6] , \nOut5_30[5] , \nOut5_30[4] , 
        \nOut5_30[3] , \nOut5_30[2] , \nOut5_30[1] , \nOut5_30[0] }), .WestIn(
        {\nOut3_30[7] , \nOut3_30[6] , \nOut3_30[5] , \nOut3_30[4] , 
        \nOut3_30[3] , \nOut3_30[2] , \nOut3_30[1] , \nOut3_30[0] }), .Out({
        \nOut4_30[7] , \nOut4_30[6] , \nOut4_30[5] , \nOut4_30[4] , 
        \nOut4_30[3] , \nOut4_30[2] , \nOut4_30[1] , \nOut4_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_268 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut269[7] , \nScanOut269[6] , 
        \nScanOut269[5] , \nScanOut269[4] , \nScanOut269[3] , \nScanOut269[2] , 
        \nScanOut269[1] , \nScanOut269[0] }), .ScanOut({\nScanOut268[7] , 
        \nScanOut268[6] , \nScanOut268[5] , \nScanOut268[4] , \nScanOut268[3] , 
        \nScanOut268[2] , \nScanOut268[1] , \nScanOut268[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_11[7] , \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , 
        \nOut8_11[3] , \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }), 
        .SouthIn({\nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }), .EastIn(
        {\nOut9_12[7] , \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , 
        \nOut9_12[3] , \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }), .WestIn(
        {\nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }), .Out({
        \nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_479 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut480[7] , \nScanOut480[6] , 
        \nScanOut480[5] , \nScanOut480[4] , \nScanOut480[3] , \nScanOut480[2] , 
        \nScanOut480[1] , \nScanOut480[0] }), .ScanOut({\nScanOut479[7] , 
        \nScanOut479[6] , \nScanOut479[5] , \nScanOut479[4] , \nScanOut479[3] , 
        \nScanOut479[2] , \nScanOut479[1] , \nScanOut479[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut14_31[7] , \nOut14_31[6] , 
        \nOut14_31[5] , \nOut14_31[4] , \nOut14_31[3] , \nOut14_31[2] , 
        \nOut14_31[1] , \nOut14_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_727 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut728[7] , \nScanOut728[6] , 
        \nScanOut728[5] , \nScanOut728[4] , \nScanOut728[3] , \nScanOut728[2] , 
        \nScanOut728[1] , \nScanOut728[0] }), .ScanOut({\nScanOut727[7] , 
        \nScanOut727[6] , \nScanOut727[5] , \nScanOut727[4] , \nScanOut727[3] , 
        \nScanOut727[2] , \nScanOut727[1] , \nScanOut727[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_22[7] , \nOut22_22[6] , \nOut22_22[5] , \nOut22_22[4] , 
        \nOut22_22[3] , \nOut22_22[2] , \nOut22_22[1] , \nOut22_22[0] }), 
        .SouthIn({\nOut22_24[7] , \nOut22_24[6] , \nOut22_24[5] , 
        \nOut22_24[4] , \nOut22_24[3] , \nOut22_24[2] , \nOut22_24[1] , 
        \nOut22_24[0] }), .EastIn({\nOut23_23[7] , \nOut23_23[6] , 
        \nOut23_23[5] , \nOut23_23[4] , \nOut23_23[3] , \nOut23_23[2] , 
        \nOut23_23[1] , \nOut23_23[0] }), .WestIn({\nOut21_23[7] , 
        \nOut21_23[6] , \nOut21_23[5] , \nOut21_23[4] , \nOut21_23[3] , 
        \nOut21_23[2] , \nOut21_23[1] , \nOut21_23[0] }), .Out({\nOut22_23[7] , 
        \nOut22_23[6] , \nOut22_23[5] , \nOut22_23[4] , \nOut22_23[3] , 
        \nOut22_23[2] , \nOut22_23[1] , \nOut22_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_749 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut750[7] , \nScanOut750[6] , 
        \nScanOut750[5] , \nScanOut750[4] , \nScanOut750[3] , \nScanOut750[2] , 
        \nScanOut750[1] , \nScanOut750[0] }), .ScanOut({\nScanOut749[7] , 
        \nScanOut749[6] , \nScanOut749[5] , \nScanOut749[4] , \nScanOut749[3] , 
        \nScanOut749[2] , \nScanOut749[1] , \nScanOut749[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_12[7] , \nOut23_12[6] , \nOut23_12[5] , \nOut23_12[4] , 
        \nOut23_12[3] , \nOut23_12[2] , \nOut23_12[1] , \nOut23_12[0] }), 
        .SouthIn({\nOut23_14[7] , \nOut23_14[6] , \nOut23_14[5] , 
        \nOut23_14[4] , \nOut23_14[3] , \nOut23_14[2] , \nOut23_14[1] , 
        \nOut23_14[0] }), .EastIn({\nOut24_13[7] , \nOut24_13[6] , 
        \nOut24_13[5] , \nOut24_13[4] , \nOut24_13[3] , \nOut24_13[2] , 
        \nOut24_13[1] , \nOut24_13[0] }), .WestIn({\nOut22_13[7] , 
        \nOut22_13[6] , \nOut22_13[5] , \nOut22_13[4] , \nOut22_13[3] , 
        \nOut22_13[2] , \nOut22_13[1] , \nOut22_13[0] }), .Out({\nOut23_13[7] , 
        \nOut23_13[6] , \nOut23_13[5] , \nOut23_13[4] , \nOut23_13[3] , 
        \nOut23_13[2] , \nOut23_13[1] , \nOut23_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_373 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut374[7] , \nScanOut374[6] , 
        \nScanOut374[5] , \nScanOut374[4] , \nScanOut374[3] , \nScanOut374[2] , 
        \nScanOut374[1] , \nScanOut374[0] }), .ScanOut({\nScanOut373[7] , 
        \nScanOut373[6] , \nScanOut373[5] , \nScanOut373[4] , \nScanOut373[3] , 
        \nScanOut373[2] , \nScanOut373[1] , \nScanOut373[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_20[7] , \nOut11_20[6] , \nOut11_20[5] , \nOut11_20[4] , 
        \nOut11_20[3] , \nOut11_20[2] , \nOut11_20[1] , \nOut11_20[0] }), 
        .SouthIn({\nOut11_22[7] , \nOut11_22[6] , \nOut11_22[5] , 
        \nOut11_22[4] , \nOut11_22[3] , \nOut11_22[2] , \nOut11_22[1] , 
        \nOut11_22[0] }), .EastIn({\nOut12_21[7] , \nOut12_21[6] , 
        \nOut12_21[5] , \nOut12_21[4] , \nOut12_21[3] , \nOut12_21[2] , 
        \nOut12_21[1] , \nOut12_21[0] }), .WestIn({\nOut10_21[7] , 
        \nOut10_21[6] , \nOut10_21[5] , \nOut10_21[4] , \nOut10_21[3] , 
        \nOut10_21[2] , \nOut10_21[1] , \nOut10_21[0] }), .Out({\nOut11_21[7] , 
        \nOut11_21[6] , \nOut11_21[5] , \nOut11_21[4] , \nOut11_21[3] , 
        \nOut11_21[2] , \nOut11_21[1] , \nOut11_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_880 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut881[7] , \nScanOut881[6] , 
        \nScanOut881[5] , \nScanOut881[4] , \nScanOut881[3] , \nScanOut881[2] , 
        \nScanOut881[1] , \nScanOut881[0] }), .ScanOut({\nScanOut880[7] , 
        \nScanOut880[6] , \nScanOut880[5] , \nScanOut880[4] , \nScanOut880[3] , 
        \nScanOut880[2] , \nScanOut880[1] , \nScanOut880[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_15[7] , \nOut27_15[6] , \nOut27_15[5] , \nOut27_15[4] , 
        \nOut27_15[3] , \nOut27_15[2] , \nOut27_15[1] , \nOut27_15[0] }), 
        .SouthIn({\nOut27_17[7] , \nOut27_17[6] , \nOut27_17[5] , 
        \nOut27_17[4] , \nOut27_17[3] , \nOut27_17[2] , \nOut27_17[1] , 
        \nOut27_17[0] }), .EastIn({\nOut28_16[7] , \nOut28_16[6] , 
        \nOut28_16[5] , \nOut28_16[4] , \nOut28_16[3] , \nOut28_16[2] , 
        \nOut28_16[1] , \nOut28_16[0] }), .WestIn({\nOut26_16[7] , 
        \nOut26_16[6] , \nOut26_16[5] , \nOut26_16[4] , \nOut26_16[3] , 
        \nOut26_16[2] , \nOut26_16[1] , \nOut26_16[0] }), .Out({\nOut27_16[7] , 
        \nOut27_16[6] , \nOut27_16[5] , \nOut27_16[4] , \nOut27_16[3] , 
        \nOut27_16[2] , \nOut27_16[1] , \nOut27_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_910 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut911[7] , \nScanOut911[6] , 
        \nScanOut911[5] , \nScanOut911[4] , \nScanOut911[3] , \nScanOut911[2] , 
        \nScanOut911[1] , \nScanOut911[0] }), .ScanOut({\nScanOut910[7] , 
        \nScanOut910[6] , \nScanOut910[5] , \nScanOut910[4] , \nScanOut910[3] , 
        \nScanOut910[2] , \nScanOut910[1] , \nScanOut910[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_13[7] , \nOut28_13[6] , \nOut28_13[5] , \nOut28_13[4] , 
        \nOut28_13[3] , \nOut28_13[2] , \nOut28_13[1] , \nOut28_13[0] }), 
        .SouthIn({\nOut28_15[7] , \nOut28_15[6] , \nOut28_15[5] , 
        \nOut28_15[4] , \nOut28_15[3] , \nOut28_15[2] , \nOut28_15[1] , 
        \nOut28_15[0] }), .EastIn({\nOut29_14[7] , \nOut29_14[6] , 
        \nOut29_14[5] , \nOut29_14[4] , \nOut29_14[3] , \nOut29_14[2] , 
        \nOut29_14[1] , \nOut29_14[0] }), .WestIn({\nOut27_14[7] , 
        \nOut27_14[6] , \nOut27_14[5] , \nOut27_14[4] , \nOut27_14[3] , 
        \nOut27_14[2] , \nOut27_14[1] , \nOut27_14[0] }), .Out({\nOut28_14[7] , 
        \nOut28_14[6] , \nOut28_14[5] , \nOut28_14[4] , \nOut28_14[3] , 
        \nOut28_14[2] , \nOut28_14[1] , \nOut28_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_562 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut563[7] , \nScanOut563[6] , 
        \nScanOut563[5] , \nScanOut563[4] , \nScanOut563[3] , \nScanOut563[2] , 
        \nScanOut563[1] , \nScanOut563[0] }), .ScanOut({\nScanOut562[7] , 
        \nScanOut562[6] , \nScanOut562[5] , \nScanOut562[4] , \nScanOut562[3] , 
        \nScanOut562[2] , \nScanOut562[1] , \nScanOut562[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_17[7] , \nOut17_17[6] , \nOut17_17[5] , \nOut17_17[4] , 
        \nOut17_17[3] , \nOut17_17[2] , \nOut17_17[1] , \nOut17_17[0] }), 
        .SouthIn({\nOut17_19[7] , \nOut17_19[6] , \nOut17_19[5] , 
        \nOut17_19[4] , \nOut17_19[3] , \nOut17_19[2] , \nOut17_19[1] , 
        \nOut17_19[0] }), .EastIn({\nOut18_18[7] , \nOut18_18[6] , 
        \nOut18_18[5] , \nOut18_18[4] , \nOut18_18[3] , \nOut18_18[2] , 
        \nOut18_18[1] , \nOut18_18[0] }), .WestIn({\nOut16_18[7] , 
        \nOut16_18[6] , \nOut16_18[5] , \nOut16_18[4] , \nOut16_18[3] , 
        \nOut16_18[2] , \nOut16_18[1] , \nOut16_18[0] }), .Out({\nOut17_18[7] , 
        \nOut17_18[6] , \nOut17_18[5] , \nOut17_18[4] , \nOut17_18[3] , 
        \nOut17_18[2] , \nOut17_18[1] , \nOut17_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_652 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut653[7] , \nScanOut653[6] , 
        \nScanOut653[5] , \nScanOut653[4] , \nScanOut653[3] , \nScanOut653[2] , 
        \nScanOut653[1] , \nScanOut653[0] }), .ScanOut({\nScanOut652[7] , 
        \nScanOut652[6] , \nScanOut652[5] , \nScanOut652[4] , \nScanOut652[3] , 
        \nScanOut652[2] , \nScanOut652[1] , \nScanOut652[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_11[7] , \nOut20_11[6] , \nOut20_11[5] , \nOut20_11[4] , 
        \nOut20_11[3] , \nOut20_11[2] , \nOut20_11[1] , \nOut20_11[0] }), 
        .SouthIn({\nOut20_13[7] , \nOut20_13[6] , \nOut20_13[5] , 
        \nOut20_13[4] , \nOut20_13[3] , \nOut20_13[2] , \nOut20_13[1] , 
        \nOut20_13[0] }), .EastIn({\nOut21_12[7] , \nOut21_12[6] , 
        \nOut21_12[5] , \nOut21_12[4] , \nOut21_12[3] , \nOut21_12[2] , 
        \nOut21_12[1] , \nOut21_12[0] }), .WestIn({\nOut19_12[7] , 
        \nOut19_12[6] , \nOut19_12[5] , \nOut19_12[4] , \nOut19_12[3] , 
        \nOut19_12[2] , \nOut19_12[1] , \nOut19_12[0] }), .Out({\nOut20_12[7] , 
        \nOut20_12[6] , \nOut20_12[5] , \nOut20_12[4] , \nOut20_12[3] , 
        \nOut20_12[2] , \nOut20_12[1] , \nOut20_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_6 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut7[7] , \nScanOut7[6] , 
        \nScanOut7[5] , \nScanOut7[4] , \nScanOut7[3] , \nScanOut7[2] , 
        \nScanOut7[1] , \nScanOut7[0] }), .ScanOut({\nScanOut6[7] , 
        \nScanOut6[6] , \nScanOut6[5] , \nScanOut6[4] , \nScanOut6[3] , 
        \nScanOut6[2] , \nScanOut6[1] , \nScanOut6[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_6[7] , \nOut0_6[6] , 
        \nOut0_6[5] , \nOut0_6[4] , \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , 
        \nOut0_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_8 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut9[7] , \nScanOut9[6] , 
        \nScanOut9[5] , \nScanOut9[4] , \nScanOut9[3] , \nScanOut9[2] , 
        \nScanOut9[1] , \nScanOut9[0] }), .ScanOut({\nScanOut8[7] , 
        \nScanOut8[6] , \nScanOut8[5] , \nScanOut8[4] , \nScanOut8[3] , 
        \nScanOut8[2] , \nScanOut8[1] , \nScanOut8[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_8[7] , \nOut0_8[6] , 
        \nOut0_8[5] , \nOut0_8[4] , \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , 
        \nOut0_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_15 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut16[7] , \nScanOut16[6] , 
        \nScanOut16[5] , \nScanOut16[4] , \nScanOut16[3] , \nScanOut16[2] , 
        \nScanOut16[1] , \nScanOut16[0] }), .ScanOut({\nScanOut15[7] , 
        \nScanOut15[6] , \nScanOut15[5] , \nScanOut15[4] , \nScanOut15[3] , 
        \nScanOut15[2] , \nScanOut15[1] , \nScanOut15[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_15[7] , \nOut0_15[6] , 
        \nOut0_15[5] , \nOut0_15[4] , \nOut0_15[3] , \nOut0_15[2] , 
        \nOut0_15[1] , \nOut0_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_32 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut33[7] , \nScanOut33[6] , 
        \nScanOut33[5] , \nScanOut33[4] , \nScanOut33[3] , \nScanOut33[2] , 
        \nScanOut33[1] , \nScanOut33[0] }), .ScanOut({\nScanOut32[7] , 
        \nScanOut32[6] , \nScanOut32[5] , \nScanOut32[4] , \nScanOut32[3] , 
        \nScanOut32[2] , \nScanOut32[1] , \nScanOut32[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut1_0[7] , \nOut1_0[6] , 
        \nOut1_0[5] , \nOut1_0[4] , \nOut1_0[3] , \nOut1_0[2] , \nOut1_0[1] , 
        \nOut1_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_47 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut48[7] , \nScanOut48[6] , 
        \nScanOut48[5] , \nScanOut48[4] , \nScanOut48[3] , \nScanOut48[2] , 
        \nScanOut48[1] , \nScanOut48[0] }), .ScanOut({\nScanOut47[7] , 
        \nScanOut47[6] , \nScanOut47[5] , \nScanOut47[4] , \nScanOut47[3] , 
        \nScanOut47[2] , \nScanOut47[1] , \nScanOut47[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), 
        .SouthIn({\nOut1_16[7] , \nOut1_16[6] , \nOut1_16[5] , \nOut1_16[4] , 
        \nOut1_16[3] , \nOut1_16[2] , \nOut1_16[1] , \nOut1_16[0] }), .EastIn(
        {\nOut2_15[7] , \nOut2_15[6] , \nOut2_15[5] , \nOut2_15[4] , 
        \nOut2_15[3] , \nOut2_15[2] , \nOut2_15[1] , \nOut2_15[0] }), .WestIn(
        {\nOut0_15[7] , \nOut0_15[6] , \nOut0_15[5] , \nOut0_15[4] , 
        \nOut0_15[3] , \nOut0_15[2] , \nOut0_15[1] , \nOut0_15[0] }), .Out({
        \nOut1_15[7] , \nOut1_15[6] , \nOut1_15[5] , \nOut1_15[4] , 
        \nOut1_15[3] , \nOut1_15[2] , \nOut1_15[1] , \nOut1_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_60 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut61[7] , \nScanOut61[6] , 
        \nScanOut61[5] , \nScanOut61[4] , \nScanOut61[3] , \nScanOut61[2] , 
        \nScanOut61[1] , \nScanOut61[0] }), .ScanOut({\nScanOut60[7] , 
        \nScanOut60[6] , \nScanOut60[5] , \nScanOut60[4] , \nScanOut60[3] , 
        \nScanOut60[2] , \nScanOut60[1] , \nScanOut60[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_27[7] , \nOut1_27[6] , \nOut1_27[5] , \nOut1_27[4] , 
        \nOut1_27[3] , \nOut1_27[2] , \nOut1_27[1] , \nOut1_27[0] }), 
        .SouthIn({\nOut1_29[7] , \nOut1_29[6] , \nOut1_29[5] , \nOut1_29[4] , 
        \nOut1_29[3] , \nOut1_29[2] , \nOut1_29[1] , \nOut1_29[0] }), .EastIn(
        {\nOut2_28[7] , \nOut2_28[6] , \nOut2_28[5] , \nOut2_28[4] , 
        \nOut2_28[3] , \nOut2_28[2] , \nOut2_28[1] , \nOut2_28[0] }), .WestIn(
        {\nOut0_28[7] , \nOut0_28[6] , \nOut0_28[5] , \nOut0_28[4] , 
        \nOut0_28[3] , \nOut0_28[2] , \nOut0_28[1] , \nOut0_28[0] }), .Out({
        \nOut1_28[7] , \nOut1_28[6] , \nOut1_28[5] , \nOut1_28[4] , 
        \nOut1_28[3] , \nOut1_28[2] , \nOut1_28[1] , \nOut1_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_675 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut676[7] , \nScanOut676[6] , 
        \nScanOut676[5] , \nScanOut676[4] , \nScanOut676[3] , \nScanOut676[2] , 
        \nScanOut676[1] , \nScanOut676[0] }), .ScanOut({\nScanOut675[7] , 
        \nScanOut675[6] , \nScanOut675[5] , \nScanOut675[4] , \nScanOut675[3] , 
        \nScanOut675[2] , \nScanOut675[1] , \nScanOut675[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_2[7] , \nOut21_2[6] , \nOut21_2[5] , \nOut21_2[4] , 
        \nOut21_2[3] , \nOut21_2[2] , \nOut21_2[1] , \nOut21_2[0] }), 
        .SouthIn({\nOut21_4[7] , \nOut21_4[6] , \nOut21_4[5] , \nOut21_4[4] , 
        \nOut21_4[3] , \nOut21_4[2] , \nOut21_4[1] , \nOut21_4[0] }), .EastIn(
        {\nOut22_3[7] , \nOut22_3[6] , \nOut22_3[5] , \nOut22_3[4] , 
        \nOut22_3[3] , \nOut22_3[2] , \nOut22_3[1] , \nOut22_3[0] }), .WestIn(
        {\nOut20_3[7] , \nOut20_3[6] , \nOut20_3[5] , \nOut20_3[4] , 
        \nOut20_3[3] , \nOut20_3[2] , \nOut20_3[1] , \nOut20_3[0] }), .Out({
        \nOut21_3[7] , \nOut21_3[6] , \nOut21_3[5] , \nOut21_3[4] , 
        \nOut21_3[3] , \nOut21_3[2] , \nOut21_3[1] , \nOut21_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_143 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut144[7] , \nScanOut144[6] , 
        \nScanOut144[5] , \nScanOut144[4] , \nScanOut144[3] , \nScanOut144[2] , 
        \nScanOut144[1] , \nScanOut144[0] }), .ScanOut({\nScanOut143[7] , 
        \nScanOut143[6] , \nScanOut143[5] , \nScanOut143[4] , \nScanOut143[3] , 
        \nScanOut143[2] , \nScanOut143[1] , \nScanOut143[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }), 
        .SouthIn({\nOut4_16[7] , \nOut4_16[6] , \nOut4_16[5] , \nOut4_16[4] , 
        \nOut4_16[3] , \nOut4_16[2] , \nOut4_16[1] , \nOut4_16[0] }), .EastIn(
        {\nOut5_15[7] , \nOut5_15[6] , \nOut5_15[5] , \nOut5_15[4] , 
        \nOut5_15[3] , \nOut5_15[2] , \nOut5_15[1] , \nOut5_15[0] }), .WestIn(
        {\nOut3_15[7] , \nOut3_15[6] , \nOut3_15[5] , \nOut3_15[4] , 
        \nOut3_15[3] , \nOut3_15[2] , \nOut3_15[1] , \nOut3_15[0] }), .Out({
        \nOut4_15[7] , \nOut4_15[6] , \nOut4_15[5] , \nOut4_15[4] , 
        \nOut4_15[3] , \nOut4_15[2] , \nOut4_15[1] , \nOut4_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_164 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut165[7] , \nScanOut165[6] , 
        \nScanOut165[5] , \nScanOut165[4] , \nScanOut165[3] , \nScanOut165[2] , 
        \nScanOut165[1] , \nScanOut165[0] }), .ScanOut({\nScanOut164[7] , 
        \nScanOut164[6] , \nScanOut164[5] , \nScanOut164[4] , \nScanOut164[3] , 
        \nScanOut164[2] , \nScanOut164[1] , \nScanOut164[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_3[7] , \nOut5_3[6] , \nOut5_3[5] , \nOut5_3[4] , \nOut5_3[3] , 
        \nOut5_3[2] , \nOut5_3[1] , \nOut5_3[0] }), .SouthIn({\nOut5_5[7] , 
        \nOut5_5[6] , \nOut5_5[5] , \nOut5_5[4] , \nOut5_5[3] , \nOut5_5[2] , 
        \nOut5_5[1] , \nOut5_5[0] }), .EastIn({\nOut6_4[7] , \nOut6_4[6] , 
        \nOut6_4[5] , \nOut6_4[4] , \nOut6_4[3] , \nOut6_4[2] , \nOut6_4[1] , 
        \nOut6_4[0] }), .WestIn({\nOut4_4[7] , \nOut4_4[6] , \nOut4_4[5] , 
        \nOut4_4[4] , \nOut4_4[3] , \nOut4_4[2] , \nOut4_4[1] , \nOut4_4[0] }), 
        .Out({\nOut5_4[7] , \nOut5_4[6] , \nOut5_4[5] , \nOut5_4[4] , 
        \nOut5_4[3] , \nOut5_4[2] , \nOut5_4[1] , \nOut5_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_254 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut255[7] , \nScanOut255[6] , 
        \nScanOut255[5] , \nScanOut255[4] , \nScanOut255[3] , \nScanOut255[2] , 
        \nScanOut255[1] , \nScanOut255[0] }), .ScanOut({\nScanOut254[7] , 
        \nScanOut254[6] , \nScanOut254[5] , \nScanOut254[4] , \nScanOut254[3] , 
        \nScanOut254[2] , \nScanOut254[1] , \nScanOut254[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_29[7] , \nOut7_29[6] , \nOut7_29[5] , \nOut7_29[4] , 
        \nOut7_29[3] , \nOut7_29[2] , \nOut7_29[1] , \nOut7_29[0] }), 
        .SouthIn({\nOut7_31[7] , \nOut7_31[6] , \nOut7_31[5] , \nOut7_31[4] , 
        \nOut7_31[3] , \nOut7_31[2] , \nOut7_31[1] , \nOut7_31[0] }), .EastIn(
        {\nOut8_30[7] , \nOut8_30[6] , \nOut8_30[5] , \nOut8_30[4] , 
        \nOut8_30[3] , \nOut8_30[2] , \nOut8_30[1] , \nOut8_30[0] }), .WestIn(
        {\nOut6_30[7] , \nOut6_30[6] , \nOut6_30[5] , \nOut6_30[4] , 
        \nOut6_30[3] , \nOut6_30[2] , \nOut6_30[1] , \nOut6_30[0] }), .Out({
        \nOut7_30[7] , \nOut7_30[6] , \nOut7_30[5] , \nOut7_30[4] , 
        \nOut7_30[3] , \nOut7_30[2] , \nOut7_30[1] , \nOut7_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_354 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut355[7] , \nScanOut355[6] , 
        \nScanOut355[5] , \nScanOut355[4] , \nScanOut355[3] , \nScanOut355[2] , 
        \nScanOut355[1] , \nScanOut355[0] }), .ScanOut({\nScanOut354[7] , 
        \nScanOut354[6] , \nScanOut354[5] , \nScanOut354[4] , \nScanOut354[3] , 
        \nScanOut354[2] , \nScanOut354[1] , \nScanOut354[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_1[7] , \nOut11_1[6] , \nOut11_1[5] , \nOut11_1[4] , 
        \nOut11_1[3] , \nOut11_1[2] , \nOut11_1[1] , \nOut11_1[0] }), 
        .SouthIn({\nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }), .EastIn(
        {\nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }), .WestIn(
        {\nOut10_2[7] , \nOut10_2[6] , \nOut10_2[5] , \nOut10_2[4] , 
        \nOut10_2[3] , \nOut10_2[2] , \nOut10_2[1] , \nOut10_2[0] }), .Out({
        \nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_545 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut546[7] , \nScanOut546[6] , 
        \nScanOut546[5] , \nScanOut546[4] , \nScanOut546[3] , \nScanOut546[2] , 
        \nScanOut546[1] , \nScanOut546[0] }), .ScanOut({\nScanOut545[7] , 
        \nScanOut545[6] , \nScanOut545[5] , \nScanOut545[4] , \nScanOut545[3] , 
        \nScanOut545[2] , \nScanOut545[1] , \nScanOut545[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_0[7] , \nOut17_0[6] , \nOut17_0[5] , \nOut17_0[4] , 
        \nOut17_0[3] , \nOut17_0[2] , \nOut17_0[1] , \nOut17_0[0] }), 
        .SouthIn({\nOut17_2[7] , \nOut17_2[6] , \nOut17_2[5] , \nOut17_2[4] , 
        \nOut17_2[3] , \nOut17_2[2] , \nOut17_2[1] , \nOut17_2[0] }), .EastIn(
        {\nOut18_1[7] , \nOut18_1[6] , \nOut18_1[5] , \nOut18_1[4] , 
        \nOut18_1[3] , \nOut18_1[2] , \nOut18_1[1] , \nOut18_1[0] }), .WestIn(
        {\nOut16_1[7] , \nOut16_1[6] , \nOut16_1[5] , \nOut16_1[4] , 
        \nOut16_1[3] , \nOut16_1[2] , \nOut16_1[1] , \nOut16_1[0] }), .Out({
        \nOut17_1[7] , \nOut17_1[6] , \nOut17_1[5] , \nOut17_1[4] , 
        \nOut17_1[3] , \nOut17_1[2] , \nOut17_1[1] , \nOut17_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_937 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut938[7] , \nScanOut938[6] , 
        \nScanOut938[5] , \nScanOut938[4] , \nScanOut938[3] , \nScanOut938[2] , 
        \nScanOut938[1] , \nScanOut938[0] }), .ScanOut({\nScanOut937[7] , 
        \nScanOut937[6] , \nScanOut937[5] , \nScanOut937[4] , \nScanOut937[3] , 
        \nScanOut937[2] , \nScanOut937[1] , \nScanOut937[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_8[7] , \nOut29_8[6] , \nOut29_8[5] , \nOut29_8[4] , 
        \nOut29_8[3] , \nOut29_8[2] , \nOut29_8[1] , \nOut29_8[0] }), 
        .SouthIn({\nOut29_10[7] , \nOut29_10[6] , \nOut29_10[5] , 
        \nOut29_10[4] , \nOut29_10[3] , \nOut29_10[2] , \nOut29_10[1] , 
        \nOut29_10[0] }), .EastIn({\nOut30_9[7] , \nOut30_9[6] , \nOut30_9[5] , 
        \nOut30_9[4] , \nOut30_9[3] , \nOut30_9[2] , \nOut30_9[1] , 
        \nOut30_9[0] }), .WestIn({\nOut28_9[7] , \nOut28_9[6] , \nOut28_9[5] , 
        \nOut28_9[4] , \nOut28_9[3] , \nOut28_9[2] , \nOut28_9[1] , 
        \nOut28_9[0] }), .Out({\nOut29_9[7] , \nOut29_9[6] , \nOut29_9[5] , 
        \nOut29_9[4] , \nOut29_9[3] , \nOut29_9[2] , \nOut29_9[1] , 
        \nOut29_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_368 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut369[7] , \nScanOut369[6] , 
        \nScanOut369[5] , \nScanOut369[4] , \nScanOut369[3] , \nScanOut369[2] , 
        \nScanOut369[1] , \nScanOut369[0] }), .ScanOut({\nScanOut368[7] , 
        \nScanOut368[6] , \nScanOut368[5] , \nScanOut368[4] , \nScanOut368[3] , 
        \nScanOut368[2] , \nScanOut368[1] , \nScanOut368[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_15[7] , \nOut11_15[6] , \nOut11_15[5] , \nOut11_15[4] , 
        \nOut11_15[3] , \nOut11_15[2] , \nOut11_15[1] , \nOut11_15[0] }), 
        .SouthIn({\nOut11_17[7] , \nOut11_17[6] , \nOut11_17[5] , 
        \nOut11_17[4] , \nOut11_17[3] , \nOut11_17[2] , \nOut11_17[1] , 
        \nOut11_17[0] }), .EastIn({\nOut12_16[7] , \nOut12_16[6] , 
        \nOut12_16[5] , \nOut12_16[4] , \nOut12_16[3] , \nOut12_16[2] , 
        \nOut12_16[1] , \nOut12_16[0] }), .WestIn({\nOut10_16[7] , 
        \nOut10_16[6] , \nOut10_16[5] , \nOut10_16[4] , \nOut10_16[3] , 
        \nOut10_16[2] , \nOut10_16[1] , \nOut10_16[0] }), .Out({\nOut11_16[7] , 
        \nOut11_16[6] , \nOut11_16[5] , \nOut11_16[4] , \nOut11_16[3] , 
        \nOut11_16[2] , \nOut11_16[1] , \nOut11_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_649 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut650[7] , \nScanOut650[6] , 
        \nScanOut650[5] , \nScanOut650[4] , \nScanOut650[3] , \nScanOut650[2] , 
        \nScanOut650[1] , \nScanOut650[0] }), .ScanOut({\nScanOut649[7] , 
        \nScanOut649[6] , \nScanOut649[5] , \nScanOut649[4] , \nScanOut649[3] , 
        \nScanOut649[2] , \nScanOut649[1] , \nScanOut649[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_8[7] , \nOut20_8[6] , \nOut20_8[5] , \nOut20_8[4] , 
        \nOut20_8[3] , \nOut20_8[2] , \nOut20_8[1] , \nOut20_8[0] }), 
        .SouthIn({\nOut20_10[7] , \nOut20_10[6] , \nOut20_10[5] , 
        \nOut20_10[4] , \nOut20_10[3] , \nOut20_10[2] , \nOut20_10[1] , 
        \nOut20_10[0] }), .EastIn({\nOut21_9[7] , \nOut21_9[6] , \nOut21_9[5] , 
        \nOut21_9[4] , \nOut21_9[3] , \nOut21_9[2] , \nOut21_9[1] , 
        \nOut21_9[0] }), .WestIn({\nOut19_9[7] , \nOut19_9[6] , \nOut19_9[5] , 
        \nOut19_9[4] , \nOut19_9[3] , \nOut19_9[2] , \nOut19_9[1] , 
        \nOut19_9[0] }), .Out({\nOut20_9[7] , \nOut20_9[6] , \nOut20_9[5] , 
        \nOut20_9[4] , \nOut20_9[3] , \nOut20_9[2] , \nOut20_9[1] , 
        \nOut20_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_579 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut580[7] , \nScanOut580[6] , 
        \nScanOut580[5] , \nScanOut580[4] , \nScanOut580[3] , \nScanOut580[2] , 
        \nScanOut580[1] , \nScanOut580[0] }), .ScanOut({\nScanOut579[7] , 
        \nScanOut579[6] , \nScanOut579[5] , \nScanOut579[4] , \nScanOut579[3] , 
        \nScanOut579[2] , \nScanOut579[1] , \nScanOut579[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_2[7] , \nOut18_2[6] , \nOut18_2[5] , \nOut18_2[4] , 
        \nOut18_2[3] , \nOut18_2[2] , \nOut18_2[1] , \nOut18_2[0] }), 
        .SouthIn({\nOut18_4[7] , \nOut18_4[6] , \nOut18_4[5] , \nOut18_4[4] , 
        \nOut18_4[3] , \nOut18_4[2] , \nOut18_4[1] , \nOut18_4[0] }), .EastIn(
        {\nOut19_3[7] , \nOut19_3[6] , \nOut19_3[5] , \nOut19_3[4] , 
        \nOut19_3[3] , \nOut19_3[2] , \nOut19_3[1] , \nOut19_3[0] }), .WestIn(
        {\nOut17_3[7] , \nOut17_3[6] , \nOut17_3[5] , \nOut17_3[4] , 
        \nOut17_3[3] , \nOut17_3[2] , \nOut17_3[1] , \nOut17_3[0] }), .Out({
        \nOut18_3[7] , \nOut18_3[6] , \nOut18_3[5] , \nOut18_3[4] , 
        \nOut18_3[3] , \nOut18_3[2] , \nOut18_3[1] , \nOut18_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_837 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut838[7] , \nScanOut838[6] , 
        \nScanOut838[5] , \nScanOut838[4] , \nScanOut838[3] , \nScanOut838[2] , 
        \nScanOut838[1] , \nScanOut838[0] }), .ScanOut({\nScanOut837[7] , 
        \nScanOut837[6] , \nScanOut837[5] , \nScanOut837[4] , \nScanOut837[3] , 
        \nScanOut837[2] , \nScanOut837[1] , \nScanOut837[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_4[7] , \nOut26_4[6] , \nOut26_4[5] , \nOut26_4[4] , 
        \nOut26_4[3] , \nOut26_4[2] , \nOut26_4[1] , \nOut26_4[0] }), 
        .SouthIn({\nOut26_6[7] , \nOut26_6[6] , \nOut26_6[5] , \nOut26_6[4] , 
        \nOut26_6[3] , \nOut26_6[2] , \nOut26_6[1] , \nOut26_6[0] }), .EastIn(
        {\nOut27_5[7] , \nOut27_5[6] , \nOut27_5[5] , \nOut27_5[4] , 
        \nOut27_5[3] , \nOut27_5[2] , \nOut27_5[1] , \nOut27_5[0] }), .WestIn(
        {\nOut25_5[7] , \nOut25_5[6] , \nOut25_5[5] , \nOut25_5[4] , 
        \nOut25_5[3] , \nOut25_5[2] , \nOut25_5[1] , \nOut25_5[0] }), .Out({
        \nOut26_5[7] , \nOut26_5[6] , \nOut26_5[5] , \nOut26_5[4] , 
        \nOut26_5[3] , \nOut26_5[2] , \nOut26_5[1] , \nOut26_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_445 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut446[7] , \nScanOut446[6] , 
        \nScanOut446[5] , \nScanOut446[4] , \nScanOut446[3] , \nScanOut446[2] , 
        \nScanOut446[1] , \nScanOut446[0] }), .ScanOut({\nScanOut445[7] , 
        \nScanOut445[6] , \nScanOut445[5] , \nScanOut445[4] , \nScanOut445[3] , 
        \nScanOut445[2] , \nScanOut445[1] , \nScanOut445[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_28[7] , \nOut13_28[6] , \nOut13_28[5] , \nOut13_28[4] , 
        \nOut13_28[3] , \nOut13_28[2] , \nOut13_28[1] , \nOut13_28[0] }), 
        .SouthIn({\nOut13_30[7] , \nOut13_30[6] , \nOut13_30[5] , 
        \nOut13_30[4] , \nOut13_30[3] , \nOut13_30[2] , \nOut13_30[1] , 
        \nOut13_30[0] }), .EastIn({\nOut14_29[7] , \nOut14_29[6] , 
        \nOut14_29[5] , \nOut14_29[4] , \nOut14_29[3] , \nOut14_29[2] , 
        \nOut14_29[1] , \nOut14_29[0] }), .WestIn({\nOut12_29[7] , 
        \nOut12_29[6] , \nOut12_29[5] , \nOut12_29[4] , \nOut12_29[3] , 
        \nOut12_29[2] , \nOut12_29[1] , \nOut12_29[0] }), .Out({\nOut13_29[7] , 
        \nOut13_29[6] , \nOut13_29[5] , \nOut13_29[4] , \nOut13_29[3] , 
        \nOut13_29[2] , \nOut13_29[1] , \nOut13_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_752 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut753[7] , \nScanOut753[6] , 
        \nScanOut753[5] , \nScanOut753[4] , \nScanOut753[3] , \nScanOut753[2] , 
        \nScanOut753[1] , \nScanOut753[0] }), .ScanOut({\nScanOut752[7] , 
        \nScanOut752[6] , \nScanOut752[5] , \nScanOut752[4] , \nScanOut752[3] , 
        \nScanOut752[2] , \nScanOut752[1] , \nScanOut752[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_15[7] , \nOut23_15[6] , \nOut23_15[5] , \nOut23_15[4] , 
        \nOut23_15[3] , \nOut23_15[2] , \nOut23_15[1] , \nOut23_15[0] }), 
        .SouthIn({\nOut23_17[7] , \nOut23_17[6] , \nOut23_17[5] , 
        \nOut23_17[4] , \nOut23_17[3] , \nOut23_17[2] , \nOut23_17[1] , 
        \nOut23_17[0] }), .EastIn({\nOut24_16[7] , \nOut24_16[6] , 
        \nOut24_16[5] , \nOut24_16[4] , \nOut24_16[3] , \nOut24_16[2] , 
        \nOut24_16[1] , \nOut24_16[0] }), .WestIn({\nOut22_16[7] , 
        \nOut22_16[6] , \nOut22_16[5] , \nOut22_16[4] , \nOut22_16[3] , 
        \nOut22_16[2] , \nOut22_16[1] , \nOut22_16[0] }), .Out({\nOut23_16[7] , 
        \nOut23_16[6] , \nOut23_16[5] , \nOut23_16[4] , \nOut23_16[3] , 
        \nOut23_16[2] , \nOut23_16[1] , \nOut23_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_775 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut776[7] , \nScanOut776[6] , 
        \nScanOut776[5] , \nScanOut776[4] , \nScanOut776[3] , \nScanOut776[2] , 
        \nScanOut776[1] , \nScanOut776[0] }), .ScanOut({\nScanOut775[7] , 
        \nScanOut775[6] , \nScanOut775[5] , \nScanOut775[4] , \nScanOut775[3] , 
        \nScanOut775[2] , \nScanOut775[1] , \nScanOut775[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_6[7] , \nOut24_6[6] , \nOut24_6[5] , \nOut24_6[4] , 
        \nOut24_6[3] , \nOut24_6[2] , \nOut24_6[1] , \nOut24_6[0] }), 
        .SouthIn({\nOut24_8[7] , \nOut24_8[6] , \nOut24_8[5] , \nOut24_8[4] , 
        \nOut24_8[3] , \nOut24_8[2] , \nOut24_8[1] , \nOut24_8[0] }), .EastIn(
        {\nOut25_7[7] , \nOut25_7[6] , \nOut25_7[5] , \nOut25_7[4] , 
        \nOut25_7[3] , \nOut25_7[2] , \nOut25_7[1] , \nOut25_7[0] }), .WestIn(
        {\nOut23_7[7] , \nOut23_7[6] , \nOut23_7[5] , \nOut23_7[4] , 
        \nOut23_7[3] , \nOut23_7[2] , \nOut23_7[1] , \nOut23_7[0] }), .Out({
        \nOut24_7[7] , \nOut24_7[6] , \nOut24_7[5] , \nOut24_7[4] , 
        \nOut24_7[3] , \nOut24_7[2] , \nOut24_7[1] , \nOut24_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_273 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut274[7] , \nScanOut274[6] , 
        \nScanOut274[5] , \nScanOut274[4] , \nScanOut274[3] , \nScanOut274[2] , 
        \nScanOut274[1] , \nScanOut274[0] }), .ScanOut({\nScanOut273[7] , 
        \nScanOut273[6] , \nScanOut273[5] , \nScanOut273[4] , \nScanOut273[3] , 
        \nScanOut273[2] , \nScanOut273[1] , \nScanOut273[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_16[7] , \nOut8_16[6] , \nOut8_16[5] , \nOut8_16[4] , 
        \nOut8_16[3] , \nOut8_16[2] , \nOut8_16[1] , \nOut8_16[0] }), 
        .SouthIn({\nOut8_18[7] , \nOut8_18[6] , \nOut8_18[5] , \nOut8_18[4] , 
        \nOut8_18[3] , \nOut8_18[2] , \nOut8_18[1] , \nOut8_18[0] }), .EastIn(
        {\nOut9_17[7] , \nOut9_17[6] , \nOut9_17[5] , \nOut9_17[4] , 
        \nOut9_17[3] , \nOut9_17[2] , \nOut9_17[1] , \nOut9_17[0] }), .WestIn(
        {\nOut7_17[7] , \nOut7_17[6] , \nOut7_17[5] , \nOut7_17[4] , 
        \nOut7_17[3] , \nOut7_17[2] , \nOut7_17[1] , \nOut7_17[0] }), .Out({
        \nOut8_17[7] , \nOut8_17[6] , \nOut8_17[5] , \nOut8_17[4] , 
        \nOut8_17[3] , \nOut8_17[2] , \nOut8_17[1] , \nOut8_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_462 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut463[7] , \nScanOut463[6] , 
        \nScanOut463[5] , \nScanOut463[4] , \nScanOut463[3] , \nScanOut463[2] , 
        \nScanOut463[1] , \nScanOut463[0] }), .ScanOut({\nScanOut462[7] , 
        \nScanOut462[6] , \nScanOut462[5] , \nScanOut462[4] , \nScanOut462[3] , 
        \nScanOut462[2] , \nScanOut462[1] , \nScanOut462[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_13[7] , \nOut14_13[6] , \nOut14_13[5] , \nOut14_13[4] , 
        \nOut14_13[3] , \nOut14_13[2] , \nOut14_13[1] , \nOut14_13[0] }), 
        .SouthIn({\nOut14_15[7] , \nOut14_15[6] , \nOut14_15[5] , 
        \nOut14_15[4] , \nOut14_15[3] , \nOut14_15[2] , \nOut14_15[1] , 
        \nOut14_15[0] }), .EastIn({\nOut15_14[7] , \nOut15_14[6] , 
        \nOut15_14[5] , \nOut15_14[4] , \nOut15_14[3] , \nOut15_14[2] , 
        \nOut15_14[1] , \nOut15_14[0] }), .WestIn({\nOut13_14[7] , 
        \nOut13_14[6] , \nOut13_14[5] , \nOut13_14[4] , \nOut13_14[3] , 
        \nOut13_14[2] , \nOut13_14[1] , \nOut13_14[0] }), .Out({\nOut14_14[7] , 
        \nOut14_14[6] , \nOut14_14[5] , \nOut14_14[4] , \nOut14_14[3] , 
        \nOut14_14[2] , \nOut14_14[1] , \nOut14_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_810 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut811[7] , \nScanOut811[6] , 
        \nScanOut811[5] , \nScanOut811[4] , \nScanOut811[3] , \nScanOut811[2] , 
        \nScanOut811[1] , \nScanOut811[0] }), .ScanOut({\nScanOut810[7] , 
        \nScanOut810[6] , \nScanOut810[5] , \nScanOut810[4] , \nScanOut810[3] , 
        \nScanOut810[2] , \nScanOut810[1] , \nScanOut810[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_9[7] , \nOut25_9[6] , \nOut25_9[5] , \nOut25_9[4] , 
        \nOut25_9[3] , \nOut25_9[2] , \nOut25_9[1] , \nOut25_9[0] }), 
        .SouthIn({\nOut25_11[7] , \nOut25_11[6] , \nOut25_11[5] , 
        \nOut25_11[4] , \nOut25_11[3] , \nOut25_11[2] , \nOut25_11[1] , 
        \nOut25_11[0] }), .EastIn({\nOut26_10[7] , \nOut26_10[6] , 
        \nOut26_10[5] , \nOut26_10[4] , \nOut26_10[3] , \nOut26_10[2] , 
        \nOut26_10[1] , \nOut26_10[0] }), .WestIn({\nOut24_10[7] , 
        \nOut24_10[6] , \nOut24_10[5] , \nOut24_10[4] , \nOut24_10[3] , 
        \nOut24_10[2] , \nOut24_10[1] , \nOut24_10[0] }), .Out({\nOut25_10[7] , 
        \nOut25_10[6] , \nOut25_10[5] , \nOut25_10[4] , \nOut25_10[3] , 
        \nOut25_10[2] , \nOut25_10[1] , \nOut25_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_980 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut981[7] , \nScanOut981[6] , 
        \nScanOut981[5] , \nScanOut981[4] , \nScanOut981[3] , \nScanOut981[2] , 
        \nScanOut981[1] , \nScanOut981[0] }), .ScanOut({\nScanOut980[7] , 
        \nScanOut980[6] , \nScanOut980[5] , \nScanOut980[4] , \nScanOut980[3] , 
        \nScanOut980[2] , \nScanOut980[1] , \nScanOut980[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_19[7] , \nOut30_19[6] , \nOut30_19[5] , \nOut30_19[4] , 
        \nOut30_19[3] , \nOut30_19[2] , \nOut30_19[1] , \nOut30_19[0] }), 
        .SouthIn({\nOut30_21[7] , \nOut30_21[6] , \nOut30_21[5] , 
        \nOut30_21[4] , \nOut30_21[3] , \nOut30_21[2] , \nOut30_21[1] , 
        \nOut30_21[0] }), .EastIn({\nOut31_20[7] , \nOut31_20[6] , 
        \nOut31_20[5] , \nOut31_20[4] , \nOut31_20[3] , \nOut31_20[2] , 
        \nOut31_20[1] , \nOut31_20[0] }), .WestIn({\nOut29_20[7] , 
        \nOut29_20[6] , \nOut29_20[5] , \nOut29_20[4] , \nOut29_20[3] , 
        \nOut29_20[2] , \nOut29_20[1] , \nOut29_20[0] }), .Out({\nOut30_20[7] , 
        \nOut30_20[6] , \nOut30_20[5] , \nOut30_20[4] , \nOut30_20[3] , 
        \nOut30_20[2] , \nOut30_20[1] , \nOut30_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_859 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut860[7] , \nScanOut860[6] , 
        \nScanOut860[5] , \nScanOut860[4] , \nScanOut860[3] , \nScanOut860[2] , 
        \nScanOut860[1] , \nScanOut860[0] }), .ScanOut({\nScanOut859[7] , 
        \nScanOut859[6] , \nScanOut859[5] , \nScanOut859[4] , \nScanOut859[3] , 
        \nScanOut859[2] , \nScanOut859[1] , \nScanOut859[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_26[7] , \nOut26_26[6] , \nOut26_26[5] , \nOut26_26[4] , 
        \nOut26_26[3] , \nOut26_26[2] , \nOut26_26[1] , \nOut26_26[0] }), 
        .SouthIn({\nOut26_28[7] , \nOut26_28[6] , \nOut26_28[5] , 
        \nOut26_28[4] , \nOut26_28[3] , \nOut26_28[2] , \nOut26_28[1] , 
        \nOut26_28[0] }), .EastIn({\nOut27_27[7] , \nOut27_27[6] , 
        \nOut27_27[5] , \nOut27_27[4] , \nOut27_27[3] , \nOut27_27[2] , 
        \nOut27_27[1] , \nOut27_27[0] }), .WestIn({\nOut25_27[7] , 
        \nOut25_27[6] , \nOut25_27[5] , \nOut25_27[4] , \nOut25_27[3] , 
        \nOut25_27[2] , \nOut25_27[1] , \nOut25_27[0] }), .Out({\nOut26_27[7] , 
        \nOut26_27[6] , \nOut26_27[5] , \nOut26_27[4] , \nOut26_27[3] , 
        \nOut26_27[2] , \nOut26_27[1] , \nOut26_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_296 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut297[7] , \nScanOut297[6] , 
        \nScanOut297[5] , \nScanOut297[4] , \nScanOut297[3] , \nScanOut297[2] , 
        \nScanOut297[1] , \nScanOut297[0] }), .ScanOut({\nScanOut296[7] , 
        \nScanOut296[6] , \nScanOut296[5] , \nScanOut296[4] , \nScanOut296[3] , 
        \nScanOut296[2] , \nScanOut296[1] , \nScanOut296[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_7[7] , \nOut9_7[6] , \nOut9_7[5] , \nOut9_7[4] , \nOut9_7[3] , 
        \nOut9_7[2] , \nOut9_7[1] , \nOut9_7[0] }), .SouthIn({\nOut9_9[7] , 
        \nOut9_9[6] , \nOut9_9[5] , \nOut9_9[4] , \nOut9_9[3] , \nOut9_9[2] , 
        \nOut9_9[1] , \nOut9_9[0] }), .EastIn({\nOut10_8[7] , \nOut10_8[6] , 
        \nOut10_8[5] , \nOut10_8[4] , \nOut10_8[3] , \nOut10_8[2] , 
        \nOut10_8[1] , \nOut10_8[0] }), .WestIn({\nOut8_8[7] , \nOut8_8[6] , 
        \nOut8_8[5] , \nOut8_8[4] , \nOut8_8[3] , \nOut8_8[2] , \nOut8_8[1] , 
        \nOut8_8[0] }), .Out({\nOut9_8[7] , \nOut9_8[6] , \nOut9_8[5] , 
        \nOut9_8[4] , \nOut9_8[3] , \nOut9_8[2] , \nOut9_8[1] , \nOut9_8[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_627 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut628[7] , \nScanOut628[6] , 
        \nScanOut628[5] , \nScanOut628[4] , \nScanOut628[3] , \nScanOut628[2] , 
        \nScanOut628[1] , \nScanOut628[0] }), .ScanOut({\nScanOut627[7] , 
        \nScanOut627[6] , \nScanOut627[5] , \nScanOut627[4] , \nScanOut627[3] , 
        \nScanOut627[2] , \nScanOut627[1] , \nScanOut627[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_18[7] , \nOut19_18[6] , \nOut19_18[5] , \nOut19_18[4] , 
        \nOut19_18[3] , \nOut19_18[2] , \nOut19_18[1] , \nOut19_18[0] }), 
        .SouthIn({\nOut19_20[7] , \nOut19_20[6] , \nOut19_20[5] , 
        \nOut19_20[4] , \nOut19_20[3] , \nOut19_20[2] , \nOut19_20[1] , 
        \nOut19_20[0] }), .EastIn({\nOut20_19[7] , \nOut20_19[6] , 
        \nOut20_19[5] , \nOut20_19[4] , \nOut20_19[3] , \nOut20_19[2] , 
        \nOut20_19[1] , \nOut20_19[0] }), .WestIn({\nOut18_19[7] , 
        \nOut18_19[6] , \nOut18_19[5] , \nOut18_19[4] , \nOut18_19[3] , 
        \nOut18_19[2] , \nOut18_19[1] , \nOut18_19[0] }), .Out({\nOut19_19[7] , 
        \nOut19_19[6] , \nOut19_19[5] , \nOut19_19[4] , \nOut19_19[3] , 
        \nOut19_19[2] , \nOut19_19[1] , \nOut19_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_965 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut966[7] , \nScanOut966[6] , 
        \nScanOut966[5] , \nScanOut966[4] , \nScanOut966[3] , \nScanOut966[2] , 
        \nScanOut966[1] , \nScanOut966[0] }), .ScanOut({\nScanOut965[7] , 
        \nScanOut965[6] , \nScanOut965[5] , \nScanOut965[4] , \nScanOut965[3] , 
        \nScanOut965[2] , \nScanOut965[1] , \nScanOut965[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_4[7] , \nOut30_4[6] , \nOut30_4[5] , \nOut30_4[4] , 
        \nOut30_4[3] , \nOut30_4[2] , \nOut30_4[1] , \nOut30_4[0] }), 
        .SouthIn({\nOut30_6[7] , \nOut30_6[6] , \nOut30_6[5] , \nOut30_6[4] , 
        \nOut30_6[3] , \nOut30_6[2] , \nOut30_6[1] , \nOut30_6[0] }), .EastIn(
        {\nOut31_5[7] , \nOut31_5[6] , \nOut31_5[5] , \nOut31_5[4] , 
        \nOut31_5[3] , \nOut31_5[2] , \nOut31_5[1] , \nOut31_5[0] }), .WestIn(
        {\nOut29_5[7] , \nOut29_5[6] , \nOut29_5[5] , \nOut29_5[4] , 
        \nOut29_5[3] , \nOut29_5[2] , \nOut29_5[1] , \nOut29_5[0] }), .Out({
        \nOut30_5[7] , \nOut30_5[6] , \nOut30_5[5] , \nOut30_5[4] , 
        \nOut30_5[3] , \nOut30_5[2] , \nOut30_5[1] , \nOut30_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_306 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut307[7] , \nScanOut307[6] , 
        \nScanOut307[5] , \nScanOut307[4] , \nScanOut307[3] , \nScanOut307[2] , 
        \nScanOut307[1] , \nScanOut307[0] }), .ScanOut({\nScanOut306[7] , 
        \nScanOut306[6] , \nScanOut306[5] , \nScanOut306[4] , \nScanOut306[3] , 
        \nScanOut306[2] , \nScanOut306[1] , \nScanOut306[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_17[7] , \nOut9_17[6] , \nOut9_17[5] , \nOut9_17[4] , 
        \nOut9_17[3] , \nOut9_17[2] , \nOut9_17[1] , \nOut9_17[0] }), 
        .SouthIn({\nOut9_19[7] , \nOut9_19[6] , \nOut9_19[5] , \nOut9_19[4] , 
        \nOut9_19[3] , \nOut9_19[2] , \nOut9_19[1] , \nOut9_19[0] }), .EastIn(
        {\nOut10_18[7] , \nOut10_18[6] , \nOut10_18[5] , \nOut10_18[4] , 
        \nOut10_18[3] , \nOut10_18[2] , \nOut10_18[1] , \nOut10_18[0] }), 
        .WestIn({\nOut8_18[7] , \nOut8_18[6] , \nOut8_18[5] , \nOut8_18[4] , 
        \nOut8_18[3] , \nOut8_18[2] , \nOut8_18[1] , \nOut8_18[0] }), .Out({
        \nOut9_18[7] , \nOut9_18[6] , \nOut9_18[5] , \nOut9_18[4] , 
        \nOut9_18[3] , \nOut9_18[2] , \nOut9_18[1] , \nOut9_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_517 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut518[7] , \nScanOut518[6] , 
        \nScanOut518[5] , \nScanOut518[4] , \nScanOut518[3] , \nScanOut518[2] , 
        \nScanOut518[1] , \nScanOut518[0] }), .ScanOut({\nScanOut517[7] , 
        \nScanOut517[6] , \nScanOut517[5] , \nScanOut517[4] , \nScanOut517[3] , 
        \nScanOut517[2] , \nScanOut517[1] , \nScanOut517[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_4[7] , \nOut16_4[6] , \nOut16_4[5] , \nOut16_4[4] , 
        \nOut16_4[3] , \nOut16_4[2] , \nOut16_4[1] , \nOut16_4[0] }), 
        .SouthIn({\nOut16_6[7] , \nOut16_6[6] , \nOut16_6[5] , \nOut16_6[4] , 
        \nOut16_6[3] , \nOut16_6[2] , \nOut16_6[1] , \nOut16_6[0] }), .EastIn(
        {\nOut17_5[7] , \nOut17_5[6] , \nOut17_5[5] , \nOut17_5[4] , 
        \nOut17_5[3] , \nOut17_5[2] , \nOut17_5[1] , \nOut17_5[0] }), .WestIn(
        {\nOut15_5[7] , \nOut15_5[6] , \nOut15_5[5] , \nOut15_5[4] , 
        \nOut15_5[3] , \nOut15_5[2] , \nOut15_5[1] , \nOut15_5[0] }), .Out({
        \nOut16_5[7] , \nOut16_5[6] , \nOut16_5[5] , \nOut16_5[4] , 
        \nOut16_5[3] , \nOut16_5[2] , \nOut16_5[1] , \nOut16_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_321 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut322[7] , \nScanOut322[6] , 
        \nScanOut322[5] , \nScanOut322[4] , \nScanOut322[3] , \nScanOut322[2] , 
        \nScanOut322[1] , \nScanOut322[0] }), .ScanOut({\nScanOut321[7] , 
        \nScanOut321[6] , \nScanOut321[5] , \nScanOut321[4] , \nScanOut321[3] , 
        \nScanOut321[2] , \nScanOut321[1] , \nScanOut321[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_0[7] , \nOut10_0[6] , \nOut10_0[5] , \nOut10_0[4] , 
        \nOut10_0[3] , \nOut10_0[2] , \nOut10_0[1] , \nOut10_0[0] }), 
        .SouthIn({\nOut10_2[7] , \nOut10_2[6] , \nOut10_2[5] , \nOut10_2[4] , 
        \nOut10_2[3] , \nOut10_2[2] , \nOut10_2[1] , \nOut10_2[0] }), .EastIn(
        {\nOut11_1[7] , \nOut11_1[6] , \nOut11_1[5] , \nOut11_1[4] , 
        \nOut11_1[3] , \nOut11_1[2] , \nOut11_1[1] , \nOut11_1[0] }), .WestIn(
        {\nOut9_1[7] , \nOut9_1[6] , \nOut9_1[5] , \nOut9_1[4] , \nOut9_1[3] , 
        \nOut9_1[2] , \nOut9_1[1] , \nOut9_1[0] }), .Out({\nOut10_1[7] , 
        \nOut10_1[6] , \nOut10_1[5] , \nOut10_1[4] , \nOut10_1[3] , 
        \nOut10_1[2] , \nOut10_1[1] , \nOut10_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_487 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut488[7] , \nScanOut488[6] , 
        \nScanOut488[5] , \nScanOut488[4] , \nScanOut488[3] , \nScanOut488[2] , 
        \nScanOut488[1] , \nScanOut488[0] }), .ScanOut({\nScanOut487[7] , 
        \nScanOut487[6] , \nScanOut487[5] , \nScanOut487[4] , \nScanOut487[3] , 
        \nScanOut487[2] , \nScanOut487[1] , \nScanOut487[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_6[7] , \nOut15_6[6] , \nOut15_6[5] , \nOut15_6[4] , 
        \nOut15_6[3] , \nOut15_6[2] , \nOut15_6[1] , \nOut15_6[0] }), 
        .SouthIn({\nOut15_8[7] , \nOut15_8[6] , \nOut15_8[5] , \nOut15_8[4] , 
        \nOut15_8[3] , \nOut15_8[2] , \nOut15_8[1] , \nOut15_8[0] }), .EastIn(
        {\nOut16_7[7] , \nOut16_7[6] , \nOut16_7[5] , \nOut16_7[4] , 
        \nOut16_7[3] , \nOut16_7[2] , \nOut16_7[1] , \nOut16_7[0] }), .WestIn(
        {\nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }), .Out({
        \nOut15_7[7] , \nOut15_7[6] , \nOut15_7[5] , \nOut15_7[4] , 
        \nOut15_7[3] , \nOut15_7[2] , \nOut15_7[1] , \nOut15_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_942 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut943[7] , \nScanOut943[6] , 
        \nScanOut943[5] , \nScanOut943[4] , \nScanOut943[3] , \nScanOut943[2] , 
        \nScanOut943[1] , \nScanOut943[0] }), .ScanOut({\nScanOut942[7] , 
        \nScanOut942[6] , \nScanOut942[5] , \nScanOut942[4] , \nScanOut942[3] , 
        \nScanOut942[2] , \nScanOut942[1] , \nScanOut942[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_13[7] , \nOut29_13[6] , \nOut29_13[5] , \nOut29_13[4] , 
        \nOut29_13[3] , \nOut29_13[2] , \nOut29_13[1] , \nOut29_13[0] }), 
        .SouthIn({\nOut29_15[7] , \nOut29_15[6] , \nOut29_15[5] , 
        \nOut29_15[4] , \nOut29_15[3] , \nOut29_15[2] , \nOut29_15[1] , 
        \nOut29_15[0] }), .EastIn({\nOut30_14[7] , \nOut30_14[6] , 
        \nOut30_14[5] , \nOut30_14[4] , \nOut30_14[3] , \nOut30_14[2] , 
        \nOut30_14[1] , \nOut30_14[0] }), .WestIn({\nOut28_14[7] , 
        \nOut28_14[6] , \nOut28_14[5] , \nOut28_14[4] , \nOut28_14[3] , 
        \nOut28_14[2] , \nOut28_14[1] , \nOut28_14[0] }), .Out({\nOut29_14[7] , 
        \nOut29_14[6] , \nOut29_14[5] , \nOut29_14[4] , \nOut29_14[3] , 
        \nOut29_14[2] , \nOut29_14[1] , \nOut29_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_530 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut531[7] , \nScanOut531[6] , 
        \nScanOut531[5] , \nScanOut531[4] , \nScanOut531[3] , \nScanOut531[2] , 
        \nScanOut531[1] , \nScanOut531[0] }), .ScanOut({\nScanOut530[7] , 
        \nScanOut530[6] , \nScanOut530[5] , \nScanOut530[4] , \nScanOut530[3] , 
        \nScanOut530[2] , \nScanOut530[1] , \nScanOut530[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_17[7] , \nOut16_17[6] , \nOut16_17[5] , \nOut16_17[4] , 
        \nOut16_17[3] , \nOut16_17[2] , \nOut16_17[1] , \nOut16_17[0] }), 
        .SouthIn({\nOut16_19[7] , \nOut16_19[6] , \nOut16_19[5] , 
        \nOut16_19[4] , \nOut16_19[3] , \nOut16_19[2] , \nOut16_19[1] , 
        \nOut16_19[0] }), .EastIn({\nOut17_18[7] , \nOut17_18[6] , 
        \nOut17_18[5] , \nOut17_18[4] , \nOut17_18[3] , \nOut17_18[2] , 
        \nOut17_18[1] , \nOut17_18[0] }), .WestIn({\nOut15_18[7] , 
        \nOut15_18[6] , \nOut15_18[5] , \nOut15_18[4] , \nOut15_18[3] , 
        \nOut15_18[2] , \nOut15_18[1] , \nOut15_18[0] }), .Out({\nOut16_18[7] , 
        \nOut16_18[6] , \nOut16_18[5] , \nOut16_18[4] , \nOut16_18[3] , 
        \nOut16_18[2] , \nOut16_18[1] , \nOut16_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_20 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut21[7] , \nScanOut21[6] , 
        \nScanOut21[5] , \nScanOut21[4] , \nScanOut21[3] , \nScanOut21[2] , 
        \nScanOut21[1] , \nScanOut21[0] }), .ScanOut({\nScanOut20[7] , 
        \nScanOut20[6] , \nScanOut20[5] , \nScanOut20[4] , \nScanOut20[3] , 
        \nScanOut20[2] , \nScanOut20[1] , \nScanOut20[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_20[7] , \nOut0_20[6] , 
        \nOut0_20[5] , \nOut0_20[4] , \nOut0_20[3] , \nOut0_20[2] , 
        \nOut0_20[1] , \nOut0_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_181 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut182[7] , \nScanOut182[6] , 
        \nScanOut182[5] , \nScanOut182[4] , \nScanOut182[3] , \nScanOut182[2] , 
        \nScanOut182[1] , \nScanOut182[0] }), .ScanOut({\nScanOut181[7] , 
        \nScanOut181[6] , \nScanOut181[5] , \nScanOut181[4] , \nScanOut181[3] , 
        \nScanOut181[2] , \nScanOut181[1] , \nScanOut181[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_20[7] , \nOut5_20[6] , \nOut5_20[5] , \nOut5_20[4] , 
        \nOut5_20[3] , \nOut5_20[2] , \nOut5_20[1] , \nOut5_20[0] }), 
        .SouthIn({\nOut5_22[7] , \nOut5_22[6] , \nOut5_22[5] , \nOut5_22[4] , 
        \nOut5_22[3] , \nOut5_22[2] , \nOut5_22[1] , \nOut5_22[0] }), .EastIn(
        {\nOut6_21[7] , \nOut6_21[6] , \nOut6_21[5] , \nOut6_21[4] , 
        \nOut6_21[3] , \nOut6_21[2] , \nOut6_21[1] , \nOut6_21[0] }), .WestIn(
        {\nOut4_21[7] , \nOut4_21[6] , \nOut4_21[5] , \nOut4_21[4] , 
        \nOut4_21[3] , \nOut4_21[2] , \nOut4_21[1] , \nOut4_21[0] }), .Out({
        \nOut5_21[7] , \nOut5_21[6] , \nOut5_21[5] , \nOut5_21[4] , 
        \nOut5_21[3] , \nOut5_21[2] , \nOut5_21[1] , \nOut5_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_600 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut601[7] , \nScanOut601[6] , 
        \nScanOut601[5] , \nScanOut601[4] , \nScanOut601[3] , \nScanOut601[2] , 
        \nScanOut601[1] , \nScanOut601[0] }), .ScanOut({\nScanOut600[7] , 
        \nScanOut600[6] , \nScanOut600[5] , \nScanOut600[4] , \nScanOut600[3] , 
        \nScanOut600[2] , \nScanOut600[1] , \nScanOut600[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_23[7] , \nOut18_23[6] , \nOut18_23[5] , \nOut18_23[4] , 
        \nOut18_23[3] , \nOut18_23[2] , \nOut18_23[1] , \nOut18_23[0] }), 
        .SouthIn({\nOut18_25[7] , \nOut18_25[6] , \nOut18_25[5] , 
        \nOut18_25[4] , \nOut18_25[3] , \nOut18_25[2] , \nOut18_25[1] , 
        \nOut18_25[0] }), .EastIn({\nOut19_24[7] , \nOut19_24[6] , 
        \nOut19_24[5] , \nOut19_24[4] , \nOut19_24[3] , \nOut19_24[2] , 
        \nOut19_24[1] , \nOut19_24[0] }), .WestIn({\nOut17_24[7] , 
        \nOut17_24[6] , \nOut17_24[5] , \nOut17_24[4] , \nOut17_24[3] , 
        \nOut17_24[2] , \nOut17_24[1] , \nOut17_24[0] }), .Out({\nOut18_24[7] , 
        \nOut18_24[6] , \nOut18_24[5] , \nOut18_24[4] , \nOut18_24[3] , 
        \nOut18_24[2] , \nOut18_24[1] , \nOut18_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_790 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut791[7] , \nScanOut791[6] , 
        \nScanOut791[5] , \nScanOut791[4] , \nScanOut791[3] , \nScanOut791[2] , 
        \nScanOut791[1] , \nScanOut791[0] }), .ScanOut({\nScanOut790[7] , 
        \nScanOut790[6] , \nScanOut790[5] , \nScanOut790[4] , \nScanOut790[3] , 
        \nScanOut790[2] , \nScanOut790[1] , \nScanOut790[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_21[7] , \nOut24_21[6] , \nOut24_21[5] , \nOut24_21[4] , 
        \nOut24_21[3] , \nOut24_21[2] , \nOut24_21[1] , \nOut24_21[0] }), 
        .SouthIn({\nOut24_23[7] , \nOut24_23[6] , \nOut24_23[5] , 
        \nOut24_23[4] , \nOut24_23[3] , \nOut24_23[2] , \nOut24_23[1] , 
        \nOut24_23[0] }), .EastIn({\nOut25_22[7] , \nOut25_22[6] , 
        \nOut25_22[5] , \nOut25_22[4] , \nOut25_22[3] , \nOut25_22[2] , 
        \nOut25_22[1] , \nOut25_22[0] }), .WestIn({\nOut23_22[7] , 
        \nOut23_22[6] , \nOut23_22[5] , \nOut23_22[4] , \nOut23_22[3] , 
        \nOut23_22[2] , \nOut23_22[1] , \nOut23_22[0] }), .Out({\nOut24_22[7] , 
        \nOut24_22[6] , \nOut24_22[5] , \nOut24_22[4] , \nOut24_22[3] , 
        \nOut24_22[2] , \nOut24_22[1] , \nOut24_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_69 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut70[7] , \nScanOut70[6] , 
        \nScanOut70[5] , \nScanOut70[4] , \nScanOut70[3] , \nScanOut70[2] , 
        \nScanOut70[1] , \nScanOut70[0] }), .ScanOut({\nScanOut69[7] , 
        \nScanOut69[6] , \nScanOut69[5] , \nScanOut69[4] , \nScanOut69[3] , 
        \nScanOut69[2] , \nScanOut69[1] , \nScanOut69[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_4[7] , \nOut2_4[6] , \nOut2_4[5] , \nOut2_4[4] , \nOut2_4[3] , 
        \nOut2_4[2] , \nOut2_4[1] , \nOut2_4[0] }), .SouthIn({\nOut2_6[7] , 
        \nOut2_6[6] , \nOut2_6[5] , \nOut2_6[4] , \nOut2_6[3] , \nOut2_6[2] , 
        \nOut2_6[1] , \nOut2_6[0] }), .EastIn({\nOut3_5[7] , \nOut3_5[6] , 
        \nOut3_5[5] , \nOut3_5[4] , \nOut3_5[3] , \nOut3_5[2] , \nOut3_5[1] , 
        \nOut3_5[0] }), .WestIn({\nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , 
        \nOut1_5[4] , \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }), 
        .Out({\nOut2_5[7] , \nOut2_5[6] , \nOut2_5[5] , \nOut2_5[4] , 
        \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , \nOut2_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_118 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut119[7] , \nScanOut119[6] , 
        \nScanOut119[5] , \nScanOut119[4] , \nScanOut119[3] , \nScanOut119[2] , 
        \nScanOut119[1] , \nScanOut119[0] }), .ScanOut({\nScanOut118[7] , 
        \nScanOut118[6] , \nScanOut118[5] , \nScanOut118[4] , \nScanOut118[3] , 
        \nScanOut118[2] , \nScanOut118[1] , \nScanOut118[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_21[7] , \nOut3_21[6] , \nOut3_21[5] , \nOut3_21[4] , 
        \nOut3_21[3] , \nOut3_21[2] , \nOut3_21[1] , \nOut3_21[0] }), 
        .SouthIn({\nOut3_23[7] , \nOut3_23[6] , \nOut3_23[5] , \nOut3_23[4] , 
        \nOut3_23[3] , \nOut3_23[2] , \nOut3_23[1] , \nOut3_23[0] }), .EastIn(
        {\nOut4_22[7] , \nOut4_22[6] , \nOut4_22[5] , \nOut4_22[4] , 
        \nOut4_22[3] , \nOut4_22[2] , \nOut4_22[1] , \nOut4_22[0] }), .WestIn(
        {\nOut2_22[7] , \nOut2_22[6] , \nOut2_22[5] , \nOut2_22[4] , 
        \nOut2_22[3] , \nOut2_22[2] , \nOut2_22[1] , \nOut2_22[0] }), .Out({
        \nOut3_22[7] , \nOut3_22[6] , \nOut3_22[5] , \nOut3_22[4] , 
        \nOut3_22[3] , \nOut3_22[2] , \nOut3_22[1] , \nOut3_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_193 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut194[7] , \nScanOut194[6] , 
        \nScanOut194[5] , \nScanOut194[4] , \nScanOut194[3] , \nScanOut194[2] , 
        \nScanOut194[1] , \nScanOut194[0] }), .ScanOut({\nScanOut193[7] , 
        \nScanOut193[6] , \nScanOut193[5] , \nScanOut193[4] , \nScanOut193[3] , 
        \nScanOut193[2] , \nScanOut193[1] , \nScanOut193[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_0[7] , \nOut6_0[6] , \nOut6_0[5] , \nOut6_0[4] , \nOut6_0[3] , 
        \nOut6_0[2] , \nOut6_0[1] , \nOut6_0[0] }), .SouthIn({\nOut6_2[7] , 
        \nOut6_2[6] , \nOut6_2[5] , \nOut6_2[4] , \nOut6_2[3] , \nOut6_2[2] , 
        \nOut6_2[1] , \nOut6_2[0] }), .EastIn({\nOut7_1[7] , \nOut7_1[6] , 
        \nOut7_1[5] , \nOut7_1[4] , \nOut7_1[3] , \nOut7_1[2] , \nOut7_1[1] , 
        \nOut7_1[0] }), .WestIn({\nOut5_1[7] , \nOut5_1[6] , \nOut5_1[5] , 
        \nOut5_1[4] , \nOut5_1[3] , \nOut5_1[2] , \nOut5_1[1] , \nOut5_1[0] }), 
        .Out({\nOut6_1[7] , \nOut6_1[6] , \nOut6_1[5] , \nOut6_1[4] , 
        \nOut6_1[3] , \nOut6_1[2] , \nOut6_1[1] , \nOut6_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_284 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut285[7] , \nScanOut285[6] , 
        \nScanOut285[5] , \nScanOut285[4] , \nScanOut285[3] , \nScanOut285[2] , 
        \nScanOut285[1] , \nScanOut285[0] }), .ScanOut({\nScanOut284[7] , 
        \nScanOut284[6] , \nScanOut284[5] , \nScanOut284[4] , \nScanOut284[3] , 
        \nScanOut284[2] , \nScanOut284[1] , \nScanOut284[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_27[7] , \nOut8_27[6] , \nOut8_27[5] , \nOut8_27[4] , 
        \nOut8_27[3] , \nOut8_27[2] , \nOut8_27[1] , \nOut8_27[0] }), 
        .SouthIn({\nOut8_29[7] , \nOut8_29[6] , \nOut8_29[5] , \nOut8_29[4] , 
        \nOut8_29[3] , \nOut8_29[2] , \nOut8_29[1] , \nOut8_29[0] }), .EastIn(
        {\nOut9_28[7] , \nOut9_28[6] , \nOut9_28[5] , \nOut9_28[4] , 
        \nOut9_28[3] , \nOut9_28[2] , \nOut9_28[1] , \nOut9_28[0] }), .WestIn(
        {\nOut7_28[7] , \nOut7_28[6] , \nOut7_28[5] , \nOut7_28[4] , 
        \nOut7_28[3] , \nOut7_28[2] , \nOut7_28[1] , \nOut7_28[0] }), .Out({
        \nOut8_28[7] , \nOut8_28[6] , \nOut8_28[5] , \nOut8_28[4] , 
        \nOut8_28[3] , \nOut8_28[2] , \nOut8_28[1] , \nOut8_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_314 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut315[7] , \nScanOut315[6] , 
        \nScanOut315[5] , \nScanOut315[4] , \nScanOut315[3] , \nScanOut315[2] , 
        \nScanOut315[1] , \nScanOut315[0] }), .ScanOut({\nScanOut314[7] , 
        \nScanOut314[6] , \nScanOut314[5] , \nScanOut314[4] , \nScanOut314[3] , 
        \nScanOut314[2] , \nScanOut314[1] , \nScanOut314[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_25[7] , \nOut9_25[6] , \nOut9_25[5] , \nOut9_25[4] , 
        \nOut9_25[3] , \nOut9_25[2] , \nOut9_25[1] , \nOut9_25[0] }), 
        .SouthIn({\nOut9_27[7] , \nOut9_27[6] , \nOut9_27[5] , \nOut9_27[4] , 
        \nOut9_27[3] , \nOut9_27[2] , \nOut9_27[1] , \nOut9_27[0] }), .EastIn(
        {\nOut10_26[7] , \nOut10_26[6] , \nOut10_26[5] , \nOut10_26[4] , 
        \nOut10_26[3] , \nOut10_26[2] , \nOut10_26[1] , \nOut10_26[0] }), 
        .WestIn({\nOut8_26[7] , \nOut8_26[6] , \nOut8_26[5] , \nOut8_26[4] , 
        \nOut8_26[3] , \nOut8_26[2] , \nOut8_26[1] , \nOut8_26[0] }), .Out({
        \nOut9_26[7] , \nOut9_26[6] , \nOut9_26[5] , \nOut9_26[4] , 
        \nOut9_26[3] , \nOut9_26[2] , \nOut9_26[1] , \nOut9_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_635 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut636[7] , \nScanOut636[6] , 
        \nScanOut636[5] , \nScanOut636[4] , \nScanOut636[3] , \nScanOut636[2] , 
        \nScanOut636[1] , \nScanOut636[0] }), .ScanOut({\nScanOut635[7] , 
        \nScanOut635[6] , \nScanOut635[5] , \nScanOut635[4] , \nScanOut635[3] , 
        \nScanOut635[2] , \nScanOut635[1] , \nScanOut635[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_26[7] , \nOut19_26[6] , \nOut19_26[5] , \nOut19_26[4] , 
        \nOut19_26[3] , \nOut19_26[2] , \nOut19_26[1] , \nOut19_26[0] }), 
        .SouthIn({\nOut19_28[7] , \nOut19_28[6] , \nOut19_28[5] , 
        \nOut19_28[4] , \nOut19_28[3] , \nOut19_28[2] , \nOut19_28[1] , 
        \nOut19_28[0] }), .EastIn({\nOut20_27[7] , \nOut20_27[6] , 
        \nOut20_27[5] , \nOut20_27[4] , \nOut20_27[3] , \nOut20_27[2] , 
        \nOut20_27[1] , \nOut20_27[0] }), .WestIn({\nOut18_27[7] , 
        \nOut18_27[6] , \nOut18_27[5] , \nOut18_27[4] , \nOut18_27[3] , 
        \nOut18_27[2] , \nOut18_27[1] , \nOut18_27[0] }), .Out({\nOut19_27[7] , 
        \nOut19_27[6] , \nOut19_27[5] , \nOut19_27[4] , \nOut19_27[3] , 
        \nOut19_27[2] , \nOut19_27[1] , \nOut19_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_495 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut496[7] , \nScanOut496[6] , 
        \nScanOut496[5] , \nScanOut496[4] , \nScanOut496[3] , \nScanOut496[2] , 
        \nScanOut496[1] , \nScanOut496[0] }), .ScanOut({\nScanOut495[7] , 
        \nScanOut495[6] , \nScanOut495[5] , \nScanOut495[4] , \nScanOut495[3] , 
        \nScanOut495[2] , \nScanOut495[1] , \nScanOut495[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_14[7] , \nOut15_14[6] , \nOut15_14[5] , \nOut15_14[4] , 
        \nOut15_14[3] , \nOut15_14[2] , \nOut15_14[1] , \nOut15_14[0] }), 
        .SouthIn({\nOut15_16[7] , \nOut15_16[6] , \nOut15_16[5] , 
        \nOut15_16[4] , \nOut15_16[3] , \nOut15_16[2] , \nOut15_16[1] , 
        \nOut15_16[0] }), .EastIn({\nOut16_15[7] , \nOut16_15[6] , 
        \nOut16_15[5] , \nOut16_15[4] , \nOut16_15[3] , \nOut16_15[2] , 
        \nOut16_15[1] , \nOut16_15[0] }), .WestIn({\nOut14_15[7] , 
        \nOut14_15[6] , \nOut14_15[5] , \nOut14_15[4] , \nOut14_15[3] , 
        \nOut14_15[2] , \nOut14_15[1] , \nOut14_15[0] }), .Out({\nOut15_15[7] , 
        \nOut15_15[6] , \nOut15_15[5] , \nOut15_15[4] , \nOut15_15[3] , 
        \nOut15_15[2] , \nOut15_15[1] , \nOut15_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_333 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut334[7] , \nScanOut334[6] , 
        \nScanOut334[5] , \nScanOut334[4] , \nScanOut334[3] , \nScanOut334[2] , 
        \nScanOut334[1] , \nScanOut334[0] }), .ScanOut({\nScanOut333[7] , 
        \nScanOut333[6] , \nScanOut333[5] , \nScanOut333[4] , \nScanOut333[3] , 
        \nScanOut333[2] , \nScanOut333[1] , \nScanOut333[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_12[7] , \nOut10_12[6] , \nOut10_12[5] , \nOut10_12[4] , 
        \nOut10_12[3] , \nOut10_12[2] , \nOut10_12[1] , \nOut10_12[0] }), 
        .SouthIn({\nOut10_14[7] , \nOut10_14[6] , \nOut10_14[5] , 
        \nOut10_14[4] , \nOut10_14[3] , \nOut10_14[2] , \nOut10_14[1] , 
        \nOut10_14[0] }), .EastIn({\nOut11_13[7] , \nOut11_13[6] , 
        \nOut11_13[5] , \nOut11_13[4] , \nOut11_13[3] , \nOut11_13[2] , 
        \nOut11_13[1] , \nOut11_13[0] }), .WestIn({\nOut9_13[7] , 
        \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , \nOut9_13[3] , 
        \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }), .Out({\nOut10_13[7] , 
        \nOut10_13[6] , \nOut10_13[5] , \nOut10_13[4] , \nOut10_13[3] , 
        \nOut10_13[2] , \nOut10_13[1] , \nOut10_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_505 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut506[7] , \nScanOut506[6] , 
        \nScanOut506[5] , \nScanOut506[4] , \nScanOut506[3] , \nScanOut506[2] , 
        \nScanOut506[1] , \nScanOut506[0] }), .ScanOut({\nScanOut505[7] , 
        \nScanOut505[6] , \nScanOut505[5] , \nScanOut505[4] , \nScanOut505[3] , 
        \nScanOut505[2] , \nScanOut505[1] , \nScanOut505[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_24[7] , \nOut15_24[6] , \nOut15_24[5] , \nOut15_24[4] , 
        \nOut15_24[3] , \nOut15_24[2] , \nOut15_24[1] , \nOut15_24[0] }), 
        .SouthIn({\nOut15_26[7] , \nOut15_26[6] , \nOut15_26[5] , 
        \nOut15_26[4] , \nOut15_26[3] , \nOut15_26[2] , \nOut15_26[1] , 
        \nOut15_26[0] }), .EastIn({\nOut16_25[7] , \nOut16_25[6] , 
        \nOut16_25[5] , \nOut16_25[4] , \nOut16_25[3] , \nOut16_25[2] , 
        \nOut16_25[1] , \nOut16_25[0] }), .WestIn({\nOut14_25[7] , 
        \nOut14_25[6] , \nOut14_25[5] , \nOut14_25[4] , \nOut14_25[3] , 
        \nOut14_25[2] , \nOut14_25[1] , \nOut14_25[0] }), .Out({\nOut15_25[7] , 
        \nOut15_25[6] , \nOut15_25[5] , \nOut15_25[4] , \nOut15_25[3] , 
        \nOut15_25[2] , \nOut15_25[1] , \nOut15_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_522 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut523[7] , \nScanOut523[6] , 
        \nScanOut523[5] , \nScanOut523[4] , \nScanOut523[3] , \nScanOut523[2] , 
        \nScanOut523[1] , \nScanOut523[0] }), .ScanOut({\nScanOut522[7] , 
        \nScanOut522[6] , \nScanOut522[5] , \nScanOut522[4] , \nScanOut522[3] , 
        \nScanOut522[2] , \nScanOut522[1] , \nScanOut522[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_9[7] , \nOut16_9[6] , \nOut16_9[5] , \nOut16_9[4] , 
        \nOut16_9[3] , \nOut16_9[2] , \nOut16_9[1] , \nOut16_9[0] }), 
        .SouthIn({\nOut16_11[7] , \nOut16_11[6] , \nOut16_11[5] , 
        \nOut16_11[4] , \nOut16_11[3] , \nOut16_11[2] , \nOut16_11[1] , 
        \nOut16_11[0] }), .EastIn({\nOut17_10[7] , \nOut17_10[6] , 
        \nOut17_10[5] , \nOut17_10[4] , \nOut17_10[3] , \nOut17_10[2] , 
        \nOut17_10[1] , \nOut17_10[0] }), .WestIn({\nOut15_10[7] , 
        \nOut15_10[6] , \nOut15_10[5] , \nOut15_10[4] , \nOut15_10[3] , 
        \nOut15_10[2] , \nOut15_10[1] , \nOut15_10[0] }), .Out({\nOut16_10[7] , 
        \nOut16_10[6] , \nOut16_10[5] , \nOut16_10[4] , \nOut16_10[3] , 
        \nOut16_10[2] , \nOut16_10[1] , \nOut16_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_977 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut978[7] , \nScanOut978[6] , 
        \nScanOut978[5] , \nScanOut978[4] , \nScanOut978[3] , \nScanOut978[2] , 
        \nScanOut978[1] , \nScanOut978[0] }), .ScanOut({\nScanOut977[7] , 
        \nScanOut977[6] , \nScanOut977[5] , \nScanOut977[4] , \nScanOut977[3] , 
        \nScanOut977[2] , \nScanOut977[1] , \nScanOut977[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_16[7] , \nOut30_16[6] , \nOut30_16[5] , \nOut30_16[4] , 
        \nOut30_16[3] , \nOut30_16[2] , \nOut30_16[1] , \nOut30_16[0] }), 
        .SouthIn({\nOut30_18[7] , \nOut30_18[6] , \nOut30_18[5] , 
        \nOut30_18[4] , \nOut30_18[3] , \nOut30_18[2] , \nOut30_18[1] , 
        \nOut30_18[0] }), .EastIn({\nOut31_17[7] , \nOut31_17[6] , 
        \nOut31_17[5] , \nOut31_17[4] , \nOut31_17[3] , \nOut31_17[2] , 
        \nOut31_17[1] , \nOut31_17[0] }), .WestIn({\nOut29_17[7] , 
        \nOut29_17[6] , \nOut29_17[5] , \nOut29_17[4] , \nOut29_17[3] , 
        \nOut29_17[2] , \nOut29_17[1] , \nOut29_17[0] }), .Out({\nOut30_17[7] , 
        \nOut30_17[6] , \nOut30_17[5] , \nOut30_17[4] , \nOut30_17[3] , 
        \nOut30_17[2] , \nOut30_17[1] , \nOut30_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_612 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut613[7] , \nScanOut613[6] , 
        \nScanOut613[5] , \nScanOut613[4] , \nScanOut613[3] , \nScanOut613[2] , 
        \nScanOut613[1] , \nScanOut613[0] }), .ScanOut({\nScanOut612[7] , 
        \nScanOut612[6] , \nScanOut612[5] , \nScanOut612[4] , \nScanOut612[3] , 
        \nScanOut612[2] , \nScanOut612[1] , \nScanOut612[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_3[7] , \nOut19_3[6] , \nOut19_3[5] , \nOut19_3[4] , 
        \nOut19_3[3] , \nOut19_3[2] , \nOut19_3[1] , \nOut19_3[0] }), 
        .SouthIn({\nOut19_5[7] , \nOut19_5[6] , \nOut19_5[5] , \nOut19_5[4] , 
        \nOut19_5[3] , \nOut19_5[2] , \nOut19_5[1] , \nOut19_5[0] }), .EastIn(
        {\nOut20_4[7] , \nOut20_4[6] , \nOut20_4[5] , \nOut20_4[4] , 
        \nOut20_4[3] , \nOut20_4[2] , \nOut20_4[1] , \nOut20_4[0] }), .WestIn(
        {\nOut18_4[7] , \nOut18_4[6] , \nOut18_4[5] , \nOut18_4[4] , 
        \nOut18_4[3] , \nOut18_4[2] , \nOut18_4[1] , \nOut18_4[0] }), .Out({
        \nOut19_4[7] , \nOut19_4[6] , \nOut19_4[5] , \nOut19_4[4] , 
        \nOut19_4[3] , \nOut19_4[2] , \nOut19_4[1] , \nOut19_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_950 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut951[7] , \nScanOut951[6] , 
        \nScanOut951[5] , \nScanOut951[4] , \nScanOut951[3] , \nScanOut951[2] , 
        \nScanOut951[1] , \nScanOut951[0] }), .ScanOut({\nScanOut950[7] , 
        \nScanOut950[6] , \nScanOut950[5] , \nScanOut950[4] , \nScanOut950[3] , 
        \nScanOut950[2] , \nScanOut950[1] , \nScanOut950[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_21[7] , \nOut29_21[6] , \nOut29_21[5] , \nOut29_21[4] , 
        \nOut29_21[3] , \nOut29_21[2] , \nOut29_21[1] , \nOut29_21[0] }), 
        .SouthIn({\nOut29_23[7] , \nOut29_23[6] , \nOut29_23[5] , 
        \nOut29_23[4] , \nOut29_23[3] , \nOut29_23[2] , \nOut29_23[1] , 
        \nOut29_23[0] }), .EastIn({\nOut30_22[7] , \nOut30_22[6] , 
        \nOut30_22[5] , \nOut30_22[4] , \nOut30_22[3] , \nOut30_22[2] , 
        \nOut30_22[1] , \nOut30_22[0] }), .WestIn({\nOut28_22[7] , 
        \nOut28_22[6] , \nOut28_22[5] , \nOut28_22[4] , \nOut28_22[3] , 
        \nOut28_22[2] , \nOut28_22[1] , \nOut28_22[0] }), .Out({\nOut29_22[7] , 
        \nOut29_22[6] , \nOut29_22[5] , \nOut29_22[4] , \nOut29_22[3] , 
        \nOut29_22[2] , \nOut29_22[1] , \nOut29_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_228 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut229[7] , \nScanOut229[6] , 
        \nScanOut229[5] , \nScanOut229[4] , \nScanOut229[3] , \nScanOut229[2] , 
        \nScanOut229[1] , \nScanOut229[0] }), .ScanOut({\nScanOut228[7] , 
        \nScanOut228[6] , \nScanOut228[5] , \nScanOut228[4] , \nScanOut228[3] , 
        \nScanOut228[2] , \nScanOut228[1] , \nScanOut228[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_3[7] , \nOut7_3[6] , \nOut7_3[5] , \nOut7_3[4] , \nOut7_3[3] , 
        \nOut7_3[2] , \nOut7_3[1] , \nOut7_3[0] }), .SouthIn({\nOut7_5[7] , 
        \nOut7_5[6] , \nOut7_5[5] , \nOut7_5[4] , \nOut7_5[3] , \nOut7_5[2] , 
        \nOut7_5[1] , \nOut7_5[0] }), .EastIn({\nOut8_4[7] , \nOut8_4[6] , 
        \nOut8_4[5] , \nOut8_4[4] , \nOut8_4[3] , \nOut8_4[2] , \nOut8_4[1] , 
        \nOut8_4[0] }), .WestIn({\nOut6_4[7] , \nOut6_4[6] , \nOut6_4[5] , 
        \nOut6_4[4] , \nOut6_4[3] , \nOut6_4[2] , \nOut6_4[1] , \nOut6_4[0] }), 
        .Out({\nOut7_4[7] , \nOut7_4[6] , \nOut7_4[5] , \nOut7_4[4] , 
        \nOut7_4[3] , \nOut7_4[2] , \nOut7_4[1] , \nOut7_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_782 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut783[7] , \nScanOut783[6] , 
        \nScanOut783[5] , \nScanOut783[4] , \nScanOut783[3] , \nScanOut783[2] , 
        \nScanOut783[1] , \nScanOut783[0] }), .ScanOut({\nScanOut782[7] , 
        \nScanOut782[6] , \nScanOut782[5] , \nScanOut782[4] , \nScanOut782[3] , 
        \nScanOut782[2] , \nScanOut782[1] , \nScanOut782[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_13[7] , \nOut24_13[6] , \nOut24_13[5] , \nOut24_13[4] , 
        \nOut24_13[3] , \nOut24_13[2] , \nOut24_13[1] , \nOut24_13[0] }), 
        .SouthIn({\nOut24_15[7] , \nOut24_15[6] , \nOut24_15[5] , 
        \nOut24_15[4] , \nOut24_15[3] , \nOut24_15[2] , \nOut24_15[1] , 
        \nOut24_15[0] }), .EastIn({\nOut25_14[7] , \nOut25_14[6] , 
        \nOut25_14[5] , \nOut25_14[4] , \nOut25_14[3] , \nOut25_14[2] , 
        \nOut25_14[1] , \nOut25_14[0] }), .WestIn({\nOut23_14[7] , 
        \nOut23_14[6] , \nOut23_14[5] , \nOut23_14[4] , \nOut23_14[3] , 
        \nOut23_14[2] , \nOut23_14[1] , \nOut23_14[0] }), .Out({\nOut24_14[7] , 
        \nOut24_14[6] , \nOut24_14[5] , \nOut24_14[4] , \nOut24_14[3] , 
        \nOut24_14[2] , \nOut24_14[1] , \nOut24_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_439 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut440[7] , \nScanOut440[6] , 
        \nScanOut440[5] , \nScanOut440[4] , \nScanOut440[3] , \nScanOut440[2] , 
        \nScanOut440[1] , \nScanOut440[0] }), .ScanOut({\nScanOut439[7] , 
        \nScanOut439[6] , \nScanOut439[5] , \nScanOut439[4] , \nScanOut439[3] , 
        \nScanOut439[2] , \nScanOut439[1] , \nScanOut439[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_22[7] , \nOut13_22[6] , \nOut13_22[5] , \nOut13_22[4] , 
        \nOut13_22[3] , \nOut13_22[2] , \nOut13_22[1] , \nOut13_22[0] }), 
        .SouthIn({\nOut13_24[7] , \nOut13_24[6] , \nOut13_24[5] , 
        \nOut13_24[4] , \nOut13_24[3] , \nOut13_24[2] , \nOut13_24[1] , 
        \nOut13_24[0] }), .EastIn({\nOut14_23[7] , \nOut14_23[6] , 
        \nOut14_23[5] , \nOut14_23[4] , \nOut14_23[3] , \nOut14_23[2] , 
        \nOut14_23[1] , \nOut14_23[0] }), .WestIn({\nOut12_23[7] , 
        \nOut12_23[6] , \nOut12_23[5] , \nOut12_23[4] , \nOut12_23[3] , 
        \nOut12_23[2] , \nOut12_23[1] , \nOut12_23[0] }), .Out({\nOut13_23[7] , 
        \nOut13_23[6] , \nOut13_23[5] , \nOut13_23[4] , \nOut13_23[3] , 
        \nOut13_23[2] , \nOut13_23[1] , \nOut13_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_699 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut700[7] , \nScanOut700[6] , 
        \nScanOut700[5] , \nScanOut700[4] , \nScanOut700[3] , \nScanOut700[2] , 
        \nScanOut700[1] , \nScanOut700[0] }), .ScanOut({\nScanOut699[7] , 
        \nScanOut699[6] , \nScanOut699[5] , \nScanOut699[4] , \nScanOut699[3] , 
        \nScanOut699[2] , \nScanOut699[1] , \nScanOut699[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_26[7] , \nOut21_26[6] , \nOut21_26[5] , \nOut21_26[4] , 
        \nOut21_26[3] , \nOut21_26[2] , \nOut21_26[1] , \nOut21_26[0] }), 
        .SouthIn({\nOut21_28[7] , \nOut21_28[6] , \nOut21_28[5] , 
        \nOut21_28[4] , \nOut21_28[3] , \nOut21_28[2] , \nOut21_28[1] , 
        \nOut21_28[0] }), .EastIn({\nOut22_27[7] , \nOut22_27[6] , 
        \nOut22_27[5] , \nOut22_27[4] , \nOut22_27[3] , \nOut22_27[2] , 
        \nOut22_27[1] , \nOut22_27[0] }), .WestIn({\nOut20_27[7] , 
        \nOut20_27[6] , \nOut20_27[5] , \nOut20_27[4] , \nOut20_27[3] , 
        \nOut20_27[2] , \nOut20_27[1] , \nOut20_27[0] }), .Out({\nOut21_27[7] , 
        \nOut21_27[6] , \nOut21_27[5] , \nOut21_27[4] , \nOut21_27[3] , 
        \nOut21_27[2] , \nOut21_27[1] , \nOut21_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_151 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut152[7] , \nScanOut152[6] , 
        \nScanOut152[5] , \nScanOut152[4] , \nScanOut152[3] , \nScanOut152[2] , 
        \nScanOut152[1] , \nScanOut152[0] }), .ScanOut({\nScanOut151[7] , 
        \nScanOut151[6] , \nScanOut151[5] , \nScanOut151[4] , \nScanOut151[3] , 
        \nScanOut151[2] , \nScanOut151[1] , \nScanOut151[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_22[7] , \nOut4_22[6] , \nOut4_22[5] , \nOut4_22[4] , 
        \nOut4_22[3] , \nOut4_22[2] , \nOut4_22[1] , \nOut4_22[0] }), 
        .SouthIn({\nOut4_24[7] , \nOut4_24[6] , \nOut4_24[5] , \nOut4_24[4] , 
        \nOut4_24[3] , \nOut4_24[2] , \nOut4_24[1] , \nOut4_24[0] }), .EastIn(
        {\nOut5_23[7] , \nOut5_23[6] , \nOut5_23[5] , \nOut5_23[4] , 
        \nOut5_23[3] , \nOut5_23[2] , \nOut5_23[1] , \nOut5_23[0] }), .WestIn(
        {\nOut3_23[7] , \nOut3_23[6] , \nOut3_23[5] , \nOut3_23[4] , 
        \nOut3_23[3] , \nOut3_23[2] , \nOut3_23[1] , \nOut3_23[0] }), .Out({
        \nOut4_23[7] , \nOut4_23[6] , \nOut4_23[5] , \nOut4_23[4] , 
        \nOut4_23[3] , \nOut4_23[2] , \nOut4_23[1] , \nOut4_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_176 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut177[7] , \nScanOut177[6] , 
        \nScanOut177[5] , \nScanOut177[4] , \nScanOut177[3] , \nScanOut177[2] , 
        \nScanOut177[1] , \nScanOut177[0] }), .ScanOut({\nScanOut176[7] , 
        \nScanOut176[6] , \nScanOut176[5] , \nScanOut176[4] , \nScanOut176[3] , 
        \nScanOut176[2] , \nScanOut176[1] , \nScanOut176[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_15[7] , \nOut5_15[6] , \nOut5_15[5] , \nOut5_15[4] , 
        \nOut5_15[3] , \nOut5_15[2] , \nOut5_15[1] , \nOut5_15[0] }), 
        .SouthIn({\nOut5_17[7] , \nOut5_17[6] , \nOut5_17[5] , \nOut5_17[4] , 
        \nOut5_17[3] , \nOut5_17[2] , \nOut5_17[1] , \nOut5_17[0] }), .EastIn(
        {\nOut6_16[7] , \nOut6_16[6] , \nOut6_16[5] , \nOut6_16[4] , 
        \nOut6_16[3] , \nOut6_16[2] , \nOut6_16[1] , \nOut6_16[0] }), .WestIn(
        {\nOut4_16[7] , \nOut4_16[6] , \nOut4_16[5] , \nOut4_16[4] , 
        \nOut4_16[3] , \nOut4_16[2] , \nOut4_16[1] , \nOut4_16[0] }), .Out({
        \nOut5_16[7] , \nOut5_16[6] , \nOut5_16[5] , \nOut5_16[4] , 
        \nOut5_16[3] , \nOut5_16[2] , \nOut5_16[1] , \nOut5_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_246 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut247[7] , \nScanOut247[6] , 
        \nScanOut247[5] , \nScanOut247[4] , \nScanOut247[3] , \nScanOut247[2] , 
        \nScanOut247[1] , \nScanOut247[0] }), .ScanOut({\nScanOut246[7] , 
        \nScanOut246[6] , \nScanOut246[5] , \nScanOut246[4] , \nScanOut246[3] , 
        \nScanOut246[2] , \nScanOut246[1] , \nScanOut246[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_21[7] , \nOut7_21[6] , \nOut7_21[5] , \nOut7_21[4] , 
        \nOut7_21[3] , \nOut7_21[2] , \nOut7_21[1] , \nOut7_21[0] }), 
        .SouthIn({\nOut7_23[7] , \nOut7_23[6] , \nOut7_23[5] , \nOut7_23[4] , 
        \nOut7_23[3] , \nOut7_23[2] , \nOut7_23[1] , \nOut7_23[0] }), .EastIn(
        {\nOut8_22[7] , \nOut8_22[6] , \nOut8_22[5] , \nOut8_22[4] , 
        \nOut8_22[3] , \nOut8_22[2] , \nOut8_22[1] , \nOut8_22[0] }), .WestIn(
        {\nOut6_22[7] , \nOut6_22[6] , \nOut6_22[5] , \nOut6_22[4] , 
        \nOut6_22[3] , \nOut6_22[2] , \nOut6_22[1] , \nOut6_22[0] }), .Out({
        \nOut7_22[7] , \nOut7_22[6] , \nOut7_22[5] , \nOut7_22[4] , 
        \nOut7_22[3] , \nOut7_22[2] , \nOut7_22[1] , \nOut7_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_457 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut458[7] , \nScanOut458[6] , 
        \nScanOut458[5] , \nScanOut458[4] , \nScanOut458[3] , \nScanOut458[2] , 
        \nScanOut458[1] , \nScanOut458[0] }), .ScanOut({\nScanOut457[7] , 
        \nScanOut457[6] , \nScanOut457[5] , \nScanOut457[4] , \nScanOut457[3] , 
        \nScanOut457[2] , \nScanOut457[1] , \nScanOut457[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }), 
        .SouthIn({\nOut14_10[7] , \nOut14_10[6] , \nOut14_10[5] , 
        \nOut14_10[4] , \nOut14_10[3] , \nOut14_10[2] , \nOut14_10[1] , 
        \nOut14_10[0] }), .EastIn({\nOut15_9[7] , \nOut15_9[6] , \nOut15_9[5] , 
        \nOut15_9[4] , \nOut15_9[3] , \nOut15_9[2] , \nOut15_9[1] , 
        \nOut15_9[0] }), .WestIn({\nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , 
        \nOut13_9[4] , \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , 
        \nOut13_9[0] }), .Out({\nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , 
        \nOut14_9[4] , \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , 
        \nOut14_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_709 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut710[7] , \nScanOut710[6] , 
        \nScanOut710[5] , \nScanOut710[4] , \nScanOut710[3] , \nScanOut710[2] , 
        \nScanOut710[1] , \nScanOut710[0] }), .ScanOut({\nScanOut709[7] , 
        \nScanOut709[6] , \nScanOut709[5] , \nScanOut709[4] , \nScanOut709[3] , 
        \nScanOut709[2] , \nScanOut709[1] , \nScanOut709[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_4[7] , \nOut22_4[6] , \nOut22_4[5] , \nOut22_4[4] , 
        \nOut22_4[3] , \nOut22_4[2] , \nOut22_4[1] , \nOut22_4[0] }), 
        .SouthIn({\nOut22_6[7] , \nOut22_6[6] , \nOut22_6[5] , \nOut22_6[4] , 
        \nOut22_6[3] , \nOut22_6[2] , \nOut22_6[1] , \nOut22_6[0] }), .EastIn(
        {\nOut23_5[7] , \nOut23_5[6] , \nOut23_5[5] , \nOut23_5[4] , 
        \nOut23_5[3] , \nOut23_5[2] , \nOut23_5[1] , \nOut23_5[0] }), .WestIn(
        {\nOut21_5[7] , \nOut21_5[6] , \nOut21_5[5] , \nOut21_5[4] , 
        \nOut21_5[3] , \nOut21_5[2] , \nOut21_5[1] , \nOut21_5[0] }), .Out({
        \nOut22_5[7] , \nOut22_5[6] , \nOut22_5[5] , \nOut22_5[4] , 
        \nOut22_5[3] , \nOut22_5[2] , \nOut22_5[1] , \nOut22_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_767 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut768[7] , \nScanOut768[6] , 
        \nScanOut768[5] , \nScanOut768[4] , \nScanOut768[3] , \nScanOut768[2] , 
        \nScanOut768[1] , \nScanOut768[0] }), .ScanOut({\nScanOut767[7] , 
        \nScanOut767[6] , \nScanOut767[5] , \nScanOut767[4] , \nScanOut767[3] , 
        \nScanOut767[2] , \nScanOut767[1] , \nScanOut767[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut23_31[7] , \nOut23_31[6] , 
        \nOut23_31[5] , \nOut23_31[4] , \nOut23_31[3] , \nOut23_31[2] , 
        \nOut23_31[1] , \nOut23_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_825 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut826[7] , \nScanOut826[6] , 
        \nScanOut826[5] , \nScanOut826[4] , \nScanOut826[3] , \nScanOut826[2] , 
        \nScanOut826[1] , \nScanOut826[0] }), .ScanOut({\nScanOut825[7] , 
        \nScanOut825[6] , \nScanOut825[5] , \nScanOut825[4] , \nScanOut825[3] , 
        \nScanOut825[2] , \nScanOut825[1] , \nScanOut825[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_24[7] , \nOut25_24[6] , \nOut25_24[5] , \nOut25_24[4] , 
        \nOut25_24[3] , \nOut25_24[2] , \nOut25_24[1] , \nOut25_24[0] }), 
        .SouthIn({\nOut25_26[7] , \nOut25_26[6] , \nOut25_26[5] , 
        \nOut25_26[4] , \nOut25_26[3] , \nOut25_26[2] , \nOut25_26[1] , 
        \nOut25_26[0] }), .EastIn({\nOut26_25[7] , \nOut26_25[6] , 
        \nOut26_25[5] , \nOut26_25[4] , \nOut26_25[3] , \nOut26_25[2] , 
        \nOut26_25[1] , \nOut26_25[0] }), .WestIn({\nOut24_25[7] , 
        \nOut24_25[6] , \nOut24_25[5] , \nOut24_25[4] , \nOut24_25[3] , 
        \nOut24_25[2] , \nOut24_25[1] , \nOut24_25[0] }), .Out({\nOut25_25[7] , 
        \nOut25_25[6] , \nOut25_25[5] , \nOut25_25[4] , \nOut25_25[3] , 
        \nOut25_25[2] , \nOut25_25[1] , \nOut25_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_261 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut262[7] , \nScanOut262[6] , 
        \nScanOut262[5] , \nScanOut262[4] , \nScanOut262[3] , \nScanOut262[2] , 
        \nScanOut262[1] , \nScanOut262[0] }), .ScanOut({\nScanOut261[7] , 
        \nScanOut261[6] , \nScanOut261[5] , \nScanOut261[4] , \nScanOut261[3] , 
        \nScanOut261[2] , \nScanOut261[1] , \nScanOut261[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_4[7] , \nOut8_4[6] , \nOut8_4[5] , \nOut8_4[4] , \nOut8_4[3] , 
        \nOut8_4[2] , \nOut8_4[1] , \nOut8_4[0] }), .SouthIn({\nOut8_6[7] , 
        \nOut8_6[6] , \nOut8_6[5] , \nOut8_6[4] , \nOut8_6[3] , \nOut8_6[2] , 
        \nOut8_6[1] , \nOut8_6[0] }), .EastIn({\nOut9_5[7] , \nOut9_5[6] , 
        \nOut9_5[5] , \nOut9_5[4] , \nOut9_5[3] , \nOut9_5[2] , \nOut9_5[1] , 
        \nOut9_5[0] }), .WestIn({\nOut7_5[7] , \nOut7_5[6] , \nOut7_5[5] , 
        \nOut7_5[4] , \nOut7_5[3] , \nOut7_5[2] , \nOut7_5[1] , \nOut7_5[0] }), 
        .Out({\nOut8_5[7] , \nOut8_5[6] , \nOut8_5[5] , \nOut8_5[4] , 
        \nOut8_5[3] , \nOut8_5[2] , \nOut8_5[1] , \nOut8_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_740 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut741[7] , \nScanOut741[6] , 
        \nScanOut741[5] , \nScanOut741[4] , \nScanOut741[3] , \nScanOut741[2] , 
        \nScanOut741[1] , \nScanOut741[0] }), .ScanOut({\nScanOut740[7] , 
        \nScanOut740[6] , \nScanOut740[5] , \nScanOut740[4] , \nScanOut740[3] , 
        \nScanOut740[2] , \nScanOut740[1] , \nScanOut740[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_3[7] , \nOut23_3[6] , \nOut23_3[5] , \nOut23_3[4] , 
        \nOut23_3[3] , \nOut23_3[2] , \nOut23_3[1] , \nOut23_3[0] }), 
        .SouthIn({\nOut23_5[7] , \nOut23_5[6] , \nOut23_5[5] , \nOut23_5[4] , 
        \nOut23_5[3] , \nOut23_5[2] , \nOut23_5[1] , \nOut23_5[0] }), .EastIn(
        {\nOut24_4[7] , \nOut24_4[6] , \nOut24_4[5] , \nOut24_4[4] , 
        \nOut24_4[3] , \nOut24_4[2] , \nOut24_4[1] , \nOut24_4[0] }), .WestIn(
        {\nOut22_4[7] , \nOut22_4[6] , \nOut22_4[5] , \nOut22_4[4] , 
        \nOut22_4[3] , \nOut22_4[2] , \nOut22_4[1] , \nOut22_4[0] }), .Out({
        \nOut23_4[7] , \nOut23_4[6] , \nOut23_4[5] , \nOut23_4[4] , 
        \nOut23_4[3] , \nOut23_4[2] , \nOut23_4[1] , \nOut23_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_470 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut471[7] , \nScanOut471[6] , 
        \nScanOut471[5] , \nScanOut471[4] , \nScanOut471[3] , \nScanOut471[2] , 
        \nScanOut471[1] , \nScanOut471[0] }), .ScanOut({\nScanOut470[7] , 
        \nScanOut470[6] , \nScanOut470[5] , \nScanOut470[4] , \nScanOut470[3] , 
        \nScanOut470[2] , \nScanOut470[1] , \nScanOut470[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_21[7] , \nOut14_21[6] , \nOut14_21[5] , \nOut14_21[4] , 
        \nOut14_21[3] , \nOut14_21[2] , \nOut14_21[1] , \nOut14_21[0] }), 
        .SouthIn({\nOut14_23[7] , \nOut14_23[6] , \nOut14_23[5] , 
        \nOut14_23[4] , \nOut14_23[3] , \nOut14_23[2] , \nOut14_23[1] , 
        \nOut14_23[0] }), .EastIn({\nOut15_22[7] , \nOut15_22[6] , 
        \nOut15_22[5] , \nOut15_22[4] , \nOut15_22[3] , \nOut15_22[2] , 
        \nOut15_22[1] , \nOut15_22[0] }), .WestIn({\nOut13_22[7] , 
        \nOut13_22[6] , \nOut13_22[5] , \nOut13_22[4] , \nOut13_22[3] , 
        \nOut13_22[2] , \nOut13_22[1] , \nOut13_22[0] }), .Out({\nOut14_22[7] , 
        \nOut14_22[6] , \nOut14_22[5] , \nOut14_22[4] , \nOut14_22[3] , 
        \nOut14_22[2] , \nOut14_22[1] , \nOut14_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_802 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut803[7] , \nScanOut803[6] , 
        \nScanOut803[5] , \nScanOut803[4] , \nScanOut803[3] , \nScanOut803[2] , 
        \nScanOut803[1] , \nScanOut803[0] }), .ScanOut({\nScanOut802[7] , 
        \nScanOut802[6] , \nScanOut802[5] , \nScanOut802[4] , \nScanOut802[3] , 
        \nScanOut802[2] , \nScanOut802[1] , \nScanOut802[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_1[7] , \nOut25_1[6] , \nOut25_1[5] , \nOut25_1[4] , 
        \nOut25_1[3] , \nOut25_1[2] , \nOut25_1[1] , \nOut25_1[0] }), 
        .SouthIn({\nOut25_3[7] , \nOut25_3[6] , \nOut25_3[5] , \nOut25_3[4] , 
        \nOut25_3[3] , \nOut25_3[2] , \nOut25_3[1] , \nOut25_3[0] }), .EastIn(
        {\nOut26_2[7] , \nOut26_2[6] , \nOut26_2[5] , \nOut26_2[4] , 
        \nOut26_2[3] , \nOut26_2[2] , \nOut26_2[1] , \nOut26_2[0] }), .WestIn(
        {\nOut24_2[7] , \nOut24_2[6] , \nOut24_2[5] , \nOut24_2[4] , 
        \nOut24_2[3] , \nOut24_2[2] , \nOut24_2[1] , \nOut24_2[0] }), .Out({
        \nOut25_2[7] , \nOut25_2[6] , \nOut25_2[5] , \nOut25_2[4] , 
        \nOut25_2[3] , \nOut25_2[2] , \nOut25_2[1] , \nOut25_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_992 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut993[7] , \nScanOut993[6] , 
        \nScanOut993[5] , \nScanOut993[4] , \nScanOut993[3] , \nScanOut993[2] , 
        \nScanOut993[1] , \nScanOut993[0] }), .ScanOut({\nScanOut992[7] , 
        \nScanOut992[6] , \nScanOut992[5] , \nScanOut992[4] , \nScanOut992[3] , 
        \nScanOut992[2] , \nScanOut992[1] , \nScanOut992[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_12 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut13[7] , \nScanOut13[6] , 
        \nScanOut13[5] , \nScanOut13[4] , \nScanOut13[3] , \nScanOut13[2] , 
        \nScanOut13[1] , \nScanOut13[0] }), .ScanOut({\nScanOut12[7] , 
        \nScanOut12[6] , \nScanOut12[5] , \nScanOut12[4] , \nScanOut12[3] , 
        \nScanOut12[2] , \nScanOut12[1] , \nScanOut12[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_12[7] , \nOut0_12[6] , 
        \nOut0_12[5] , \nOut0_12[4] , \nOut0_12[3] , \nOut0_12[2] , 
        \nOut0_12[1] , \nOut0_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_27 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut28[7] , \nScanOut28[6] , 
        \nScanOut28[5] , \nScanOut28[4] , \nScanOut28[3] , \nScanOut28[2] , 
        \nScanOut28[1] , \nScanOut28[0] }), .ScanOut({\nScanOut27[7] , 
        \nScanOut27[6] , \nScanOut27[5] , \nScanOut27[4] , \nScanOut27[3] , 
        \nScanOut27[2] , \nScanOut27[1] , \nScanOut27[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_27[7] , \nOut0_27[6] , 
        \nOut0_27[5] , \nOut0_27[4] , \nOut0_27[3] , \nOut0_27[2] , 
        \nOut0_27[1] , \nOut0_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_49 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut50[7] , \nScanOut50[6] , 
        \nScanOut50[5] , \nScanOut50[4] , \nScanOut50[3] , \nScanOut50[2] , 
        \nScanOut50[1] , \nScanOut50[0] }), .ScanOut({\nScanOut49[7] , 
        \nScanOut49[6] , \nScanOut49[5] , \nScanOut49[4] , \nScanOut49[3] , 
        \nScanOut49[2] , \nScanOut49[1] , \nScanOut49[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_16[7] , \nOut1_16[6] , \nOut1_16[5] , \nOut1_16[4] , 
        \nOut1_16[3] , \nOut1_16[2] , \nOut1_16[1] , \nOut1_16[0] }), 
        .SouthIn({\nOut1_18[7] , \nOut1_18[6] , \nOut1_18[5] , \nOut1_18[4] , 
        \nOut1_18[3] , \nOut1_18[2] , \nOut1_18[1] , \nOut1_18[0] }), .EastIn(
        {\nOut2_17[7] , \nOut2_17[6] , \nOut2_17[5] , \nOut2_17[4] , 
        \nOut2_17[3] , \nOut2_17[2] , \nOut2_17[1] , \nOut2_17[0] }), .WestIn(
        {\nOut0_17[7] , \nOut0_17[6] , \nOut0_17[5] , \nOut0_17[4] , 
        \nOut0_17[3] , \nOut0_17[2] , \nOut0_17[1] , \nOut0_17[0] }), .Out({
        \nOut1_17[7] , \nOut1_17[6] , \nOut1_17[5] , \nOut1_17[4] , 
        \nOut1_17[3] , \nOut1_17[2] , \nOut1_17[1] , \nOut1_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_52 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut53[7] , \nScanOut53[6] , 
        \nScanOut53[5] , \nScanOut53[4] , \nScanOut53[3] , \nScanOut53[2] , 
        \nScanOut53[1] , \nScanOut53[0] }), .ScanOut({\nScanOut52[7] , 
        \nScanOut52[6] , \nScanOut52[5] , \nScanOut52[4] , \nScanOut52[3] , 
        \nScanOut52[2] , \nScanOut52[1] , \nScanOut52[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_19[7] , \nOut1_19[6] , \nOut1_19[5] , \nOut1_19[4] , 
        \nOut1_19[3] , \nOut1_19[2] , \nOut1_19[1] , \nOut1_19[0] }), 
        .SouthIn({\nOut1_21[7] , \nOut1_21[6] , \nOut1_21[5] , \nOut1_21[4] , 
        \nOut1_21[3] , \nOut1_21[2] , \nOut1_21[1] , \nOut1_21[0] }), .EastIn(
        {\nOut2_20[7] , \nOut2_20[6] , \nOut2_20[5] , \nOut2_20[4] , 
        \nOut2_20[3] , \nOut2_20[2] , \nOut2_20[1] , \nOut2_20[0] }), .WestIn(
        {\nOut0_20[7] , \nOut0_20[6] , \nOut0_20[5] , \nOut0_20[4] , 
        \nOut0_20[3] , \nOut0_20[2] , \nOut0_20[1] , \nOut0_20[0] }), .Out({
        \nOut1_20[7] , \nOut1_20[6] , \nOut1_20[5] , \nOut1_20[4] , 
        \nOut1_20[3] , \nOut1_20[2] , \nOut1_20[1] , \nOut1_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_55 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut56[7] , \nScanOut56[6] , 
        \nScanOut56[5] , \nScanOut56[4] , \nScanOut56[3] , \nScanOut56[2] , 
        \nScanOut56[1] , \nScanOut56[0] }), .ScanOut({\nScanOut55[7] , 
        \nScanOut55[6] , \nScanOut55[5] , \nScanOut55[4] , \nScanOut55[3] , 
        \nScanOut55[2] , \nScanOut55[1] , \nScanOut55[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_22[7] , \nOut1_22[6] , \nOut1_22[5] , \nOut1_22[4] , 
        \nOut1_22[3] , \nOut1_22[2] , \nOut1_22[1] , \nOut1_22[0] }), 
        .SouthIn({\nOut1_24[7] , \nOut1_24[6] , \nOut1_24[5] , \nOut1_24[4] , 
        \nOut1_24[3] , \nOut1_24[2] , \nOut1_24[1] , \nOut1_24[0] }), .EastIn(
        {\nOut2_23[7] , \nOut2_23[6] , \nOut2_23[5] , \nOut2_23[4] , 
        \nOut2_23[3] , \nOut2_23[2] , \nOut2_23[1] , \nOut2_23[0] }), .WestIn(
        {\nOut0_23[7] , \nOut0_23[6] , \nOut0_23[5] , \nOut0_23[4] , 
        \nOut0_23[3] , \nOut0_23[2] , \nOut0_23[1] , \nOut0_23[0] }), .Out({
        \nOut1_23[7] , \nOut1_23[6] , \nOut1_23[5] , \nOut1_23[4] , 
        \nOut1_23[3] , \nOut1_23[2] , \nOut1_23[1] , \nOut1_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_361 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut362[7] , \nScanOut362[6] , 
        \nScanOut362[5] , \nScanOut362[4] , \nScanOut362[3] , \nScanOut362[2] , 
        \nScanOut362[1] , \nScanOut362[0] }), .ScanOut({\nScanOut361[7] , 
        \nScanOut361[6] , \nScanOut361[5] , \nScanOut361[4] , \nScanOut361[3] , 
        \nScanOut361[2] , \nScanOut361[1] , \nScanOut361[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }), 
        .SouthIn({\nOut11_10[7] , \nOut11_10[6] , \nOut11_10[5] , 
        \nOut11_10[4] , \nOut11_10[3] , \nOut11_10[2] , \nOut11_10[1] , 
        \nOut11_10[0] }), .EastIn({\nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , 
        \nOut12_9[4] , \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , 
        \nOut12_9[0] }), .WestIn({\nOut10_9[7] , \nOut10_9[6] , \nOut10_9[5] , 
        \nOut10_9[4] , \nOut10_9[3] , \nOut10_9[2] , \nOut10_9[1] , 
        \nOut10_9[0] }), .Out({\nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , 
        \nOut11_9[4] , \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , 
        \nOut11_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_570 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut571[7] , \nScanOut571[6] , 
        \nScanOut571[5] , \nScanOut571[4] , \nScanOut571[3] , \nScanOut571[2] , 
        \nScanOut571[1] , \nScanOut571[0] }), .ScanOut({\nScanOut570[7] , 
        \nScanOut570[6] , \nScanOut570[5] , \nScanOut570[4] , \nScanOut570[3] , 
        \nScanOut570[2] , \nScanOut570[1] , \nScanOut570[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_25[7] , \nOut17_25[6] , \nOut17_25[5] , \nOut17_25[4] , 
        \nOut17_25[3] , \nOut17_25[2] , \nOut17_25[1] , \nOut17_25[0] }), 
        .SouthIn({\nOut17_27[7] , \nOut17_27[6] , \nOut17_27[5] , 
        \nOut17_27[4] , \nOut17_27[3] , \nOut17_27[2] , \nOut17_27[1] , 
        \nOut17_27[0] }), .EastIn({\nOut18_26[7] , \nOut18_26[6] , 
        \nOut18_26[5] , \nOut18_26[4] , \nOut18_26[3] , \nOut18_26[2] , 
        \nOut18_26[1] , \nOut18_26[0] }), .WestIn({\nOut16_26[7] , 
        \nOut16_26[6] , \nOut16_26[5] , \nOut16_26[4] , \nOut16_26[3] , 
        \nOut16_26[2] , \nOut16_26[1] , \nOut16_26[0] }), .Out({\nOut17_26[7] , 
        \nOut17_26[6] , \nOut17_26[5] , \nOut17_26[4] , \nOut17_26[3] , 
        \nOut17_26[2] , \nOut17_26[1] , \nOut17_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_889 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut890[7] , \nScanOut890[6] , 
        \nScanOut890[5] , \nScanOut890[4] , \nScanOut890[3] , \nScanOut890[2] , 
        \nScanOut890[1] , \nScanOut890[0] }), .ScanOut({\nScanOut889[7] , 
        \nScanOut889[6] , \nScanOut889[5] , \nScanOut889[4] , \nScanOut889[3] , 
        \nScanOut889[2] , \nScanOut889[1] , \nScanOut889[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_24[7] , \nOut27_24[6] , \nOut27_24[5] , \nOut27_24[4] , 
        \nOut27_24[3] , \nOut27_24[2] , \nOut27_24[1] , \nOut27_24[0] }), 
        .SouthIn({\nOut27_26[7] , \nOut27_26[6] , \nOut27_26[5] , 
        \nOut27_26[4] , \nOut27_26[3] , \nOut27_26[2] , \nOut27_26[1] , 
        \nOut27_26[0] }), .EastIn({\nOut28_25[7] , \nOut28_25[6] , 
        \nOut28_25[5] , \nOut28_25[4] , \nOut28_25[3] , \nOut28_25[2] , 
        \nOut28_25[1] , \nOut28_25[0] }), .WestIn({\nOut26_25[7] , 
        \nOut26_25[6] , \nOut26_25[5] , \nOut26_25[4] , \nOut26_25[3] , 
        \nOut26_25[2] , \nOut26_25[1] , \nOut26_25[0] }), .Out({\nOut27_25[7] , 
        \nOut27_25[6] , \nOut27_25[5] , \nOut27_25[4] , \nOut27_25[3] , 
        \nOut27_25[2] , \nOut27_25[1] , \nOut27_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_919 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut920[7] , \nScanOut920[6] , 
        \nScanOut920[5] , \nScanOut920[4] , \nScanOut920[3] , \nScanOut920[2] , 
        \nScanOut920[1] , \nScanOut920[0] }), .ScanOut({\nScanOut919[7] , 
        \nScanOut919[6] , \nScanOut919[5] , \nScanOut919[4] , \nScanOut919[3] , 
        \nScanOut919[2] , \nScanOut919[1] , \nScanOut919[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_22[7] , \nOut28_22[6] , \nOut28_22[5] , \nOut28_22[4] , 
        \nOut28_22[3] , \nOut28_22[2] , \nOut28_22[1] , \nOut28_22[0] }), 
        .SouthIn({\nOut28_24[7] , \nOut28_24[6] , \nOut28_24[5] , 
        \nOut28_24[4] , \nOut28_24[3] , \nOut28_24[2] , \nOut28_24[1] , 
        \nOut28_24[0] }), .EastIn({\nOut29_23[7] , \nOut29_23[6] , 
        \nOut29_23[5] , \nOut29_23[4] , \nOut29_23[3] , \nOut29_23[2] , 
        \nOut29_23[1] , \nOut29_23[0] }), .WestIn({\nOut27_23[7] , 
        \nOut27_23[6] , \nOut27_23[5] , \nOut27_23[4] , \nOut27_23[3] , 
        \nOut27_23[2] , \nOut27_23[1] , \nOut27_23[0] }), .Out({\nOut28_23[7] , 
        \nOut28_23[6] , \nOut28_23[5] , \nOut28_23[4] , \nOut28_23[3] , 
        \nOut28_23[2] , \nOut28_23[1] , \nOut28_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_640 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut641[7] , \nScanOut641[6] , 
        \nScanOut641[5] , \nScanOut641[4] , \nScanOut641[3] , \nScanOut641[2] , 
        \nScanOut641[1] , \nScanOut641[0] }), .ScanOut({\nScanOut640[7] , 
        \nScanOut640[6] , \nScanOut640[5] , \nScanOut640[4] , \nScanOut640[3] , 
        \nScanOut640[2] , \nScanOut640[1] , \nScanOut640[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut20_0[7] , \nOut20_0[6] , 
        \nOut20_0[5] , \nOut20_0[4] , \nOut20_0[3] , \nOut20_0[2] , 
        \nOut20_0[1] , \nOut20_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_892 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut893[7] , \nScanOut893[6] , 
        \nScanOut893[5] , \nScanOut893[4] , \nScanOut893[3] , \nScanOut893[2] , 
        \nScanOut893[1] , \nScanOut893[0] }), .ScanOut({\nScanOut892[7] , 
        \nScanOut892[6] , \nScanOut892[5] , \nScanOut892[4] , \nScanOut892[3] , 
        \nScanOut892[2] , \nScanOut892[1] , \nScanOut892[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_27[7] , \nOut27_27[6] , \nOut27_27[5] , \nOut27_27[4] , 
        \nOut27_27[3] , \nOut27_27[2] , \nOut27_27[1] , \nOut27_27[0] }), 
        .SouthIn({\nOut27_29[7] , \nOut27_29[6] , \nOut27_29[5] , 
        \nOut27_29[4] , \nOut27_29[3] , \nOut27_29[2] , \nOut27_29[1] , 
        \nOut27_29[0] }), .EastIn({\nOut28_28[7] , \nOut28_28[6] , 
        \nOut28_28[5] , \nOut28_28[4] , \nOut28_28[3] , \nOut28_28[2] , 
        \nOut28_28[1] , \nOut28_28[0] }), .WestIn({\nOut26_28[7] , 
        \nOut26_28[6] , \nOut26_28[5] , \nOut26_28[4] , \nOut26_28[3] , 
        \nOut26_28[2] , \nOut26_28[1] , \nOut26_28[0] }), .Out({\nOut27_28[7] , 
        \nOut27_28[6] , \nOut27_28[5] , \nOut27_28[4] , \nOut27_28[3] , 
        \nOut27_28[2] , \nOut27_28[1] , \nOut27_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_902 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut903[7] , \nScanOut903[6] , 
        \nScanOut903[5] , \nScanOut903[4] , \nScanOut903[3] , \nScanOut903[2] , 
        \nScanOut903[1] , \nScanOut903[0] }), .ScanOut({\nScanOut902[7] , 
        \nScanOut902[6] , \nScanOut902[5] , \nScanOut902[4] , \nScanOut902[3] , 
        \nScanOut902[2] , \nScanOut902[1] , \nScanOut902[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_5[7] , \nOut28_5[6] , \nOut28_5[5] , \nOut28_5[4] , 
        \nOut28_5[3] , \nOut28_5[2] , \nOut28_5[1] , \nOut28_5[0] }), 
        .SouthIn({\nOut28_7[7] , \nOut28_7[6] , \nOut28_7[5] , \nOut28_7[4] , 
        \nOut28_7[3] , \nOut28_7[2] , \nOut28_7[1] , \nOut28_7[0] }), .EastIn(
        {\nOut29_6[7] , \nOut29_6[6] , \nOut29_6[5] , \nOut29_6[4] , 
        \nOut29_6[3] , \nOut29_6[2] , \nOut29_6[1] , \nOut29_6[0] }), .WestIn(
        {\nOut27_6[7] , \nOut27_6[6] , \nOut27_6[5] , \nOut27_6[4] , 
        \nOut27_6[3] , \nOut27_6[2] , \nOut27_6[1] , \nOut27_6[0] }), .Out({
        \nOut28_6[7] , \nOut28_6[6] , \nOut28_6[5] , \nOut28_6[4] , 
        \nOut28_6[3] , \nOut28_6[2] , \nOut28_6[1] , \nOut28_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_72 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut73[7] , \nScanOut73[6] , 
        \nScanOut73[5] , \nScanOut73[4] , \nScanOut73[3] , \nScanOut73[2] , 
        \nScanOut73[1] , \nScanOut73[0] }), .ScanOut({\nScanOut72[7] , 
        \nScanOut72[6] , \nScanOut72[5] , \nScanOut72[4] , \nScanOut72[3] , 
        \nScanOut72[2] , \nScanOut72[1] , \nScanOut72[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_7[7] , \nOut2_7[6] , \nOut2_7[5] , \nOut2_7[4] , \nOut2_7[3] , 
        \nOut2_7[2] , \nOut2_7[1] , \nOut2_7[0] }), .SouthIn({\nOut2_9[7] , 
        \nOut2_9[6] , \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , 
        \nOut2_9[1] , \nOut2_9[0] }), .EastIn({\nOut3_8[7] , \nOut3_8[6] , 
        \nOut3_8[5] , \nOut3_8[4] , \nOut3_8[3] , \nOut3_8[2] , \nOut3_8[1] , 
        \nOut3_8[0] }), .WestIn({\nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , 
        \nOut1_8[4] , \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }), 
        .Out({\nOut2_8[7] , \nOut2_8[6] , \nOut2_8[5] , \nOut2_8[4] , 
        \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , \nOut2_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_667 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut668[7] , \nScanOut668[6] , 
        \nScanOut668[5] , \nScanOut668[4] , \nScanOut668[3] , \nScanOut668[2] , 
        \nScanOut668[1] , \nScanOut668[0] }), .ScanOut({\nScanOut667[7] , 
        \nScanOut667[6] , \nScanOut667[5] , \nScanOut667[4] , \nScanOut667[3] , 
        \nScanOut667[2] , \nScanOut667[1] , \nScanOut667[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_26[7] , \nOut20_26[6] , \nOut20_26[5] , \nOut20_26[4] , 
        \nOut20_26[3] , \nOut20_26[2] , \nOut20_26[1] , \nOut20_26[0] }), 
        .SouthIn({\nOut20_28[7] , \nOut20_28[6] , \nOut20_28[5] , 
        \nOut20_28[4] , \nOut20_28[3] , \nOut20_28[2] , \nOut20_28[1] , 
        \nOut20_28[0] }), .EastIn({\nOut21_27[7] , \nOut21_27[6] , 
        \nOut21_27[5] , \nOut21_27[4] , \nOut21_27[3] , \nOut21_27[2] , 
        \nOut21_27[1] , \nOut21_27[0] }), .WestIn({\nOut19_27[7] , 
        \nOut19_27[6] , \nOut19_27[5] , \nOut19_27[4] , \nOut19_27[3] , 
        \nOut19_27[2] , \nOut19_27[1] , \nOut19_27[0] }), .Out({\nOut20_27[7] , 
        \nOut20_27[6] , \nOut20_27[5] , \nOut20_27[4] , \nOut20_27[3] , 
        \nOut20_27[2] , \nOut20_27[1] , \nOut20_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_75 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut76[7] , \nScanOut76[6] , 
        \nScanOut76[5] , \nScanOut76[4] , \nScanOut76[3] , \nScanOut76[2] , 
        \nScanOut76[1] , \nScanOut76[0] }), .ScanOut({\nScanOut75[7] , 
        \nScanOut75[6] , \nScanOut75[5] , \nScanOut75[4] , \nScanOut75[3] , 
        \nScanOut75[2] , \nScanOut75[1] , \nScanOut75[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_10[7] , \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , 
        \nOut2_10[3] , \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), 
        .SouthIn({\nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), .EastIn(
        {\nOut3_11[7] , \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , 
        \nOut3_11[3] , \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }), .WestIn(
        {\nOut1_11[7] , \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , 
        \nOut1_11[3] , \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), .Out({
        \nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_90 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut91[7] , \nScanOut91[6] , 
        \nScanOut91[5] , \nScanOut91[4] , \nScanOut91[3] , \nScanOut91[2] , 
        \nScanOut91[1] , \nScanOut91[0] }), .ScanOut({\nScanOut90[7] , 
        \nScanOut90[6] , \nScanOut90[5] , \nScanOut90[4] , \nScanOut90[3] , 
        \nScanOut90[2] , \nScanOut90[1] , \nScanOut90[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_25[7] , \nOut2_25[6] , \nOut2_25[5] , \nOut2_25[4] , 
        \nOut2_25[3] , \nOut2_25[2] , \nOut2_25[1] , \nOut2_25[0] }), 
        .SouthIn({\nOut2_27[7] , \nOut2_27[6] , \nOut2_27[5] , \nOut2_27[4] , 
        \nOut2_27[3] , \nOut2_27[2] , \nOut2_27[1] , \nOut2_27[0] }), .EastIn(
        {\nOut3_26[7] , \nOut3_26[6] , \nOut3_26[5] , \nOut3_26[4] , 
        \nOut3_26[3] , \nOut3_26[2] , \nOut3_26[1] , \nOut3_26[0] }), .WestIn(
        {\nOut1_26[7] , \nOut1_26[6] , \nOut1_26[5] , \nOut1_26[4] , 
        \nOut1_26[3] , \nOut1_26[2] , \nOut1_26[1] , \nOut1_26[0] }), .Out({
        \nOut2_26[7] , \nOut2_26[6] , \nOut2_26[5] , \nOut2_26[4] , 
        \nOut2_26[3] , \nOut2_26[2] , \nOut2_26[1] , \nOut2_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_97 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut98[7] , \nScanOut98[6] , 
        \nScanOut98[5] , \nScanOut98[4] , \nScanOut98[3] , \nScanOut98[2] , 
        \nScanOut98[1] , \nScanOut98[0] }), .ScanOut({\nScanOut97[7] , 
        \nScanOut97[6] , \nScanOut97[5] , \nScanOut97[4] , \nScanOut97[3] , 
        \nScanOut97[2] , \nScanOut97[1] , \nScanOut97[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_0[7] , \nOut3_0[6] , \nOut3_0[5] , \nOut3_0[4] , \nOut3_0[3] , 
        \nOut3_0[2] , \nOut3_0[1] , \nOut3_0[0] }), .SouthIn({\nOut3_2[7] , 
        \nOut3_2[6] , \nOut3_2[5] , \nOut3_2[4] , \nOut3_2[3] , \nOut3_2[2] , 
        \nOut3_2[1] , \nOut3_2[0] }), .EastIn({\nOut4_1[7] , \nOut4_1[6] , 
        \nOut4_1[5] , \nOut4_1[4] , \nOut4_1[3] , \nOut4_1[2] , \nOut4_1[1] , 
        \nOut4_1[0] }), .WestIn({\nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , 
        \nOut2_1[4] , \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }), 
        .Out({\nOut3_1[7] , \nOut3_1[6] , \nOut3_1[5] , \nOut3_1[4] , 
        \nOut3_1[3] , \nOut3_1[2] , \nOut3_1[1] , \nOut3_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_346 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut347[7] , \nScanOut347[6] , 
        \nScanOut347[5] , \nScanOut347[4] , \nScanOut347[3] , \nScanOut347[2] , 
        \nScanOut347[1] , \nScanOut347[0] }), .ScanOut({\nScanOut346[7] , 
        \nScanOut346[6] , \nScanOut346[5] , \nScanOut346[4] , \nScanOut346[3] , 
        \nScanOut346[2] , \nScanOut346[1] , \nScanOut346[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_25[7] , \nOut10_25[6] , \nOut10_25[5] , \nOut10_25[4] , 
        \nOut10_25[3] , \nOut10_25[2] , \nOut10_25[1] , \nOut10_25[0] }), 
        .SouthIn({\nOut10_27[7] , \nOut10_27[6] , \nOut10_27[5] , 
        \nOut10_27[4] , \nOut10_27[3] , \nOut10_27[2] , \nOut10_27[1] , 
        \nOut10_27[0] }), .EastIn({\nOut11_26[7] , \nOut11_26[6] , 
        \nOut11_26[5] , \nOut11_26[4] , \nOut11_26[3] , \nOut11_26[2] , 
        \nOut11_26[1] , \nOut11_26[0] }), .WestIn({\nOut9_26[7] , 
        \nOut9_26[6] , \nOut9_26[5] , \nOut9_26[4] , \nOut9_26[3] , 
        \nOut9_26[2] , \nOut9_26[1] , \nOut9_26[0] }), .Out({\nOut10_26[7] , 
        \nOut10_26[6] , \nOut10_26[5] , \nOut10_26[4] , \nOut10_26[3] , 
        \nOut10_26[2] , \nOut10_26[1] , \nOut10_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_557 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut558[7] , \nScanOut558[6] , 
        \nScanOut558[5] , \nScanOut558[4] , \nScanOut558[3] , \nScanOut558[2] , 
        \nScanOut558[1] , \nScanOut558[0] }), .ScanOut({\nScanOut557[7] , 
        \nScanOut557[6] , \nScanOut557[5] , \nScanOut557[4] , \nScanOut557[3] , 
        \nScanOut557[2] , \nScanOut557[1] , \nScanOut557[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_12[7] , \nOut17_12[6] , \nOut17_12[5] , \nOut17_12[4] , 
        \nOut17_12[3] , \nOut17_12[2] , \nOut17_12[1] , \nOut17_12[0] }), 
        .SouthIn({\nOut17_14[7] , \nOut17_14[6] , \nOut17_14[5] , 
        \nOut17_14[4] , \nOut17_14[3] , \nOut17_14[2] , \nOut17_14[1] , 
        \nOut17_14[0] }), .EastIn({\nOut18_13[7] , \nOut18_13[6] , 
        \nOut18_13[5] , \nOut18_13[4] , \nOut18_13[3] , \nOut18_13[2] , 
        \nOut18_13[1] , \nOut18_13[0] }), .WestIn({\nOut16_13[7] , 
        \nOut16_13[6] , \nOut16_13[5] , \nOut16_13[4] , \nOut16_13[3] , 
        \nOut16_13[2] , \nOut16_13[1] , \nOut16_13[0] }), .Out({\nOut17_13[7] , 
        \nOut17_13[6] , \nOut17_13[5] , \nOut17_13[4] , \nOut17_13[3] , 
        \nOut17_13[2] , \nOut17_13[1] , \nOut17_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_819 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut820[7] , \nScanOut820[6] , 
        \nScanOut820[5] , \nScanOut820[4] , \nScanOut820[3] , \nScanOut820[2] , 
        \nScanOut820[1] , \nScanOut820[0] }), .ScanOut({\nScanOut819[7] , 
        \nScanOut819[6] , \nScanOut819[5] , \nScanOut819[4] , \nScanOut819[3] , 
        \nScanOut819[2] , \nScanOut819[1] , \nScanOut819[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_18[7] , \nOut25_18[6] , \nOut25_18[5] , \nOut25_18[4] , 
        \nOut25_18[3] , \nOut25_18[2] , \nOut25_18[1] , \nOut25_18[0] }), 
        .SouthIn({\nOut25_20[7] , \nOut25_20[6] , \nOut25_20[5] , 
        \nOut25_20[4] , \nOut25_20[3] , \nOut25_20[2] , \nOut25_20[1] , 
        \nOut25_20[0] }), .EastIn({\nOut26_19[7] , \nOut26_19[6] , 
        \nOut26_19[5] , \nOut26_19[4] , \nOut26_19[3] , \nOut26_19[2] , 
        \nOut26_19[1] , \nOut26_19[0] }), .WestIn({\nOut24_19[7] , 
        \nOut24_19[6] , \nOut24_19[5] , \nOut24_19[4] , \nOut24_19[3] , 
        \nOut24_19[2] , \nOut24_19[1] , \nOut24_19[0] }), .Out({\nOut25_19[7] , 
        \nOut25_19[6] , \nOut25_19[5] , \nOut25_19[4] , \nOut25_19[3] , 
        \nOut25_19[2] , \nOut25_19[1] , \nOut25_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_925 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut926[7] , \nScanOut926[6] , 
        \nScanOut926[5] , \nScanOut926[4] , \nScanOut926[3] , \nScanOut926[2] , 
        \nScanOut926[1] , \nScanOut926[0] }), .ScanOut({\nScanOut925[7] , 
        \nScanOut925[6] , \nScanOut925[5] , \nScanOut925[4] , \nScanOut925[3] , 
        \nScanOut925[2] , \nScanOut925[1] , \nScanOut925[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_28[7] , \nOut28_28[6] , \nOut28_28[5] , \nOut28_28[4] , 
        \nOut28_28[3] , \nOut28_28[2] , \nOut28_28[1] , \nOut28_28[0] }), 
        .SouthIn({\nOut28_30[7] , \nOut28_30[6] , \nOut28_30[5] , 
        \nOut28_30[4] , \nOut28_30[3] , \nOut28_30[2] , \nOut28_30[1] , 
        \nOut28_30[0] }), .EastIn({\nOut29_29[7] , \nOut29_29[6] , 
        \nOut29_29[5] , \nOut29_29[4] , \nOut29_29[3] , \nOut29_29[2] , 
        \nOut29_29[1] , \nOut29_29[0] }), .WestIn({\nOut27_29[7] , 
        \nOut27_29[6] , \nOut27_29[5] , \nOut27_29[4] , \nOut27_29[3] , 
        \nOut27_29[2] , \nOut27_29[1] , \nOut27_29[0] }), .Out({\nOut28_29[7] , 
        \nOut28_29[6] , \nOut28_29[5] , \nOut28_29[4] , \nOut28_29[3] , 
        \nOut28_29[2] , \nOut28_29[1] , \nOut28_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_989 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut990[7] , \nScanOut990[6] , 
        \nScanOut990[5] , \nScanOut990[4] , \nScanOut990[3] , \nScanOut990[2] , 
        \nScanOut990[1] , \nScanOut990[0] }), .ScanOut({\nScanOut989[7] , 
        \nScanOut989[6] , \nScanOut989[5] , \nScanOut989[4] , \nScanOut989[3] , 
        \nScanOut989[2] , \nScanOut989[1] , \nScanOut989[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_28[7] , \nOut30_28[6] , \nOut30_28[5] , \nOut30_28[4] , 
        \nOut30_28[3] , \nOut30_28[2] , \nOut30_28[1] , \nOut30_28[0] }), 
        .SouthIn({\nOut30_30[7] , \nOut30_30[6] , \nOut30_30[5] , 
        \nOut30_30[4] , \nOut30_30[3] , \nOut30_30[2] , \nOut30_30[1] , 
        \nOut30_30[0] }), .EastIn({\nOut31_29[7] , \nOut31_29[6] , 
        \nOut31_29[5] , \nOut31_29[4] , \nOut31_29[3] , \nOut31_29[2] , 
        \nOut31_29[1] , \nOut31_29[0] }), .WestIn({\nOut29_29[7] , 
        \nOut29_29[6] , \nOut29_29[5] , \nOut29_29[4] , \nOut29_29[3] , 
        \nOut29_29[2] , \nOut29_29[1] , \nOut29_29[0] }), .Out({\nOut30_29[7] , 
        \nOut30_29[6] , \nOut30_29[5] , \nOut30_29[4] , \nOut30_29[3] , 
        \nOut30_29[2] , \nOut30_29[1] , \nOut30_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_103 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut104[7] , \nScanOut104[6] , 
        \nScanOut104[5] , \nScanOut104[4] , \nScanOut104[3] , \nScanOut104[2] , 
        \nScanOut104[1] , \nScanOut104[0] }), .ScanOut({\nScanOut103[7] , 
        \nScanOut103[6] , \nScanOut103[5] , \nScanOut103[4] , \nScanOut103[3] , 
        \nScanOut103[2] , \nScanOut103[1] , \nScanOut103[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_6[7] , \nOut3_6[6] , \nOut3_6[5] , \nOut3_6[4] , \nOut3_6[3] , 
        \nOut3_6[2] , \nOut3_6[1] , \nOut3_6[0] }), .SouthIn({\nOut3_8[7] , 
        \nOut3_8[6] , \nOut3_8[5] , \nOut3_8[4] , \nOut3_8[3] , \nOut3_8[2] , 
        \nOut3_8[1] , \nOut3_8[0] }), .EastIn({\nOut4_7[7] , \nOut4_7[6] , 
        \nOut4_7[5] , \nOut4_7[4] , \nOut4_7[3] , \nOut4_7[2] , \nOut4_7[1] , 
        \nOut4_7[0] }), .WestIn({\nOut2_7[7] , \nOut2_7[6] , \nOut2_7[5] , 
        \nOut2_7[4] , \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , \nOut2_7[0] }), 
        .Out({\nOut3_7[7] , \nOut3_7[6] , \nOut3_7[5] , \nOut3_7[4] , 
        \nOut3_7[3] , \nOut3_7[2] , \nOut3_7[1] , \nOut3_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_682 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut683[7] , \nScanOut683[6] , 
        \nScanOut683[5] , \nScanOut683[4] , \nScanOut683[3] , \nScanOut683[2] , 
        \nScanOut683[1] , \nScanOut683[0] }), .ScanOut({\nScanOut682[7] , 
        \nScanOut682[6] , \nScanOut682[5] , \nScanOut682[4] , \nScanOut682[3] , 
        \nScanOut682[2] , \nScanOut682[1] , \nScanOut682[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_9[7] , \nOut21_9[6] , \nOut21_9[5] , \nOut21_9[4] , 
        \nOut21_9[3] , \nOut21_9[2] , \nOut21_9[1] , \nOut21_9[0] }), 
        .SouthIn({\nOut21_11[7] , \nOut21_11[6] , \nOut21_11[5] , 
        \nOut21_11[4] , \nOut21_11[3] , \nOut21_11[2] , \nOut21_11[1] , 
        \nOut21_11[0] }), .EastIn({\nOut22_10[7] , \nOut22_10[6] , 
        \nOut22_10[5] , \nOut22_10[4] , \nOut22_10[3] , \nOut22_10[2] , 
        \nOut22_10[1] , \nOut22_10[0] }), .WestIn({\nOut20_10[7] , 
        \nOut20_10[6] , \nOut20_10[5] , \nOut20_10[4] , \nOut20_10[3] , 
        \nOut20_10[2] , \nOut20_10[1] , \nOut20_10[0] }), .Out({\nOut21_10[7] , 
        \nOut21_10[6] , \nOut21_10[5] , \nOut21_10[4] , \nOut21_10[3] , 
        \nOut21_10[2] , \nOut21_10[1] , \nOut21_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1014 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1015[7] , \nScanOut1015[6] , 
        \nScanOut1015[5] , \nScanOut1015[4] , \nScanOut1015[3] , 
        \nScanOut1015[2] , \nScanOut1015[1] , \nScanOut1015[0] }), .ScanOut({
        \nScanOut1014[7] , \nScanOut1014[6] , \nScanOut1014[5] , 
        \nScanOut1014[4] , \nScanOut1014[3] , \nScanOut1014[2] , 
        \nScanOut1014[1] , \nScanOut1014[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_22[7] , \nOut31_22[6] , \nOut31_22[5] , 
        \nOut31_22[4] , \nOut31_22[3] , \nOut31_22[2] , \nOut31_22[1] , 
        \nOut31_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_104 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut105[7] , \nScanOut105[6] , 
        \nScanOut105[5] , \nScanOut105[4] , \nScanOut105[3] , \nScanOut105[2] , 
        \nScanOut105[1] , \nScanOut105[0] }), .ScanOut({\nScanOut104[7] , 
        \nScanOut104[6] , \nScanOut104[5] , \nScanOut104[4] , \nScanOut104[3] , 
        \nScanOut104[2] , \nScanOut104[1] , \nScanOut104[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_7[7] , \nOut3_7[6] , \nOut3_7[5] , \nOut3_7[4] , \nOut3_7[3] , 
        \nOut3_7[2] , \nOut3_7[1] , \nOut3_7[0] }), .SouthIn({\nOut3_9[7] , 
        \nOut3_9[6] , \nOut3_9[5] , \nOut3_9[4] , \nOut3_9[3] , \nOut3_9[2] , 
        \nOut3_9[1] , \nOut3_9[0] }), .EastIn({\nOut4_8[7] , \nOut4_8[6] , 
        \nOut4_8[5] , \nOut4_8[4] , \nOut4_8[3] , \nOut4_8[2] , \nOut4_8[1] , 
        \nOut4_8[0] }), .WestIn({\nOut2_8[7] , \nOut2_8[6] , \nOut2_8[5] , 
        \nOut2_8[4] , \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , \nOut2_8[0] }), 
        .Out({\nOut3_8[7] , \nOut3_8[6] , \nOut3_8[5] , \nOut3_8[4] , 
        \nOut3_8[3] , \nOut3_8[2] , \nOut3_8[1] , \nOut3_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_123 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut124[7] , \nScanOut124[6] , 
        \nScanOut124[5] , \nScanOut124[4] , \nScanOut124[3] , \nScanOut124[2] , 
        \nScanOut124[1] , \nScanOut124[0] }), .ScanOut({\nScanOut123[7] , 
        \nScanOut123[6] , \nScanOut123[5] , \nScanOut123[4] , \nScanOut123[3] , 
        \nScanOut123[2] , \nScanOut123[1] , \nScanOut123[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_26[7] , \nOut3_26[6] , \nOut3_26[5] , \nOut3_26[4] , 
        \nOut3_26[3] , \nOut3_26[2] , \nOut3_26[1] , \nOut3_26[0] }), 
        .SouthIn({\nOut3_28[7] , \nOut3_28[6] , \nOut3_28[5] , \nOut3_28[4] , 
        \nOut3_28[3] , \nOut3_28[2] , \nOut3_28[1] , \nOut3_28[0] }), .EastIn(
        {\nOut4_27[7] , \nOut4_27[6] , \nOut4_27[5] , \nOut4_27[4] , 
        \nOut4_27[3] , \nOut4_27[2] , \nOut4_27[1] , \nOut4_27[0] }), .WestIn(
        {\nOut2_27[7] , \nOut2_27[6] , \nOut2_27[5] , \nOut2_27[4] , 
        \nOut2_27[3] , \nOut2_27[2] , \nOut2_27[1] , \nOut2_27[0] }), .Out({
        \nOut3_27[7] , \nOut3_27[6] , \nOut3_27[5] , \nOut3_27[4] , 
        \nOut3_27[3] , \nOut3_27[2] , \nOut3_27[1] , \nOut3_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_124 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut125[7] , \nScanOut125[6] , 
        \nScanOut125[5] , \nScanOut125[4] , \nScanOut125[3] , \nScanOut125[2] , 
        \nScanOut125[1] , \nScanOut125[0] }), .ScanOut({\nScanOut124[7] , 
        \nScanOut124[6] , \nScanOut124[5] , \nScanOut124[4] , \nScanOut124[3] , 
        \nScanOut124[2] , \nScanOut124[1] , \nScanOut124[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_27[7] , \nOut3_27[6] , \nOut3_27[5] , \nOut3_27[4] , 
        \nOut3_27[3] , \nOut3_27[2] , \nOut3_27[1] , \nOut3_27[0] }), 
        .SouthIn({\nOut3_29[7] , \nOut3_29[6] , \nOut3_29[5] , \nOut3_29[4] , 
        \nOut3_29[3] , \nOut3_29[2] , \nOut3_29[1] , \nOut3_29[0] }), .EastIn(
        {\nOut4_28[7] , \nOut4_28[6] , \nOut4_28[5] , \nOut4_28[4] , 
        \nOut4_28[3] , \nOut4_28[2] , \nOut4_28[1] , \nOut4_28[0] }), .WestIn(
        {\nOut2_28[7] , \nOut2_28[6] , \nOut2_28[5] , \nOut2_28[4] , 
        \nOut2_28[3] , \nOut2_28[2] , \nOut2_28[1] , \nOut2_28[0] }), .Out({
        \nOut3_28[7] , \nOut3_28[6] , \nOut3_28[5] , \nOut3_28[4] , 
        \nOut3_28[3] , \nOut3_28[2] , \nOut3_28[1] , \nOut3_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_214 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut215[7] , \nScanOut215[6] , 
        \nScanOut215[5] , \nScanOut215[4] , \nScanOut215[3] , \nScanOut215[2] , 
        \nScanOut215[1] , \nScanOut215[0] }), .ScanOut({\nScanOut214[7] , 
        \nScanOut214[6] , \nScanOut214[5] , \nScanOut214[4] , \nScanOut214[3] , 
        \nScanOut214[2] , \nScanOut214[1] , \nScanOut214[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_21[7] , \nOut6_21[6] , \nOut6_21[5] , \nOut6_21[4] , 
        \nOut6_21[3] , \nOut6_21[2] , \nOut6_21[1] , \nOut6_21[0] }), 
        .SouthIn({\nOut6_23[7] , \nOut6_23[6] , \nOut6_23[5] , \nOut6_23[4] , 
        \nOut6_23[3] , \nOut6_23[2] , \nOut6_23[1] , \nOut6_23[0] }), .EastIn(
        {\nOut7_22[7] , \nOut7_22[6] , \nOut7_22[5] , \nOut7_22[4] , 
        \nOut7_22[3] , \nOut7_22[2] , \nOut7_22[1] , \nOut7_22[0] }), .WestIn(
        {\nOut5_22[7] , \nOut5_22[6] , \nOut5_22[5] , \nOut5_22[4] , 
        \nOut5_22[3] , \nOut5_22[2] , \nOut5_22[1] , \nOut5_22[0] }), .Out({
        \nOut6_22[7] , \nOut6_22[6] , \nOut6_22[5] , \nOut6_22[4] , 
        \nOut6_22[3] , \nOut6_22[2] , \nOut6_22[1] , \nOut6_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_233 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut234[7] , \nScanOut234[6] , 
        \nScanOut234[5] , \nScanOut234[4] , \nScanOut234[3] , \nScanOut234[2] , 
        \nScanOut234[1] , \nScanOut234[0] }), .ScanOut({\nScanOut233[7] , 
        \nScanOut233[6] , \nScanOut233[5] , \nScanOut233[4] , \nScanOut233[3] , 
        \nScanOut233[2] , \nScanOut233[1] , \nScanOut233[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_8[7] , \nOut7_8[6] , \nOut7_8[5] , \nOut7_8[4] , \nOut7_8[3] , 
        \nOut7_8[2] , \nOut7_8[1] , \nOut7_8[0] }), .SouthIn({\nOut7_10[7] , 
        \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , \nOut7_10[3] , 
        \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }), .EastIn({\nOut8_9[7] , 
        \nOut8_9[6] , \nOut8_9[5] , \nOut8_9[4] , \nOut8_9[3] , \nOut8_9[2] , 
        \nOut8_9[1] , \nOut8_9[0] }), .WestIn({\nOut6_9[7] , \nOut6_9[6] , 
        \nOut6_9[5] , \nOut6_9[4] , \nOut6_9[3] , \nOut6_9[2] , \nOut6_9[1] , 
        \nOut6_9[0] }), .Out({\nOut7_9[7] , \nOut7_9[6] , \nOut7_9[5] , 
        \nOut7_9[4] , \nOut7_9[3] , \nOut7_9[2] , \nOut7_9[1] , \nOut7_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_712 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut713[7] , \nScanOut713[6] , 
        \nScanOut713[5] , \nScanOut713[4] , \nScanOut713[3] , \nScanOut713[2] , 
        \nScanOut713[1] , \nScanOut713[0] }), .ScanOut({\nScanOut712[7] , 
        \nScanOut712[6] , \nScanOut712[5] , \nScanOut712[4] , \nScanOut712[3] , 
        \nScanOut712[2] , \nScanOut712[1] , \nScanOut712[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_7[7] , \nOut22_7[6] , \nOut22_7[5] , \nOut22_7[4] , 
        \nOut22_7[3] , \nOut22_7[2] , \nOut22_7[1] , \nOut22_7[0] }), 
        .SouthIn({\nOut22_9[7] , \nOut22_9[6] , \nOut22_9[5] , \nOut22_9[4] , 
        \nOut22_9[3] , \nOut22_9[2] , \nOut22_9[1] , \nOut22_9[0] }), .EastIn(
        {\nOut23_8[7] , \nOut23_8[6] , \nOut23_8[5] , \nOut23_8[4] , 
        \nOut23_8[3] , \nOut23_8[2] , \nOut23_8[1] , \nOut23_8[0] }), .WestIn(
        {\nOut21_8[7] , \nOut21_8[6] , \nOut21_8[5] , \nOut21_8[4] , 
        \nOut21_8[3] , \nOut21_8[2] , \nOut21_8[1] , \nOut21_8[0] }), .Out({
        \nOut22_8[7] , \nOut22_8[6] , \nOut22_8[5] , \nOut22_8[4] , 
        \nOut22_8[3] , \nOut22_8[2] , \nOut22_8[1] , \nOut22_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_384 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut385[7] , \nScanOut385[6] , 
        \nScanOut385[5] , \nScanOut385[4] , \nScanOut385[3] , \nScanOut385[2] , 
        \nScanOut385[1] , \nScanOut385[0] }), .ScanOut({\nScanOut384[7] , 
        \nScanOut384[6] , \nScanOut384[5] , \nScanOut384[4] , \nScanOut384[3] , 
        \nScanOut384[2] , \nScanOut384[1] , \nScanOut384[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut12_0[7] , \nOut12_0[6] , 
        \nOut12_0[5] , \nOut12_0[4] , \nOut12_0[3] , \nOut12_0[2] , 
        \nOut12_0[1] , \nOut12_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_422 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut423[7] , \nScanOut423[6] , 
        \nScanOut423[5] , \nScanOut423[4] , \nScanOut423[3] , \nScanOut423[2] , 
        \nScanOut423[1] , \nScanOut423[0] }), .ScanOut({\nScanOut422[7] , 
        \nScanOut422[6] , \nScanOut422[5] , \nScanOut422[4] , \nScanOut422[3] , 
        \nScanOut422[2] , \nScanOut422[1] , \nScanOut422[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }), 
        .SouthIn({\nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }), .EastIn(
        {\nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }), .WestIn(
        {\nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }), .Out({
        \nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_850 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut851[7] , \nScanOut851[6] , 
        \nScanOut851[5] , \nScanOut851[4] , \nScanOut851[3] , \nScanOut851[2] , 
        \nScanOut851[1] , \nScanOut851[0] }), .ScanOut({\nScanOut850[7] , 
        \nScanOut850[6] , \nScanOut850[5] , \nScanOut850[4] , \nScanOut850[3] , 
        \nScanOut850[2] , \nScanOut850[1] , \nScanOut850[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_17[7] , \nOut26_17[6] , \nOut26_17[5] , \nOut26_17[4] , 
        \nOut26_17[3] , \nOut26_17[2] , \nOut26_17[1] , \nOut26_17[0] }), 
        .SouthIn({\nOut26_19[7] , \nOut26_19[6] , \nOut26_19[5] , 
        \nOut26_19[4] , \nOut26_19[3] , \nOut26_19[2] , \nOut26_19[1] , 
        \nOut26_19[0] }), .EastIn({\nOut27_18[7] , \nOut27_18[6] , 
        \nOut27_18[5] , \nOut27_18[4] , \nOut27_18[3] , \nOut27_18[2] , 
        \nOut27_18[1] , \nOut27_18[0] }), .WestIn({\nOut25_18[7] , 
        \nOut25_18[6] , \nOut25_18[5] , \nOut25_18[4] , \nOut25_18[3] , 
        \nOut25_18[2] , \nOut25_18[1] , \nOut25_18[0] }), .Out({\nOut26_18[7] , 
        \nOut26_18[6] , \nOut26_18[5] , \nOut26_18[4] , \nOut26_18[3] , 
        \nOut26_18[2] , \nOut26_18[1] , \nOut26_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_405 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut406[7] , \nScanOut406[6] , 
        \nScanOut406[5] , \nScanOut406[4] , \nScanOut406[3] , \nScanOut406[2] , 
        \nScanOut406[1] , \nScanOut406[0] }), .ScanOut({\nScanOut405[7] , 
        \nScanOut405[6] , \nScanOut405[5] , \nScanOut405[4] , \nScanOut405[3] , 
        \nScanOut405[2] , \nScanOut405[1] , \nScanOut405[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_20[7] , \nOut12_20[6] , \nOut12_20[5] , \nOut12_20[4] , 
        \nOut12_20[3] , \nOut12_20[2] , \nOut12_20[1] , \nOut12_20[0] }), 
        .SouthIn({\nOut12_22[7] , \nOut12_22[6] , \nOut12_22[5] , 
        \nOut12_22[4] , \nOut12_22[3] , \nOut12_22[2] , \nOut12_22[1] , 
        \nOut12_22[0] }), .EastIn({\nOut13_21[7] , \nOut13_21[6] , 
        \nOut13_21[5] , \nOut13_21[4] , \nOut13_21[3] , \nOut13_21[2] , 
        \nOut13_21[1] , \nOut13_21[0] }), .WestIn({\nOut11_21[7] , 
        \nOut11_21[6] , \nOut11_21[5] , \nOut11_21[4] , \nOut11_21[3] , 
        \nOut11_21[2] , \nOut11_21[1] , \nOut11_21[0] }), .Out({\nOut12_21[7] , 
        \nOut12_21[6] , \nOut12_21[5] , \nOut12_21[4] , \nOut12_21[3] , 
        \nOut12_21[2] , \nOut12_21[1] , \nOut12_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_595 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut596[7] , \nScanOut596[6] , 
        \nScanOut596[5] , \nScanOut596[4] , \nScanOut596[3] , \nScanOut596[2] , 
        \nScanOut596[1] , \nScanOut596[0] }), .ScanOut({\nScanOut595[7] , 
        \nScanOut595[6] , \nScanOut595[5] , \nScanOut595[4] , \nScanOut595[3] , 
        \nScanOut595[2] , \nScanOut595[1] , \nScanOut595[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_18[7] , \nOut18_18[6] , \nOut18_18[5] , \nOut18_18[4] , 
        \nOut18_18[3] , \nOut18_18[2] , \nOut18_18[1] , \nOut18_18[0] }), 
        .SouthIn({\nOut18_20[7] , \nOut18_20[6] , \nOut18_20[5] , 
        \nOut18_20[4] , \nOut18_20[3] , \nOut18_20[2] , \nOut18_20[1] , 
        \nOut18_20[0] }), .EastIn({\nOut19_19[7] , \nOut19_19[6] , 
        \nOut19_19[5] , \nOut19_19[4] , \nOut19_19[3] , \nOut19_19[2] , 
        \nOut19_19[1] , \nOut19_19[0] }), .WestIn({\nOut17_19[7] , 
        \nOut17_19[6] , \nOut17_19[5] , \nOut17_19[4] , \nOut17_19[3] , 
        \nOut17_19[2] , \nOut17_19[1] , \nOut17_19[0] }), .Out({\nOut18_19[7] , 
        \nOut18_19[6] , \nOut18_19[5] , \nOut18_19[4] , \nOut18_19[3] , 
        \nOut18_19[2] , \nOut18_19[1] , \nOut18_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_735 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut736[7] , \nScanOut736[6] , 
        \nScanOut736[5] , \nScanOut736[4] , \nScanOut736[3] , \nScanOut736[2] , 
        \nScanOut736[1] , \nScanOut736[0] }), .ScanOut({\nScanOut735[7] , 
        \nScanOut735[6] , \nScanOut735[5] , \nScanOut735[4] , \nScanOut735[3] , 
        \nScanOut735[2] , \nScanOut735[1] , \nScanOut735[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut22_31[7] , \nOut22_31[6] , 
        \nOut22_31[5] , \nOut22_31[4] , \nOut22_31[3] , \nOut22_31[2] , 
        \nOut22_31[1] , \nOut22_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_877 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut878[7] , \nScanOut878[6] , 
        \nScanOut878[5] , \nScanOut878[4] , \nScanOut878[3] , \nScanOut878[2] , 
        \nScanOut878[1] , \nScanOut878[0] }), .ScanOut({\nScanOut877[7] , 
        \nScanOut877[6] , \nScanOut877[5] , \nScanOut877[4] , \nScanOut877[3] , 
        \nScanOut877[2] , \nScanOut877[1] , \nScanOut877[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_12[7] , \nOut27_12[6] , \nOut27_12[5] , \nOut27_12[4] , 
        \nOut27_12[3] , \nOut27_12[2] , \nOut27_12[1] , \nOut27_12[0] }), 
        .SouthIn({\nOut27_14[7] , \nOut27_14[6] , \nOut27_14[5] , 
        \nOut27_14[4] , \nOut27_14[3] , \nOut27_14[2] , \nOut27_14[1] , 
        \nOut27_14[0] }), .EastIn({\nOut28_13[7] , \nOut28_13[6] , 
        \nOut28_13[5] , \nOut28_13[4] , \nOut28_13[3] , \nOut28_13[2] , 
        \nOut28_13[1] , \nOut28_13[0] }), .WestIn({\nOut26_13[7] , 
        \nOut26_13[6] , \nOut26_13[5] , \nOut26_13[4] , \nOut26_13[3] , 
        \nOut26_13[2] , \nOut26_13[1] , \nOut26_13[0] }), .Out({\nOut27_13[7] , 
        \nOut27_13[6] , \nOut27_13[5] , \nOut27_13[4] , \nOut27_13[3] , 
        \nOut27_13[2] , \nOut27_13[1] , \nOut27_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_188 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut189[7] , \nScanOut189[6] , 
        \nScanOut189[5] , \nScanOut189[4] , \nScanOut189[3] , \nScanOut189[2] , 
        \nScanOut189[1] , \nScanOut189[0] }), .ScanOut({\nScanOut188[7] , 
        \nScanOut188[6] , \nScanOut188[5] , \nScanOut188[4] , \nScanOut188[3] , 
        \nScanOut188[2] , \nScanOut188[1] , \nScanOut188[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_27[7] , \nOut5_27[6] , \nOut5_27[5] , \nOut5_27[4] , 
        \nOut5_27[3] , \nOut5_27[2] , \nOut5_27[1] , \nOut5_27[0] }), 
        .SouthIn({\nOut5_29[7] , \nOut5_29[6] , \nOut5_29[5] , \nOut5_29[4] , 
        \nOut5_29[3] , \nOut5_29[2] , \nOut5_29[1] , \nOut5_29[0] }), .EastIn(
        {\nOut6_28[7] , \nOut6_28[6] , \nOut6_28[5] , \nOut6_28[4] , 
        \nOut6_28[3] , \nOut6_28[2] , \nOut6_28[1] , \nOut6_28[0] }), .WestIn(
        {\nOut4_28[7] , \nOut4_28[6] , \nOut4_28[5] , \nOut4_28[4] , 
        \nOut4_28[3] , \nOut4_28[2] , \nOut4_28[1] , \nOut4_28[0] }), .Out({
        \nOut5_28[7] , \nOut5_28[6] , \nOut5_28[5] , \nOut5_28[4] , 
        \nOut5_28[3] , \nOut5_28[2] , \nOut5_28[1] , \nOut5_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_609 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut610[7] , \nScanOut610[6] , 
        \nScanOut610[5] , \nScanOut610[4] , \nScanOut610[3] , \nScanOut610[2] , 
        \nScanOut610[1] , \nScanOut610[0] }), .ScanOut({\nScanOut609[7] , 
        \nScanOut609[6] , \nScanOut609[5] , \nScanOut609[4] , \nScanOut609[3] , 
        \nScanOut609[2] , \nScanOut609[1] , \nScanOut609[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_0[7] , \nOut19_0[6] , \nOut19_0[5] , \nOut19_0[4] , 
        \nOut19_0[3] , \nOut19_0[2] , \nOut19_0[1] , \nOut19_0[0] }), 
        .SouthIn({\nOut19_2[7] , \nOut19_2[6] , \nOut19_2[5] , \nOut19_2[4] , 
        \nOut19_2[3] , \nOut19_2[2] , \nOut19_2[1] , \nOut19_2[0] }), .EastIn(
        {\nOut20_1[7] , \nOut20_1[6] , \nOut20_1[5] , \nOut20_1[4] , 
        \nOut20_1[3] , \nOut20_1[2] , \nOut20_1[1] , \nOut20_1[0] }), .WestIn(
        {\nOut18_1[7] , \nOut18_1[6] , \nOut18_1[5] , \nOut18_1[4] , 
        \nOut18_1[3] , \nOut18_1[2] , \nOut18_1[1] , \nOut18_1[0] }), .Out({
        \nOut19_1[7] , \nOut19_1[6] , \nOut19_1[5] , \nOut19_1[4] , 
        \nOut19_1[3] , \nOut19_1[2] , \nOut19_1[1] , \nOut19_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_328 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut329[7] , \nScanOut329[6] , 
        \nScanOut329[5] , \nScanOut329[4] , \nScanOut329[3] , \nScanOut329[2] , 
        \nScanOut329[1] , \nScanOut329[0] }), .ScanOut({\nScanOut328[7] , 
        \nScanOut328[6] , \nScanOut328[5] , \nScanOut328[4] , \nScanOut328[3] , 
        \nScanOut328[2] , \nScanOut328[1] , \nScanOut328[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_7[7] , \nOut10_7[6] , \nOut10_7[5] , \nOut10_7[4] , 
        \nOut10_7[3] , \nOut10_7[2] , \nOut10_7[1] , \nOut10_7[0] }), 
        .SouthIn({\nOut10_9[7] , \nOut10_9[6] , \nOut10_9[5] , \nOut10_9[4] , 
        \nOut10_9[3] , \nOut10_9[2] , \nOut10_9[1] , \nOut10_9[0] }), .EastIn(
        {\nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }), .WestIn(
        {\nOut9_8[7] , \nOut9_8[6] , \nOut9_8[5] , \nOut9_8[4] , \nOut9_8[3] , 
        \nOut9_8[2] , \nOut9_8[1] , \nOut9_8[0] }), .Out({\nOut10_8[7] , 
        \nOut10_8[6] , \nOut10_8[5] , \nOut10_8[4] , \nOut10_8[3] , 
        \nOut10_8[2] , \nOut10_8[1] , \nOut10_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_539 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut540[7] , \nScanOut540[6] , 
        \nScanOut540[5] , \nScanOut540[4] , \nScanOut540[3] , \nScanOut540[2] , 
        \nScanOut540[1] , \nScanOut540[0] }), .ScanOut({\nScanOut539[7] , 
        \nScanOut539[6] , \nScanOut539[5] , \nScanOut539[4] , \nScanOut539[3] , 
        \nScanOut539[2] , \nScanOut539[1] , \nScanOut539[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_26[7] , \nOut16_26[6] , \nOut16_26[5] , \nOut16_26[4] , 
        \nOut16_26[3] , \nOut16_26[2] , \nOut16_26[1] , \nOut16_26[0] }), 
        .SouthIn({\nOut16_28[7] , \nOut16_28[6] , \nOut16_28[5] , 
        \nOut16_28[4] , \nOut16_28[3] , \nOut16_28[2] , \nOut16_28[1] , 
        \nOut16_28[0] }), .EastIn({\nOut17_27[7] , \nOut17_27[6] , 
        \nOut17_27[5] , \nOut17_27[4] , \nOut17_27[3] , \nOut17_27[2] , 
        \nOut17_27[1] , \nOut17_27[0] }), .WestIn({\nOut15_27[7] , 
        \nOut15_27[6] , \nOut15_27[5] , \nOut15_27[4] , \nOut15_27[3] , 
        \nOut15_27[2] , \nOut15_27[1] , \nOut15_27[0] }), .Out({\nOut16_27[7] , 
        \nOut16_27[6] , \nOut16_27[5] , \nOut16_27[4] , \nOut16_27[3] , 
        \nOut16_27[2] , \nOut16_27[1] , \nOut16_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_799 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut800[7] , \nScanOut800[6] , 
        \nScanOut800[5] , \nScanOut800[4] , \nScanOut800[3] , \nScanOut800[2] , 
        \nScanOut800[1] , \nScanOut800[0] }), .ScanOut({\nScanOut799[7] , 
        \nScanOut799[6] , \nScanOut799[5] , \nScanOut799[4] , \nScanOut799[3] , 
        \nScanOut799[2] , \nScanOut799[1] , \nScanOut799[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut24_31[7] , \nOut24_31[6] , 
        \nOut24_31[5] , \nOut24_31[4] , \nOut24_31[3] , \nOut24_31[2] , 
        \nOut24_31[1] , \nOut24_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_213 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut214[7] , \nScanOut214[6] , 
        \nScanOut214[5] , \nScanOut214[4] , \nScanOut214[3] , \nScanOut214[2] , 
        \nScanOut214[1] , \nScanOut214[0] }), .ScanOut({\nScanOut213[7] , 
        \nScanOut213[6] , \nScanOut213[5] , \nScanOut213[4] , \nScanOut213[3] , 
        \nScanOut213[2] , \nScanOut213[1] , \nScanOut213[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_20[7] , \nOut6_20[6] , \nOut6_20[5] , \nOut6_20[4] , 
        \nOut6_20[3] , \nOut6_20[2] , \nOut6_20[1] , \nOut6_20[0] }), 
        .SouthIn({\nOut6_22[7] , \nOut6_22[6] , \nOut6_22[5] , \nOut6_22[4] , 
        \nOut6_22[3] , \nOut6_22[2] , \nOut6_22[1] , \nOut6_22[0] }), .EastIn(
        {\nOut7_21[7] , \nOut7_21[6] , \nOut7_21[5] , \nOut7_21[4] , 
        \nOut7_21[3] , \nOut7_21[2] , \nOut7_21[1] , \nOut7_21[0] }), .WestIn(
        {\nOut5_21[7] , \nOut5_21[6] , \nOut5_21[5] , \nOut5_21[4] , 
        \nOut5_21[3] , \nOut5_21[2] , \nOut5_21[1] , \nOut5_21[0] }), .Out({
        \nOut6_21[7] , \nOut6_21[6] , \nOut6_21[5] , \nOut6_21[4] , 
        \nOut6_21[3] , \nOut6_21[2] , \nOut6_21[1] , \nOut6_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_592 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut593[7] , \nScanOut593[6] , 
        \nScanOut593[5] , \nScanOut593[4] , \nScanOut593[3] , \nScanOut593[2] , 
        \nScanOut593[1] , \nScanOut593[0] }), .ScanOut({\nScanOut592[7] , 
        \nScanOut592[6] , \nScanOut592[5] , \nScanOut592[4] , \nScanOut592[3] , 
        \nScanOut592[2] , \nScanOut592[1] , \nScanOut592[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_15[7] , \nOut18_15[6] , \nOut18_15[5] , \nOut18_15[4] , 
        \nOut18_15[3] , \nOut18_15[2] , \nOut18_15[1] , \nOut18_15[0] }), 
        .SouthIn({\nOut18_17[7] , \nOut18_17[6] , \nOut18_17[5] , 
        \nOut18_17[4] , \nOut18_17[3] , \nOut18_17[2] , \nOut18_17[1] , 
        \nOut18_17[0] }), .EastIn({\nOut19_16[7] , \nOut19_16[6] , 
        \nOut19_16[5] , \nOut19_16[4] , \nOut19_16[3] , \nOut19_16[2] , 
        \nOut19_16[1] , \nOut19_16[0] }), .WestIn({\nOut17_16[7] , 
        \nOut17_16[6] , \nOut17_16[5] , \nOut17_16[4] , \nOut17_16[3] , 
        \nOut17_16[2] , \nOut17_16[1] , \nOut17_16[0] }), .Out({\nOut18_16[7] , 
        \nOut18_16[6] , \nOut18_16[5] , \nOut18_16[4] , \nOut18_16[3] , 
        \nOut18_16[2] , \nOut18_16[1] , \nOut18_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_732 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut733[7] , \nScanOut733[6] , 
        \nScanOut733[5] , \nScanOut733[4] , \nScanOut733[3] , \nScanOut733[2] , 
        \nScanOut733[1] , \nScanOut733[0] }), .ScanOut({\nScanOut732[7] , 
        \nScanOut732[6] , \nScanOut732[5] , \nScanOut732[4] , \nScanOut732[3] , 
        \nScanOut732[2] , \nScanOut732[1] , \nScanOut732[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_27[7] , \nOut22_27[6] , \nOut22_27[5] , \nOut22_27[4] , 
        \nOut22_27[3] , \nOut22_27[2] , \nOut22_27[1] , \nOut22_27[0] }), 
        .SouthIn({\nOut22_29[7] , \nOut22_29[6] , \nOut22_29[5] , 
        \nOut22_29[4] , \nOut22_29[3] , \nOut22_29[2] , \nOut22_29[1] , 
        \nOut22_29[0] }), .EastIn({\nOut23_28[7] , \nOut23_28[6] , 
        \nOut23_28[5] , \nOut23_28[4] , \nOut23_28[3] , \nOut23_28[2] , 
        \nOut23_28[1] , \nOut23_28[0] }), .WestIn({\nOut21_28[7] , 
        \nOut21_28[6] , \nOut21_28[5] , \nOut21_28[4] , \nOut21_28[3] , 
        \nOut21_28[2] , \nOut21_28[1] , \nOut21_28[0] }), .Out({\nOut22_28[7] , 
        \nOut22_28[6] , \nOut22_28[5] , \nOut22_28[4] , \nOut22_28[3] , 
        \nOut22_28[2] , \nOut22_28[1] , \nOut22_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_870 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut871[7] , \nScanOut871[6] , 
        \nScanOut871[5] , \nScanOut871[4] , \nScanOut871[3] , \nScanOut871[2] , 
        \nScanOut871[1] , \nScanOut871[0] }), .ScanOut({\nScanOut870[7] , 
        \nScanOut870[6] , \nScanOut870[5] , \nScanOut870[4] , \nScanOut870[3] , 
        \nScanOut870[2] , \nScanOut870[1] , \nScanOut870[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_5[7] , \nOut27_5[6] , \nOut27_5[5] , \nOut27_5[4] , 
        \nOut27_5[3] , \nOut27_5[2] , \nOut27_5[1] , \nOut27_5[0] }), 
        .SouthIn({\nOut27_7[7] , \nOut27_7[6] , \nOut27_7[5] , \nOut27_7[4] , 
        \nOut27_7[3] , \nOut27_7[2] , \nOut27_7[1] , \nOut27_7[0] }), .EastIn(
        {\nOut28_6[7] , \nOut28_6[6] , \nOut28_6[5] , \nOut28_6[4] , 
        \nOut28_6[3] , \nOut28_6[2] , \nOut28_6[1] , \nOut28_6[0] }), .WestIn(
        {\nOut26_6[7] , \nOut26_6[6] , \nOut26_6[5] , \nOut26_6[4] , 
        \nOut26_6[3] , \nOut26_6[2] , \nOut26_6[1] , \nOut26_6[0] }), .Out({
        \nOut27_6[7] , \nOut27_6[6] , \nOut27_6[5] , \nOut27_6[4] , 
        \nOut27_6[3] , \nOut27_6[2] , \nOut27_6[1] , \nOut27_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_234 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut235[7] , \nScanOut235[6] , 
        \nScanOut235[5] , \nScanOut235[4] , \nScanOut235[3] , \nScanOut235[2] , 
        \nScanOut235[1] , \nScanOut235[0] }), .ScanOut({\nScanOut234[7] , 
        \nScanOut234[6] , \nScanOut234[5] , \nScanOut234[4] , \nScanOut234[3] , 
        \nScanOut234[2] , \nScanOut234[1] , \nScanOut234[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_9[7] , \nOut7_9[6] , \nOut7_9[5] , \nOut7_9[4] , \nOut7_9[3] , 
        \nOut7_9[2] , \nOut7_9[1] , \nOut7_9[0] }), .SouthIn({\nOut7_11[7] , 
        \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , \nOut7_11[3] , 
        \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }), .EastIn({\nOut8_10[7] , 
        \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , \nOut8_10[3] , 
        \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }), .WestIn({\nOut6_10[7] , 
        \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , \nOut6_10[3] , 
        \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }), .Out({\nOut7_10[7] , 
        \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , \nOut7_10[3] , 
        \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_383 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut384[7] , \nScanOut384[6] , 
        \nScanOut384[5] , \nScanOut384[4] , \nScanOut384[3] , \nScanOut384[2] , 
        \nScanOut384[1] , \nScanOut384[0] }), .ScanOut({\nScanOut383[7] , 
        \nScanOut383[6] , \nScanOut383[5] , \nScanOut383[4] , \nScanOut383[3] , 
        \nScanOut383[2] , \nScanOut383[1] , \nScanOut383[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut11_31[7] , \nOut11_31[6] , 
        \nOut11_31[5] , \nOut11_31[4] , \nOut11_31[3] , \nOut11_31[2] , 
        \nOut11_31[1] , \nOut11_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_402 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut403[7] , \nScanOut403[6] , 
        \nScanOut403[5] , \nScanOut403[4] , \nScanOut403[3] , \nScanOut403[2] , 
        \nScanOut403[1] , \nScanOut403[0] }), .ScanOut({\nScanOut402[7] , 
        \nScanOut402[6] , \nScanOut402[5] , \nScanOut402[4] , \nScanOut402[3] , 
        \nScanOut402[2] , \nScanOut402[1] , \nScanOut402[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_17[7] , \nOut12_17[6] , \nOut12_17[5] , \nOut12_17[4] , 
        \nOut12_17[3] , \nOut12_17[2] , \nOut12_17[1] , \nOut12_17[0] }), 
        .SouthIn({\nOut12_19[7] , \nOut12_19[6] , \nOut12_19[5] , 
        \nOut12_19[4] , \nOut12_19[3] , \nOut12_19[2] , \nOut12_19[1] , 
        \nOut12_19[0] }), .EastIn({\nOut13_18[7] , \nOut13_18[6] , 
        \nOut13_18[5] , \nOut13_18[4] , \nOut13_18[3] , \nOut13_18[2] , 
        \nOut13_18[1] , \nOut13_18[0] }), .WestIn({\nOut11_18[7] , 
        \nOut11_18[6] , \nOut11_18[5] , \nOut11_18[4] , \nOut11_18[3] , 
        \nOut11_18[2] , \nOut11_18[1] , \nOut11_18[0] }), .Out({\nOut12_18[7] , 
        \nOut12_18[6] , \nOut12_18[5] , \nOut12_18[4] , \nOut12_18[3] , 
        \nOut12_18[2] , \nOut12_18[1] , \nOut12_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_425 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut426[7] , \nScanOut426[6] , 
        \nScanOut426[5] , \nScanOut426[4] , \nScanOut426[3] , \nScanOut426[2] , 
        \nScanOut426[1] , \nScanOut426[0] }), .ScanOut({\nScanOut425[7] , 
        \nScanOut425[6] , \nScanOut425[5] , \nScanOut425[4] , \nScanOut425[3] , 
        \nScanOut425[2] , \nScanOut425[1] , \nScanOut425[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }), 
        .SouthIn({\nOut13_10[7] , \nOut13_10[6] , \nOut13_10[5] , 
        \nOut13_10[4] , \nOut13_10[3] , \nOut13_10[2] , \nOut13_10[1] , 
        \nOut13_10[0] }), .EastIn({\nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , 
        \nOut14_9[4] , \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , 
        \nOut14_9[0] }), .WestIn({\nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , 
        \nOut12_9[4] , \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , 
        \nOut12_9[0] }), .Out({\nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , 
        \nOut13_9[4] , \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , 
        \nOut13_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_857 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut858[7] , \nScanOut858[6] , 
        \nScanOut858[5] , \nScanOut858[4] , \nScanOut858[3] , \nScanOut858[2] , 
        \nScanOut858[1] , \nScanOut858[0] }), .ScanOut({\nScanOut857[7] , 
        \nScanOut857[6] , \nScanOut857[5] , \nScanOut857[4] , \nScanOut857[3] , 
        \nScanOut857[2] , \nScanOut857[1] , \nScanOut857[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_24[7] , \nOut26_24[6] , \nOut26_24[5] , \nOut26_24[4] , 
        \nOut26_24[3] , \nOut26_24[2] , \nOut26_24[1] , \nOut26_24[0] }), 
        .SouthIn({\nOut26_26[7] , \nOut26_26[6] , \nOut26_26[5] , 
        \nOut26_26[4] , \nOut26_26[3] , \nOut26_26[2] , \nOut26_26[1] , 
        \nOut26_26[0] }), .EastIn({\nOut27_25[7] , \nOut27_25[6] , 
        \nOut27_25[5] , \nOut27_25[4] , \nOut27_25[3] , \nOut27_25[2] , 
        \nOut27_25[1] , \nOut27_25[0] }), .WestIn({\nOut25_25[7] , 
        \nOut25_25[6] , \nOut25_25[5] , \nOut25_25[4] , \nOut25_25[3] , 
        \nOut25_25[2] , \nOut25_25[1] , \nOut25_25[0] }), .Out({\nOut26_25[7] , 
        \nOut26_25[6] , \nOut26_25[5] , \nOut26_25[4] , \nOut26_25[3] , 
        \nOut26_25[2] , \nOut26_25[1] , \nOut26_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_715 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut716[7] , \nScanOut716[6] , 
        \nScanOut716[5] , \nScanOut716[4] , \nScanOut716[3] , \nScanOut716[2] , 
        \nScanOut716[1] , \nScanOut716[0] }), .ScanOut({\nScanOut715[7] , 
        \nScanOut715[6] , \nScanOut715[5] , \nScanOut715[4] , \nScanOut715[3] , 
        \nScanOut715[2] , \nScanOut715[1] , \nScanOut715[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_10[7] , \nOut22_10[6] , \nOut22_10[5] , \nOut22_10[4] , 
        \nOut22_10[3] , \nOut22_10[2] , \nOut22_10[1] , \nOut22_10[0] }), 
        .SouthIn({\nOut22_12[7] , \nOut22_12[6] , \nOut22_12[5] , 
        \nOut22_12[4] , \nOut22_12[3] , \nOut22_12[2] , \nOut22_12[1] , 
        \nOut22_12[0] }), .EastIn({\nOut23_11[7] , \nOut23_11[6] , 
        \nOut23_11[5] , \nOut23_11[4] , \nOut23_11[3] , \nOut23_11[2] , 
        \nOut23_11[1] , \nOut23_11[0] }), .WestIn({\nOut21_11[7] , 
        \nOut21_11[6] , \nOut21_11[5] , \nOut21_11[4] , \nOut21_11[3] , 
        \nOut21_11[2] , \nOut21_11[1] , \nOut21_11[0] }), .Out({\nOut22_11[7] , 
        \nOut22_11[6] , \nOut22_11[5] , \nOut22_11[4] , \nOut22_11[3] , 
        \nOut22_11[2] , \nOut22_11[1] , \nOut22_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_685 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut686[7] , \nScanOut686[6] , 
        \nScanOut686[5] , \nScanOut686[4] , \nScanOut686[3] , \nScanOut686[2] , 
        \nScanOut686[1] , \nScanOut686[0] }), .ScanOut({\nScanOut685[7] , 
        \nScanOut685[6] , \nScanOut685[5] , \nScanOut685[4] , \nScanOut685[3] , 
        \nScanOut685[2] , \nScanOut685[1] , \nScanOut685[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_12[7] , \nOut21_12[6] , \nOut21_12[5] , \nOut21_12[4] , 
        \nOut21_12[3] , \nOut21_12[2] , \nOut21_12[1] , \nOut21_12[0] }), 
        .SouthIn({\nOut21_14[7] , \nOut21_14[6] , \nOut21_14[5] , 
        \nOut21_14[4] , \nOut21_14[3] , \nOut21_14[2] , \nOut21_14[1] , 
        \nOut21_14[0] }), .EastIn({\nOut22_13[7] , \nOut22_13[6] , 
        \nOut22_13[5] , \nOut22_13[4] , \nOut22_13[3] , \nOut22_13[2] , 
        \nOut22_13[1] , \nOut22_13[0] }), .WestIn({\nOut20_13[7] , 
        \nOut20_13[6] , \nOut20_13[5] , \nOut20_13[4] , \nOut20_13[3] , 
        \nOut20_13[2] , \nOut20_13[1] , \nOut20_13[0] }), .Out({\nOut21_13[7] , 
        \nOut21_13[6] , \nOut21_13[5] , \nOut21_13[4] , \nOut21_13[3] , 
        \nOut21_13[2] , \nOut21_13[1] , \nOut21_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1013 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1014[7] , \nScanOut1014[6] , 
        \nScanOut1014[5] , \nScanOut1014[4] , \nScanOut1014[3] , 
        \nScanOut1014[2] , \nScanOut1014[1] , \nScanOut1014[0] }), .ScanOut({
        \nScanOut1013[7] , \nScanOut1013[6] , \nScanOut1013[5] , 
        \nScanOut1013[4] , \nScanOut1013[3] , \nScanOut1013[2] , 
        \nScanOut1013[1] , \nScanOut1013[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_21[7] , \nOut31_21[6] , \nOut31_21[5] , 
        \nOut31_21[4] , \nOut31_21[3] , \nOut31_21[2] , \nOut31_21[1] , 
        \nOut31_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_298 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut299[7] , \nScanOut299[6] , 
        \nScanOut299[5] , \nScanOut299[4] , \nScanOut299[3] , \nScanOut299[2] , 
        \nScanOut299[1] , \nScanOut299[0] }), .ScanOut({\nScanOut298[7] , 
        \nScanOut298[6] , \nScanOut298[5] , \nScanOut298[4] , \nScanOut298[3] , 
        \nScanOut298[2] , \nScanOut298[1] , \nScanOut298[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_9[7] , \nOut9_9[6] , \nOut9_9[5] , \nOut9_9[4] , \nOut9_9[3] , 
        \nOut9_9[2] , \nOut9_9[1] , \nOut9_9[0] }), .SouthIn({\nOut9_11[7] , 
        \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , \nOut9_11[3] , 
        \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }), .EastIn({\nOut10_10[7] , 
        \nOut10_10[6] , \nOut10_10[5] , \nOut10_10[4] , \nOut10_10[3] , 
        \nOut10_10[2] , \nOut10_10[1] , \nOut10_10[0] }), .WestIn({
        \nOut8_10[7] , \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , 
        \nOut8_10[3] , \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }), .Out({
        \nOut9_10[7] , \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , 
        \nOut9_10[3] , \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_519 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut520[7] , \nScanOut520[6] , 
        \nScanOut520[5] , \nScanOut520[4] , \nScanOut520[3] , \nScanOut520[2] , 
        \nScanOut520[1] , \nScanOut520[0] }), .ScanOut({\nScanOut519[7] , 
        \nScanOut519[6] , \nScanOut519[5] , \nScanOut519[4] , \nScanOut519[3] , 
        \nScanOut519[2] , \nScanOut519[1] , \nScanOut519[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_6[7] , \nOut16_6[6] , \nOut16_6[5] , \nOut16_6[4] , 
        \nOut16_6[3] , \nOut16_6[2] , \nOut16_6[1] , \nOut16_6[0] }), 
        .SouthIn({\nOut16_8[7] , \nOut16_8[6] , \nOut16_8[5] , \nOut16_8[4] , 
        \nOut16_8[3] , \nOut16_8[2] , \nOut16_8[1] , \nOut16_8[0] }), .EastIn(
        {\nOut17_7[7] , \nOut17_7[6] , \nOut17_7[5] , \nOut17_7[4] , 
        \nOut17_7[3] , \nOut17_7[2] , \nOut17_7[1] , \nOut17_7[0] }), .WestIn(
        {\nOut15_7[7] , \nOut15_7[6] , \nOut15_7[5] , \nOut15_7[4] , 
        \nOut15_7[3] , \nOut15_7[2] , \nOut15_7[1] , \nOut15_7[0] }), .Out({
        \nOut16_7[7] , \nOut16_7[6] , \nOut16_7[5] , \nOut16_7[4] , 
        \nOut16_7[3] , \nOut16_7[2] , \nOut16_7[1] , \nOut16_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_629 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut630[7] , \nScanOut630[6] , 
        \nScanOut630[5] , \nScanOut630[4] , \nScanOut630[3] , \nScanOut630[2] , 
        \nScanOut630[1] , \nScanOut630[0] }), .ScanOut({\nScanOut629[7] , 
        \nScanOut629[6] , \nScanOut629[5] , \nScanOut629[4] , \nScanOut629[3] , 
        \nScanOut629[2] , \nScanOut629[1] , \nScanOut629[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_20[7] , \nOut19_20[6] , \nOut19_20[5] , \nOut19_20[4] , 
        \nOut19_20[3] , \nOut19_20[2] , \nOut19_20[1] , \nOut19_20[0] }), 
        .SouthIn({\nOut19_22[7] , \nOut19_22[6] , \nOut19_22[5] , 
        \nOut19_22[4] , \nOut19_22[3] , \nOut19_22[2] , \nOut19_22[1] , 
        \nOut19_22[0] }), .EastIn({\nOut20_21[7] , \nOut20_21[6] , 
        \nOut20_21[5] , \nOut20_21[4] , \nOut20_21[3] , \nOut20_21[2] , 
        \nOut20_21[1] , \nOut20_21[0] }), .WestIn({\nOut18_21[7] , 
        \nOut18_21[6] , \nOut18_21[5] , \nOut18_21[4] , \nOut18_21[3] , 
        \nOut18_21[2] , \nOut18_21[1] , \nOut18_21[0] }), .Out({\nOut19_21[7] , 
        \nOut19_21[6] , \nOut19_21[5] , \nOut19_21[4] , \nOut19_21[3] , 
        \nOut19_21[2] , \nOut19_21[1] , \nOut19_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_308 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut309[7] , \nScanOut309[6] , 
        \nScanOut309[5] , \nScanOut309[4] , \nScanOut309[3] , \nScanOut309[2] , 
        \nScanOut309[1] , \nScanOut309[0] }), .ScanOut({\nScanOut308[7] , 
        \nScanOut308[6] , \nScanOut308[5] , \nScanOut308[4] , \nScanOut308[3] , 
        \nScanOut308[2] , \nScanOut308[1] , \nScanOut308[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_19[7] , \nOut9_19[6] , \nOut9_19[5] , \nOut9_19[4] , 
        \nOut9_19[3] , \nOut9_19[2] , \nOut9_19[1] , \nOut9_19[0] }), 
        .SouthIn({\nOut9_21[7] , \nOut9_21[6] , \nOut9_21[5] , \nOut9_21[4] , 
        \nOut9_21[3] , \nOut9_21[2] , \nOut9_21[1] , \nOut9_21[0] }), .EastIn(
        {\nOut10_20[7] , \nOut10_20[6] , \nOut10_20[5] , \nOut10_20[4] , 
        \nOut10_20[3] , \nOut10_20[2] , \nOut10_20[1] , \nOut10_20[0] }), 
        .WestIn({\nOut8_20[7] , \nOut8_20[6] , \nOut8_20[5] , \nOut8_20[4] , 
        \nOut8_20[3] , \nOut8_20[2] , \nOut8_20[1] , \nOut8_20[0] }), .Out({
        \nOut9_20[7] , \nOut9_20[6] , \nOut9_20[5] , \nOut9_20[4] , 
        \nOut9_20[3] , \nOut9_20[2] , \nOut9_20[1] , \nOut9_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_489 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut490[7] , \nScanOut490[6] , 
        \nScanOut490[5] , \nScanOut490[4] , \nScanOut490[3] , \nScanOut490[2] , 
        \nScanOut490[1] , \nScanOut490[0] }), .ScanOut({\nScanOut489[7] , 
        \nScanOut489[6] , \nScanOut489[5] , \nScanOut489[4] , \nScanOut489[3] , 
        \nScanOut489[2] , \nScanOut489[1] , \nScanOut489[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_8[7] , \nOut15_8[6] , \nOut15_8[5] , \nOut15_8[4] , 
        \nOut15_8[3] , \nOut15_8[2] , \nOut15_8[1] , \nOut15_8[0] }), 
        .SouthIn({\nOut15_10[7] , \nOut15_10[6] , \nOut15_10[5] , 
        \nOut15_10[4] , \nOut15_10[3] , \nOut15_10[2] , \nOut15_10[1] , 
        \nOut15_10[0] }), .EastIn({\nOut16_9[7] , \nOut16_9[6] , \nOut16_9[5] , 
        \nOut16_9[4] , \nOut16_9[3] , \nOut16_9[2] , \nOut16_9[1] , 
        \nOut16_9[0] }), .WestIn({\nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , 
        \nOut14_9[4] , \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , 
        \nOut14_9[0] }), .Out({\nOut15_9[7] , \nOut15_9[6] , \nOut15_9[5] , 
        \nOut15_9[4] , \nOut15_9[3] , \nOut15_9[2] , \nOut15_9[1] , 
        \nOut15_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_341 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut342[7] , \nScanOut342[6] , 
        \nScanOut342[5] , \nScanOut342[4] , \nScanOut342[3] , \nScanOut342[2] , 
        \nScanOut342[1] , \nScanOut342[0] }), .ScanOut({\nScanOut341[7] , 
        \nScanOut341[6] , \nScanOut341[5] , \nScanOut341[4] , \nScanOut341[3] , 
        \nScanOut341[2] , \nScanOut341[1] , \nScanOut341[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_20[7] , \nOut10_20[6] , \nOut10_20[5] , \nOut10_20[4] , 
        \nOut10_20[3] , \nOut10_20[2] , \nOut10_20[1] , \nOut10_20[0] }), 
        .SouthIn({\nOut10_22[7] , \nOut10_22[6] , \nOut10_22[5] , 
        \nOut10_22[4] , \nOut10_22[3] , \nOut10_22[2] , \nOut10_22[1] , 
        \nOut10_22[0] }), .EastIn({\nOut11_21[7] , \nOut11_21[6] , 
        \nOut11_21[5] , \nOut11_21[4] , \nOut11_21[3] , \nOut11_21[2] , 
        \nOut11_21[1] , \nOut11_21[0] }), .WestIn({\nOut9_21[7] , 
        \nOut9_21[6] , \nOut9_21[5] , \nOut9_21[4] , \nOut9_21[3] , 
        \nOut9_21[2] , \nOut9_21[1] , \nOut9_21[0] }), .Out({\nOut10_21[7] , 
        \nOut10_21[6] , \nOut10_21[5] , \nOut10_21[4] , \nOut10_21[3] , 
        \nOut10_21[2] , \nOut10_21[1] , \nOut10_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_550 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut551[7] , \nScanOut551[6] , 
        \nScanOut551[5] , \nScanOut551[4] , \nScanOut551[3] , \nScanOut551[2] , 
        \nScanOut551[1] , \nScanOut551[0] }), .ScanOut({\nScanOut550[7] , 
        \nScanOut550[6] , \nScanOut550[5] , \nScanOut550[4] , \nScanOut550[3] , 
        \nScanOut550[2] , \nScanOut550[1] , \nScanOut550[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_5[7] , \nOut17_5[6] , \nOut17_5[5] , \nOut17_5[4] , 
        \nOut17_5[3] , \nOut17_5[2] , \nOut17_5[1] , \nOut17_5[0] }), 
        .SouthIn({\nOut17_7[7] , \nOut17_7[6] , \nOut17_7[5] , \nOut17_7[4] , 
        \nOut17_7[3] , \nOut17_7[2] , \nOut17_7[1] , \nOut17_7[0] }), .EastIn(
        {\nOut18_6[7] , \nOut18_6[6] , \nOut18_6[5] , \nOut18_6[4] , 
        \nOut18_6[3] , \nOut18_6[2] , \nOut18_6[1] , \nOut18_6[0] }), .WestIn(
        {\nOut16_6[7] , \nOut16_6[6] , \nOut16_6[5] , \nOut16_6[4] , 
        \nOut16_6[3] , \nOut16_6[2] , \nOut16_6[1] , \nOut16_6[0] }), .Out({
        \nOut17_6[7] , \nOut17_6[6] , \nOut17_6[5] , \nOut17_6[4] , 
        \nOut17_6[3] , \nOut17_6[2] , \nOut17_6[1] , \nOut17_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_922 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut923[7] , \nScanOut923[6] , 
        \nScanOut923[5] , \nScanOut923[4] , \nScanOut923[3] , \nScanOut923[2] , 
        \nScanOut923[1] , \nScanOut923[0] }), .ScanOut({\nScanOut922[7] , 
        \nScanOut922[6] , \nScanOut922[5] , \nScanOut922[4] , \nScanOut922[3] , 
        \nScanOut922[2] , \nScanOut922[1] , \nScanOut922[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_25[7] , \nOut28_25[6] , \nOut28_25[5] , \nOut28_25[4] , 
        \nOut28_25[3] , \nOut28_25[2] , \nOut28_25[1] , \nOut28_25[0] }), 
        .SouthIn({\nOut28_27[7] , \nOut28_27[6] , \nOut28_27[5] , 
        \nOut28_27[4] , \nOut28_27[3] , \nOut28_27[2] , \nOut28_27[1] , 
        \nOut28_27[0] }), .EastIn({\nOut29_26[7] , \nOut29_26[6] , 
        \nOut29_26[5] , \nOut29_26[4] , \nOut29_26[3] , \nOut29_26[2] , 
        \nOut29_26[1] , \nOut29_26[0] }), .WestIn({\nOut27_26[7] , 
        \nOut27_26[6] , \nOut27_26[5] , \nOut27_26[4] , \nOut27_26[3] , 
        \nOut27_26[2] , \nOut27_26[1] , \nOut27_26[0] }), .Out({\nOut28_26[7] , 
        \nOut28_26[6] , \nOut28_26[5] , \nOut28_26[4] , \nOut28_26[3] , 
        \nOut28_26[2] , \nOut28_26[1] , \nOut28_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_660 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut661[7] , \nScanOut661[6] , 
        \nScanOut661[5] , \nScanOut661[4] , \nScanOut661[3] , \nScanOut661[2] , 
        \nScanOut661[1] , \nScanOut661[0] }), .ScanOut({\nScanOut660[7] , 
        \nScanOut660[6] , \nScanOut660[5] , \nScanOut660[4] , \nScanOut660[3] , 
        \nScanOut660[2] , \nScanOut660[1] , \nScanOut660[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_19[7] , \nOut20_19[6] , \nOut20_19[5] , \nOut20_19[4] , 
        \nOut20_19[3] , \nOut20_19[2] , \nOut20_19[1] , \nOut20_19[0] }), 
        .SouthIn({\nOut20_21[7] , \nOut20_21[6] , \nOut20_21[5] , 
        \nOut20_21[4] , \nOut20_21[3] , \nOut20_21[2] , \nOut20_21[1] , 
        \nOut20_21[0] }), .EastIn({\nOut21_20[7] , \nOut21_20[6] , 
        \nOut21_20[5] , \nOut21_20[4] , \nOut21_20[3] , \nOut21_20[2] , 
        \nOut21_20[1] , \nOut21_20[0] }), .WestIn({\nOut19_20[7] , 
        \nOut19_20[6] , \nOut19_20[5] , \nOut19_20[4] , \nOut19_20[3] , 
        \nOut19_20[2] , \nOut19_20[1] , \nOut19_20[0] }), .Out({\nOut20_20[7] , 
        \nOut20_20[6] , \nOut20_20[5] , \nOut20_20[4] , \nOut20_20[3] , 
        \nOut20_20[2] , \nOut20_20[1] , \nOut20_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_156 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut157[7] , \nScanOut157[6] , 
        \nScanOut157[5] , \nScanOut157[4] , \nScanOut157[3] , \nScanOut157[2] , 
        \nScanOut157[1] , \nScanOut157[0] }), .ScanOut({\nScanOut156[7] , 
        \nScanOut156[6] , \nScanOut156[5] , \nScanOut156[4] , \nScanOut156[3] , 
        \nScanOut156[2] , \nScanOut156[1] , \nScanOut156[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_27[7] , \nOut4_27[6] , \nOut4_27[5] , \nOut4_27[4] , 
        \nOut4_27[3] , \nOut4_27[2] , \nOut4_27[1] , \nOut4_27[0] }), 
        .SouthIn({\nOut4_29[7] , \nOut4_29[6] , \nOut4_29[5] , \nOut4_29[4] , 
        \nOut4_29[3] , \nOut4_29[2] , \nOut4_29[1] , \nOut4_29[0] }), .EastIn(
        {\nOut5_28[7] , \nOut5_28[6] , \nOut5_28[5] , \nOut5_28[4] , 
        \nOut5_28[3] , \nOut5_28[2] , \nOut5_28[1] , \nOut5_28[0] }), .WestIn(
        {\nOut3_28[7] , \nOut3_28[6] , \nOut3_28[5] , \nOut3_28[4] , 
        \nOut3_28[3] , \nOut3_28[2] , \nOut3_28[1] , \nOut3_28[0] }), .Out({
        \nOut4_28[7] , \nOut4_28[6] , \nOut4_28[5] , \nOut4_28[4] , 
        \nOut4_28[3] , \nOut4_28[2] , \nOut4_28[1] , \nOut4_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_266 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut267[7] , \nScanOut267[6] , 
        \nScanOut267[5] , \nScanOut267[4] , \nScanOut267[3] , \nScanOut267[2] , 
        \nScanOut267[1] , \nScanOut267[0] }), .ScanOut({\nScanOut266[7] , 
        \nScanOut266[6] , \nScanOut266[5] , \nScanOut266[4] , \nScanOut266[3] , 
        \nScanOut266[2] , \nScanOut266[1] , \nScanOut266[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_9[7] , \nOut8_9[6] , \nOut8_9[5] , \nOut8_9[4] , \nOut8_9[3] , 
        \nOut8_9[2] , \nOut8_9[1] , \nOut8_9[0] }), .SouthIn({\nOut8_11[7] , 
        \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , \nOut8_11[3] , 
        \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }), .EastIn({\nOut9_10[7] , 
        \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , \nOut9_10[3] , 
        \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }), .WestIn({\nOut7_10[7] , 
        \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , \nOut7_10[3] , 
        \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }), .Out({\nOut8_10[7] , 
        \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , \nOut8_10[3] , 
        \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_366 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut367[7] , \nScanOut367[6] , 
        \nScanOut367[5] , \nScanOut367[4] , \nScanOut367[3] , \nScanOut367[2] , 
        \nScanOut367[1] , \nScanOut367[0] }), .ScanOut({\nScanOut366[7] , 
        \nScanOut366[6] , \nScanOut366[5] , \nScanOut366[4] , \nScanOut366[3] , 
        \nScanOut366[2] , \nScanOut366[1] , \nScanOut366[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_13[7] , \nOut11_13[6] , \nOut11_13[5] , \nOut11_13[4] , 
        \nOut11_13[3] , \nOut11_13[2] , \nOut11_13[1] , \nOut11_13[0] }), 
        .SouthIn({\nOut11_15[7] , \nOut11_15[6] , \nOut11_15[5] , 
        \nOut11_15[4] , \nOut11_15[3] , \nOut11_15[2] , \nOut11_15[1] , 
        \nOut11_15[0] }), .EastIn({\nOut12_14[7] , \nOut12_14[6] , 
        \nOut12_14[5] , \nOut12_14[4] , \nOut12_14[3] , \nOut12_14[2] , 
        \nOut12_14[1] , \nOut12_14[0] }), .WestIn({\nOut10_14[7] , 
        \nOut10_14[6] , \nOut10_14[5] , \nOut10_14[4] , \nOut10_14[3] , 
        \nOut10_14[2] , \nOut10_14[1] , \nOut10_14[0] }), .Out({\nOut11_14[7] , 
        \nOut11_14[6] , \nOut11_14[5] , \nOut11_14[4] , \nOut11_14[3] , 
        \nOut11_14[2] , \nOut11_14[1] , \nOut11_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_647 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut648[7] , \nScanOut648[6] , 
        \nScanOut648[5] , \nScanOut648[4] , \nScanOut648[3] , \nScanOut648[2] , 
        \nScanOut648[1] , \nScanOut648[0] }), .ScanOut({\nScanOut647[7] , 
        \nScanOut647[6] , \nScanOut647[5] , \nScanOut647[4] , \nScanOut647[3] , 
        \nScanOut647[2] , \nScanOut647[1] , \nScanOut647[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_6[7] , \nOut20_6[6] , \nOut20_6[5] , \nOut20_6[4] , 
        \nOut20_6[3] , \nOut20_6[2] , \nOut20_6[1] , \nOut20_6[0] }), 
        .SouthIn({\nOut20_8[7] , \nOut20_8[6] , \nOut20_8[5] , \nOut20_8[4] , 
        \nOut20_8[3] , \nOut20_8[2] , \nOut20_8[1] , \nOut20_8[0] }), .EastIn(
        {\nOut21_7[7] , \nOut21_7[6] , \nOut21_7[5] , \nOut21_7[4] , 
        \nOut21_7[3] , \nOut21_7[2] , \nOut21_7[1] , \nOut21_7[0] }), .WestIn(
        {\nOut19_7[7] , \nOut19_7[6] , \nOut19_7[5] , \nOut19_7[4] , 
        \nOut19_7[3] , \nOut19_7[2] , \nOut19_7[1] , \nOut19_7[0] }), .Out({
        \nOut20_7[7] , \nOut20_7[6] , \nOut20_7[5] , \nOut20_7[4] , 
        \nOut20_7[3] , \nOut20_7[2] , \nOut20_7[1] , \nOut20_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_895 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut896[7] , \nScanOut896[6] , 
        \nScanOut896[5] , \nScanOut896[4] , \nScanOut896[3] , \nScanOut896[2] , 
        \nScanOut896[1] , \nScanOut896[0] }), .ScanOut({\nScanOut895[7] , 
        \nScanOut895[6] , \nScanOut895[5] , \nScanOut895[4] , \nScanOut895[3] , 
        \nScanOut895[2] , \nScanOut895[1] , \nScanOut895[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut27_31[7] , \nOut27_31[6] , 
        \nOut27_31[5] , \nOut27_31[4] , \nOut27_31[3] , \nOut27_31[2] , 
        \nOut27_31[1] , \nOut27_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_905 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut906[7] , \nScanOut906[6] , 
        \nScanOut906[5] , \nScanOut906[4] , \nScanOut906[3] , \nScanOut906[2] , 
        \nScanOut906[1] , \nScanOut906[0] }), .ScanOut({\nScanOut905[7] , 
        \nScanOut905[6] , \nScanOut905[5] , \nScanOut905[4] , \nScanOut905[3] , 
        \nScanOut905[2] , \nScanOut905[1] , \nScanOut905[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_8[7] , \nOut28_8[6] , \nOut28_8[5] , \nOut28_8[4] , 
        \nOut28_8[3] , \nOut28_8[2] , \nOut28_8[1] , \nOut28_8[0] }), 
        .SouthIn({\nOut28_10[7] , \nOut28_10[6] , \nOut28_10[5] , 
        \nOut28_10[4] , \nOut28_10[3] , \nOut28_10[2] , \nOut28_10[1] , 
        \nOut28_10[0] }), .EastIn({\nOut29_9[7] , \nOut29_9[6] , \nOut29_9[5] , 
        \nOut29_9[4] , \nOut29_9[3] , \nOut29_9[2] , \nOut29_9[1] , 
        \nOut29_9[0] }), .WestIn({\nOut27_9[7] , \nOut27_9[6] , \nOut27_9[5] , 
        \nOut27_9[4] , \nOut27_9[3] , \nOut27_9[2] , \nOut27_9[1] , 
        \nOut27_9[0] }), .Out({\nOut28_9[7] , \nOut28_9[6] , \nOut28_9[5] , 
        \nOut28_9[4] , \nOut28_9[3] , \nOut28_9[2] , \nOut28_9[1] , 
        \nOut28_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_477 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut478[7] , \nScanOut478[6] , 
        \nScanOut478[5] , \nScanOut478[4] , \nScanOut478[3] , \nScanOut478[2] , 
        \nScanOut478[1] , \nScanOut478[0] }), .ScanOut({\nScanOut477[7] , 
        \nScanOut477[6] , \nScanOut477[5] , \nScanOut477[4] , \nScanOut477[3] , 
        \nScanOut477[2] , \nScanOut477[1] , \nScanOut477[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_28[7] , \nOut14_28[6] , \nOut14_28[5] , \nOut14_28[4] , 
        \nOut14_28[3] , \nOut14_28[2] , \nOut14_28[1] , \nOut14_28[0] }), 
        .SouthIn({\nOut14_30[7] , \nOut14_30[6] , \nOut14_30[5] , 
        \nOut14_30[4] , \nOut14_30[3] , \nOut14_30[2] , \nOut14_30[1] , 
        \nOut14_30[0] }), .EastIn({\nOut15_29[7] , \nOut15_29[6] , 
        \nOut15_29[5] , \nOut15_29[4] , \nOut15_29[3] , \nOut15_29[2] , 
        \nOut15_29[1] , \nOut15_29[0] }), .WestIn({\nOut13_29[7] , 
        \nOut13_29[6] , \nOut13_29[5] , \nOut13_29[4] , \nOut13_29[3] , 
        \nOut13_29[2] , \nOut13_29[1] , \nOut13_29[0] }), .Out({\nOut14_29[7] , 
        \nOut14_29[6] , \nOut14_29[5] , \nOut14_29[4] , \nOut14_29[3] , 
        \nOut14_29[2] , \nOut14_29[1] , \nOut14_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_577 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut578[7] , \nScanOut578[6] , 
        \nScanOut578[5] , \nScanOut578[4] , \nScanOut578[3] , \nScanOut578[2] , 
        \nScanOut578[1] , \nScanOut578[0] }), .ScanOut({\nScanOut577[7] , 
        \nScanOut577[6] , \nScanOut577[5] , \nScanOut577[4] , \nScanOut577[3] , 
        \nScanOut577[2] , \nScanOut577[1] , \nScanOut577[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_0[7] , \nOut18_0[6] , \nOut18_0[5] , \nOut18_0[4] , 
        \nOut18_0[3] , \nOut18_0[2] , \nOut18_0[1] , \nOut18_0[0] }), 
        .SouthIn({\nOut18_2[7] , \nOut18_2[6] , \nOut18_2[5] , \nOut18_2[4] , 
        \nOut18_2[3] , \nOut18_2[2] , \nOut18_2[1] , \nOut18_2[0] }), .EastIn(
        {\nOut19_1[7] , \nOut19_1[6] , \nOut19_1[5] , \nOut19_1[4] , 
        \nOut19_1[3] , \nOut19_1[2] , \nOut19_1[1] , \nOut19_1[0] }), .WestIn(
        {\nOut17_1[7] , \nOut17_1[6] , \nOut17_1[5] , \nOut17_1[4] , 
        \nOut17_1[3] , \nOut17_1[2] , \nOut17_1[1] , \nOut17_1[0] }), .Out({
        \nOut18_1[7] , \nOut18_1[6] , \nOut18_1[5] , \nOut18_1[4] , 
        \nOut18_1[3] , \nOut18_1[2] , \nOut18_1[1] , \nOut18_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_805 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut806[7] , \nScanOut806[6] , 
        \nScanOut806[5] , \nScanOut806[4] , \nScanOut806[3] , \nScanOut806[2] , 
        \nScanOut806[1] , \nScanOut806[0] }), .ScanOut({\nScanOut805[7] , 
        \nScanOut805[6] , \nScanOut805[5] , \nScanOut805[4] , \nScanOut805[3] , 
        \nScanOut805[2] , \nScanOut805[1] , \nScanOut805[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_4[7] , \nOut25_4[6] , \nOut25_4[5] , \nOut25_4[4] , 
        \nOut25_4[3] , \nOut25_4[2] , \nOut25_4[1] , \nOut25_4[0] }), 
        .SouthIn({\nOut25_6[7] , \nOut25_6[6] , \nOut25_6[5] , \nOut25_6[4] , 
        \nOut25_6[3] , \nOut25_6[2] , \nOut25_6[1] , \nOut25_6[0] }), .EastIn(
        {\nOut26_5[7] , \nOut26_5[6] , \nOut26_5[5] , \nOut26_5[4] , 
        \nOut26_5[3] , \nOut26_5[2] , \nOut26_5[1] , \nOut26_5[0] }), .WestIn(
        {\nOut24_5[7] , \nOut24_5[6] , \nOut24_5[5] , \nOut24_5[4] , 
        \nOut24_5[3] , \nOut24_5[2] , \nOut24_5[1] , \nOut24_5[0] }), .Out({
        \nOut25_5[7] , \nOut25_5[6] , \nOut25_5[5] , \nOut25_5[4] , 
        \nOut25_5[3] , \nOut25_5[2] , \nOut25_5[1] , \nOut25_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_839 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut840[7] , \nScanOut840[6] , 
        \nScanOut840[5] , \nScanOut840[4] , \nScanOut840[3] , \nScanOut840[2] , 
        \nScanOut840[1] , \nScanOut840[0] }), .ScanOut({\nScanOut839[7] , 
        \nScanOut839[6] , \nScanOut839[5] , \nScanOut839[4] , \nScanOut839[3] , 
        \nScanOut839[2] , \nScanOut839[1] , \nScanOut839[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_6[7] , \nOut26_6[6] , \nOut26_6[5] , \nOut26_6[4] , 
        \nOut26_6[3] , \nOut26_6[2] , \nOut26_6[1] , \nOut26_6[0] }), 
        .SouthIn({\nOut26_8[7] , \nOut26_8[6] , \nOut26_8[5] , \nOut26_8[4] , 
        \nOut26_8[3] , \nOut26_8[2] , \nOut26_8[1] , \nOut26_8[0] }), .EastIn(
        {\nOut27_7[7] , \nOut27_7[6] , \nOut27_7[5] , \nOut27_7[4] , 
        \nOut27_7[3] , \nOut27_7[2] , \nOut27_7[1] , \nOut27_7[0] }), .WestIn(
        {\nOut25_7[7] , \nOut25_7[6] , \nOut25_7[5] , \nOut25_7[4] , 
        \nOut25_7[3] , \nOut25_7[2] , \nOut25_7[1] , \nOut25_7[0] }), .Out({
        \nOut26_7[7] , \nOut26_7[6] , \nOut26_7[5] , \nOut26_7[4] , 
        \nOut26_7[3] , \nOut26_7[2] , \nOut26_7[1] , \nOut26_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_995 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut996[7] , \nScanOut996[6] , 
        \nScanOut996[5] , \nScanOut996[4] , \nScanOut996[3] , \nScanOut996[2] , 
        \nScanOut996[1] , \nScanOut996[0] }), .ScanOut({\nScanOut995[7] , 
        \nScanOut995[6] , \nScanOut995[5] , \nScanOut995[4] , \nScanOut995[3] , 
        \nScanOut995[2] , \nScanOut995[1] , \nScanOut995[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut31_3[7] , \nOut31_3[6] , 
        \nOut31_3[5] , \nOut31_3[4] , \nOut31_3[3] , \nOut31_3[2] , 
        \nOut31_3[1] , \nOut31_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_747 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut748[7] , \nScanOut748[6] , 
        \nScanOut748[5] , \nScanOut748[4] , \nScanOut748[3] , \nScanOut748[2] , 
        \nScanOut748[1] , \nScanOut748[0] }), .ScanOut({\nScanOut747[7] , 
        \nScanOut747[6] , \nScanOut747[5] , \nScanOut747[4] , \nScanOut747[3] , 
        \nScanOut747[2] , \nScanOut747[1] , \nScanOut747[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_10[7] , \nOut23_10[6] , \nOut23_10[5] , \nOut23_10[4] , 
        \nOut23_10[3] , \nOut23_10[2] , \nOut23_10[1] , \nOut23_10[0] }), 
        .SouthIn({\nOut23_12[7] , \nOut23_12[6] , \nOut23_12[5] , 
        \nOut23_12[4] , \nOut23_12[3] , \nOut23_12[2] , \nOut23_12[1] , 
        \nOut23_12[0] }), .EastIn({\nOut24_11[7] , \nOut24_11[6] , 
        \nOut24_11[5] , \nOut24_11[4] , \nOut24_11[3] , \nOut24_11[2] , 
        \nOut24_11[1] , \nOut24_11[0] }), .WestIn({\nOut22_11[7] , 
        \nOut22_11[6] , \nOut22_11[5] , \nOut22_11[4] , \nOut22_11[3] , 
        \nOut22_11[2] , \nOut22_11[1] , \nOut22_11[0] }), .Out({\nOut23_11[7] , 
        \nOut23_11[6] , \nOut23_11[5] , \nOut23_11[4] , \nOut23_11[3] , 
        \nOut23_11[2] , \nOut23_11[1] , \nOut23_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_171 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut172[7] , \nScanOut172[6] , 
        \nScanOut172[5] , \nScanOut172[4] , \nScanOut172[3] , \nScanOut172[2] , 
        \nScanOut172[1] , \nScanOut172[0] }), .ScanOut({\nScanOut171[7] , 
        \nScanOut171[6] , \nScanOut171[5] , \nScanOut171[4] , \nScanOut171[3] , 
        \nScanOut171[2] , \nScanOut171[1] , \nScanOut171[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_10[7] , \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , 
        \nOut5_10[3] , \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }), 
        .SouthIn({\nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }), .EastIn(
        {\nOut6_11[7] , \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , 
        \nOut6_11[3] , \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }), .WestIn(
        {\nOut4_11[7] , \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , 
        \nOut4_11[3] , \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }), .Out({
        \nOut5_11[7] , \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , 
        \nOut5_11[3] , \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_241 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut242[7] , \nScanOut242[6] , 
        \nScanOut242[5] , \nScanOut242[4] , \nScanOut242[3] , \nScanOut242[2] , 
        \nScanOut242[1] , \nScanOut242[0] }), .ScanOut({\nScanOut241[7] , 
        \nScanOut241[6] , \nScanOut241[5] , \nScanOut241[4] , \nScanOut241[3] , 
        \nScanOut241[2] , \nScanOut241[1] , \nScanOut241[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_16[7] , \nOut7_16[6] , \nOut7_16[5] , \nOut7_16[4] , 
        \nOut7_16[3] , \nOut7_16[2] , \nOut7_16[1] , \nOut7_16[0] }), 
        .SouthIn({\nOut7_18[7] , \nOut7_18[6] , \nOut7_18[5] , \nOut7_18[4] , 
        \nOut7_18[3] , \nOut7_18[2] , \nOut7_18[1] , \nOut7_18[0] }), .EastIn(
        {\nOut8_17[7] , \nOut8_17[6] , \nOut8_17[5] , \nOut8_17[4] , 
        \nOut8_17[3] , \nOut8_17[2] , \nOut8_17[1] , \nOut8_17[0] }), .WestIn(
        {\nOut6_17[7] , \nOut6_17[6] , \nOut6_17[5] , \nOut6_17[4] , 
        \nOut6_17[3] , \nOut6_17[2] , \nOut6_17[1] , \nOut6_17[0] }), .Out({
        \nOut7_17[7] , \nOut7_17[6] , \nOut7_17[5] , \nOut7_17[4] , 
        \nOut7_17[3] , \nOut7_17[2] , \nOut7_17[1] , \nOut7_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_760 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut761[7] , \nScanOut761[6] , 
        \nScanOut761[5] , \nScanOut761[4] , \nScanOut761[3] , \nScanOut761[2] , 
        \nScanOut761[1] , \nScanOut761[0] }), .ScanOut({\nScanOut760[7] , 
        \nScanOut760[6] , \nScanOut760[5] , \nScanOut760[4] , \nScanOut760[3] , 
        \nScanOut760[2] , \nScanOut760[1] , \nScanOut760[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_23[7] , \nOut23_23[6] , \nOut23_23[5] , \nOut23_23[4] , 
        \nOut23_23[3] , \nOut23_23[2] , \nOut23_23[1] , \nOut23_23[0] }), 
        .SouthIn({\nOut23_25[7] , \nOut23_25[6] , \nOut23_25[5] , 
        \nOut23_25[4] , \nOut23_25[3] , \nOut23_25[2] , \nOut23_25[1] , 
        \nOut23_25[0] }), .EastIn({\nOut24_24[7] , \nOut24_24[6] , 
        \nOut24_24[5] , \nOut24_24[4] , \nOut24_24[3] , \nOut24_24[2] , 
        \nOut24_24[1] , \nOut24_24[0] }), .WestIn({\nOut22_24[7] , 
        \nOut22_24[6] , \nOut22_24[5] , \nOut22_24[4] , \nOut22_24[3] , 
        \nOut22_24[2] , \nOut22_24[1] , \nOut22_24[0] }), .Out({\nOut23_24[7] , 
        \nOut23_24[6] , \nOut23_24[5] , \nOut23_24[4] , \nOut23_24[3] , 
        \nOut23_24[2] , \nOut23_24[1] , \nOut23_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_822 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut823[7] , \nScanOut823[6] , 
        \nScanOut823[5] , \nScanOut823[4] , \nScanOut823[3] , \nScanOut823[2] , 
        \nScanOut823[1] , \nScanOut823[0] }), .ScanOut({\nScanOut822[7] , 
        \nScanOut822[6] , \nScanOut822[5] , \nScanOut822[4] , \nScanOut822[3] , 
        \nScanOut822[2] , \nScanOut822[1] , \nScanOut822[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_21[7] , \nOut25_21[6] , \nOut25_21[5] , \nOut25_21[4] , 
        \nOut25_21[3] , \nOut25_21[2] , \nOut25_21[1] , \nOut25_21[0] }), 
        .SouthIn({\nOut25_23[7] , \nOut25_23[6] , \nOut25_23[5] , 
        \nOut25_23[4] , \nOut25_23[3] , \nOut25_23[2] , \nOut25_23[1] , 
        \nOut25_23[0] }), .EastIn({\nOut26_22[7] , \nOut26_22[6] , 
        \nOut26_22[5] , \nOut26_22[4] , \nOut26_22[3] , \nOut26_22[2] , 
        \nOut26_22[1] , \nOut26_22[0] }), .WestIn({\nOut24_22[7] , 
        \nOut24_22[6] , \nOut24_22[5] , \nOut24_22[4] , \nOut24_22[3] , 
        \nOut24_22[2] , \nOut24_22[1] , \nOut24_22[0] }), .Out({\nOut25_22[7] , 
        \nOut25_22[6] , \nOut25_22[5] , \nOut25_22[4] , \nOut25_22[3] , 
        \nOut25_22[2] , \nOut25_22[1] , \nOut25_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_450 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut451[7] , \nScanOut451[6] , 
        \nScanOut451[5] , \nScanOut451[4] , \nScanOut451[3] , \nScanOut451[2] , 
        \nScanOut451[1] , \nScanOut451[0] }), .ScanOut({\nScanOut450[7] , 
        \nScanOut450[6] , \nScanOut450[5] , \nScanOut450[4] , \nScanOut450[3] , 
        \nScanOut450[2] , \nScanOut450[1] , \nScanOut450[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_1[7] , \nOut14_1[6] , \nOut14_1[5] , \nOut14_1[4] , 
        \nOut14_1[3] , \nOut14_1[2] , \nOut14_1[1] , \nOut14_1[0] }), 
        .SouthIn({\nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }), .EastIn(
        {\nOut15_2[7] , \nOut15_2[6] , \nOut15_2[5] , \nOut15_2[4] , 
        \nOut15_2[3] , \nOut15_2[2] , \nOut15_2[1] , \nOut15_2[0] }), .WestIn(
        {\nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }), .Out({
        \nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_194 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut195[7] , \nScanOut195[6] , 
        \nScanOut195[5] , \nScanOut195[4] , \nScanOut195[3] , \nScanOut195[2] , 
        \nScanOut195[1] , \nScanOut195[0] }), .ScanOut({\nScanOut194[7] , 
        \nScanOut194[6] , \nScanOut194[5] , \nScanOut194[4] , \nScanOut194[3] , 
        \nScanOut194[2] , \nScanOut194[1] , \nScanOut194[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_1[7] , \nOut6_1[6] , \nOut6_1[5] , \nOut6_1[4] , \nOut6_1[3] , 
        \nOut6_1[2] , \nOut6_1[1] , \nOut6_1[0] }), .SouthIn({\nOut6_3[7] , 
        \nOut6_3[6] , \nOut6_3[5] , \nOut6_3[4] , \nOut6_3[3] , \nOut6_3[2] , 
        \nOut6_3[1] , \nOut6_3[0] }), .EastIn({\nOut7_2[7] , \nOut7_2[6] , 
        \nOut7_2[5] , \nOut7_2[4] , \nOut7_2[3] , \nOut7_2[2] , \nOut7_2[1] , 
        \nOut7_2[0] }), .WestIn({\nOut5_2[7] , \nOut5_2[6] , \nOut5_2[5] , 
        \nOut5_2[4] , \nOut5_2[3] , \nOut5_2[2] , \nOut5_2[1] , \nOut5_2[0] }), 
        .Out({\nOut6_2[7] , \nOut6_2[6] , \nOut6_2[5] , \nOut6_2[4] , 
        \nOut6_2[3] , \nOut6_2[2] , \nOut6_2[1] , \nOut6_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_785 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut786[7] , \nScanOut786[6] , 
        \nScanOut786[5] , \nScanOut786[4] , \nScanOut786[3] , \nScanOut786[2] , 
        \nScanOut786[1] , \nScanOut786[0] }), .ScanOut({\nScanOut785[7] , 
        \nScanOut785[6] , \nScanOut785[5] , \nScanOut785[4] , \nScanOut785[3] , 
        \nScanOut785[2] , \nScanOut785[1] , \nScanOut785[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_16[7] , \nOut24_16[6] , \nOut24_16[5] , \nOut24_16[4] , 
        \nOut24_16[3] , \nOut24_16[2] , \nOut24_16[1] , \nOut24_16[0] }), 
        .SouthIn({\nOut24_18[7] , \nOut24_18[6] , \nOut24_18[5] , 
        \nOut24_18[4] , \nOut24_18[3] , \nOut24_18[2] , \nOut24_18[1] , 
        \nOut24_18[0] }), .EastIn({\nOut25_17[7] , \nOut25_17[6] , 
        \nOut25_17[5] , \nOut25_17[4] , \nOut25_17[3] , \nOut25_17[2] , 
        \nOut25_17[1] , \nOut25_17[0] }), .WestIn({\nOut23_17[7] , 
        \nOut23_17[6] , \nOut23_17[5] , \nOut23_17[4] , \nOut23_17[3] , 
        \nOut23_17[2] , \nOut23_17[1] , \nOut23_17[0] }), .Out({\nOut24_17[7] , 
        \nOut24_17[6] , \nOut24_17[5] , \nOut24_17[4] , \nOut24_17[3] , 
        \nOut24_17[2] , \nOut24_17[1] , \nOut24_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_939 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut940[7] , \nScanOut940[6] , 
        \nScanOut940[5] , \nScanOut940[4] , \nScanOut940[3] , \nScanOut940[2] , 
        \nScanOut940[1] , \nScanOut940[0] }), .ScanOut({\nScanOut939[7] , 
        \nScanOut939[6] , \nScanOut939[5] , \nScanOut939[4] , \nScanOut939[3] , 
        \nScanOut939[2] , \nScanOut939[1] , \nScanOut939[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_10[7] , \nOut29_10[6] , \nOut29_10[5] , \nOut29_10[4] , 
        \nOut29_10[3] , \nOut29_10[2] , \nOut29_10[1] , \nOut29_10[0] }), 
        .SouthIn({\nOut29_12[7] , \nOut29_12[6] , \nOut29_12[5] , 
        \nOut29_12[4] , \nOut29_12[3] , \nOut29_12[2] , \nOut29_12[1] , 
        \nOut29_12[0] }), .EastIn({\nOut30_11[7] , \nOut30_11[6] , 
        \nOut30_11[5] , \nOut30_11[4] , \nOut30_11[3] , \nOut30_11[2] , 
        \nOut30_11[1] , \nOut30_11[0] }), .WestIn({\nOut28_11[7] , 
        \nOut28_11[6] , \nOut28_11[5] , \nOut28_11[4] , \nOut28_11[3] , 
        \nOut28_11[2] , \nOut28_11[1] , \nOut28_11[0] }), .Out({\nOut29_11[7] , 
        \nOut29_11[6] , \nOut29_11[5] , \nOut29_11[4] , \nOut29_11[3] , 
        \nOut29_11[2] , \nOut29_11[1] , \nOut29_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_283 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut284[7] , \nScanOut284[6] , 
        \nScanOut284[5] , \nScanOut284[4] , \nScanOut284[3] , \nScanOut284[2] , 
        \nScanOut284[1] , \nScanOut284[0] }), .ScanOut({\nScanOut283[7] , 
        \nScanOut283[6] , \nScanOut283[5] , \nScanOut283[4] , \nScanOut283[3] , 
        \nScanOut283[2] , \nScanOut283[1] , \nScanOut283[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_26[7] , \nOut8_26[6] , \nOut8_26[5] , \nOut8_26[4] , 
        \nOut8_26[3] , \nOut8_26[2] , \nOut8_26[1] , \nOut8_26[0] }), 
        .SouthIn({\nOut8_28[7] , \nOut8_28[6] , \nOut8_28[5] , \nOut8_28[4] , 
        \nOut8_28[3] , \nOut8_28[2] , \nOut8_28[1] , \nOut8_28[0] }), .EastIn(
        {\nOut9_27[7] , \nOut9_27[6] , \nOut9_27[5] , \nOut9_27[4] , 
        \nOut9_27[3] , \nOut9_27[2] , \nOut9_27[1] , \nOut9_27[0] }), .WestIn(
        {\nOut7_27[7] , \nOut7_27[6] , \nOut7_27[5] , \nOut7_27[4] , 
        \nOut7_27[3] , \nOut7_27[2] , \nOut7_27[1] , \nOut7_27[0] }), .Out({
        \nOut8_27[7] , \nOut8_27[6] , \nOut8_27[5] , \nOut8_27[4] , 
        \nOut8_27[3] , \nOut8_27[2] , \nOut8_27[1] , \nOut8_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_334 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut335[7] , \nScanOut335[6] , 
        \nScanOut335[5] , \nScanOut335[4] , \nScanOut335[3] , \nScanOut335[2] , 
        \nScanOut335[1] , \nScanOut335[0] }), .ScanOut({\nScanOut334[7] , 
        \nScanOut334[6] , \nScanOut334[5] , \nScanOut334[4] , \nScanOut334[3] , 
        \nScanOut334[2] , \nScanOut334[1] , \nScanOut334[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_13[7] , \nOut10_13[6] , \nOut10_13[5] , \nOut10_13[4] , 
        \nOut10_13[3] , \nOut10_13[2] , \nOut10_13[1] , \nOut10_13[0] }), 
        .SouthIn({\nOut10_15[7] , \nOut10_15[6] , \nOut10_15[5] , 
        \nOut10_15[4] , \nOut10_15[3] , \nOut10_15[2] , \nOut10_15[1] , 
        \nOut10_15[0] }), .EastIn({\nOut11_14[7] , \nOut11_14[6] , 
        \nOut11_14[5] , \nOut11_14[4] , \nOut11_14[3] , \nOut11_14[2] , 
        \nOut11_14[1] , \nOut11_14[0] }), .WestIn({\nOut9_14[7] , 
        \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , \nOut9_14[3] , 
        \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }), .Out({\nOut10_14[7] , 
        \nOut10_14[6] , \nOut10_14[5] , \nOut10_14[4] , \nOut10_14[3] , 
        \nOut10_14[2] , \nOut10_14[1] , \nOut10_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_615 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut616[7] , \nScanOut616[6] , 
        \nScanOut616[5] , \nScanOut616[4] , \nScanOut616[3] , \nScanOut616[2] , 
        \nScanOut616[1] , \nScanOut616[0] }), .ScanOut({\nScanOut615[7] , 
        \nScanOut615[6] , \nScanOut615[5] , \nScanOut615[4] , \nScanOut615[3] , 
        \nScanOut615[2] , \nScanOut615[1] , \nScanOut615[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_6[7] , \nOut19_6[6] , \nOut19_6[5] , \nOut19_6[4] , 
        \nOut19_6[3] , \nOut19_6[2] , \nOut19_6[1] , \nOut19_6[0] }), 
        .SouthIn({\nOut19_8[7] , \nOut19_8[6] , \nOut19_8[5] , \nOut19_8[4] , 
        \nOut19_8[3] , \nOut19_8[2] , \nOut19_8[1] , \nOut19_8[0] }), .EastIn(
        {\nOut20_7[7] , \nOut20_7[6] , \nOut20_7[5] , \nOut20_7[4] , 
        \nOut20_7[3] , \nOut20_7[2] , \nOut20_7[1] , \nOut20_7[0] }), .WestIn(
        {\nOut18_7[7] , \nOut18_7[6] , \nOut18_7[5] , \nOut18_7[4] , 
        \nOut18_7[3] , \nOut18_7[2] , \nOut18_7[1] , \nOut18_7[0] }), .Out({
        \nOut19_7[7] , \nOut19_7[6] , \nOut19_7[5] , \nOut19_7[4] , 
        \nOut19_7[3] , \nOut19_7[2] , \nOut19_7[1] , \nOut19_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_957 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut958[7] , \nScanOut958[6] , 
        \nScanOut958[5] , \nScanOut958[4] , \nScanOut958[3] , \nScanOut958[2] , 
        \nScanOut958[1] , \nScanOut958[0] }), .ScanOut({\nScanOut957[7] , 
        \nScanOut957[6] , \nScanOut957[5] , \nScanOut957[4] , \nScanOut957[3] , 
        \nScanOut957[2] , \nScanOut957[1] , \nScanOut957[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_28[7] , \nOut29_28[6] , \nOut29_28[5] , \nOut29_28[4] , 
        \nOut29_28[3] , \nOut29_28[2] , \nOut29_28[1] , \nOut29_28[0] }), 
        .SouthIn({\nOut29_30[7] , \nOut29_30[6] , \nOut29_30[5] , 
        \nOut29_30[4] , \nOut29_30[3] , \nOut29_30[2] , \nOut29_30[1] , 
        \nOut29_30[0] }), .EastIn({\nOut30_29[7] , \nOut30_29[6] , 
        \nOut30_29[5] , \nOut30_29[4] , \nOut30_29[3] , \nOut30_29[2] , 
        \nOut30_29[1] , \nOut30_29[0] }), .WestIn({\nOut28_29[7] , 
        \nOut28_29[6] , \nOut28_29[5] , \nOut28_29[4] , \nOut28_29[3] , 
        \nOut28_29[2] , \nOut28_29[1] , \nOut28_29[0] }), .Out({\nOut29_29[7] , 
        \nOut29_29[6] , \nOut29_29[5] , \nOut29_29[4] , \nOut29_29[3] , 
        \nOut29_29[2] , \nOut29_29[1] , \nOut29_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_502 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut503[7] , \nScanOut503[6] , 
        \nScanOut503[5] , \nScanOut503[4] , \nScanOut503[3] , \nScanOut503[2] , 
        \nScanOut503[1] , \nScanOut503[0] }), .ScanOut({\nScanOut502[7] , 
        \nScanOut502[6] , \nScanOut502[5] , \nScanOut502[4] , \nScanOut502[3] , 
        \nScanOut502[2] , \nScanOut502[1] , \nScanOut502[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_21[7] , \nOut15_21[6] , \nOut15_21[5] , \nOut15_21[4] , 
        \nOut15_21[3] , \nOut15_21[2] , \nOut15_21[1] , \nOut15_21[0] }), 
        .SouthIn({\nOut15_23[7] , \nOut15_23[6] , \nOut15_23[5] , 
        \nOut15_23[4] , \nOut15_23[3] , \nOut15_23[2] , \nOut15_23[1] , 
        \nOut15_23[0] }), .EastIn({\nOut16_22[7] , \nOut16_22[6] , 
        \nOut16_22[5] , \nOut16_22[4] , \nOut16_22[3] , \nOut16_22[2] , 
        \nOut16_22[1] , \nOut16_22[0] }), .WestIn({\nOut14_22[7] , 
        \nOut14_22[6] , \nOut14_22[5] , \nOut14_22[4] , \nOut14_22[3] , 
        \nOut14_22[2] , \nOut14_22[1] , \nOut14_22[0] }), .Out({\nOut15_22[7] , 
        \nOut15_22[6] , \nOut15_22[5] , \nOut15_22[4] , \nOut15_22[3] , 
        \nOut15_22[2] , \nOut15_22[1] , \nOut15_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_525 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut526[7] , \nScanOut526[6] , 
        \nScanOut526[5] , \nScanOut526[4] , \nScanOut526[3] , \nScanOut526[2] , 
        \nScanOut526[1] , \nScanOut526[0] }), .ScanOut({\nScanOut525[7] , 
        \nScanOut525[6] , \nScanOut525[5] , \nScanOut525[4] , \nScanOut525[3] , 
        \nScanOut525[2] , \nScanOut525[1] , \nScanOut525[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_12[7] , \nOut16_12[6] , \nOut16_12[5] , \nOut16_12[4] , 
        \nOut16_12[3] , \nOut16_12[2] , \nOut16_12[1] , \nOut16_12[0] }), 
        .SouthIn({\nOut16_14[7] , \nOut16_14[6] , \nOut16_14[5] , 
        \nOut16_14[4] , \nOut16_14[3] , \nOut16_14[2] , \nOut16_14[1] , 
        \nOut16_14[0] }), .EastIn({\nOut17_13[7] , \nOut17_13[6] , 
        \nOut17_13[5] , \nOut17_13[4] , \nOut17_13[3] , \nOut17_13[2] , 
        \nOut17_13[1] , \nOut17_13[0] }), .WestIn({\nOut15_13[7] , 
        \nOut15_13[6] , \nOut15_13[5] , \nOut15_13[4] , \nOut15_13[3] , 
        \nOut15_13[2] , \nOut15_13[1] , \nOut15_13[0] }), .Out({\nOut16_13[7] , 
        \nOut16_13[6] , \nOut16_13[5] , \nOut16_13[4] , \nOut16_13[3] , 
        \nOut16_13[2] , \nOut16_13[1] , \nOut16_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_970 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut971[7] , \nScanOut971[6] , 
        \nScanOut971[5] , \nScanOut971[4] , \nScanOut971[3] , \nScanOut971[2] , 
        \nScanOut971[1] , \nScanOut971[0] }), .ScanOut({\nScanOut970[7] , 
        \nScanOut970[6] , \nScanOut970[5] , \nScanOut970[4] , \nScanOut970[3] , 
        \nScanOut970[2] , \nScanOut970[1] , \nScanOut970[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_9[7] , \nOut30_9[6] , \nOut30_9[5] , \nOut30_9[4] , 
        \nOut30_9[3] , \nOut30_9[2] , \nOut30_9[1] , \nOut30_9[0] }), 
        .SouthIn({\nOut30_11[7] , \nOut30_11[6] , \nOut30_11[5] , 
        \nOut30_11[4] , \nOut30_11[3] , \nOut30_11[2] , \nOut30_11[1] , 
        \nOut30_11[0] }), .EastIn({\nOut31_10[7] , \nOut31_10[6] , 
        \nOut31_10[5] , \nOut31_10[4] , \nOut31_10[3] , \nOut31_10[2] , 
        \nOut31_10[1] , \nOut31_10[0] }), .WestIn({\nOut29_10[7] , 
        \nOut29_10[6] , \nOut29_10[5] , \nOut29_10[4] , \nOut29_10[3] , 
        \nOut29_10[2] , \nOut29_10[1] , \nOut29_10[0] }), .Out({\nOut30_10[7] , 
        \nOut30_10[6] , \nOut30_10[5] , \nOut30_10[4] , \nOut30_10[3] , 
        \nOut30_10[2] , \nOut30_10[1] , \nOut30_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_313 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut314[7] , \nScanOut314[6] , 
        \nScanOut314[5] , \nScanOut314[4] , \nScanOut314[3] , \nScanOut314[2] , 
        \nScanOut314[1] , \nScanOut314[0] }), .ScanOut({\nScanOut313[7] , 
        \nScanOut313[6] , \nScanOut313[5] , \nScanOut313[4] , \nScanOut313[3] , 
        \nScanOut313[2] , \nScanOut313[1] , \nScanOut313[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_24[7] , \nOut9_24[6] , \nOut9_24[5] , \nOut9_24[4] , 
        \nOut9_24[3] , \nOut9_24[2] , \nOut9_24[1] , \nOut9_24[0] }), 
        .SouthIn({\nOut9_26[7] , \nOut9_26[6] , \nOut9_26[5] , \nOut9_26[4] , 
        \nOut9_26[3] , \nOut9_26[2] , \nOut9_26[1] , \nOut9_26[0] }), .EastIn(
        {\nOut10_25[7] , \nOut10_25[6] , \nOut10_25[5] , \nOut10_25[4] , 
        \nOut10_25[3] , \nOut10_25[2] , \nOut10_25[1] , \nOut10_25[0] }), 
        .WestIn({\nOut8_25[7] , \nOut8_25[6] , \nOut8_25[5] , \nOut8_25[4] , 
        \nOut8_25[3] , \nOut8_25[2] , \nOut8_25[1] , \nOut8_25[0] }), .Out({
        \nOut9_25[7] , \nOut9_25[6] , \nOut9_25[5] , \nOut9_25[4] , 
        \nOut9_25[3] , \nOut9_25[2] , \nOut9_25[1] , \nOut9_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_492 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut493[7] , \nScanOut493[6] , 
        \nScanOut493[5] , \nScanOut493[4] , \nScanOut493[3] , \nScanOut493[2] , 
        \nScanOut493[1] , \nScanOut493[0] }), .ScanOut({\nScanOut492[7] , 
        \nScanOut492[6] , \nScanOut492[5] , \nScanOut492[4] , \nScanOut492[3] , 
        \nScanOut492[2] , \nScanOut492[1] , \nScanOut492[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_11[7] , \nOut15_11[6] , \nOut15_11[5] , \nOut15_11[4] , 
        \nOut15_11[3] , \nOut15_11[2] , \nOut15_11[1] , \nOut15_11[0] }), 
        .SouthIn({\nOut15_13[7] , \nOut15_13[6] , \nOut15_13[5] , 
        \nOut15_13[4] , \nOut15_13[3] , \nOut15_13[2] , \nOut15_13[1] , 
        \nOut15_13[0] }), .EastIn({\nOut16_12[7] , \nOut16_12[6] , 
        \nOut16_12[5] , \nOut16_12[4] , \nOut16_12[3] , \nOut16_12[2] , 
        \nOut16_12[1] , \nOut16_12[0] }), .WestIn({\nOut14_12[7] , 
        \nOut14_12[6] , \nOut14_12[5] , \nOut14_12[4] , \nOut14_12[3] , 
        \nOut14_12[2] , \nOut14_12[1] , \nOut14_12[0] }), .Out({\nOut15_12[7] , 
        \nOut15_12[6] , \nOut15_12[5] , \nOut15_12[4] , \nOut15_12[3] , 
        \nOut15_12[2] , \nOut15_12[1] , \nOut15_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_632 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut633[7] , \nScanOut633[6] , 
        \nScanOut633[5] , \nScanOut633[4] , \nScanOut633[3] , \nScanOut633[2] , 
        \nScanOut633[1] , \nScanOut633[0] }), .ScanOut({\nScanOut632[7] , 
        \nScanOut632[6] , \nScanOut632[5] , \nScanOut632[4] , \nScanOut632[3] , 
        \nScanOut632[2] , \nScanOut632[1] , \nScanOut632[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_23[7] , \nOut19_23[6] , \nOut19_23[5] , \nOut19_23[4] , 
        \nOut19_23[3] , \nOut19_23[2] , \nOut19_23[1] , \nOut19_23[0] }), 
        .SouthIn({\nOut19_25[7] , \nOut19_25[6] , \nOut19_25[5] , 
        \nOut19_25[4] , \nOut19_25[3] , \nOut19_25[2] , \nOut19_25[1] , 
        \nOut19_25[0] }), .EastIn({\nOut20_24[7] , \nOut20_24[6] , 
        \nOut20_24[5] , \nOut20_24[4] , \nOut20_24[3] , \nOut20_24[2] , 
        \nOut20_24[1] , \nOut20_24[0] }), .WestIn({\nOut18_24[7] , 
        \nOut18_24[6] , \nOut18_24[5] , \nOut18_24[4] , \nOut18_24[3] , 
        \nOut18_24[2] , \nOut18_24[1] , \nOut18_24[0] }), .Out({\nOut19_24[7] , 
        \nOut19_24[6] , \nOut19_24[5] , \nOut19_24[4] , \nOut19_24[3] , 
        \nOut19_24[2] , \nOut19_24[1] , \nOut19_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_99 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut100[7] , \nScanOut100[6] , 
        \nScanOut100[5] , \nScanOut100[4] , \nScanOut100[3] , \nScanOut100[2] , 
        \nScanOut100[1] , \nScanOut100[0] }), .ScanOut({\nScanOut99[7] , 
        \nScanOut99[6] , \nScanOut99[5] , \nScanOut99[4] , \nScanOut99[3] , 
        \nScanOut99[2] , \nScanOut99[1] , \nScanOut99[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_2[7] , \nOut3_2[6] , \nOut3_2[5] , \nOut3_2[4] , \nOut3_2[3] , 
        \nOut3_2[2] , \nOut3_2[1] , \nOut3_2[0] }), .SouthIn({\nOut3_4[7] , 
        \nOut3_4[6] , \nOut3_4[5] , \nOut3_4[4] , \nOut3_4[3] , \nOut3_4[2] , 
        \nOut3_4[1] , \nOut3_4[0] }), .EastIn({\nOut4_3[7] , \nOut4_3[6] , 
        \nOut4_3[5] , \nOut4_3[4] , \nOut4_3[3] , \nOut4_3[2] , \nOut4_3[1] , 
        \nOut4_3[0] }), .WestIn({\nOut2_3[7] , \nOut2_3[6] , \nOut2_3[5] , 
        \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , \nOut2_3[0] }), 
        .Out({\nOut3_3[7] , \nOut3_3[6] , \nOut3_3[5] , \nOut3_3[4] , 
        \nOut3_3[3] , \nOut3_3[2] , \nOut3_3[1] , \nOut3_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_138 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut139[7] , \nScanOut139[6] , 
        \nScanOut139[5] , \nScanOut139[4] , \nScanOut139[3] , \nScanOut139[2] , 
        \nScanOut139[1] , \nScanOut139[0] }), .ScanOut({\nScanOut138[7] , 
        \nScanOut138[6] , \nScanOut138[5] , \nScanOut138[4] , \nScanOut138[3] , 
        \nScanOut138[2] , \nScanOut138[1] , \nScanOut138[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_9[7] , \nOut4_9[6] , \nOut4_9[5] , \nOut4_9[4] , \nOut4_9[3] , 
        \nOut4_9[2] , \nOut4_9[1] , \nOut4_9[0] }), .SouthIn({\nOut4_11[7] , 
        \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , \nOut4_11[3] , 
        \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }), .EastIn({\nOut5_10[7] , 
        \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , \nOut5_10[3] , 
        \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }), .WestIn({\nOut3_10[7] , 
        \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , \nOut3_10[3] , 
        \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }), .Out({\nOut4_10[7] , 
        \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , \nOut4_10[3] , 
        \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_208 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut209[7] , \nScanOut209[6] , 
        \nScanOut209[5] , \nScanOut209[4] , \nScanOut209[3] , \nScanOut209[2] , 
        \nScanOut209[1] , \nScanOut209[0] }), .ScanOut({\nScanOut208[7] , 
        \nScanOut208[6] , \nScanOut208[5] , \nScanOut208[4] , \nScanOut208[3] , 
        \nScanOut208[2] , \nScanOut208[1] , \nScanOut208[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_15[7] , \nOut6_15[6] , \nOut6_15[5] , \nOut6_15[4] , 
        \nOut6_15[3] , \nOut6_15[2] , \nOut6_15[1] , \nOut6_15[0] }), 
        .SouthIn({\nOut6_17[7] , \nOut6_17[6] , \nOut6_17[5] , \nOut6_17[4] , 
        \nOut6_17[3] , \nOut6_17[2] , \nOut6_17[1] , \nOut6_17[0] }), .EastIn(
        {\nOut7_16[7] , \nOut7_16[6] , \nOut7_16[5] , \nOut7_16[4] , 
        \nOut7_16[3] , \nOut7_16[2] , \nOut7_16[1] , \nOut7_16[0] }), .WestIn(
        {\nOut5_16[7] , \nOut5_16[6] , \nOut5_16[5] , \nOut5_16[4] , 
        \nOut5_16[3] , \nOut5_16[2] , \nOut5_16[1] , \nOut5_16[0] }), .Out({
        \nOut6_16[7] , \nOut6_16[6] , \nOut6_16[5] , \nOut6_16[4] , 
        \nOut6_16[3] , \nOut6_16[2] , \nOut6_16[1] , \nOut6_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_589 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut590[7] , \nScanOut590[6] , 
        \nScanOut590[5] , \nScanOut590[4] , \nScanOut590[3] , \nScanOut590[2] , 
        \nScanOut590[1] , \nScanOut590[0] }), .ScanOut({\nScanOut589[7] , 
        \nScanOut589[6] , \nScanOut589[5] , \nScanOut589[4] , \nScanOut589[3] , 
        \nScanOut589[2] , \nScanOut589[1] , \nScanOut589[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_12[7] , \nOut18_12[6] , \nOut18_12[5] , \nOut18_12[4] , 
        \nOut18_12[3] , \nOut18_12[2] , \nOut18_12[1] , \nOut18_12[0] }), 
        .SouthIn({\nOut18_14[7] , \nOut18_14[6] , \nOut18_14[5] , 
        \nOut18_14[4] , \nOut18_14[3] , \nOut18_14[2] , \nOut18_14[1] , 
        \nOut18_14[0] }), .EastIn({\nOut19_13[7] , \nOut19_13[6] , 
        \nOut19_13[5] , \nOut19_13[4] , \nOut19_13[3] , \nOut19_13[2] , 
        \nOut19_13[1] , \nOut19_13[0] }), .WestIn({\nOut17_13[7] , 
        \nOut17_13[6] , \nOut17_13[5] , \nOut17_13[4] , \nOut17_13[3] , 
        \nOut17_13[2] , \nOut17_13[1] , \nOut17_13[0] }), .Out({\nOut18_13[7] , 
        \nOut18_13[6] , \nOut18_13[5] , \nOut18_13[4] , \nOut18_13[3] , 
        \nOut18_13[2] , \nOut18_13[1] , \nOut18_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1008 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1009[7] , \nScanOut1009[6] , 
        \nScanOut1009[5] , \nScanOut1009[4] , \nScanOut1009[3] , 
        \nScanOut1009[2] , \nScanOut1009[1] , \nScanOut1009[0] }), .ScanOut({
        \nScanOut1008[7] , \nScanOut1008[6] , \nScanOut1008[5] , 
        \nScanOut1008[4] , \nScanOut1008[3] , \nScanOut1008[2] , 
        \nScanOut1008[1] , \nScanOut1008[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_16[7] , \nOut31_16[6] , \nOut31_16[5] , 
        \nOut31_16[4] , \nOut31_16[3] , \nOut31_16[2] , \nOut31_16[1] , 
        \nOut31_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_398 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut399[7] , \nScanOut399[6] , 
        \nScanOut399[5] , \nScanOut399[4] , \nScanOut399[3] , \nScanOut399[2] , 
        \nScanOut399[1] , \nScanOut399[0] }), .ScanOut({\nScanOut398[7] , 
        \nScanOut398[6] , \nScanOut398[5] , \nScanOut398[4] , \nScanOut398[3] , 
        \nScanOut398[2] , \nScanOut398[1] , \nScanOut398[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_13[7] , \nOut12_13[6] , \nOut12_13[5] , \nOut12_13[4] , 
        \nOut12_13[3] , \nOut12_13[2] , \nOut12_13[1] , \nOut12_13[0] }), 
        .SouthIn({\nOut12_15[7] , \nOut12_15[6] , \nOut12_15[5] , 
        \nOut12_15[4] , \nOut12_15[3] , \nOut12_15[2] , \nOut12_15[1] , 
        \nOut12_15[0] }), .EastIn({\nOut13_14[7] , \nOut13_14[6] , 
        \nOut13_14[5] , \nOut13_14[4] , \nOut13_14[3] , \nOut13_14[2] , 
        \nOut13_14[1] , \nOut13_14[0] }), .WestIn({\nOut11_14[7] , 
        \nOut11_14[6] , \nOut11_14[5] , \nOut11_14[4] , \nOut11_14[3] , 
        \nOut11_14[2] , \nOut11_14[1] , \nOut11_14[0] }), .Out({\nOut12_14[7] , 
        \nOut12_14[6] , \nOut12_14[5] , \nOut12_14[4] , \nOut12_14[3] , 
        \nOut12_14[2] , \nOut12_14[1] , \nOut12_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_419 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut420[7] , \nScanOut420[6] , 
        \nScanOut420[5] , \nScanOut420[4] , \nScanOut420[3] , \nScanOut420[2] , 
        \nScanOut420[1] , \nScanOut420[0] }), .ScanOut({\nScanOut419[7] , 
        \nScanOut419[6] , \nScanOut419[5] , \nScanOut419[4] , \nScanOut419[3] , 
        \nScanOut419[2] , \nScanOut419[1] , \nScanOut419[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }), 
        .SouthIn({\nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }), .EastIn(
        {\nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }), .WestIn(
        {\nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }), .Out({
        \nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_729 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut730[7] , \nScanOut730[6] , 
        \nScanOut730[5] , \nScanOut730[4] , \nScanOut730[3] , \nScanOut730[2] , 
        \nScanOut730[1] , \nScanOut730[0] }), .ScanOut({\nScanOut729[7] , 
        \nScanOut729[6] , \nScanOut729[5] , \nScanOut729[4] , \nScanOut729[3] , 
        \nScanOut729[2] , \nScanOut729[1] , \nScanOut729[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_24[7] , \nOut22_24[6] , \nOut22_24[5] , \nOut22_24[4] , 
        \nOut22_24[3] , \nOut22_24[2] , \nOut22_24[1] , \nOut22_24[0] }), 
        .SouthIn({\nOut22_26[7] , \nOut22_26[6] , \nOut22_26[5] , 
        \nOut22_26[4] , \nOut22_26[3] , \nOut22_26[2] , \nOut22_26[1] , 
        \nOut22_26[0] }), .EastIn({\nOut23_25[7] , \nOut23_25[6] , 
        \nOut23_25[5] , \nOut23_25[4] , \nOut23_25[3] , \nOut23_25[2] , 
        \nOut23_25[1] , \nOut23_25[0] }), .WestIn({\nOut21_25[7] , 
        \nOut21_25[6] , \nOut21_25[5] , \nOut21_25[4] , \nOut21_25[3] , 
        \nOut21_25[2] , \nOut21_25[1] , \nOut21_25[0] }), .Out({\nOut22_25[7] , 
        \nOut22_25[6] , \nOut22_25[5] , \nOut22_25[4] , \nOut22_25[3] , 
        \nOut22_25[2] , \nOut22_25[1] , \nOut22_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_186 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut187[7] , \nScanOut187[6] , 
        \nScanOut187[5] , \nScanOut187[4] , \nScanOut187[3] , \nScanOut187[2] , 
        \nScanOut187[1] , \nScanOut187[0] }), .ScanOut({\nScanOut186[7] , 
        \nScanOut186[6] , \nScanOut186[5] , \nScanOut186[4] , \nScanOut186[3] , 
        \nScanOut186[2] , \nScanOut186[1] , \nScanOut186[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_25[7] , \nOut5_25[6] , \nOut5_25[5] , \nOut5_25[4] , 
        \nOut5_25[3] , \nOut5_25[2] , \nOut5_25[1] , \nOut5_25[0] }), 
        .SouthIn({\nOut5_27[7] , \nOut5_27[6] , \nOut5_27[5] , \nOut5_27[4] , 
        \nOut5_27[3] , \nOut5_27[2] , \nOut5_27[1] , \nOut5_27[0] }), .EastIn(
        {\nOut6_26[7] , \nOut6_26[6] , \nOut6_26[5] , \nOut6_26[4] , 
        \nOut6_26[3] , \nOut6_26[2] , \nOut6_26[1] , \nOut6_26[0] }), .WestIn(
        {\nOut4_26[7] , \nOut4_26[6] , \nOut4_26[5] , \nOut4_26[4] , 
        \nOut4_26[3] , \nOut4_26[2] , \nOut4_26[1] , \nOut4_26[0] }), .Out({
        \nOut5_26[7] , \nOut5_26[6] , \nOut5_26[5] , \nOut5_26[4] , 
        \nOut5_26[3] , \nOut5_26[2] , \nOut5_26[1] , \nOut5_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_879 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut880[7] , \nScanOut880[6] , 
        \nScanOut880[5] , \nScanOut880[4] , \nScanOut880[3] , \nScanOut880[2] , 
        \nScanOut880[1] , \nScanOut880[0] }), .ScanOut({\nScanOut879[7] , 
        \nScanOut879[6] , \nScanOut879[5] , \nScanOut879[4] , \nScanOut879[3] , 
        \nScanOut879[2] , \nScanOut879[1] , \nScanOut879[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_14[7] , \nOut27_14[6] , \nOut27_14[5] , \nOut27_14[4] , 
        \nOut27_14[3] , \nOut27_14[2] , \nOut27_14[1] , \nOut27_14[0] }), 
        .SouthIn({\nOut27_16[7] , \nOut27_16[6] , \nOut27_16[5] , 
        \nOut27_16[4] , \nOut27_16[3] , \nOut27_16[2] , \nOut27_16[1] , 
        \nOut27_16[0] }), .EastIn({\nOut28_15[7] , \nOut28_15[6] , 
        \nOut28_15[5] , \nOut28_15[4] , \nOut28_15[3] , \nOut28_15[2] , 
        \nOut28_15[1] , \nOut28_15[0] }), .WestIn({\nOut26_15[7] , 
        \nOut26_15[6] , \nOut26_15[5] , \nOut26_15[4] , \nOut26_15[3] , 
        \nOut26_15[2] , \nOut26_15[1] , \nOut26_15[0] }), .Out({\nOut27_15[7] , 
        \nOut27_15[6] , \nOut27_15[5] , \nOut27_15[4] , \nOut27_15[3] , 
        \nOut27_15[2] , \nOut27_15[1] , \nOut27_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_607 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut608[7] , \nScanOut608[6] , 
        \nScanOut608[5] , \nScanOut608[4] , \nScanOut608[3] , \nScanOut608[2] , 
        \nScanOut608[1] , \nScanOut608[0] }), .ScanOut({\nScanOut607[7] , 
        \nScanOut607[6] , \nScanOut607[5] , \nScanOut607[4] , \nScanOut607[3] , 
        \nScanOut607[2] , \nScanOut607[1] , \nScanOut607[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut18_31[7] , \nOut18_31[6] , 
        \nOut18_31[5] , \nOut18_31[4] , \nOut18_31[3] , \nOut18_31[2] , 
        \nOut18_31[1] , \nOut18_31[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_797 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut798[7] , \nScanOut798[6] , 
        \nScanOut798[5] , \nScanOut798[4] , \nScanOut798[3] , \nScanOut798[2] , 
        \nScanOut798[1] , \nScanOut798[0] }), .ScanOut({\nScanOut797[7] , 
        \nScanOut797[6] , \nScanOut797[5] , \nScanOut797[4] , \nScanOut797[3] , 
        \nScanOut797[2] , \nScanOut797[1] , \nScanOut797[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_28[7] , \nOut24_28[6] , \nOut24_28[5] , \nOut24_28[4] , 
        \nOut24_28[3] , \nOut24_28[2] , \nOut24_28[1] , \nOut24_28[0] }), 
        .SouthIn({\nOut24_30[7] , \nOut24_30[6] , \nOut24_30[5] , 
        \nOut24_30[4] , \nOut24_30[3] , \nOut24_30[2] , \nOut24_30[1] , 
        \nOut24_30[0] }), .EastIn({\nOut25_29[7] , \nOut25_29[6] , 
        \nOut25_29[5] , \nOut25_29[4] , \nOut25_29[3] , \nOut25_29[2] , 
        \nOut25_29[1] , \nOut25_29[0] }), .WestIn({\nOut23_29[7] , 
        \nOut23_29[6] , \nOut23_29[5] , \nOut23_29[4] , \nOut23_29[3] , 
        \nOut23_29[2] , \nOut23_29[1] , \nOut23_29[0] }), .Out({\nOut24_29[7] , 
        \nOut24_29[6] , \nOut24_29[5] , \nOut24_29[4] , \nOut24_29[3] , 
        \nOut24_29[2] , \nOut24_29[1] , \nOut24_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_35 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut36[7] , \nScanOut36[6] , 
        \nScanOut36[5] , \nScanOut36[4] , \nScanOut36[3] , \nScanOut36[2] , 
        \nScanOut36[1] , \nScanOut36[0] }), .ScanOut({\nScanOut35[7] , 
        \nScanOut35[6] , \nScanOut35[5] , \nScanOut35[4] , \nScanOut35[3] , 
        \nScanOut35[2] , \nScanOut35[1] , \nScanOut35[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , \nOut1_2[3] , 
        \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), .SouthIn({\nOut1_4[7] , 
        \nOut1_4[6] , \nOut1_4[5] , \nOut1_4[4] , \nOut1_4[3] , \nOut1_4[2] , 
        \nOut1_4[1] , \nOut1_4[0] }), .EastIn({\nOut2_3[7] , \nOut2_3[6] , 
        \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , 
        \nOut2_3[0] }), .WestIn({\nOut0_3[7] , \nOut0_3[6] , \nOut0_3[5] , 
        \nOut0_3[4] , \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , \nOut0_3[0] }), 
        .Out({\nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , 
        \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_291 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut292[7] , \nScanOut292[6] , 
        \nScanOut292[5] , \nScanOut292[4] , \nScanOut292[3] , \nScanOut292[2] , 
        \nScanOut292[1] , \nScanOut292[0] }), .ScanOut({\nScanOut291[7] , 
        \nScanOut291[6] , \nScanOut291[5] , \nScanOut291[4] , \nScanOut291[3] , 
        \nScanOut291[2] , \nScanOut291[1] , \nScanOut291[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_2[7] , \nOut9_2[6] , \nOut9_2[5] , \nOut9_2[4] , \nOut9_2[3] , 
        \nOut9_2[2] , \nOut9_2[1] , \nOut9_2[0] }), .SouthIn({\nOut9_4[7] , 
        \nOut9_4[6] , \nOut9_4[5] , \nOut9_4[4] , \nOut9_4[3] , \nOut9_4[2] , 
        \nOut9_4[1] , \nOut9_4[0] }), .EastIn({\nOut10_3[7] , \nOut10_3[6] , 
        \nOut10_3[5] , \nOut10_3[4] , \nOut10_3[3] , \nOut10_3[2] , 
        \nOut10_3[1] , \nOut10_3[0] }), .WestIn({\nOut8_3[7] , \nOut8_3[6] , 
        \nOut8_3[5] , \nOut8_3[4] , \nOut8_3[3] , \nOut8_3[2] , \nOut8_3[1] , 
        \nOut8_3[0] }), .Out({\nOut9_3[7] , \nOut9_3[6] , \nOut9_3[5] , 
        \nOut9_3[4] , \nOut9_3[3] , \nOut9_3[2] , \nOut9_3[1] , \nOut9_3[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_301 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut302[7] , \nScanOut302[6] , 
        \nScanOut302[5] , \nScanOut302[4] , \nScanOut302[3] , \nScanOut302[2] , 
        \nScanOut302[1] , \nScanOut302[0] }), .ScanOut({\nScanOut301[7] , 
        \nScanOut301[6] , \nScanOut301[5] , \nScanOut301[4] , \nScanOut301[3] , 
        \nScanOut301[2] , \nScanOut301[1] , \nScanOut301[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_12[7] , \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , 
        \nOut9_12[3] , \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }), 
        .SouthIn({\nOut9_14[7] , \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , 
        \nOut9_14[3] , \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }), .EastIn(
        {\nOut10_13[7] , \nOut10_13[6] , \nOut10_13[5] , \nOut10_13[4] , 
        \nOut10_13[3] , \nOut10_13[2] , \nOut10_13[1] , \nOut10_13[0] }), 
        .WestIn({\nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }), .Out({
        \nOut9_13[7] , \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , 
        \nOut9_13[3] , \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_326 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut327[7] , \nScanOut327[6] , 
        \nScanOut327[5] , \nScanOut327[4] , \nScanOut327[3] , \nScanOut327[2] , 
        \nScanOut327[1] , \nScanOut327[0] }), .ScanOut({\nScanOut326[7] , 
        \nScanOut326[6] , \nScanOut326[5] , \nScanOut326[4] , \nScanOut326[3] , 
        \nScanOut326[2] , \nScanOut326[1] , \nScanOut326[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_5[7] , \nOut10_5[6] , \nOut10_5[5] , \nOut10_5[4] , 
        \nOut10_5[3] , \nOut10_5[2] , \nOut10_5[1] , \nOut10_5[0] }), 
        .SouthIn({\nOut10_7[7] , \nOut10_7[6] , \nOut10_7[5] , \nOut10_7[4] , 
        \nOut10_7[3] , \nOut10_7[2] , \nOut10_7[1] , \nOut10_7[0] }), .EastIn(
        {\nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }), .WestIn(
        {\nOut9_6[7] , \nOut9_6[6] , \nOut9_6[5] , \nOut9_6[4] , \nOut9_6[3] , 
        \nOut9_6[2] , \nOut9_6[1] , \nOut9_6[0] }), .Out({\nOut10_6[7] , 
        \nOut10_6[6] , \nOut10_6[5] , \nOut10_6[4] , \nOut10_6[3] , 
        \nOut10_6[2] , \nOut10_6[1] , \nOut10_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_537 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut538[7] , \nScanOut538[6] , 
        \nScanOut538[5] , \nScanOut538[4] , \nScanOut538[3] , \nScanOut538[2] , 
        \nScanOut538[1] , \nScanOut538[0] }), .ScanOut({\nScanOut537[7] , 
        \nScanOut537[6] , \nScanOut537[5] , \nScanOut537[4] , \nScanOut537[3] , 
        \nScanOut537[2] , \nScanOut537[1] , \nScanOut537[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_24[7] , \nOut16_24[6] , \nOut16_24[5] , \nOut16_24[4] , 
        \nOut16_24[3] , \nOut16_24[2] , \nOut16_24[1] , \nOut16_24[0] }), 
        .SouthIn({\nOut16_26[7] , \nOut16_26[6] , \nOut16_26[5] , 
        \nOut16_26[4] , \nOut16_26[3] , \nOut16_26[2] , \nOut16_26[1] , 
        \nOut16_26[0] }), .EastIn({\nOut17_25[7] , \nOut17_25[6] , 
        \nOut17_25[5] , \nOut17_25[4] , \nOut17_25[3] , \nOut17_25[2] , 
        \nOut17_25[1] , \nOut17_25[0] }), .WestIn({\nOut15_25[7] , 
        \nOut15_25[6] , \nOut15_25[5] , \nOut15_25[4] , \nOut15_25[3] , 
        \nOut15_25[2] , \nOut15_25[1] , \nOut15_25[0] }), .Out({\nOut16_25[7] , 
        \nOut16_25[6] , \nOut16_25[5] , \nOut16_25[4] , \nOut16_25[3] , 
        \nOut16_25[2] , \nOut16_25[1] , \nOut16_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_480 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut481[7] , \nScanOut481[6] , 
        \nScanOut481[5] , \nScanOut481[4] , \nScanOut481[3] , \nScanOut481[2] , 
        \nScanOut481[1] , \nScanOut481[0] }), .ScanOut({\nScanOut480[7] , 
        \nScanOut480[6] , \nScanOut480[5] , \nScanOut480[4] , \nScanOut480[3] , 
        \nScanOut480[2] , \nScanOut480[1] , \nScanOut480[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_0[7] , \nOut15_0[6] , 
        \nOut15_0[5] , \nOut15_0[4] , \nOut15_0[3] , \nOut15_0[2] , 
        \nOut15_0[1] , \nOut15_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_945 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut946[7] , \nScanOut946[6] , 
        \nScanOut946[5] , \nScanOut946[4] , \nScanOut946[3] , \nScanOut946[2] , 
        \nScanOut946[1] , \nScanOut946[0] }), .ScanOut({\nScanOut945[7] , 
        \nScanOut945[6] , \nScanOut945[5] , \nScanOut945[4] , \nScanOut945[3] , 
        \nScanOut945[2] , \nScanOut945[1] , \nScanOut945[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_16[7] , \nOut29_16[6] , \nOut29_16[5] , \nOut29_16[4] , 
        \nOut29_16[3] , \nOut29_16[2] , \nOut29_16[1] , \nOut29_16[0] }), 
        .SouthIn({\nOut29_18[7] , \nOut29_18[6] , \nOut29_18[5] , 
        \nOut29_18[4] , \nOut29_18[3] , \nOut29_18[2] , \nOut29_18[1] , 
        \nOut29_18[0] }), .EastIn({\nOut30_17[7] , \nOut30_17[6] , 
        \nOut30_17[5] , \nOut30_17[4] , \nOut30_17[3] , \nOut30_17[2] , 
        \nOut30_17[1] , \nOut30_17[0] }), .WestIn({\nOut28_17[7] , 
        \nOut28_17[6] , \nOut28_17[5] , \nOut28_17[4] , \nOut28_17[3] , 
        \nOut28_17[2] , \nOut28_17[1] , \nOut28_17[0] }), .Out({\nOut29_17[7] , 
        \nOut29_17[6] , \nOut29_17[5] , \nOut29_17[4] , \nOut29_17[3] , 
        \nOut29_17[2] , \nOut29_17[1] , \nOut29_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_510 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut511[7] , \nScanOut511[6] , 
        \nScanOut511[5] , \nScanOut511[4] , \nScanOut511[3] , \nScanOut511[2] , 
        \nScanOut511[1] , \nScanOut511[0] }), .ScanOut({\nScanOut510[7] , 
        \nScanOut510[6] , \nScanOut510[5] , \nScanOut510[4] , \nScanOut510[3] , 
        \nScanOut510[2] , \nScanOut510[1] , \nScanOut510[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut15_29[7] , \nOut15_29[6] , \nOut15_29[5] , \nOut15_29[4] , 
        \nOut15_29[3] , \nOut15_29[2] , \nOut15_29[1] , \nOut15_29[0] }), 
        .SouthIn({\nOut15_31[7] , \nOut15_31[6] , \nOut15_31[5] , 
        \nOut15_31[4] , \nOut15_31[3] , \nOut15_31[2] , \nOut15_31[1] , 
        \nOut15_31[0] }), .EastIn({\nOut16_30[7] , \nOut16_30[6] , 
        \nOut16_30[5] , \nOut16_30[4] , \nOut16_30[3] , \nOut16_30[2] , 
        \nOut16_30[1] , \nOut16_30[0] }), .WestIn({\nOut14_30[7] , 
        \nOut14_30[6] , \nOut14_30[5] , \nOut14_30[4] , \nOut14_30[3] , 
        \nOut14_30[2] , \nOut14_30[1] , \nOut14_30[0] }), .Out({\nOut15_30[7] , 
        \nOut15_30[6] , \nOut15_30[5] , \nOut15_30[4] , \nOut15_30[3] , 
        \nOut15_30[2] , \nOut15_30[1] , \nOut15_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_620 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut621[7] , \nScanOut621[6] , 
        \nScanOut621[5] , \nScanOut621[4] , \nScanOut621[3] , \nScanOut621[2] , 
        \nScanOut621[1] , \nScanOut621[0] }), .ScanOut({\nScanOut620[7] , 
        \nScanOut620[6] , \nScanOut620[5] , \nScanOut620[4] , \nScanOut620[3] , 
        \nScanOut620[2] , \nScanOut620[1] , \nScanOut620[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut19_11[7] , \nOut19_11[6] , \nOut19_11[5] , \nOut19_11[4] , 
        \nOut19_11[3] , \nOut19_11[2] , \nOut19_11[1] , \nOut19_11[0] }), 
        .SouthIn({\nOut19_13[7] , \nOut19_13[6] , \nOut19_13[5] , 
        \nOut19_13[4] , \nOut19_13[3] , \nOut19_13[2] , \nOut19_13[1] , 
        \nOut19_13[0] }), .EastIn({\nOut20_12[7] , \nOut20_12[6] , 
        \nOut20_12[5] , \nOut20_12[4] , \nOut20_12[3] , \nOut20_12[2] , 
        \nOut20_12[1] , \nOut20_12[0] }), .WestIn({\nOut18_12[7] , 
        \nOut18_12[6] , \nOut18_12[5] , \nOut18_12[4] , \nOut18_12[3] , 
        \nOut18_12[2] , \nOut18_12[1] , \nOut18_12[0] }), .Out({\nOut19_12[7] , 
        \nOut19_12[6] , \nOut19_12[5] , \nOut19_12[4] , \nOut19_12[3] , 
        \nOut19_12[2] , \nOut19_12[1] , \nOut19_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_962 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut963[7] , \nScanOut963[6] , 
        \nScanOut963[5] , \nScanOut963[4] , \nScanOut963[3] , \nScanOut963[2] , 
        \nScanOut963[1] , \nScanOut963[0] }), .ScanOut({\nScanOut962[7] , 
        \nScanOut962[6] , \nScanOut962[5] , \nScanOut962[4] , \nScanOut962[3] , 
        \nScanOut962[2] , \nScanOut962[1] , \nScanOut962[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_1[7] , \nOut30_1[6] , \nOut30_1[5] , \nOut30_1[4] , 
        \nOut30_1[3] , \nOut30_1[2] , \nOut30_1[1] , \nOut30_1[0] }), 
        .SouthIn({\nOut30_3[7] , \nOut30_3[6] , \nOut30_3[5] , \nOut30_3[4] , 
        \nOut30_3[3] , \nOut30_3[2] , \nOut30_3[1] , \nOut30_3[0] }), .EastIn(
        {\nOut31_2[7] , \nOut31_2[6] , \nOut31_2[5] , \nOut31_2[4] , 
        \nOut31_2[3] , \nOut31_2[2] , \nOut31_2[1] , \nOut31_2[0] }), .WestIn(
        {\nOut29_2[7] , \nOut29_2[6] , \nOut29_2[5] , \nOut29_2[4] , 
        \nOut29_2[3] , \nOut29_2[2] , \nOut29_2[1] , \nOut29_2[0] }), .Out({
        \nOut30_2[7] , \nOut30_2[6] , \nOut30_2[5] , \nOut30_2[4] , 
        \nOut30_2[3] , \nOut30_2[2] , \nOut30_2[1] , \nOut30_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_40 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut41[7] , \nScanOut41[6] , 
        \nScanOut41[5] , \nScanOut41[4] , \nScanOut41[3] , \nScanOut41[2] , 
        \nScanOut41[1] , \nScanOut41[0] }), .ScanOut({\nScanOut40[7] , 
        \nScanOut40[6] , \nScanOut40[5] , \nScanOut40[4] , \nScanOut40[3] , 
        \nScanOut40[2] , \nScanOut40[1] , \nScanOut40[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , \nOut1_7[4] , \nOut1_7[3] , 
        \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }), .SouthIn({\nOut1_9[7] , 
        \nOut1_9[6] , \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , 
        \nOut1_9[1] , \nOut1_9[0] }), .EastIn({\nOut2_8[7] , \nOut2_8[6] , 
        \nOut2_8[5] , \nOut2_8[4] , \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , 
        \nOut2_8[0] }), .WestIn({\nOut0_8[7] , \nOut0_8[6] , \nOut0_8[5] , 
        \nOut0_8[4] , \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , \nOut0_8[0] }), 
        .Out({\nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , \nOut1_8[4] , 
        \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_67 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut68[7] , \nScanOut68[6] , 
        \nScanOut68[5] , \nScanOut68[4] , \nScanOut68[3] , \nScanOut68[2] , 
        \nScanOut68[1] , \nScanOut68[0] }), .ScanOut({\nScanOut67[7] , 
        \nScanOut67[6] , \nScanOut67[5] , \nScanOut67[4] , \nScanOut67[3] , 
        \nScanOut67[2] , \nScanOut67[1] , \nScanOut67[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , 
        \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }), .SouthIn({\nOut2_4[7] , 
        \nOut2_4[6] , \nOut2_4[5] , \nOut2_4[4] , \nOut2_4[3] , \nOut2_4[2] , 
        \nOut2_4[1] , \nOut2_4[0] }), .EastIn({\nOut3_3[7] , \nOut3_3[6] , 
        \nOut3_3[5] , \nOut3_3[4] , \nOut3_3[3] , \nOut3_3[2] , \nOut3_3[1] , 
        \nOut3_3[0] }), .WestIn({\nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , 
        \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }), 
        .Out({\nOut2_3[7] , \nOut2_3[6] , \nOut2_3[5] , \nOut2_3[4] , 
        \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , \nOut2_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_144 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut145[7] , \nScanOut145[6] , 
        \nScanOut145[5] , \nScanOut145[4] , \nScanOut145[3] , \nScanOut145[2] , 
        \nScanOut145[1] , \nScanOut145[0] }), .ScanOut({\nScanOut144[7] , 
        \nScanOut144[6] , \nScanOut144[5] , \nScanOut144[4] , \nScanOut144[3] , 
        \nScanOut144[2] , \nScanOut144[1] , \nScanOut144[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_15[7] , \nOut4_15[6] , \nOut4_15[5] , \nOut4_15[4] , 
        \nOut4_15[3] , \nOut4_15[2] , \nOut4_15[1] , \nOut4_15[0] }), 
        .SouthIn({\nOut4_17[7] , \nOut4_17[6] , \nOut4_17[5] , \nOut4_17[4] , 
        \nOut4_17[3] , \nOut4_17[2] , \nOut4_17[1] , \nOut4_17[0] }), .EastIn(
        {\nOut5_16[7] , \nOut5_16[6] , \nOut5_16[5] , \nOut5_16[4] , 
        \nOut5_16[3] , \nOut5_16[2] , \nOut5_16[1] , \nOut5_16[0] }), .WestIn(
        {\nOut3_16[7] , \nOut3_16[6] , \nOut3_16[5] , \nOut3_16[4] , 
        \nOut3_16[3] , \nOut3_16[2] , \nOut3_16[1] , \nOut3_16[0] }), .Out({
        \nOut4_16[7] , \nOut4_16[6] , \nOut4_16[5] , \nOut4_16[4] , 
        \nOut4_16[3] , \nOut4_16[2] , \nOut4_16[1] , \nOut4_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_274 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut275[7] , \nScanOut275[6] , 
        \nScanOut275[5] , \nScanOut275[4] , \nScanOut275[3] , \nScanOut275[2] , 
        \nScanOut275[1] , \nScanOut275[0] }), .ScanOut({\nScanOut274[7] , 
        \nScanOut274[6] , \nScanOut274[5] , \nScanOut274[4] , \nScanOut274[3] , 
        \nScanOut274[2] , \nScanOut274[1] , \nScanOut274[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_17[7] , \nOut8_17[6] , \nOut8_17[5] , \nOut8_17[4] , 
        \nOut8_17[3] , \nOut8_17[2] , \nOut8_17[1] , \nOut8_17[0] }), 
        .SouthIn({\nOut8_19[7] , \nOut8_19[6] , \nOut8_19[5] , \nOut8_19[4] , 
        \nOut8_19[3] , \nOut8_19[2] , \nOut8_19[1] , \nOut8_19[0] }), .EastIn(
        {\nOut9_18[7] , \nOut9_18[6] , \nOut9_18[5] , \nOut9_18[4] , 
        \nOut9_18[3] , \nOut9_18[2] , \nOut9_18[1] , \nOut9_18[0] }), .WestIn(
        {\nOut7_18[7] , \nOut7_18[6] , \nOut7_18[5] , \nOut7_18[4] , 
        \nOut7_18[3] , \nOut7_18[2] , \nOut7_18[1] , \nOut7_18[0] }), .Out({
        \nOut8_18[7] , \nOut8_18[6] , \nOut8_18[5] , \nOut8_18[4] , 
        \nOut8_18[3] , \nOut8_18[2] , \nOut8_18[1] , \nOut8_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_348 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut349[7] , \nScanOut349[6] , 
        \nScanOut349[5] , \nScanOut349[4] , \nScanOut349[3] , \nScanOut349[2] , 
        \nScanOut349[1] , \nScanOut349[0] }), .ScanOut({\nScanOut348[7] , 
        \nScanOut348[6] , \nScanOut348[5] , \nScanOut348[4] , \nScanOut348[3] , 
        \nScanOut348[2] , \nScanOut348[1] , \nScanOut348[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_27[7] , \nOut10_27[6] , \nOut10_27[5] , \nOut10_27[4] , 
        \nOut10_27[3] , \nOut10_27[2] , \nOut10_27[1] , \nOut10_27[0] }), 
        .SouthIn({\nOut10_29[7] , \nOut10_29[6] , \nOut10_29[5] , 
        \nOut10_29[4] , \nOut10_29[3] , \nOut10_29[2] , \nOut10_29[1] , 
        \nOut10_29[0] }), .EastIn({\nOut11_28[7] , \nOut11_28[6] , 
        \nOut11_28[5] , \nOut11_28[4] , \nOut11_28[3] , \nOut11_28[2] , 
        \nOut11_28[1] , \nOut11_28[0] }), .WestIn({\nOut9_28[7] , 
        \nOut9_28[6] , \nOut9_28[5] , \nOut9_28[4] , \nOut9_28[3] , 
        \nOut9_28[2] , \nOut9_28[1] , \nOut9_28[0] }), .Out({\nOut10_28[7] , 
        \nOut10_28[6] , \nOut10_28[5] , \nOut10_28[4] , \nOut10_28[3] , 
        \nOut10_28[2] , \nOut10_28[1] , \nOut10_28[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_669 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut670[7] , \nScanOut670[6] , 
        \nScanOut670[5] , \nScanOut670[4] , \nScanOut670[3] , \nScanOut670[2] , 
        \nScanOut670[1] , \nScanOut670[0] }), .ScanOut({\nScanOut669[7] , 
        \nScanOut669[6] , \nScanOut669[5] , \nScanOut669[4] , \nScanOut669[3] , 
        \nScanOut669[2] , \nScanOut669[1] , \nScanOut669[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_28[7] , \nOut20_28[6] , \nOut20_28[5] , \nOut20_28[4] , 
        \nOut20_28[3] , \nOut20_28[2] , \nOut20_28[1] , \nOut20_28[0] }), 
        .SouthIn({\nOut20_30[7] , \nOut20_30[6] , \nOut20_30[5] , 
        \nOut20_30[4] , \nOut20_30[3] , \nOut20_30[2] , \nOut20_30[1] , 
        \nOut20_30[0] }), .EastIn({\nOut21_29[7] , \nOut21_29[6] , 
        \nOut21_29[5] , \nOut21_29[4] , \nOut21_29[3] , \nOut21_29[2] , 
        \nOut21_29[1] , \nOut21_29[0] }), .WestIn({\nOut19_29[7] , 
        \nOut19_29[6] , \nOut19_29[5] , \nOut19_29[4] , \nOut19_29[3] , 
        \nOut19_29[2] , \nOut19_29[1] , \nOut19_29[0] }), .Out({\nOut20_29[7] , 
        \nOut20_29[6] , \nOut20_29[5] , \nOut20_29[4] , \nOut20_29[3] , 
        \nOut20_29[2] , \nOut20_29[1] , \nOut20_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_559 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut560[7] , \nScanOut560[6] , 
        \nScanOut560[5] , \nScanOut560[4] , \nScanOut560[3] , \nScanOut560[2] , 
        \nScanOut560[1] , \nScanOut560[0] }), .ScanOut({\nScanOut559[7] , 
        \nScanOut559[6] , \nScanOut559[5] , \nScanOut559[4] , \nScanOut559[3] , 
        \nScanOut559[2] , \nScanOut559[1] , \nScanOut559[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_14[7] , \nOut17_14[6] , \nOut17_14[5] , \nOut17_14[4] , 
        \nOut17_14[3] , \nOut17_14[2] , \nOut17_14[1] , \nOut17_14[0] }), 
        .SouthIn({\nOut17_16[7] , \nOut17_16[6] , \nOut17_16[5] , 
        \nOut17_16[4] , \nOut17_16[3] , \nOut17_16[2] , \nOut17_16[1] , 
        \nOut17_16[0] }), .EastIn({\nOut18_15[7] , \nOut18_15[6] , 
        \nOut18_15[5] , \nOut18_15[4] , \nOut18_15[3] , \nOut18_15[2] , 
        \nOut18_15[1] , \nOut18_15[0] }), .WestIn({\nOut16_15[7] , 
        \nOut16_15[6] , \nOut16_15[5] , \nOut16_15[4] , \nOut16_15[3] , 
        \nOut16_15[2] , \nOut16_15[1] , \nOut16_15[0] }), .Out({\nOut17_15[7] , 
        \nOut17_15[6] , \nOut17_15[5] , \nOut17_15[4] , \nOut17_15[3] , 
        \nOut17_15[2] , \nOut17_15[1] , \nOut17_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_465 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut466[7] , \nScanOut466[6] , 
        \nScanOut466[5] , \nScanOut466[4] , \nScanOut466[3] , \nScanOut466[2] , 
        \nScanOut466[1] , \nScanOut466[0] }), .ScanOut({\nScanOut465[7] , 
        \nScanOut465[6] , \nScanOut465[5] , \nScanOut465[4] , \nScanOut465[3] , 
        \nScanOut465[2] , \nScanOut465[1] , \nScanOut465[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_16[7] , \nOut14_16[6] , \nOut14_16[5] , \nOut14_16[4] , 
        \nOut14_16[3] , \nOut14_16[2] , \nOut14_16[1] , \nOut14_16[0] }), 
        .SouthIn({\nOut14_18[7] , \nOut14_18[6] , \nOut14_18[5] , 
        \nOut14_18[4] , \nOut14_18[3] , \nOut14_18[2] , \nOut14_18[1] , 
        \nOut14_18[0] }), .EastIn({\nOut15_17[7] , \nOut15_17[6] , 
        \nOut15_17[5] , \nOut15_17[4] , \nOut15_17[3] , \nOut15_17[2] , 
        \nOut15_17[1] , \nOut15_17[0] }), .WestIn({\nOut13_17[7] , 
        \nOut13_17[6] , \nOut13_17[5] , \nOut13_17[4] , \nOut13_17[3] , 
        \nOut13_17[2] , \nOut13_17[1] , \nOut13_17[0] }), .Out({\nOut14_17[7] , 
        \nOut14_17[6] , \nOut14_17[5] , \nOut14_17[4] , \nOut14_17[3] , 
        \nOut14_17[2] , \nOut14_17[1] , \nOut14_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_817 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut818[7] , \nScanOut818[6] , 
        \nScanOut818[5] , \nScanOut818[4] , \nScanOut818[3] , \nScanOut818[2] , 
        \nScanOut818[1] , \nScanOut818[0] }), .ScanOut({\nScanOut817[7] , 
        \nScanOut817[6] , \nScanOut817[5] , \nScanOut817[4] , \nScanOut817[3] , 
        \nScanOut817[2] , \nScanOut817[1] , \nScanOut817[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_16[7] , \nOut25_16[6] , \nOut25_16[5] , \nOut25_16[4] , 
        \nOut25_16[3] , \nOut25_16[2] , \nOut25_16[1] , \nOut25_16[0] }), 
        .SouthIn({\nOut25_18[7] , \nOut25_18[6] , \nOut25_18[5] , 
        \nOut25_18[4] , \nOut25_18[3] , \nOut25_18[2] , \nOut25_18[1] , 
        \nOut25_18[0] }), .EastIn({\nOut26_17[7] , \nOut26_17[6] , 
        \nOut26_17[5] , \nOut26_17[4] , \nOut26_17[3] , \nOut26_17[2] , 
        \nOut26_17[1] , \nOut26_17[0] }), .WestIn({\nOut24_17[7] , 
        \nOut24_17[6] , \nOut24_17[5] , \nOut24_17[4] , \nOut24_17[3] , 
        \nOut24_17[2] , \nOut24_17[1] , \nOut24_17[0] }), .Out({\nOut25_17[7] , 
        \nOut25_17[6] , \nOut25_17[5] , \nOut25_17[4] , \nOut25_17[3] , 
        \nOut25_17[2] , \nOut25_17[1] , \nOut25_17[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_987 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut988[7] , \nScanOut988[6] , 
        \nScanOut988[5] , \nScanOut988[4] , \nScanOut988[3] , \nScanOut988[2] , 
        \nScanOut988[1] , \nScanOut988[0] }), .ScanOut({\nScanOut987[7] , 
        \nScanOut987[6] , \nScanOut987[5] , \nScanOut987[4] , \nScanOut987[3] , 
        \nScanOut987[2] , \nScanOut987[1] , \nScanOut987[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_26[7] , \nOut30_26[6] , \nOut30_26[5] , \nOut30_26[4] , 
        \nOut30_26[3] , \nOut30_26[2] , \nOut30_26[1] , \nOut30_26[0] }), 
        .SouthIn({\nOut30_28[7] , \nOut30_28[6] , \nOut30_28[5] , 
        \nOut30_28[4] , \nOut30_28[3] , \nOut30_28[2] , \nOut30_28[1] , 
        \nOut30_28[0] }), .EastIn({\nOut31_27[7] , \nOut31_27[6] , 
        \nOut31_27[5] , \nOut31_27[4] , \nOut31_27[3] , \nOut31_27[2] , 
        \nOut31_27[1] , \nOut31_27[0] }), .WestIn({\nOut29_27[7] , 
        \nOut29_27[6] , \nOut29_27[5] , \nOut29_27[4] , \nOut29_27[3] , 
        \nOut29_27[2] , \nOut29_27[1] , \nOut29_27[0] }), .Out({\nOut30_27[7] , 
        \nOut30_27[6] , \nOut30_27[5] , \nOut30_27[4] , \nOut30_27[3] , 
        \nOut30_27[2] , \nOut30_27[1] , \nOut30_27[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_163 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut164[7] , \nScanOut164[6] , 
        \nScanOut164[5] , \nScanOut164[4] , \nScanOut164[3] , \nScanOut164[2] , 
        \nScanOut164[1] , \nScanOut164[0] }), .ScanOut({\nScanOut163[7] , 
        \nScanOut163[6] , \nScanOut163[5] , \nScanOut163[4] , \nScanOut163[3] , 
        \nScanOut163[2] , \nScanOut163[1] , \nScanOut163[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_2[7] , \nOut5_2[6] , \nOut5_2[5] , \nOut5_2[4] , \nOut5_2[3] , 
        \nOut5_2[2] , \nOut5_2[1] , \nOut5_2[0] }), .SouthIn({\nOut5_4[7] , 
        \nOut5_4[6] , \nOut5_4[5] , \nOut5_4[4] , \nOut5_4[3] , \nOut5_4[2] , 
        \nOut5_4[1] , \nOut5_4[0] }), .EastIn({\nOut6_3[7] , \nOut6_3[6] , 
        \nOut6_3[5] , \nOut6_3[4] , \nOut6_3[3] , \nOut6_3[2] , \nOut6_3[1] , 
        \nOut6_3[0] }), .WestIn({\nOut4_3[7] , \nOut4_3[6] , \nOut4_3[5] , 
        \nOut4_3[4] , \nOut4_3[3] , \nOut4_3[2] , \nOut4_3[1] , \nOut4_3[0] }), 
        .Out({\nOut5_3[7] , \nOut5_3[6] , \nOut5_3[5] , \nOut5_3[4] , 
        \nOut5_3[3] , \nOut5_3[2] , \nOut5_3[1] , \nOut5_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_755 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut756[7] , \nScanOut756[6] , 
        \nScanOut756[5] , \nScanOut756[4] , \nScanOut756[3] , \nScanOut756[2] , 
        \nScanOut756[1] , \nScanOut756[0] }), .ScanOut({\nScanOut755[7] , 
        \nScanOut755[6] , \nScanOut755[5] , \nScanOut755[4] , \nScanOut755[3] , 
        \nScanOut755[2] , \nScanOut755[1] , \nScanOut755[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut23_18[7] , \nOut23_18[6] , \nOut23_18[5] , \nOut23_18[4] , 
        \nOut23_18[3] , \nOut23_18[2] , \nOut23_18[1] , \nOut23_18[0] }), 
        .SouthIn({\nOut23_20[7] , \nOut23_20[6] , \nOut23_20[5] , 
        \nOut23_20[4] , \nOut23_20[3] , \nOut23_20[2] , \nOut23_20[1] , 
        \nOut23_20[0] }), .EastIn({\nOut24_19[7] , \nOut24_19[6] , 
        \nOut24_19[5] , \nOut24_19[4] , \nOut24_19[3] , \nOut24_19[2] , 
        \nOut24_19[1] , \nOut24_19[0] }), .WestIn({\nOut22_19[7] , 
        \nOut22_19[6] , \nOut22_19[5] , \nOut22_19[4] , \nOut22_19[3] , 
        \nOut22_19[2] , \nOut22_19[1] , \nOut22_19[0] }), .Out({\nOut23_19[7] , 
        \nOut23_19[6] , \nOut23_19[5] , \nOut23_19[4] , \nOut23_19[3] , 
        \nOut23_19[2] , \nOut23_19[1] , \nOut23_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_772 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut773[7] , \nScanOut773[6] , 
        \nScanOut773[5] , \nScanOut773[4] , \nScanOut773[3] , \nScanOut773[2] , 
        \nScanOut773[1] , \nScanOut773[0] }), .ScanOut({\nScanOut772[7] , 
        \nScanOut772[6] , \nScanOut772[5] , \nScanOut772[4] , \nScanOut772[3] , 
        \nScanOut772[2] , \nScanOut772[1] , \nScanOut772[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_3[7] , \nOut24_3[6] , \nOut24_3[5] , \nOut24_3[4] , 
        \nOut24_3[3] , \nOut24_3[2] , \nOut24_3[1] , \nOut24_3[0] }), 
        .SouthIn({\nOut24_5[7] , \nOut24_5[6] , \nOut24_5[5] , \nOut24_5[4] , 
        \nOut24_5[3] , \nOut24_5[2] , \nOut24_5[1] , \nOut24_5[0] }), .EastIn(
        {\nOut25_4[7] , \nOut25_4[6] , \nOut25_4[5] , \nOut25_4[4] , 
        \nOut25_4[3] , \nOut25_4[2] , \nOut25_4[1] , \nOut25_4[0] }), .WestIn(
        {\nOut23_4[7] , \nOut23_4[6] , \nOut23_4[5] , \nOut23_4[4] , 
        \nOut23_4[3] , \nOut23_4[2] , \nOut23_4[1] , \nOut23_4[0] }), .Out({
        \nOut24_4[7] , \nOut24_4[6] , \nOut24_4[5] , \nOut24_4[4] , 
        \nOut24_4[3] , \nOut24_4[2] , \nOut24_4[1] , \nOut24_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_178 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut179[7] , \nScanOut179[6] , 
        \nScanOut179[5] , \nScanOut179[4] , \nScanOut179[3] , \nScanOut179[2] , 
        \nScanOut179[1] , \nScanOut179[0] }), .ScanOut({\nScanOut178[7] , 
        \nScanOut178[6] , \nScanOut178[5] , \nScanOut178[4] , \nScanOut178[3] , 
        \nScanOut178[2] , \nScanOut178[1] , \nScanOut178[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_17[7] , \nOut5_17[6] , \nOut5_17[5] , \nOut5_17[4] , 
        \nOut5_17[3] , \nOut5_17[2] , \nOut5_17[1] , \nOut5_17[0] }), 
        .SouthIn({\nOut5_19[7] , \nOut5_19[6] , \nOut5_19[5] , \nOut5_19[4] , 
        \nOut5_19[3] , \nOut5_19[2] , \nOut5_19[1] , \nOut5_19[0] }), .EastIn(
        {\nOut6_18[7] , \nOut6_18[6] , \nOut6_18[5] , \nOut6_18[4] , 
        \nOut6_18[3] , \nOut6_18[2] , \nOut6_18[1] , \nOut6_18[0] }), .WestIn(
        {\nOut4_18[7] , \nOut4_18[6] , \nOut4_18[5] , \nOut4_18[4] , 
        \nOut4_18[3] , \nOut4_18[2] , \nOut4_18[1] , \nOut4_18[0] }), .Out({
        \nOut5_18[7] , \nOut5_18[6] , \nOut5_18[5] , \nOut5_18[4] , 
        \nOut5_18[3] , \nOut5_18[2] , \nOut5_18[1] , \nOut5_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_248 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut249[7] , \nScanOut249[6] , 
        \nScanOut249[5] , \nScanOut249[4] , \nScanOut249[3] , \nScanOut249[2] , 
        \nScanOut249[1] , \nScanOut249[0] }), .ScanOut({\nScanOut248[7] , 
        \nScanOut248[6] , \nScanOut248[5] , \nScanOut248[4] , \nScanOut248[3] , 
        \nScanOut248[2] , \nScanOut248[1] , \nScanOut248[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_23[7] , \nOut7_23[6] , \nOut7_23[5] , \nOut7_23[4] , 
        \nOut7_23[3] , \nOut7_23[2] , \nOut7_23[1] , \nOut7_23[0] }), 
        .SouthIn({\nOut7_25[7] , \nOut7_25[6] , \nOut7_25[5] , \nOut7_25[4] , 
        \nOut7_25[3] , \nOut7_25[2] , \nOut7_25[1] , \nOut7_25[0] }), .EastIn(
        {\nOut8_24[7] , \nOut8_24[6] , \nOut8_24[5] , \nOut8_24[4] , 
        \nOut8_24[3] , \nOut8_24[2] , \nOut8_24[1] , \nOut8_24[0] }), .WestIn(
        {\nOut6_24[7] , \nOut6_24[6] , \nOut6_24[5] , \nOut6_24[4] , 
        \nOut6_24[3] , \nOut6_24[2] , \nOut6_24[1] , \nOut6_24[0] }), .Out({
        \nOut7_24[7] , \nOut7_24[6] , \nOut7_24[5] , \nOut7_24[4] , 
        \nOut7_24[3] , \nOut7_24[2] , \nOut7_24[1] , \nOut7_24[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_253 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut254[7] , \nScanOut254[6] , 
        \nScanOut254[5] , \nScanOut254[4] , \nScanOut254[3] , \nScanOut254[2] , 
        \nScanOut254[1] , \nScanOut254[0] }), .ScanOut({\nScanOut253[7] , 
        \nScanOut253[6] , \nScanOut253[5] , \nScanOut253[4] , \nScanOut253[3] , 
        \nScanOut253[2] , \nScanOut253[1] , \nScanOut253[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_28[7] , \nOut7_28[6] , \nOut7_28[5] , \nOut7_28[4] , 
        \nOut7_28[3] , \nOut7_28[2] , \nOut7_28[1] , \nOut7_28[0] }), 
        .SouthIn({\nOut7_30[7] , \nOut7_30[6] , \nOut7_30[5] , \nOut7_30[4] , 
        \nOut7_30[3] , \nOut7_30[2] , \nOut7_30[1] , \nOut7_30[0] }), .EastIn(
        {\nOut8_29[7] , \nOut8_29[6] , \nOut8_29[5] , \nOut8_29[4] , 
        \nOut8_29[3] , \nOut8_29[2] , \nOut8_29[1] , \nOut8_29[0] }), .WestIn(
        {\nOut6_29[7] , \nOut6_29[6] , \nOut6_29[5] , \nOut6_29[4] , 
        \nOut6_29[3] , \nOut6_29[2] , \nOut6_29[1] , \nOut6_29[0] }), .Out({
        \nOut7_29[7] , \nOut7_29[6] , \nOut7_29[5] , \nOut7_29[4] , 
        \nOut7_29[3] , \nOut7_29[2] , \nOut7_29[1] , \nOut7_29[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_442 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut443[7] , \nScanOut443[6] , 
        \nScanOut443[5] , \nScanOut443[4] , \nScanOut443[3] , \nScanOut443[2] , 
        \nScanOut443[1] , \nScanOut443[0] }), .ScanOut({\nScanOut442[7] , 
        \nScanOut442[6] , \nScanOut442[5] , \nScanOut442[4] , \nScanOut442[3] , 
        \nScanOut442[2] , \nScanOut442[1] , \nScanOut442[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_25[7] , \nOut13_25[6] , \nOut13_25[5] , \nOut13_25[4] , 
        \nOut13_25[3] , \nOut13_25[2] , \nOut13_25[1] , \nOut13_25[0] }), 
        .SouthIn({\nOut13_27[7] , \nOut13_27[6] , \nOut13_27[5] , 
        \nOut13_27[4] , \nOut13_27[3] , \nOut13_27[2] , \nOut13_27[1] , 
        \nOut13_27[0] }), .EastIn({\nOut14_26[7] , \nOut14_26[6] , 
        \nOut14_26[5] , \nOut14_26[4] , \nOut14_26[3] , \nOut14_26[2] , 
        \nOut14_26[1] , \nOut14_26[0] }), .WestIn({\nOut12_26[7] , 
        \nOut12_26[6] , \nOut12_26[5] , \nOut12_26[4] , \nOut12_26[3] , 
        \nOut12_26[2] , \nOut12_26[1] , \nOut12_26[0] }), .Out({\nOut13_26[7] , 
        \nOut13_26[6] , \nOut13_26[5] , \nOut13_26[4] , \nOut13_26[3] , 
        \nOut13_26[2] , \nOut13_26[1] , \nOut13_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_459 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut460[7] , \nScanOut460[6] , 
        \nScanOut460[5] , \nScanOut460[4] , \nScanOut460[3] , \nScanOut460[2] , 
        \nScanOut460[1] , \nScanOut460[0] }), .ScanOut({\nScanOut459[7] , 
        \nScanOut459[6] , \nScanOut459[5] , \nScanOut459[4] , \nScanOut459[3] , 
        \nScanOut459[2] , \nScanOut459[1] , \nScanOut459[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_10[7] , \nOut14_10[6] , \nOut14_10[5] , \nOut14_10[4] , 
        \nOut14_10[3] , \nOut14_10[2] , \nOut14_10[1] , \nOut14_10[0] }), 
        .SouthIn({\nOut14_12[7] , \nOut14_12[6] , \nOut14_12[5] , 
        \nOut14_12[4] , \nOut14_12[3] , \nOut14_12[2] , \nOut14_12[1] , 
        \nOut14_12[0] }), .EastIn({\nOut15_11[7] , \nOut15_11[6] , 
        \nOut15_11[5] , \nOut15_11[4] , \nOut15_11[3] , \nOut15_11[2] , 
        \nOut15_11[1] , \nOut15_11[0] }), .WestIn({\nOut13_11[7] , 
        \nOut13_11[6] , \nOut13_11[5] , \nOut13_11[4] , \nOut13_11[3] , 
        \nOut13_11[2] , \nOut13_11[1] , \nOut13_11[0] }), .Out({\nOut14_11[7] , 
        \nOut14_11[6] , \nOut14_11[5] , \nOut14_11[4] , \nOut14_11[3] , 
        \nOut14_11[2] , \nOut14_11[1] , \nOut14_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_830 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut831[7] , \nScanOut831[6] , 
        \nScanOut831[5] , \nScanOut831[4] , \nScanOut831[3] , \nScanOut831[2] , 
        \nScanOut831[1] , \nScanOut831[0] }), .ScanOut({\nScanOut830[7] , 
        \nScanOut830[6] , \nScanOut830[5] , \nScanOut830[4] , \nScanOut830[3] , 
        \nScanOut830[2] , \nScanOut830[1] , \nScanOut830[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut25_29[7] , \nOut25_29[6] , \nOut25_29[5] , \nOut25_29[4] , 
        \nOut25_29[3] , \nOut25_29[2] , \nOut25_29[1] , \nOut25_29[0] }), 
        .SouthIn({\nOut25_31[7] , \nOut25_31[6] , \nOut25_31[5] , 
        \nOut25_31[4] , \nOut25_31[3] , \nOut25_31[2] , \nOut25_31[1] , 
        \nOut25_31[0] }), .EastIn({\nOut26_30[7] , \nOut26_30[6] , 
        \nOut26_30[5] , \nOut26_30[4] , \nOut26_30[3] , \nOut26_30[2] , 
        \nOut26_30[1] , \nOut26_30[0] }), .WestIn({\nOut24_30[7] , 
        \nOut24_30[6] , \nOut24_30[5] , \nOut24_30[4] , \nOut24_30[3] , 
        \nOut24_30[2] , \nOut24_30[1] , \nOut24_30[0] }), .Out({\nOut25_30[7] , 
        \nOut25_30[6] , \nOut25_30[5] , \nOut25_30[4] , \nOut25_30[3] , 
        \nOut25_30[2] , \nOut25_30[1] , \nOut25_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_769 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut770[7] , \nScanOut770[6] , 
        \nScanOut770[5] , \nScanOut770[4] , \nScanOut770[3] , \nScanOut770[2] , 
        \nScanOut770[1] , \nScanOut770[0] }), .ScanOut({\nScanOut769[7] , 
        \nScanOut769[6] , \nScanOut769[5] , \nScanOut769[4] , \nScanOut769[3] , 
        \nScanOut769[2] , \nScanOut769[1] , \nScanOut769[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut24_0[7] , \nOut24_0[6] , \nOut24_0[5] , \nOut24_0[4] , 
        \nOut24_0[3] , \nOut24_0[2] , \nOut24_0[1] , \nOut24_0[0] }), 
        .SouthIn({\nOut24_2[7] , \nOut24_2[6] , \nOut24_2[5] , \nOut24_2[4] , 
        \nOut24_2[3] , \nOut24_2[2] , \nOut24_2[1] , \nOut24_2[0] }), .EastIn(
        {\nOut25_1[7] , \nOut25_1[6] , \nOut25_1[5] , \nOut25_1[4] , 
        \nOut25_1[3] , \nOut25_1[2] , \nOut25_1[1] , \nOut25_1[0] }), .WestIn(
        {\nOut23_1[7] , \nOut23_1[6] , \nOut23_1[5] , \nOut23_1[4] , 
        \nOut23_1[3] , \nOut23_1[2] , \nOut23_1[1] , \nOut23_1[0] }), .Out({
        \nOut24_1[7] , \nOut24_1[6] , \nOut24_1[5] , \nOut24_1[4] , 
        \nOut24_1[3] , \nOut24_1[2] , \nOut24_1[1] , \nOut24_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_353 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut354[7] , \nScanOut354[6] , 
        \nScanOut354[5] , \nScanOut354[4] , \nScanOut354[3] , \nScanOut354[2] , 
        \nScanOut354[1] , \nScanOut354[0] }), .ScanOut({\nScanOut353[7] , 
        \nScanOut353[6] , \nScanOut353[5] , \nScanOut353[4] , \nScanOut353[3] , 
        \nScanOut353[2] , \nScanOut353[1] , \nScanOut353[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_0[7] , \nOut11_0[6] , \nOut11_0[5] , \nOut11_0[4] , 
        \nOut11_0[3] , \nOut11_0[2] , \nOut11_0[1] , \nOut11_0[0] }), 
        .SouthIn({\nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }), .EastIn(
        {\nOut12_1[7] , \nOut12_1[6] , \nOut12_1[5] , \nOut12_1[4] , 
        \nOut12_1[3] , \nOut12_1[2] , \nOut12_1[1] , \nOut12_1[0] }), .WestIn(
        {\nOut10_1[7] , \nOut10_1[6] , \nOut10_1[5] , \nOut10_1[4] , 
        \nOut10_1[3] , \nOut10_1[2] , \nOut10_1[1] , \nOut10_1[0] }), .Out({
        \nOut11_1[7] , \nOut11_1[6] , \nOut11_1[5] , \nOut11_1[4] , 
        \nOut11_1[3] , \nOut11_1[2] , \nOut11_1[1] , \nOut11_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_542 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut543[7] , \nScanOut543[6] , 
        \nScanOut543[5] , \nScanOut543[4] , \nScanOut543[3] , \nScanOut543[2] , 
        \nScanOut543[1] , \nScanOut543[0] }), .ScanOut({\nScanOut542[7] , 
        \nScanOut542[6] , \nScanOut542[5] , \nScanOut542[4] , \nScanOut542[3] , 
        \nScanOut542[2] , \nScanOut542[1] , \nScanOut542[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut16_29[7] , \nOut16_29[6] , \nOut16_29[5] , \nOut16_29[4] , 
        \nOut16_29[3] , \nOut16_29[2] , \nOut16_29[1] , \nOut16_29[0] }), 
        .SouthIn({\nOut16_31[7] , \nOut16_31[6] , \nOut16_31[5] , 
        \nOut16_31[4] , \nOut16_31[3] , \nOut16_31[2] , \nOut16_31[1] , 
        \nOut16_31[0] }), .EastIn({\nOut17_30[7] , \nOut17_30[6] , 
        \nOut17_30[5] , \nOut17_30[4] , \nOut17_30[3] , \nOut17_30[2] , 
        \nOut17_30[1] , \nOut17_30[0] }), .WestIn({\nOut15_30[7] , 
        \nOut15_30[6] , \nOut15_30[5] , \nOut15_30[4] , \nOut15_30[3] , 
        \nOut15_30[2] , \nOut15_30[1] , \nOut15_30[0] }), .Out({\nOut16_30[7] , 
        \nOut16_30[6] , \nOut16_30[5] , \nOut16_30[4] , \nOut16_30[3] , 
        \nOut16_30[2] , \nOut16_30[1] , \nOut16_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_930 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut931[7] , \nScanOut931[6] , 
        \nScanOut931[5] , \nScanOut931[4] , \nScanOut931[3] , \nScanOut931[2] , 
        \nScanOut931[1] , \nScanOut931[0] }), .ScanOut({\nScanOut930[7] , 
        \nScanOut930[6] , \nScanOut930[5] , \nScanOut930[4] , \nScanOut930[3] , 
        \nScanOut930[2] , \nScanOut930[1] , \nScanOut930[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut29_1[7] , \nOut29_1[6] , \nOut29_1[5] , \nOut29_1[4] , 
        \nOut29_1[3] , \nOut29_1[2] , \nOut29_1[1] , \nOut29_1[0] }), 
        .SouthIn({\nOut29_3[7] , \nOut29_3[6] , \nOut29_3[5] , \nOut29_3[4] , 
        \nOut29_3[3] , \nOut29_3[2] , \nOut29_3[1] , \nOut29_3[0] }), .EastIn(
        {\nOut30_2[7] , \nOut30_2[6] , \nOut30_2[5] , \nOut30_2[4] , 
        \nOut30_2[3] , \nOut30_2[2] , \nOut30_2[1] , \nOut30_2[0] }), .WestIn(
        {\nOut28_2[7] , \nOut28_2[6] , \nOut28_2[5] , \nOut28_2[4] , 
        \nOut28_2[3] , \nOut28_2[2] , \nOut28_2[1] , \nOut28_2[0] }), .Out({
        \nOut29_2[7] , \nOut29_2[6] , \nOut29_2[5] , \nOut29_2[4] , 
        \nOut29_2[3] , \nOut29_2[2] , \nOut29_2[1] , \nOut29_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_672 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut673[7] , \nScanOut673[6] , 
        \nScanOut673[5] , \nScanOut673[4] , \nScanOut673[3] , \nScanOut673[2] , 
        \nScanOut673[1] , \nScanOut673[0] }), .ScanOut({\nScanOut672[7] , 
        \nScanOut672[6] , \nScanOut672[5] , \nScanOut672[4] , \nScanOut672[3] , 
        \nScanOut672[2] , \nScanOut672[1] , \nScanOut672[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut21_0[7] , \nOut21_0[6] , 
        \nOut21_0[5] , \nOut21_0[4] , \nOut21_0[3] , \nOut21_0[2] , 
        \nOut21_0[1] , \nOut21_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_82 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut83[7] , \nScanOut83[6] , 
        \nScanOut83[5] , \nScanOut83[4] , \nScanOut83[3] , \nScanOut83[2] , 
        \nScanOut83[1] , \nScanOut83[0] }), .ScanOut({\nScanOut82[7] , 
        \nScanOut82[6] , \nScanOut82[5] , \nScanOut82[4] , \nScanOut82[3] , 
        \nScanOut82[2] , \nScanOut82[1] , \nScanOut82[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_17[7] , \nOut2_17[6] , \nOut2_17[5] , \nOut2_17[4] , 
        \nOut2_17[3] , \nOut2_17[2] , \nOut2_17[1] , \nOut2_17[0] }), 
        .SouthIn({\nOut2_19[7] , \nOut2_19[6] , \nOut2_19[5] , \nOut2_19[4] , 
        \nOut2_19[3] , \nOut2_19[2] , \nOut2_19[1] , \nOut2_19[0] }), .EastIn(
        {\nOut3_18[7] , \nOut3_18[6] , \nOut3_18[5] , \nOut3_18[4] , 
        \nOut3_18[3] , \nOut3_18[2] , \nOut3_18[1] , \nOut3_18[0] }), .WestIn(
        {\nOut1_18[7] , \nOut1_18[6] , \nOut1_18[5] , \nOut1_18[4] , 
        \nOut1_18[3] , \nOut1_18[2] , \nOut1_18[1] , \nOut1_18[0] }), .Out({
        \nOut2_18[7] , \nOut2_18[6] , \nOut2_18[5] , \nOut2_18[4] , 
        \nOut2_18[3] , \nOut2_18[2] , \nOut2_18[1] , \nOut2_18[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_116 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut117[7] , \nScanOut117[6] , 
        \nScanOut117[5] , \nScanOut117[4] , \nScanOut117[3] , \nScanOut117[2] , 
        \nScanOut117[1] , \nScanOut117[0] }), .ScanOut({\nScanOut116[7] , 
        \nScanOut116[6] , \nScanOut116[5] , \nScanOut116[4] , \nScanOut116[3] , 
        \nScanOut116[2] , \nScanOut116[1] , \nScanOut116[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_19[7] , \nOut3_19[6] , \nOut3_19[5] , \nOut3_19[4] , 
        \nOut3_19[3] , \nOut3_19[2] , \nOut3_19[1] , \nOut3_19[0] }), 
        .SouthIn({\nOut3_21[7] , \nOut3_21[6] , \nOut3_21[5] , \nOut3_21[4] , 
        \nOut3_21[3] , \nOut3_21[2] , \nOut3_21[1] , \nOut3_21[0] }), .EastIn(
        {\nOut4_20[7] , \nOut4_20[6] , \nOut4_20[5] , \nOut4_20[4] , 
        \nOut4_20[3] , \nOut4_20[2] , \nOut4_20[1] , \nOut4_20[0] }), .WestIn(
        {\nOut2_20[7] , \nOut2_20[6] , \nOut2_20[5] , \nOut2_20[4] , 
        \nOut2_20[3] , \nOut2_20[2] , \nOut2_20[1] , \nOut2_20[0] }), .Out({
        \nOut3_20[7] , \nOut3_20[6] , \nOut3_20[5] , \nOut3_20[4] , 
        \nOut3_20[3] , \nOut3_20[2] , \nOut3_20[1] , \nOut3_20[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_131 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut132[7] , \nScanOut132[6] , 
        \nScanOut132[5] , \nScanOut132[4] , \nScanOut132[3] , \nScanOut132[2] , 
        \nScanOut132[1] , \nScanOut132[0] }), .ScanOut({\nScanOut131[7] , 
        \nScanOut131[6] , \nScanOut131[5] , \nScanOut131[4] , \nScanOut131[3] , 
        \nScanOut131[2] , \nScanOut131[1] , \nScanOut131[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_2[7] , \nOut4_2[6] , \nOut4_2[5] , \nOut4_2[4] , \nOut4_2[3] , 
        \nOut4_2[2] , \nOut4_2[1] , \nOut4_2[0] }), .SouthIn({\nOut4_4[7] , 
        \nOut4_4[6] , \nOut4_4[5] , \nOut4_4[4] , \nOut4_4[3] , \nOut4_4[2] , 
        \nOut4_4[1] , \nOut4_4[0] }), .EastIn({\nOut5_3[7] , \nOut5_3[6] , 
        \nOut5_3[5] , \nOut5_3[4] , \nOut5_3[3] , \nOut5_3[2] , \nOut5_3[1] , 
        \nOut5_3[0] }), .WestIn({\nOut3_3[7] , \nOut3_3[6] , \nOut3_3[5] , 
        \nOut3_3[4] , \nOut3_3[3] , \nOut3_3[2] , \nOut3_3[1] , \nOut3_3[0] }), 
        .Out({\nOut4_3[7] , \nOut4_3[6] , \nOut4_3[5] , \nOut4_3[4] , 
        \nOut4_3[3] , \nOut4_3[2] , \nOut4_3[1] , \nOut4_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_374 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut375[7] , \nScanOut375[6] , 
        \nScanOut375[5] , \nScanOut375[4] , \nScanOut375[3] , \nScanOut375[2] , 
        \nScanOut375[1] , \nScanOut375[0] }), .ScanOut({\nScanOut374[7] , 
        \nScanOut374[6] , \nScanOut374[5] , \nScanOut374[4] , \nScanOut374[3] , 
        \nScanOut374[2] , \nScanOut374[1] , \nScanOut374[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_21[7] , \nOut11_21[6] , \nOut11_21[5] , \nOut11_21[4] , 
        \nOut11_21[3] , \nOut11_21[2] , \nOut11_21[1] , \nOut11_21[0] }), 
        .SouthIn({\nOut11_23[7] , \nOut11_23[6] , \nOut11_23[5] , 
        \nOut11_23[4] , \nOut11_23[3] , \nOut11_23[2] , \nOut11_23[1] , 
        \nOut11_23[0] }), .EastIn({\nOut12_22[7] , \nOut12_22[6] , 
        \nOut12_22[5] , \nOut12_22[4] , \nOut12_22[3] , \nOut12_22[2] , 
        \nOut12_22[1] , \nOut12_22[0] }), .WestIn({\nOut10_22[7] , 
        \nOut10_22[6] , \nOut10_22[5] , \nOut10_22[4] , \nOut10_22[3] , 
        \nOut10_22[2] , \nOut10_22[1] , \nOut10_22[0] }), .Out({\nOut11_22[7] , 
        \nOut11_22[6] , \nOut11_22[5] , \nOut11_22[4] , \nOut11_22[3] , 
        \nOut11_22[2] , \nOut11_22[1] , \nOut11_22[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_565 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut566[7] , \nScanOut566[6] , 
        \nScanOut566[5] , \nScanOut566[4] , \nScanOut566[3] , \nScanOut566[2] , 
        \nScanOut566[1] , \nScanOut566[0] }), .ScanOut({\nScanOut565[7] , 
        \nScanOut565[6] , \nScanOut565[5] , \nScanOut565[4] , \nScanOut565[3] , 
        \nScanOut565[2] , \nScanOut565[1] , \nScanOut565[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut17_20[7] , \nOut17_20[6] , \nOut17_20[5] , \nOut17_20[4] , 
        \nOut17_20[3] , \nOut17_20[2] , \nOut17_20[1] , \nOut17_20[0] }), 
        .SouthIn({\nOut17_22[7] , \nOut17_22[6] , \nOut17_22[5] , 
        \nOut17_22[4] , \nOut17_22[3] , \nOut17_22[2] , \nOut17_22[1] , 
        \nOut17_22[0] }), .EastIn({\nOut18_21[7] , \nOut18_21[6] , 
        \nOut18_21[5] , \nOut18_21[4] , \nOut18_21[3] , \nOut18_21[2] , 
        \nOut18_21[1] , \nOut18_21[0] }), .WestIn({\nOut16_21[7] , 
        \nOut16_21[6] , \nOut16_21[5] , \nOut16_21[4] , \nOut16_21[3] , 
        \nOut16_21[2] , \nOut16_21[1] , \nOut16_21[0] }), .Out({\nOut17_21[7] , 
        \nOut17_21[6] , \nOut17_21[5] , \nOut17_21[4] , \nOut17_21[3] , 
        \nOut17_21[2] , \nOut17_21[1] , \nOut17_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_655 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut656[7] , \nScanOut656[6] , 
        \nScanOut656[5] , \nScanOut656[4] , \nScanOut656[3] , \nScanOut656[2] , 
        \nScanOut656[1] , \nScanOut656[0] }), .ScanOut({\nScanOut655[7] , 
        \nScanOut655[6] , \nScanOut655[5] , \nScanOut655[4] , \nScanOut655[3] , 
        \nScanOut655[2] , \nScanOut655[1] , \nScanOut655[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut20_14[7] , \nOut20_14[6] , \nOut20_14[5] , \nOut20_14[4] , 
        \nOut20_14[3] , \nOut20_14[2] , \nOut20_14[1] , \nOut20_14[0] }), 
        .SouthIn({\nOut20_16[7] , \nOut20_16[6] , \nOut20_16[5] , 
        \nOut20_16[4] , \nOut20_16[3] , \nOut20_16[2] , \nOut20_16[1] , 
        \nOut20_16[0] }), .EastIn({\nOut21_15[7] , \nOut21_15[6] , 
        \nOut21_15[5] , \nOut21_15[4] , \nOut21_15[3] , \nOut21_15[2] , 
        \nOut21_15[1] , \nOut21_15[0] }), .WestIn({\nOut19_15[7] , 
        \nOut19_15[6] , \nOut19_15[5] , \nOut19_15[4] , \nOut19_15[3] , 
        \nOut19_15[2] , \nOut19_15[1] , \nOut19_15[0] }), .Out({\nOut20_15[7] , 
        \nOut20_15[6] , \nOut20_15[5] , \nOut20_15[4] , \nOut20_15[3] , 
        \nOut20_15[2] , \nOut20_15[1] , \nOut20_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_720 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut721[7] , \nScanOut721[6] , 
        \nScanOut721[5] , \nScanOut721[4] , \nScanOut721[3] , \nScanOut721[2] , 
        \nScanOut721[1] , \nScanOut721[0] }), .ScanOut({\nScanOut720[7] , 
        \nScanOut720[6] , \nScanOut720[5] , \nScanOut720[4] , \nScanOut720[3] , 
        \nScanOut720[2] , \nScanOut720[1] , \nScanOut720[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_15[7] , \nOut22_15[6] , \nOut22_15[5] , \nOut22_15[4] , 
        \nOut22_15[3] , \nOut22_15[2] , \nOut22_15[1] , \nOut22_15[0] }), 
        .SouthIn({\nOut22_17[7] , \nOut22_17[6] , \nOut22_17[5] , 
        \nOut22_17[4] , \nOut22_17[3] , \nOut22_17[2] , \nOut22_17[1] , 
        \nOut22_17[0] }), .EastIn({\nOut23_16[7] , \nOut23_16[6] , 
        \nOut23_16[5] , \nOut23_16[4] , \nOut23_16[3] , \nOut23_16[2] , 
        \nOut23_16[1] , \nOut23_16[0] }), .WestIn({\nOut21_16[7] , 
        \nOut21_16[6] , \nOut21_16[5] , \nOut21_16[4] , \nOut21_16[3] , 
        \nOut21_16[2] , \nOut21_16[1] , \nOut21_16[0] }), .Out({\nOut22_16[7] , 
        \nOut22_16[6] , \nOut22_16[5] , \nOut22_16[4] , \nOut22_16[3] , 
        \nOut22_16[2] , \nOut22_16[1] , \nOut22_16[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_887 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut888[7] , \nScanOut888[6] , 
        \nScanOut888[5] , \nScanOut888[4] , \nScanOut888[3] , \nScanOut888[2] , 
        \nScanOut888[1] , \nScanOut888[0] }), .ScanOut({\nScanOut887[7] , 
        \nScanOut887[6] , \nScanOut887[5] , \nScanOut887[4] , \nScanOut887[3] , 
        \nScanOut887[2] , \nScanOut887[1] , \nScanOut887[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut27_22[7] , \nOut27_22[6] , \nOut27_22[5] , \nOut27_22[4] , 
        \nOut27_22[3] , \nOut27_22[2] , \nOut27_22[1] , \nOut27_22[0] }), 
        .SouthIn({\nOut27_24[7] , \nOut27_24[6] , \nOut27_24[5] , 
        \nOut27_24[4] , \nOut27_24[3] , \nOut27_24[2] , \nOut27_24[1] , 
        \nOut27_24[0] }), .EastIn({\nOut28_23[7] , \nOut28_23[6] , 
        \nOut28_23[5] , \nOut28_23[4] , \nOut28_23[3] , \nOut28_23[2] , 
        \nOut28_23[1] , \nOut28_23[0] }), .WestIn({\nOut26_23[7] , 
        \nOut26_23[6] , \nOut26_23[5] , \nOut26_23[4] , \nOut26_23[3] , 
        \nOut26_23[2] , \nOut26_23[1] , \nOut26_23[0] }), .Out({\nOut27_23[7] , 
        \nOut27_23[6] , \nOut27_23[5] , \nOut27_23[4] , \nOut27_23[3] , 
        \nOut27_23[2] , \nOut27_23[1] , \nOut27_23[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_917 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut918[7] , \nScanOut918[6] , 
        \nScanOut918[5] , \nScanOut918[4] , \nScanOut918[3] , \nScanOut918[2] , 
        \nScanOut918[1] , \nScanOut918[0] }), .ScanOut({\nScanOut917[7] , 
        \nScanOut917[6] , \nScanOut917[5] , \nScanOut917[4] , \nScanOut917[3] , 
        \nScanOut917[2] , \nScanOut917[1] , \nScanOut917[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut28_20[7] , \nOut28_20[6] , \nOut28_20[5] , \nOut28_20[4] , 
        \nOut28_20[3] , \nOut28_20[2] , \nOut28_20[1] , \nOut28_20[0] }), 
        .SouthIn({\nOut28_22[7] , \nOut28_22[6] , \nOut28_22[5] , 
        \nOut28_22[4] , \nOut28_22[3] , \nOut28_22[2] , \nOut28_22[1] , 
        \nOut28_22[0] }), .EastIn({\nOut29_21[7] , \nOut29_21[6] , 
        \nOut29_21[5] , \nOut29_21[4] , \nOut29_21[3] , \nOut29_21[2] , 
        \nOut29_21[1] , \nOut29_21[0] }), .WestIn({\nOut27_21[7] , 
        \nOut27_21[6] , \nOut27_21[5] , \nOut27_21[4] , \nOut27_21[3] , 
        \nOut27_21[2] , \nOut27_21[1] , \nOut27_21[0] }), .Out({\nOut28_21[7] , 
        \nOut28_21[6] , \nOut28_21[5] , \nOut28_21[4] , \nOut28_21[3] , 
        \nOut28_21[2] , \nOut28_21[1] , \nOut28_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_979 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut980[7] , \nScanOut980[6] , 
        \nScanOut980[5] , \nScanOut980[4] , \nScanOut980[3] , \nScanOut980[2] , 
        \nScanOut980[1] , \nScanOut980[0] }), .ScanOut({\nScanOut979[7] , 
        \nScanOut979[6] , \nScanOut979[5] , \nScanOut979[4] , \nScanOut979[3] , 
        \nScanOut979[2] , \nScanOut979[1] , \nScanOut979[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut30_18[7] , \nOut30_18[6] , \nOut30_18[5] , \nOut30_18[4] , 
        \nOut30_18[3] , \nOut30_18[2] , \nOut30_18[1] , \nOut30_18[0] }), 
        .SouthIn({\nOut30_20[7] , \nOut30_20[6] , \nOut30_20[5] , 
        \nOut30_20[4] , \nOut30_20[3] , \nOut30_20[2] , \nOut30_20[1] , 
        \nOut30_20[0] }), .EastIn({\nOut31_19[7] , \nOut31_19[6] , 
        \nOut31_19[5] , \nOut31_19[4] , \nOut31_19[3] , \nOut31_19[2] , 
        \nOut31_19[1] , \nOut31_19[0] }), .WestIn({\nOut29_19[7] , 
        \nOut29_19[6] , \nOut29_19[5] , \nOut29_19[4] , \nOut29_19[3] , 
        \nOut29_19[2] , \nOut29_19[1] , \nOut29_19[0] }), .Out({\nOut30_19[7] , 
        \nOut30_19[6] , \nOut30_19[5] , \nOut30_19[4] , \nOut30_19[3] , 
        \nOut30_19[2] , \nOut30_19[1] , \nOut30_19[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_201 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut202[7] , \nScanOut202[6] , 
        \nScanOut202[5] , \nScanOut202[4] , \nScanOut202[3] , \nScanOut202[2] , 
        \nScanOut202[1] , \nScanOut202[0] }), .ScanOut({\nScanOut201[7] , 
        \nScanOut201[6] , \nScanOut201[5] , \nScanOut201[4] , \nScanOut201[3] , 
        \nScanOut201[2] , \nScanOut201[1] , \nScanOut201[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_8[7] , \nOut6_8[6] , \nOut6_8[5] , \nOut6_8[4] , \nOut6_8[3] , 
        \nOut6_8[2] , \nOut6_8[1] , \nOut6_8[0] }), .SouthIn({\nOut6_10[7] , 
        \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , \nOut6_10[3] , 
        \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }), .EastIn({\nOut7_9[7] , 
        \nOut7_9[6] , \nOut7_9[5] , \nOut7_9[4] , \nOut7_9[3] , \nOut7_9[2] , 
        \nOut7_9[1] , \nOut7_9[0] }), .WestIn({\nOut5_9[7] , \nOut5_9[6] , 
        \nOut5_9[5] , \nOut5_9[4] , \nOut5_9[3] , \nOut5_9[2] , \nOut5_9[1] , 
        \nOut5_9[0] }), .Out({\nOut6_9[7] , \nOut6_9[6] , \nOut6_9[5] , 
        \nOut6_9[4] , \nOut6_9[3] , \nOut6_9[2] , \nOut6_9[1] , \nOut6_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_391 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut392[7] , \nScanOut392[6] , 
        \nScanOut392[5] , \nScanOut392[4] , \nScanOut392[3] , \nScanOut392[2] , 
        \nScanOut392[1] , \nScanOut392[0] }), .ScanOut({\nScanOut391[7] , 
        \nScanOut391[6] , \nScanOut391[5] , \nScanOut391[4] , \nScanOut391[3] , 
        \nScanOut391[2] , \nScanOut391[1] , \nScanOut391[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }), 
        .SouthIn({\nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }), .EastIn(
        {\nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }), .WestIn(
        {\nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }), .Out({
        \nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_410 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut411[7] , \nScanOut411[6] , 
        \nScanOut411[5] , \nScanOut411[4] , \nScanOut411[3] , \nScanOut411[2] , 
        \nScanOut411[1] , \nScanOut411[0] }), .ScanOut({\nScanOut410[7] , 
        \nScanOut410[6] , \nScanOut410[5] , \nScanOut410[4] , \nScanOut410[3] , 
        \nScanOut410[2] , \nScanOut410[1] , \nScanOut410[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_25[7] , \nOut12_25[6] , \nOut12_25[5] , \nOut12_25[4] , 
        \nOut12_25[3] , \nOut12_25[2] , \nOut12_25[1] , \nOut12_25[0] }), 
        .SouthIn({\nOut12_27[7] , \nOut12_27[6] , \nOut12_27[5] , 
        \nOut12_27[4] , \nOut12_27[3] , \nOut12_27[2] , \nOut12_27[1] , 
        \nOut12_27[0] }), .EastIn({\nOut13_26[7] , \nOut13_26[6] , 
        \nOut13_26[5] , \nOut13_26[4] , \nOut13_26[3] , \nOut13_26[2] , 
        \nOut13_26[1] , \nOut13_26[0] }), .WestIn({\nOut11_26[7] , 
        \nOut11_26[6] , \nOut11_26[5] , \nOut11_26[4] , \nOut11_26[3] , 
        \nOut11_26[2] , \nOut11_26[1] , \nOut11_26[0] }), .Out({\nOut12_26[7] , 
        \nOut12_26[6] , \nOut12_26[5] , \nOut12_26[4] , \nOut12_26[3] , 
        \nOut12_26[2] , \nOut12_26[1] , \nOut12_26[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_580 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut581[7] , \nScanOut581[6] , 
        \nScanOut581[5] , \nScanOut581[4] , \nScanOut581[3] , \nScanOut581[2] , 
        \nScanOut581[1] , \nScanOut581[0] }), .ScanOut({\nScanOut580[7] , 
        \nScanOut580[6] , \nScanOut580[5] , \nScanOut580[4] , \nScanOut580[3] , 
        \nScanOut580[2] , \nScanOut580[1] , \nScanOut580[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut18_3[7] , \nOut18_3[6] , \nOut18_3[5] , \nOut18_3[4] , 
        \nOut18_3[3] , \nOut18_3[2] , \nOut18_3[1] , \nOut18_3[0] }), 
        .SouthIn({\nOut18_5[7] , \nOut18_5[6] , \nOut18_5[5] , \nOut18_5[4] , 
        \nOut18_5[3] , \nOut18_5[2] , \nOut18_5[1] , \nOut18_5[0] }), .EastIn(
        {\nOut19_4[7] , \nOut19_4[6] , \nOut19_4[5] , \nOut19_4[4] , 
        \nOut19_4[3] , \nOut19_4[2] , \nOut19_4[1] , \nOut19_4[0] }), .WestIn(
        {\nOut17_4[7] , \nOut17_4[6] , \nOut17_4[5] , \nOut17_4[4] , 
        \nOut17_4[3] , \nOut17_4[2] , \nOut17_4[1] , \nOut17_4[0] }), .Out({
        \nOut18_4[7] , \nOut18_4[6] , \nOut18_4[5] , \nOut18_4[4] , 
        \nOut18_4[3] , \nOut18_4[2] , \nOut18_4[1] , \nOut18_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_226 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut227[7] , \nScanOut227[6] , 
        \nScanOut227[5] , \nScanOut227[4] , \nScanOut227[3] , \nScanOut227[2] , 
        \nScanOut227[1] , \nScanOut227[0] }), .ScanOut({\nScanOut226[7] , 
        \nScanOut226[6] , \nScanOut226[5] , \nScanOut226[4] , \nScanOut226[3] , 
        \nScanOut226[2] , \nScanOut226[1] , \nScanOut226[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_1[7] , \nOut7_1[6] , \nOut7_1[5] , \nOut7_1[4] , \nOut7_1[3] , 
        \nOut7_1[2] , \nOut7_1[1] , \nOut7_1[0] }), .SouthIn({\nOut7_3[7] , 
        \nOut7_3[6] , \nOut7_3[5] , \nOut7_3[4] , \nOut7_3[3] , \nOut7_3[2] , 
        \nOut7_3[1] , \nOut7_3[0] }), .EastIn({\nOut8_2[7] , \nOut8_2[6] , 
        \nOut8_2[5] , \nOut8_2[4] , \nOut8_2[3] , \nOut8_2[2] , \nOut8_2[1] , 
        \nOut8_2[0] }), .WestIn({\nOut6_2[7] , \nOut6_2[6] , \nOut6_2[5] , 
        \nOut6_2[4] , \nOut6_2[3] , \nOut6_2[2] , \nOut6_2[1] , \nOut6_2[0] }), 
        .Out({\nOut7_2[7] , \nOut7_2[6] , \nOut7_2[5] , \nOut7_2[4] , 
        \nOut7_2[3] , \nOut7_2[2] , \nOut7_2[1] , \nOut7_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_862 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut863[7] , \nScanOut863[6] , 
        \nScanOut863[5] , \nScanOut863[4] , \nScanOut863[3] , \nScanOut863[2] , 
        \nScanOut863[1] , \nScanOut863[0] }), .ScanOut({\nScanOut862[7] , 
        \nScanOut862[6] , \nScanOut862[5] , \nScanOut862[4] , \nScanOut862[3] , 
        \nScanOut862[2] , \nScanOut862[1] , \nScanOut862[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_29[7] , \nOut26_29[6] , \nOut26_29[5] , \nOut26_29[4] , 
        \nOut26_29[3] , \nOut26_29[2] , \nOut26_29[1] , \nOut26_29[0] }), 
        .SouthIn({\nOut26_31[7] , \nOut26_31[6] , \nOut26_31[5] , 
        \nOut26_31[4] , \nOut26_31[3] , \nOut26_31[2] , \nOut26_31[1] , 
        \nOut26_31[0] }), .EastIn({\nOut27_30[7] , \nOut27_30[6] , 
        \nOut27_30[5] , \nOut27_30[4] , \nOut27_30[3] , \nOut27_30[2] , 
        \nOut27_30[1] , \nOut27_30[0] }), .WestIn({\nOut25_30[7] , 
        \nOut25_30[6] , \nOut25_30[5] , \nOut25_30[4] , \nOut25_30[3] , 
        \nOut25_30[2] , \nOut25_30[1] , \nOut25_30[0] }), .Out({\nOut26_30[7] , 
        \nOut26_30[6] , \nOut26_30[5] , \nOut26_30[4] , \nOut26_30[3] , 
        \nOut26_30[2] , \nOut26_30[1] , \nOut26_30[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_437 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut438[7] , \nScanOut438[6] , 
        \nScanOut438[5] , \nScanOut438[4] , \nScanOut438[3] , \nScanOut438[2] , 
        \nScanOut438[1] , \nScanOut438[0] }), .ScanOut({\nScanOut437[7] , 
        \nScanOut437[6] , \nScanOut437[5] , \nScanOut437[4] , \nScanOut437[3] , 
        \nScanOut437[2] , \nScanOut437[1] , \nScanOut437[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_20[7] , \nOut13_20[6] , \nOut13_20[5] , \nOut13_20[4] , 
        \nOut13_20[3] , \nOut13_20[2] , \nOut13_20[1] , \nOut13_20[0] }), 
        .SouthIn({\nOut13_22[7] , \nOut13_22[6] , \nOut13_22[5] , 
        \nOut13_22[4] , \nOut13_22[3] , \nOut13_22[2] , \nOut13_22[1] , 
        \nOut13_22[0] }), .EastIn({\nOut14_21[7] , \nOut14_21[6] , 
        \nOut14_21[5] , \nOut14_21[4] , \nOut14_21[3] , \nOut14_21[2] , 
        \nOut14_21[1] , \nOut14_21[0] }), .WestIn({\nOut12_21[7] , 
        \nOut12_21[6] , \nOut12_21[5] , \nOut12_21[4] , \nOut12_21[3] , 
        \nOut12_21[2] , \nOut12_21[1] , \nOut12_21[0] }), .Out({\nOut13_21[7] , 
        \nOut13_21[6] , \nOut13_21[5] , \nOut13_21[4] , \nOut13_21[3] , 
        \nOut13_21[2] , \nOut13_21[1] , \nOut13_21[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_845 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut846[7] , \nScanOut846[6] , 
        \nScanOut846[5] , \nScanOut846[4] , \nScanOut846[3] , \nScanOut846[2] , 
        \nScanOut846[1] , \nScanOut846[0] }), .ScanOut({\nScanOut845[7] , 
        \nScanOut845[6] , \nScanOut845[5] , \nScanOut845[4] , \nScanOut845[3] , 
        \nScanOut845[2] , \nScanOut845[1] , \nScanOut845[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut26_12[7] , \nOut26_12[6] , \nOut26_12[5] , \nOut26_12[4] , 
        \nOut26_12[3] , \nOut26_12[2] , \nOut26_12[1] , \nOut26_12[0] }), 
        .SouthIn({\nOut26_14[7] , \nOut26_14[6] , \nOut26_14[5] , 
        \nOut26_14[4] , \nOut26_14[3] , \nOut26_14[2] , \nOut26_14[1] , 
        \nOut26_14[0] }), .EastIn({\nOut27_13[7] , \nOut27_13[6] , 
        \nOut27_13[5] , \nOut27_13[4] , \nOut27_13[3] , \nOut27_13[2] , 
        \nOut27_13[1] , \nOut27_13[0] }), .WestIn({\nOut25_13[7] , 
        \nOut25_13[6] , \nOut25_13[5] , \nOut25_13[4] , \nOut25_13[3] , 
        \nOut25_13[2] , \nOut25_13[1] , \nOut25_13[0] }), .Out({\nOut26_13[7] , 
        \nOut26_13[6] , \nOut26_13[5] , \nOut26_13[4] , \nOut26_13[3] , 
        \nOut26_13[2] , \nOut26_13[1] , \nOut26_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_697 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut698[7] , \nScanOut698[6] , 
        \nScanOut698[5] , \nScanOut698[4] , \nScanOut698[3] , \nScanOut698[2] , 
        \nScanOut698[1] , \nScanOut698[0] }), .ScanOut({\nScanOut697[7] , 
        \nScanOut697[6] , \nScanOut697[5] , \nScanOut697[4] , \nScanOut697[3] , 
        \nScanOut697[2] , \nScanOut697[1] , \nScanOut697[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut21_24[7] , \nOut21_24[6] , \nOut21_24[5] , \nOut21_24[4] , 
        \nOut21_24[3] , \nOut21_24[2] , \nOut21_24[1] , \nOut21_24[0] }), 
        .SouthIn({\nOut21_26[7] , \nOut21_26[6] , \nOut21_26[5] , 
        \nOut21_26[4] , \nOut21_26[3] , \nOut21_26[2] , \nOut21_26[1] , 
        \nOut21_26[0] }), .EastIn({\nOut22_25[7] , \nOut22_25[6] , 
        \nOut22_25[5] , \nOut22_25[4] , \nOut22_25[3] , \nOut22_25[2] , 
        \nOut22_25[1] , \nOut22_25[0] }), .WestIn({\nOut20_25[7] , 
        \nOut20_25[6] , \nOut20_25[5] , \nOut20_25[4] , \nOut20_25[3] , 
        \nOut20_25[2] , \nOut20_25[1] , \nOut20_25[0] }), .Out({\nOut21_25[7] , 
        \nOut21_25[6] , \nOut21_25[5] , \nOut21_25[4] , \nOut21_25[3] , 
        \nOut21_25[2] , \nOut21_25[1] , \nOut21_25[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_707 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut708[7] , \nScanOut708[6] , 
        \nScanOut708[5] , \nScanOut708[4] , \nScanOut708[3] , \nScanOut708[2] , 
        \nScanOut708[1] , \nScanOut708[0] }), .ScanOut({\nScanOut707[7] , 
        \nScanOut707[6] , \nScanOut707[5] , \nScanOut707[4] , \nScanOut707[3] , 
        \nScanOut707[2] , \nScanOut707[1] , \nScanOut707[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut22_2[7] , \nOut22_2[6] , \nOut22_2[5] , \nOut22_2[4] , 
        \nOut22_2[3] , \nOut22_2[2] , \nOut22_2[1] , \nOut22_2[0] }), 
        .SouthIn({\nOut22_4[7] , \nOut22_4[6] , \nOut22_4[5] , \nOut22_4[4] , 
        \nOut22_4[3] , \nOut22_4[2] , \nOut22_4[1] , \nOut22_4[0] }), .EastIn(
        {\nOut23_3[7] , \nOut23_3[6] , \nOut23_3[5] , \nOut23_3[4] , 
        \nOut23_3[3] , \nOut23_3[2] , \nOut23_3[1] , \nOut23_3[0] }), .WestIn(
        {\nOut21_3[7] , \nOut21_3[6] , \nOut21_3[5] , \nOut21_3[4] , 
        \nOut21_3[3] , \nOut21_3[2] , \nOut21_3[1] , \nOut21_3[0] }), .Out({
        \nOut22_3[7] , \nOut22_3[6] , \nOut22_3[5] , \nOut22_3[4] , 
        \nOut22_3[3] , \nOut22_3[2] , \nOut22_3[1] , \nOut22_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1001 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1002[7] , \nScanOut1002[6] , 
        \nScanOut1002[5] , \nScanOut1002[4] , \nScanOut1002[3] , 
        \nScanOut1002[2] , \nScanOut1002[1] , \nScanOut1002[0] }), .ScanOut({
        \nScanOut1001[7] , \nScanOut1001[6] , \nScanOut1001[5] , 
        \nScanOut1001[4] , \nScanOut1001[3] , \nScanOut1001[2] , 
        \nScanOut1001[1] , \nScanOut1001[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Out({\nOut31_9[7] , \nOut31_9[6] , \nOut31_9[5] , 
        \nOut31_9[4] , \nOut31_9[3] , \nOut31_9[2] , \nOut31_9[1] , 
        \nOut31_9[0] }) );
endmodule

