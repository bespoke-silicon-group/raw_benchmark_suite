
module BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, Out, Enable1, Enable2, In1, In2
     );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] In1;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In2;
input  Clk, Reset, RD, WR, ScanEnable, Enable1, Enable2;
    wire \ScanOut[31] , n288, \ScanOut[5]1 , \ScanOut[4]1 , n245, n287, n262, 
        n279, n217, n230, \ScanOut[10]1 , n302, n222, n305, n257, n270, n295, 
        n239, n292, \ScanOut[23]1 , \ScanOut[8]1 , n219, n225, n250, n277, 
        n289, n237, n259, \ScanOut[22]1 , \ScanOut[11]1 , n265, n242, 
        \ScanOut[9]1 , n310, n280, n224, n276, n303, n251, n293, 
        \ScanOut[19]1 , n218, n311, n281, \ScanOut[26]1 , \ScanOut[18]1 , 
        \ScanOut[1]1 , n264, \ScanOut[0]1 , n243, n258, \ScanOut[15]1 , n236, 
        n216, n231, n278, \ScanOut[27]1 , n244, \ScanOut[14]1 , n263, n316, 
        n286, n304, n294, n271, n238, n256, n223, n233, n228, n314, n284, n214, 
        n246, n261, \ScanOut[28]1 , n221, \ScanOut[3]1 , n268, \ScanOut[30]1 , 
        \ScanOut[29]1 , \ScanOut[2]1 , n254, n273, n306, n296, n301, n291, 
        \ScanOut[25]1 , \ScanOut[24]1 , \ScanOut[17]1 , n253, n248, n274, 
        \ScanOut[16]1 , n226, n234, n308, n298, n241, n313, n266, n283, 
        \ScanOut[6]1 , n227, n249, \ScanOut[7]1 , n312, n300, n252, n290, n275, 
        n282, n215, n309, n235, n240, n267, n299, \ScanOut[13]1 , n232, n247, 
        n260, \ScanOut[21]1 , n315, n285, n229, n307, n297, \ScanOut[12]1 , 
        n272, n255, n269, \ScanOut[20]1 , n220;
    assign ScanOut[31] = \ScanOut[31] ;
    assign ScanOut[30] = \ScanOut[30]1 ;
    assign ScanOut[29] = \ScanOut[29]1 ;
    assign ScanOut[28] = \ScanOut[28]1 ;
    assign ScanOut[27] = \ScanOut[27]1 ;
    assign ScanOut[26] = \ScanOut[26]1 ;
    assign ScanOut[25] = \ScanOut[25]1 ;
    assign ScanOut[24] = \ScanOut[24]1 ;
    assign ScanOut[23] = \ScanOut[23]1 ;
    assign ScanOut[22] = \ScanOut[22]1 ;
    assign ScanOut[21] = \ScanOut[21]1 ;
    assign ScanOut[20] = \ScanOut[20]1 ;
    assign ScanOut[19] = \ScanOut[19]1 ;
    assign ScanOut[18] = \ScanOut[18]1 ;
    assign ScanOut[17] = \ScanOut[17]1 ;
    assign ScanOut[16] = \ScanOut[16]1 ;
    assign ScanOut[15] = \ScanOut[15]1 ;
    assign ScanOut[14] = \ScanOut[14]1 ;
    assign ScanOut[13] = \ScanOut[13]1 ;
    assign ScanOut[12] = \ScanOut[12]1 ;
    assign ScanOut[11] = \ScanOut[11]1 ;
    assign ScanOut[10] = \ScanOut[10]1 ;
    assign ScanOut[9] = \ScanOut[9]1 ;
    assign ScanOut[8] = \ScanOut[8]1 ;
    assign ScanOut[7] = \ScanOut[7]1 ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[31] = \ScanOut[31] ;
    assign Out[30] = \ScanOut[30]1 ;
    assign Out[29] = \ScanOut[29]1 ;
    assign Out[28] = \ScanOut[28]1 ;
    assign Out[27] = \ScanOut[27]1 ;
    assign Out[26] = \ScanOut[26]1 ;
    assign Out[25] = \ScanOut[25]1 ;
    assign Out[24] = \ScanOut[24]1 ;
    assign Out[23] = \ScanOut[23]1 ;
    assign Out[22] = \ScanOut[22]1 ;
    assign Out[21] = \ScanOut[21]1 ;
    assign Out[20] = \ScanOut[20]1 ;
    assign Out[19] = \ScanOut[19]1 ;
    assign Out[18] = \ScanOut[18]1 ;
    assign Out[17] = \ScanOut[17]1 ;
    assign Out[16] = \ScanOut[16]1 ;
    assign Out[15] = \ScanOut[15]1 ;
    assign Out[14] = \ScanOut[14]1 ;
    assign Out[13] = \ScanOut[13]1 ;
    assign Out[12] = \ScanOut[12]1 ;
    assign Out[11] = \ScanOut[11]1 ;
    assign Out[10] = \ScanOut[10]1 ;
    assign Out[9] = \ScanOut[9]1 ;
    assign Out[8] = \ScanOut[8]1 ;
    assign Out[7] = \ScanOut[7]1 ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_OR2 U54 ( .A(n258), .B(n259), .Z(n294) );
    VMW_AO22 U73 ( .A(In1[7]), .B(n281), .C(In2[7]), .D(n280), .Z(n228) );
    VMW_AO22 U113 ( .A(In1[18]), .B(n281), .C(In2[18]), .D(n280), .Z(n250) );
    VMW_INV U134 ( .A(Enable1), .Z(n282) );
    VMW_NOR4 U68 ( .A(Enable1), .B(Enable2), .C(ScanEnable), .D(Reset), .Z(
        n279) );
    VMW_AO22 U96 ( .A(\ScanOut[26]1 ), .B(n279), .C(ScanIn[26]), .D(n283), .Z(
        n267) );
    VMW_AO22 U108 ( .A(\ScanOut[20]1 ), .B(n279), .C(ScanIn[20]), .D(n283), 
        .Z(n255) );
    VMW_OR2 U33 ( .A(n216), .B(n217), .Z(n315) );
    VMW_OR2 U34 ( .A(n218), .B(n219), .Z(n314) );
    VMW_OR2 U41 ( .A(n232), .B(n233), .Z(n307) );
    VMW_OR2 U46 ( .A(n242), .B(n243), .Z(n302) );
    VMW_OR2 U61 ( .A(n272), .B(n273), .Z(n287) );
    VMW_AO22 U84 ( .A(\ScanOut[31] ), .B(n279), .C(ScanIn[31]), .D(n283), .Z(
        n277) );
    VMW_AO22 U101 ( .A(In1[23]), .B(n281), .C(In2[23]), .D(n280), .Z(n260) );
    VMW_AO22 U126 ( .A(\ScanOut[12]1 ), .B(n279), .C(ScanIn[12]), .D(n283), 
        .Z(n239) );
    VMW_NOR2 U66 ( .A(n278), .B(n282), .Z(n281) );
    VMW_AO22 U106 ( .A(\ScanOut[21]1 ), .B(n279), .C(ScanIn[21]), .D(n283), 
        .Z(n257) );
    VMW_AO22 U121 ( .A(In1[14]), .B(n281), .C(In2[14]), .D(n280), .Z(n242) );
    VMW_AO22 U83 ( .A(In1[31]), .B(n281), .C(In2[31]), .D(n280), .Z(n276) );
    VMW_AO22 U98 ( .A(\ScanOut[25]1 ), .B(n279), .C(ScanIn[25]), .D(n283), .Z(
        n265) );
    VMW_OR2 U35 ( .A(n220), .B(n221), .Z(n313) );
    VMW_OR2 U48 ( .A(n246), .B(n247), .Z(n300) );
    VMW_AO22 U128 ( .A(\ScanOut[11]1 ), .B(n279), .C(ScanIn[11]), .D(n283), 
        .Z(n237) );
    VMW_OR2 U53 ( .A(n256), .B(n257), .Z(n295) );
    VMW_AO22 U91 ( .A(In1[28]), .B(n281), .C(In2[28]), .D(n280), .Z(n270) );
    VMW_AO22 U74 ( .A(\ScanOut[7]1 ), .B(n279), .C(ScanIn[7]), .D(n283), .Z(
        n229) );
    VMW_AO22 U114 ( .A(\ScanOut[18]1 ), .B(n279), .C(ScanIn[18]), .D(n283), 
        .Z(n251) );
    VMW_INV U133 ( .A(ScanEnable), .Z(n284) );
    VMW_AO22 U99 ( .A(In1[24]), .B(n281), .C(In2[24]), .D(n280), .Z(n262) );
    VMW_FD \Out_reg[25]  ( .D(n291), .CP(Clk), .Q(\ScanOut[25]1 ) );
    VMW_FD \Out_reg[16]  ( .D(n300), .CP(Clk), .Q(\ScanOut[16]1 ) );
    VMW_OR2 U32 ( .A(n214), .B(n215), .Z(n316) );
    VMW_OR2 U40 ( .A(n230), .B(n231), .Z(n308) );
    VMW_AO22 U82 ( .A(\ScanOut[3]1 ), .B(n279), .C(ScanIn[3]), .D(n283), .Z(
        n221) );
    VMW_FD \Out_reg[5]  ( .D(n311), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_OR2 U47 ( .A(n244), .B(n245), .Z(n301) );
    VMW_OR2 U49 ( .A(n248), .B(n249), .Z(n299) );
    VMW_OR2 U52 ( .A(n254), .B(n255), .Z(n296) );
    VMW_NOR2 U67 ( .A(n284), .B(Reset), .Z(n283) );
    VMW_AO22 U107 ( .A(In1[20]), .B(n281), .C(In2[20]), .D(n280), .Z(n254) );
    VMW_AO22 U120 ( .A(\ScanOut[15]1 ), .B(n279), .C(ScanIn[15]), .D(n283), 
        .Z(n245) );
    VMW_AO22 U75 ( .A(In1[6]), .B(n281), .C(In2[6]), .D(n280), .Z(n226) );
    VMW_AO22 U115 ( .A(In1[17]), .B(n281), .C(In2[17]), .D(n280), .Z(n248) );
    VMW_AO22 U132 ( .A(\ScanOut[0]1 ), .B(n279), .C(ScanIn[0]), .D(n283), .Z(
        n215) );
    VMW_FD \Out_reg[12]  ( .D(n304), .CP(Clk), .Q(\ScanOut[12]1 ) );
    VMW_AO22 U90 ( .A(\ScanOut[29]1 ), .B(n279), .C(ScanIn[29]), .D(n283), .Z(
        n273) );
    VMW_FD \Out_reg[21]  ( .D(n295), .CP(Clk), .Q(\ScanOut[21]1 ) );
    VMW_AO22 U129 ( .A(In1[10]), .B(n281), .C(In2[10]), .D(n280), .Z(n234) );
    VMW_FD \Out_reg[31]  ( .D(n285), .CP(Clk), .Q(\ScanOut[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n288), .CP(Clk), .Q(\ScanOut[28]1 ) );
    VMW_FD \Out_reg[8]  ( .D(n308), .CP(Clk), .Q(\ScanOut[8]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n315), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_OR2 U55 ( .A(n260), .B(n261), .Z(n293) );
    VMW_AO22 U69 ( .A(In1[9]), .B(n281), .C(In2[9]), .D(n280), .Z(n232) );
    VMW_AO22 U109 ( .A(In1[1]), .B(n281), .C(In2[1]), .D(n280), .Z(n216) );
    VMW_FD \Out_reg[19]  ( .D(n297), .CP(Clk), .Q(\ScanOut[19]1 ) );
    VMW_AO22 U72 ( .A(\ScanOut[8]1 ), .B(n279), .C(ScanIn[8]), .D(n283), .Z(
        n231) );
    VMW_AO22 U97 ( .A(In1[25]), .B(n281), .C(In2[25]), .D(n280), .Z(n264) );
    VMW_FD \Out_reg[3]  ( .D(n313), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_AO22 U112 ( .A(\ScanOut[19]1 ), .B(n279), .C(ScanIn[19]), .D(n283), 
        .Z(n253) );
    VMW_FD \Out_reg[23]  ( .D(n293), .CP(Clk), .Q(\ScanOut[23]1 ) );
    VMW_FD \Out_reg[10]  ( .D(n306), .CP(Clk), .Q(\ScanOut[10]1 ) );
    VMW_OR2 U60 ( .A(n270), .B(n271), .Z(n288) );
    VMW_FD \Out_reg[7]  ( .D(n309), .CP(Clk), .Q(\ScanOut[7]1 ) );
    VMW_AO22 U100 ( .A(\ScanOut[24]1 ), .B(n279), .C(ScanIn[24]), .D(n283), 
        .Z(n263) );
    VMW_AO22 U127 ( .A(In1[11]), .B(n281), .C(In2[11]), .D(n280), .Z(n236) );
    VMW_AO22 U85 ( .A(In1[30]), .B(n281), .C(In2[30]), .D(n280), .Z(n274) );
    VMW_FD \Out_reg[27]  ( .D(n289), .CP(Clk), .Q(\ScanOut[27]1 ) );
    VMW_FD \Out_reg[14]  ( .D(n302), .CP(Clk), .Q(\ScanOut[14]1 ) );
    VMW_OR2 U36 ( .A(n222), .B(n223), .Z(n312) );
    VMW_OR2 U37 ( .A(n224), .B(n225), .Z(n311) );
    VMW_OR2 U39 ( .A(n228), .B(n229), .Z(n309) );
    VMW_OR2 U57 ( .A(n264), .B(n265), .Z(n291) );
    VMW_FD \Out_reg[6]  ( .D(n310), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U70 ( .A(\ScanOut[9]1 ), .B(n279), .C(ScanIn[9]), .D(n283), .Z(
        n233) );
    VMW_AO22 U110 ( .A(\ScanOut[1]1 ), .B(n279), .C(ScanIn[1]), .D(n283), .Z(
        n217) );
    VMW_OR2 U42 ( .A(n234), .B(n235), .Z(n306) );
    VMW_OR2 U45 ( .A(n240), .B(n241), .Z(n303) );
    VMW_AO22 U79 ( .A(In1[4]), .B(n281), .C(In2[4]), .D(n280), .Z(n222) );
    VMW_AO22 U95 ( .A(In1[26]), .B(n281), .C(In2[26]), .D(n280), .Z(n266) );
    VMW_AO22 U119 ( .A(In1[15]), .B(n281), .C(In2[15]), .D(n280), .Z(n244) );
    VMW_FD \Out_reg[26]  ( .D(n290), .CP(Clk), .Q(\ScanOut[26]1 ) );
    VMW_FD \Out_reg[15]  ( .D(n301), .CP(Clk), .Q(\ScanOut[15]1 ) );
    VMW_FD \Out_reg[18]  ( .D(n298), .CP(Clk), .Q(\ScanOut[18]1 ) );
    VMW_AO22 U87 ( .A(In1[2]), .B(n281), .C(In2[2]), .D(n280), .Z(n218) );
    VMW_FD \Out_reg[2]  ( .D(n314), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_AO22 U125 ( .A(In1[12]), .B(n281), .C(In2[12]), .D(n280), .Z(n238) );
    VMW_FD \Out_reg[11]  ( .D(n305), .CP(Clk), .Q(\ScanOut[11]1 ) );
    VMW_OR2 U62 ( .A(n274), .B(n275), .Z(n286) );
    VMW_FD \Out_reg[22]  ( .D(n294), .CP(Clk), .Q(\ScanOut[22]1 ) );
    VMW_NOR2 U65 ( .A(Enable1), .B(n278), .Z(n280) );
    VMW_AO22 U102 ( .A(\ScanOut[23]1 ), .B(n279), .C(ScanIn[23]), .D(n283), 
        .Z(n261) );
    VMW_AO22 U105 ( .A(In1[21]), .B(n281), .C(In2[21]), .D(n280), .Z(n256) );
    VMW_FD \Out_reg[20]  ( .D(n296), .CP(Clk), .Q(\ScanOut[20]1 ) );
    VMW_FD \Out_reg[13]  ( .D(n303), .CP(Clk), .Q(\ScanOut[13]1 ) );
    VMW_AO22 U80 ( .A(\ScanOut[4]1 ), .B(n279), .C(ScanIn[4]), .D(n283), .Z(
        n223) );
    VMW_AO22 U122 ( .A(\ScanOut[14]1 ), .B(n279), .C(ScanIn[14]), .D(n283), 
        .Z(n243) );
    VMW_FD \Out_reg[9]  ( .D(n307), .CP(Clk), .Q(\ScanOut[9]1 ) );
    VMW_OR2 U50 ( .A(n250), .B(n251), .Z(n298) );
    VMW_OR2 U59 ( .A(n268), .B(n269), .Z(n289) );
    VMW_FD \Out_reg[30]  ( .D(n286), .CP(Clk), .Q(\ScanOut[30]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n316), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_FD \Out_reg[29]  ( .D(n287), .CP(Clk), .Q(\ScanOut[29]1 ) );
    VMW_AO22 U77 ( .A(In1[5]), .B(n281), .C(In2[5]), .D(n280), .Z(n224) );
    VMW_AO22 U89 ( .A(In1[29]), .B(n281), .C(In2[29]), .D(n280), .Z(n272) );
    VMW_AO22 U92 ( .A(\ScanOut[28]1 ), .B(n279), .C(ScanIn[28]), .D(n283), .Z(
        n271) );
    VMW_FD \Out_reg[24]  ( .D(n292), .CP(Clk), .Q(\ScanOut[24]1 ) );
    VMW_FD \Out_reg[17]  ( .D(n299), .CP(Clk), .Q(\ScanOut[17]1 ) );
    VMW_AO22 U117 ( .A(In1[16]), .B(n281), .C(In2[16]), .D(n280), .Z(n246) );
    VMW_FD \Out_reg[4]  ( .D(n312), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_OR2 U58 ( .A(n266), .B(n267), .Z(n290) );
    VMW_AO22 U130 ( .A(\ScanOut[10]1 ), .B(n279), .C(ScanIn[10]), .D(n283), 
        .Z(n235) );
    VMW_OR2 U38 ( .A(n226), .B(n227), .Z(n310) );
    VMW_OR2 U43 ( .A(n236), .B(n237), .Z(n305) );
    VMW_OR3 U64 ( .A(Reset), .B(ScanEnable), .C(n279), .Z(n278) );
    VMW_AO22 U81 ( .A(In1[3]), .B(n281), .C(In2[3]), .D(n280), .Z(n220) );
    VMW_AO22 U104 ( .A(\ScanOut[22]1 ), .B(n279), .C(ScanIn[22]), .D(n283), 
        .Z(n259) );
    VMW_OR2 U51 ( .A(n252), .B(n253), .Z(n297) );
    VMW_AO22 U76 ( .A(\ScanOut[6]1 ), .B(n279), .C(ScanIn[6]), .D(n283), .Z(
        n227) );
    VMW_AO22 U116 ( .A(\ScanOut[17]1 ), .B(n279), .C(ScanIn[17]), .D(n283), 
        .Z(n249) );
    VMW_AO22 U123 ( .A(In1[13]), .B(n281), .C(In2[13]), .D(n280), .Z(n240) );
    VMW_AO22 U88 ( .A(\ScanOut[2]1 ), .B(n279), .C(ScanIn[2]), .D(n283), .Z(
        n219) );
    VMW_AO22 U93 ( .A(In1[27]), .B(n281), .C(In2[27]), .D(n280), .Z(n268) );
    VMW_AO22 U131 ( .A(In1[0]), .B(n281), .C(In2[0]), .D(n280), .Z(n214) );
    VMW_OR2 U44 ( .A(n238), .B(n239), .Z(n304) );
    VMW_OR2 U56 ( .A(n262), .B(n263), .Z(n292) );
    VMW_AO22 U94 ( .A(\ScanOut[27]1 ), .B(n279), .C(ScanIn[27]), .D(n283), .Z(
        n269) );
    VMW_AO22 U71 ( .A(In1[8]), .B(n281), .C(In2[8]), .D(n280), .Z(n230) );
    VMW_AO22 U111 ( .A(In1[19]), .B(n281), .C(In2[19]), .D(n280), .Z(n252) );
    VMW_AO22 U124 ( .A(\ScanOut[13]1 ), .B(n279), .C(ScanIn[13]), .D(n283), 
        .Z(n241) );
    VMW_OR2 U63 ( .A(n276), .B(n277), .Z(n285) );
    VMW_AO22 U78 ( .A(\ScanOut[5]1 ), .B(n279), .C(ScanIn[5]), .D(n283), .Z(
        n225) );
    VMW_AO22 U86 ( .A(\ScanOut[30]1 ), .B(n279), .C(ScanIn[30]), .D(n283), .Z(
        n275) );
    VMW_AO22 U103 ( .A(In1[22]), .B(n281), .C(In2[22]), .D(n280), .Z(n258) );
    VMW_AO22 U118 ( .A(\ScanOut[16]1 ), .B(n279), .C(ScanIn[16]), .D(n283), 
        .Z(n247) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_3 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n112, n32, n29, n85, n47, n60, n109, 
        n40, n67, n82, n99, n27, n35, n49, n115, n107, n52, n75, n114, n34, 
        n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, n21, n46, n54, 
        n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, n113, n118, n94, 
        n23, n103, n16, n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, n58, 
        n116, n104, n18, n24, n88, n37, n51, n93, n59, n76, n117, n80, n42, 
        n65, n19, n50, n77, n89, n25, n102, n105, n22, n39, n95, n45, n57, n70, 
        n62, n87, n17, n30, n79, n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_OR2 U54 ( .A(B[26]), .B(n99), .Z(n103) );
    VMW_INV U73 ( .A(B[27]), .Z(n109) );
    VMW_INV U96 ( .A(B[31]), .Z(n15) );
    VMW_INV U68 ( .A(A[30]), .Z(n117) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n66), .C(n62), .D(n57), .Z(n65) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U34 ( .A(B[16]), .B(n64), .Z(n67) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n75), .D(n70), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_NAND2 U61 ( .A(n114), .B(A[29]), .Z(n115) );
    VMW_INV U84 ( .A(B[15]), .Z(n66) );
    VMW_INV U101 ( .A(A[6]), .Z(n32) );
    VMW_INV U66 ( .A(B[7]), .Z(n41) );
    VMW_INV U83 ( .A(A[15]), .Z(n69) );
    VMW_INV U98 ( .A(B[13]), .Z(n60) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_NAND2 U48 ( .A(n91), .B(B[24]), .Z(n89) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n69), .C(n67), .D(n65), .Z(n68) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n102), .C(n96), .D(n89), .Z(n101) );
    VMW_INV U91 ( .A(B[11]), .Z(n54) );
    VMW_INV U74 ( .A(A[3]), .Z(n30) );
    VMW_INV U99 ( .A(A[26]), .Z(n99) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U40 ( .A(n78), .B(B[20]), .Z(n77) );
    VMW_INV U82 ( .A(B[29]), .Z(n114) );
    VMW_NAND2 U52 ( .A(n99), .B(B[26]), .Z(n97) );
    VMW_INV U67 ( .A(A[7]), .Z(n44) );
    VMW_INV U75 ( .A(B[3]), .Z(n27) );
    VMW_INV U90 ( .A(A[14]), .Z(n58) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n94), .C(n88), .D(n83), .Z(n93) );
    VMW_INV U69 ( .A(B[17]), .Z(n73) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n105), .C(n103), .D(n101), .Z(n104) );
    VMW_INV U72 ( .A(A[27]), .Z(n112) );
    VMW_INV U97 ( .A(A[16]), .Z(n64) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n114), .C(n111), .D(n106), .Z(n113) );
    VMW_INV U100 ( .A(B[23]), .Z(n94) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_INV U85 ( .A(A[4]), .Z(n25) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_NAND2 U32 ( .A(n64), .B(B[16]), .Z(n63) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n76), .C(n74), .D(n72), .Z(n75) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n109), .C(n104), .D(n97), .Z(n108) );
    VMW_INV U70 ( .A(A[17]), .Z(n76) );
    VMW_INV U95 ( .A(A[1]), .Z(n21) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_INV U79 ( .A(B[19]), .Z(n80) );
    VMW_INV U87 ( .A(A[8]), .Z(n39) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n77), .Z(n85) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n117), .C(n115), .D(n113), .Z(n116) );
    VMW_INV U65 ( .A(A[12]), .Z(n52) );
    VMW_INV U102 ( .A(A[2]), .Z(n18) );
    VMW_INV U80 ( .A(A[10]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n73), .C(n68), .D(n63), .Z(n72) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n112), .C(n110), .D(n108), .Z(n111) );
    VMW_INV U89 ( .A(A[18]), .Z(n71) );
    VMW_NAND2 U50 ( .A(n94), .B(A[23]), .Z(n95) );
    VMW_INV U77 ( .A(A[25]), .Z(n105) );
    VMW_INV U92 ( .A(A[28]), .Z(n107) );
    VMW_OR2 U58 ( .A(B[28]), .B(n107), .Z(n110) );
    VMW_NAND2 U36 ( .A(n71), .B(B[18]), .Z(n70) );
    VMW_INV U81 ( .A(B[9]), .Z(n48) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n78), .C(n81), .D(n79), .Z(n82) );
    VMW_AO22 U64 ( .A(n116), .B(n118), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n91), .C(n95), .D(n93), .Z(n96) );
    VMW_INV U76 ( .A(B[25]), .Z(n102) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_INV U88 ( .A(B[21]), .Z(n86) );
    VMW_INV U93 ( .A(A[5]), .Z(n37) );
    VMW_OR2 U38 ( .A(B[18]), .B(n71), .Z(n74) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n107), .B(B[28]), .Z(n106) );
    VMW_INV U94 ( .A(B[5]), .Z(n34) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_NAND2 U63 ( .A(n117), .B(B[30]), .Z(n118) );
    VMW_INV U86 ( .A(A[24]), .Z(n91) );
    VMW_INV U103 ( .A(A[0]), .Z(n20) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_INV U78 ( .A(A[20]), .Z(n78) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_2 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n190, n149, n152, n175, n127, n217, n135, n205, n199, n140, n167, 
        n182, n120, n129, n185, n147, n160, n132, n202, n169, n210, n155, n172, 
        n197, n133, n203, n146, n161, n121, n128, n184, n218, n154, n196, n168, 
        n173, n211, n216, n126, n148, n153, n174, n183, n191, n166, n141, n134, 
        n204, n151, n193, n198, n176, n124, n214, n188, n206, n136, n143, n158, 
        n144, n164, n163, n181, n186, n178, n123, n131, n201, n213, n171, n156, 
        n130, n138, n194, n208, n179, n200, n145, n162, n187, n195, n122, n139, 
        n209, n170, n157, n125, n212, n215, n189, n150, n177, n192, n119, n142, 
        n180, n165, n159, n137, n207;
    VMW_OAI21 U3 ( .A(A[31]), .B(n119), .C(n120), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n124), .B(B[0]), .C(n125), .D(B[1]), .Z(n123) );
    VMW_OR2 U6 ( .A(B[2]), .B(n122), .Z(n126) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n152), .C(n147), .D(n142), .Z(n151) );
    VMW_OR2 U54 ( .A(B[26]), .B(n200), .Z(n203) );
    VMW_INV U73 ( .A(B[27]), .Z(n209) );
    VMW_INV U96 ( .A(B[31]), .Z(n119) );
    VMW_INV U68 ( .A(A[30]), .Z(n217) );
    VMW_NAND2 U28 ( .A(n162), .B(B[14]), .Z(n161) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n170), .C(n166), .D(n161), .Z(n169) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n125), .C(n126), .D(n123), .Z(n127) );
    VMW_NAND2 U8 ( .A(n129), .B(B[4]), .Z(n128) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n133), .D(n128), .Z(n137) );
    VMW_OR2 U34 ( .A(B[16]), .B(n168), .Z(n171) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n184), .C(n179), .D(n174), .Z(n183) );
    VMW_NAND2 U46 ( .A(n190), .B(A[21]), .Z(n191) );
    VMW_NAND2 U61 ( .A(n214), .B(A[29]), .Z(n215) );
    VMW_INV U84 ( .A(B[15]), .Z(n170) );
    VMW_INV U101 ( .A(A[6]), .Z(n136) );
    VMW_INV U66 ( .A(B[7]), .Z(n145) );
    VMW_INV U83 ( .A(A[15]), .Z(n173) );
    VMW_INV U98 ( .A(B[13]), .Z(n164) );
    VMW_NAND2 U26 ( .A(n158), .B(A[11]), .Z(n159) );
    VMW_NAND2 U48 ( .A(n194), .B(B[24]), .Z(n193) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n131), .C(n127), .D(n121), .Z(n130) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n173), .C(n171), .D(n169), .Z(n172) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n202), .C(n198), .D(n193), .Z(n201) );
    VMW_INV U91 ( .A(B[11]), .Z(n158) );
    VMW_INV U74 ( .A(A[3]), .Z(n134) );
    VMW_INV U99 ( .A(A[26]), .Z(n200) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_NAND2 U40 ( .A(n182), .B(B[20]), .Z(n181) );
    VMW_INV U82 ( .A(B[29]), .Z(n214) );
    VMW_NAND2 U52 ( .A(n200), .B(B[26]), .Z(n199) );
    VMW_INV U67 ( .A(A[7]), .Z(n148) );
    VMW_INV U75 ( .A(B[3]), .Z(n131) );
    VMW_INV U90 ( .A(A[14]), .Z(n162) );
    VMW_NAND2 U20 ( .A(n150), .B(B[10]), .Z(n149) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n196), .C(n192), .D(n187), .Z(n195) );
    VMW_INV U69 ( .A(B[17]), .Z(n177) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n188), .C(n191), .D(n189), .Z(n192) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n205), .C(n203), .D(n201), .Z(n204) );
    VMW_INV U72 ( .A(A[27]), .Z(n212) );
    VMW_INV U97 ( .A(A[16]), .Z(n168) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n214), .C(n211), .D(n206), .Z(n213) );
    VMW_INV U100 ( .A(B[23]), .Z(n196) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_INV U85 ( .A(A[4]), .Z(n129) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n145), .C(n140), .D(n135), .Z(n144) );
    VMW_NAND2 U22 ( .A(n152), .B(A[9]), .Z(n153) );
    VMW_NAND2 U32 ( .A(n168), .B(B[16]), .Z(n167) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n180), .C(n178), .D(n176), .Z(n179) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n209), .C(n204), .D(n199), .Z(n208) );
    VMW_INV U70 ( .A(A[17]), .Z(n180) );
    VMW_INV U95 ( .A(A[1]), .Z(n125) );
    VMW_NAND2 U30 ( .A(n164), .B(A[13]), .Z(n165) );
    VMW_INV U79 ( .A(B[19]), .Z(n184) );
    VMW_INV U87 ( .A(A[8]), .Z(n143) );
    VMW_OR2 U10 ( .A(B[4]), .B(n129), .Z(n132) );
    VMW_NAND2 U42 ( .A(n184), .B(A[19]), .Z(n185) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n190), .C(n186), .D(n181), .Z(n189) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n217), .C(n215), .D(n213), .Z(n216) );
    VMW_INV U65 ( .A(A[12]), .Z(n156) );
    VMW_INV U102 ( .A(A[2]), .Z(n122) );
    VMW_INV U80 ( .A(A[10]), .Z(n150) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n134), .C(n132), .D(n130), .Z(n133) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n148), .C(n146), .D(n144), .Z(n147) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n177), .C(n172), .D(n167), .Z(n176) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n212), .C(n210), .D(n208), .Z(n211) );
    VMW_INV U89 ( .A(A[18]), .Z(n175) );
    VMW_NAND2 U50 ( .A(n196), .B(A[23]), .Z(n197) );
    VMW_INV U77 ( .A(A[25]), .Z(n205) );
    VMW_INV U92 ( .A(A[28]), .Z(n207) );
    VMW_OR2 U58 ( .A(B[28]), .B(n207), .Z(n210) );
    VMW_NAND2 U36 ( .A(n175), .B(B[18]), .Z(n174) );
    VMW_INV U81 ( .A(B[9]), .Z(n152) );
    VMW_NAND2 U4 ( .A(n122), .B(B[2]), .Z(n121) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n146) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n182), .C(n185), .D(n183), .Z(n186) );
    VMW_AO22 U64 ( .A(n216), .B(n218), .C(A[31]), .D(n119), .Z(n120) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n194), .C(n197), .D(n195), .Z(n198) );
    VMW_INV U76 ( .A(B[25]), .Z(n202) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U24 ( .A(n156), .B(B[12]), .Z(n155) );
    VMW_INV U88 ( .A(B[21]), .Z(n190) );
    VMW_INV U93 ( .A(A[5]), .Z(n141) );
    VMW_OR2 U38 ( .A(B[18]), .B(n175), .Z(n178) );
    VMW_NAND2 U44 ( .A(n188), .B(B[22]), .Z(n187) );
    VMW_NAND2 U56 ( .A(n207), .B(B[28]), .Z(n206) );
    VMW_INV U94 ( .A(B[5]), .Z(n138) );
    VMW_INV U71 ( .A(A[22]), .Z(n188) );
    VMW_NAND2 U63 ( .A(n217), .B(B[30]), .Z(n218) );
    VMW_INV U86 ( .A(A[24]), .Z(n194) );
    VMW_INV U103 ( .A(A[0]), .Z(n124) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n162), .C(n165), .D(n163), .Z(n166) );
    VMW_INV U78 ( .A(A[20]), .Z(n182) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n287, n317, n245, n262, n279, n222, n230, n257, n270, n239, n295, 
        n305, n219, n292, n302, n250, n277, n225, n237, n289, n259, n265, n242, 
        n280, n310, n224, n288, n318, n276, n236, n243, n251, n264, n281, n293, 
        n303, n311, n258, n231, n238, n244, n278, n263, n286, n316, n294, n304, 
        n256, n271, n223, n228, n284, n314, n261, n246, n233, n221, n248, n253, 
        n254, n268, n273, n291, n296, n301, n306, n274, n226, n234, n298, n308, 
        n241, n266, n227, n283, n313, n249, n252, n275, n290, n300, n282, n312, 
        n240, n267, n232, n235, n299, n309, n247, n260, n229, n285, n315, n255, 
        n272, n297, n307, n269, n220;
    VMW_OAI21 U3 ( .A(A[31]), .B(n219), .C(n220), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n224), .B(B[0]), .C(n225), .D(B[1]), .Z(n223) );
    VMW_OR2 U6 ( .A(B[2]), .B(n222), .Z(n226) );
    VMW_OR2 U14 ( .A(B[6]), .B(n236), .Z(n239) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n252), .C(n247), .D(n242), .Z(n251) );
    VMW_OR2 U54 ( .A(B[26]), .B(n300), .Z(n303) );
    VMW_INV U73 ( .A(B[27]), .Z(n309) );
    VMW_INV U96 ( .A(B[31]), .Z(n219) );
    VMW_INV U68 ( .A(A[30]), .Z(n317) );
    VMW_NAND2 U28 ( .A(n262), .B(B[14]), .Z(n261) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n270), .C(n266), .D(n261), .Z(n269) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n225), .C(n226), .D(n223), .Z(n227) );
    VMW_NAND2 U8 ( .A(n229), .B(B[4]), .Z(n228) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n238), .C(n233), .D(n228), .Z(n237) );
    VMW_OR2 U34 ( .A(B[16]), .B(n268), .Z(n271) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n284), .C(n279), .D(n274), .Z(n283) );
    VMW_NAND2 U46 ( .A(n290), .B(A[21]), .Z(n291) );
    VMW_NAND2 U61 ( .A(n314), .B(A[29]), .Z(n315) );
    VMW_INV U84 ( .A(B[15]), .Z(n270) );
    VMW_INV U101 ( .A(A[6]), .Z(n236) );
    VMW_INV U66 ( .A(B[7]), .Z(n245) );
    VMW_INV U83 ( .A(A[15]), .Z(n273) );
    VMW_INV U98 ( .A(B[13]), .Z(n264) );
    VMW_NAND2 U26 ( .A(n258), .B(A[11]), .Z(n259) );
    VMW_NAND2 U48 ( .A(n294), .B(B[24]), .Z(n293) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n231), .C(n227), .D(n221), .Z(n230) );
    VMW_NAND2 U12 ( .A(n236), .B(B[6]), .Z(n235) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n273), .C(n271), .D(n269), .Z(n272) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n302), .C(n298), .D(n293), .Z(n301) );
    VMW_INV U91 ( .A(B[11]), .Z(n258) );
    VMW_INV U74 ( .A(A[3]), .Z(n234) );
    VMW_INV U99 ( .A(A[26]), .Z(n300) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n256), .C(n259), .D(n257), .Z(n260) );
    VMW_NAND2 U40 ( .A(n282), .B(B[20]), .Z(n281) );
    VMW_INV U82 ( .A(B[29]), .Z(n314) );
    VMW_NAND2 U52 ( .A(n300), .B(B[26]), .Z(n299) );
    VMW_INV U67 ( .A(A[7]), .Z(n248) );
    VMW_INV U75 ( .A(B[3]), .Z(n231) );
    VMW_INV U90 ( .A(A[14]), .Z(n262) );
    VMW_NAND2 U20 ( .A(n250), .B(B[10]), .Z(n249) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n296), .C(n292), .D(n287), .Z(n295) );
    VMW_INV U69 ( .A(B[17]), .Z(n277) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n264), .C(n260), .D(n255), .Z(n263) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n288), .C(n291), .D(n289), .Z(n292) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n305), .C(n303), .D(n301), .Z(n304) );
    VMW_INV U72 ( .A(A[27]), .Z(n312) );
    VMW_INV U97 ( .A(A[16]), .Z(n268) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n314), .C(n311), .D(n306), .Z(n313) );
    VMW_INV U100 ( .A(B[23]), .Z(n296) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n241), .C(n239), .D(n237), .Z(n240) );
    VMW_INV U85 ( .A(A[4]), .Z(n229) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n245), .C(n240), .D(n235), .Z(n244) );
    VMW_NAND2 U22 ( .A(n252), .B(A[9]), .Z(n253) );
    VMW_NAND2 U32 ( .A(n268), .B(B[16]), .Z(n267) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n280), .C(n278), .D(n276), .Z(n279) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n309), .C(n304), .D(n299), .Z(n308) );
    VMW_INV U70 ( .A(A[17]), .Z(n280) );
    VMW_INV U95 ( .A(A[1]), .Z(n225) );
    VMW_NAND2 U30 ( .A(n264), .B(A[13]), .Z(n265) );
    VMW_INV U79 ( .A(B[19]), .Z(n284) );
    VMW_INV U87 ( .A(A[8]), .Z(n243) );
    VMW_OR2 U10 ( .A(B[4]), .B(n229), .Z(n232) );
    VMW_NAND2 U42 ( .A(n284), .B(A[19]), .Z(n285) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n290), .C(n286), .D(n281), .Z(n289) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n317), .C(n315), .D(n313), .Z(n316) );
    VMW_INV U65 ( .A(A[12]), .Z(n256) );
    VMW_INV U102 ( .A(A[2]), .Z(n222) );
    VMW_INV U80 ( .A(A[10]), .Z(n250) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n234), .C(n232), .D(n230), .Z(n233) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n248), .C(n246), .D(n244), .Z(n247) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n258), .C(n254), .D(n249), .Z(n257) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n277), .C(n272), .D(n267), .Z(n276) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n312), .C(n310), .D(n308), .Z(n311) );
    VMW_INV U89 ( .A(A[18]), .Z(n275) );
    VMW_NAND2 U50 ( .A(n296), .B(A[23]), .Z(n297) );
    VMW_INV U77 ( .A(A[25]), .Z(n305) );
    VMW_INV U92 ( .A(A[28]), .Z(n307) );
    VMW_OR2 U58 ( .A(B[28]), .B(n307), .Z(n310) );
    VMW_NAND2 U36 ( .A(n275), .B(B[18]), .Z(n274) );
    VMW_INV U81 ( .A(B[9]), .Z(n252) );
    VMW_NAND2 U4 ( .A(n222), .B(B[2]), .Z(n221) );
    VMW_OR2 U18 ( .A(B[8]), .B(n243), .Z(n246) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n282), .C(n285), .D(n283), .Z(n286) );
    VMW_AO22 U64 ( .A(n316), .B(n318), .C(A[31]), .D(n219), .Z(n220) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n294), .C(n297), .D(n295), .Z(n298) );
    VMW_INV U76 ( .A(B[25]), .Z(n302) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n250), .C(n253), .D(n251), .Z(n254) );
    VMW_NAND2 U24 ( .A(n256), .B(B[12]), .Z(n255) );
    VMW_INV U88 ( .A(B[21]), .Z(n290) );
    VMW_INV U93 ( .A(A[5]), .Z(n241) );
    VMW_OR2 U38 ( .A(B[18]), .B(n275), .Z(n278) );
    VMW_NAND2 U44 ( .A(n288), .B(B[22]), .Z(n287) );
    VMW_NAND2 U56 ( .A(n307), .B(B[28]), .Z(n306) );
    VMW_INV U94 ( .A(B[5]), .Z(n238) );
    VMW_INV U71 ( .A(A[22]), .Z(n288) );
    VMW_NAND2 U63 ( .A(n317), .B(B[30]), .Z(n318) );
    VMW_INV U86 ( .A(A[24]), .Z(n294) );
    VMW_INV U103 ( .A(A[0]), .Z(n224) );
    VMW_NAND2 U16 ( .A(n243), .B(B[8]), .Z(n242) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n262), .C(n265), .D(n263), .Z(n266) );
    VMW_INV U78 ( .A(A[20]), .Z(n282) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n330, n379, n362, n339, n345, n387, n395, n406, n414, n370, n357, 
        n322, n319, n325, n389, n408, n350, n377, n392, n413, n342, n380, n401, 
        n359, n365, n337, n351, n393, n412, n376, n324, n336, n388, n409, n343, 
        n358, n364, n381, n400, n386, n407, n323, n331, n344, n363, n378, n356, 
        n371, n333, n338, n394, n415, n328, n346, n361, n384, n405, n396, n321, 
        n354, n368, n373, n326, n348, n353, n374, n383, n391, n410, n402, n341, 
        n366, n334, n390, n398, n411, n349, n352, n375, n327, n335, n399, n340, 
        n367, n329, n382, n403, n385, n404, n347, n360, n332, n320, n369, n355, 
        n372, n397, n416;
    VMW_OAI21 U3 ( .A(A[31]), .B(n319), .C(n320), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n322), .C(B[0]), .Z(n323) );
    VMW_AO22 U6 ( .A(A[2]), .B(n325), .C(n323), .D(A[0]), .Z(n324) );
    VMW_OR2 U14 ( .A(B[6]), .B(n334), .Z(n337) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n350), .C(n345), .D(n340), .Z(n349) );
    VMW_OR2 U54 ( .A(B[26]), .B(n398), .Z(n401) );
    VMW_INV U73 ( .A(B[27]), .Z(n407) );
    VMW_INV U96 ( .A(A[16]), .Z(n366) );
    VMW_INV U68 ( .A(A[30]), .Z(n415) );
    VMW_NAND2 U28 ( .A(n360), .B(B[14]), .Z(n359) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n368), .C(n364), .D(n359), .Z(n367) );
    VMW_OAI22 U7 ( .A(n321), .B(n324), .C(A[2]), .D(n325), .Z(n326) );
    VMW_NAND2 U8 ( .A(n328), .B(B[4]), .Z(n327) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n336), .C(n332), .D(n327), .Z(n335) );
    VMW_OR2 U34 ( .A(B[16]), .B(n366), .Z(n369) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n382), .C(n377), .D(n372), .Z(n381) );
    VMW_NAND2 U46 ( .A(n388), .B(A[21]), .Z(n389) );
    VMW_NAND2 U61 ( .A(n412), .B(A[29]), .Z(n413) );
    VMW_INV U84 ( .A(A[4]), .Z(n328) );
    VMW_INV U101 ( .A(B[2]), .Z(n325) );
    VMW_INV U66 ( .A(B[7]), .Z(n343) );
    VMW_INV U83 ( .A(B[15]), .Z(n368) );
    VMW_INV U98 ( .A(A[26]), .Z(n398) );
    VMW_NAND2 U26 ( .A(n356), .B(A[11]), .Z(n357) );
    VMW_NAND2 U48 ( .A(n392), .B(B[24]), .Z(n391) );
    VMW_AO21 U9 ( .A(B[3]), .B(n330), .C(n326), .Z(n329) );
    VMW_NAND2 U12 ( .A(n334), .B(B[6]), .Z(n333) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n371), .C(n369), .D(n367), .Z(n370) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n400), .C(n396), .D(n391), .Z(n399) );
    VMW_INV U91 ( .A(A[28]), .Z(n405) );
    VMW_INV U74 ( .A(A[3]), .Z(n330) );
    VMW_INV U99 ( .A(B[23]), .Z(n394) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n354), .C(n357), .D(n355), .Z(n358) );
    VMW_NAND2 U40 ( .A(n380), .B(B[20]), .Z(n379) );
    VMW_INV U82 ( .A(A[15]), .Z(n371) );
    VMW_NAND2 U52 ( .A(n398), .B(B[26]), .Z(n397) );
    VMW_INV U67 ( .A(A[7]), .Z(n346) );
    VMW_INV U75 ( .A(B[25]), .Z(n400) );
    VMW_INV U90 ( .A(B[11]), .Z(n356) );
    VMW_NAND2 U20 ( .A(n348), .B(B[10]), .Z(n347) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n394), .C(n390), .D(n385), .Z(n393) );
    VMW_INV U69 ( .A(B[17]), .Z(n375) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n362), .C(n358), .D(n353), .Z(n361) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n386), .C(n389), .D(n387), .Z(n390) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n403), .C(n401), .D(n399), .Z(n402) );
    VMW_INV U72 ( .A(A[27]), .Z(n410) );
    VMW_INV U97 ( .A(B[13]), .Z(n362) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n412), .C(n409), .D(n404), .Z(n411) );
    VMW_INV U100 ( .A(A[6]), .Z(n334) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n339), .C(n337), .D(n335), .Z(n338) );
    VMW_INV U85 ( .A(A[24]), .Z(n392) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n343), .C(n338), .D(n333), .Z(n342) );
    VMW_NAND2 U22 ( .A(n350), .B(A[9]), .Z(n351) );
    VMW_NAND2 U32 ( .A(n366), .B(B[16]), .Z(n365) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n378), .C(n376), .D(n374), .Z(n377) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n407), .C(n402), .D(n397), .Z(n406) );
    VMW_INV U70 ( .A(A[17]), .Z(n378) );
    VMW_INV U95 ( .A(B[31]), .Z(n319) );
    VMW_NAND2 U30 ( .A(n362), .B(A[13]), .Z(n363) );
    VMW_INV U79 ( .A(A[10]), .Z(n348) );
    VMW_INV U87 ( .A(B[21]), .Z(n388) );
    VMW_OR2 U10 ( .A(B[4]), .B(n328), .Z(n331) );
    VMW_NAND2 U42 ( .A(n382), .B(A[19]), .Z(n383) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n388), .C(n384), .D(n379), .Z(n387) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n415), .C(n413), .D(n411), .Z(n414) );
    VMW_INV U65 ( .A(A[12]), .Z(n354) );
    VMW_INV U80 ( .A(B[9]), .Z(n350) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n330), .C(n331), .D(n329), .Z(n332) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n346), .C(n344), .D(n342), .Z(n345) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n356), .C(n352), .D(n347), .Z(n355) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n375), .C(n370), .D(n365), .Z(n374) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n410), .C(n408), .D(n406), .Z(n409) );
    VMW_INV U89 ( .A(A[14]), .Z(n360) );
    VMW_NAND2 U50 ( .A(n394), .B(A[23]), .Z(n395) );
    VMW_INV U77 ( .A(A[20]), .Z(n380) );
    VMW_INV U92 ( .A(A[5]), .Z(n339) );
    VMW_OR2 U58 ( .A(B[28]), .B(n405), .Z(n408) );
    VMW_NAND2 U36 ( .A(n373), .B(B[18]), .Z(n372) );
    VMW_INV U81 ( .A(B[29]), .Z(n412) );
    VMW_NOR2 U4 ( .A(n322), .B(B[1]), .Z(n321) );
    VMW_OR2 U18 ( .A(B[8]), .B(n341), .Z(n344) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n380), .C(n383), .D(n381), .Z(n384) );
    VMW_AO22 U64 ( .A(n414), .B(n416), .C(A[31]), .D(n319), .Z(n320) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n392), .C(n395), .D(n393), .Z(n396) );
    VMW_INV U76 ( .A(A[25]), .Z(n403) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n348), .C(n351), .D(n349), .Z(n352) );
    VMW_NAND2 U24 ( .A(n354), .B(B[12]), .Z(n353) );
    VMW_INV U88 ( .A(A[18]), .Z(n373) );
    VMW_INV U93 ( .A(B[5]), .Z(n336) );
    VMW_OR2 U38 ( .A(B[18]), .B(n373), .Z(n376) );
    VMW_NAND2 U44 ( .A(n386), .B(B[22]), .Z(n385) );
    VMW_NAND2 U56 ( .A(n405), .B(B[28]), .Z(n404) );
    VMW_INV U94 ( .A(A[1]), .Z(n322) );
    VMW_INV U71 ( .A(A[22]), .Z(n386) );
    VMW_NAND2 U63 ( .A(n415), .B(B[30]), .Z(n416) );
    VMW_INV U86 ( .A(A[8]), .Z(n341) );
    VMW_NAND2 U16 ( .A(n341), .B(B[8]), .Z(n340) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n360), .C(n363), .D(n361), .Z(n364) );
    VMW_INV U78 ( .A(B[19]), .Z(n382) );
endmodule


module BHeap_Node_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, Enable, 
    P_WR, P_In, P_Out, L_WR, L_In, L_Out, R_WR, R_In, R_Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
output [31:0] P_Out;
output [31:0] L_Out;
input  [31:0] R_In;
input  [31:0] P_In;
input  [31:0] L_In;
output [31:0] R_Out;
input  Clk, Reset, RD, WR, Enable;
output P_WR, L_WR, R_WR;
    wire n454, n100, n421, n433, n446, n428, n441, n434, n426, n448, n90, n453, 
        n435, n449, n98, n440, n452, n427, n420, n429, n447, n439, n432, n422, 
        n417, n430, n445, n442, n437, n425, n450, n419, n436, n443, n418, n451, 
        n92, n424, n423, n438, n444, n431;
    tri \P_Out[31] , \R_Out[25]1 , \R_Out[16]1 , \R_Out[24]1 , \R_Out[17]1 , 
        \P_Out[21]1 , \P_Out[12]1 , \P_Out[20]1 , \P_Out[13]1 , \P_Out[7]1 , 
        \R_Out[2]1 , \L_Out[20]1 , \L_Out[13]1 , \L_Out[6]1 , \R_Out[3]1 , 
        \R_Out[30]1 , \R_Out[29]1 , \P_Out[6]1 , \L_Out[7]1 , \R_Out[28]1 , 
        \L_Out[21]1 , \L_Out[12]1 , \P_Out[24]1 , \P_Out[17]1 , \P_Out[25]1 , 
        \P_Out[16]1 , \L_Out[30]1 , \R_Out[20]1 , \R_Out[13]1 , \L_Out[29]1 , 
        \L_Out[28]1 , \R_Out[21]1 , \R_Out[12]1 , \L_Out[3]1 , \P_Out[2]1 , 
        \L_Out[25]1 , \L_Out[16]1 , \P_Out[3]1 , \L_Out[2]1 , \L_Out[24]1 , 
        \L_Out[17]1 , \R_Out[7]1 , \P_Out[28]1 , \P_Out[30]1 , \P_Out[29]1 , 
        \R_Out[6]1 , \P_Out[26]1 , \P_Out[15]1 , \R_Out[9]1 , \R_Out[8]1 , 
        \P_Out[27]1 , \P_Out[14]1 , \L_Out[18]1 , \R_Out[22]1 , \R_Out[11]1 , 
        \P_Out[0]1 , \L_Out[27]1 , \L_Out[19]1 , \R_Out[23]1 , \R_Out[10]1 , 
        \L_Out[1]1 , \L_Out[14]1 , \L_Out[0]1 , \P_Out[1]1 , \L_Out[26]1 , 
        \L_Out[15]1 , \R_Out[5]1 , \P_Out[19]1 , \P_Out[18]1 , \L_Out[31] , 
        \P_Out[9]1 , \L_Out[8]1 , \R_Out[4]1 , \R_Out[27]1 , \R_Out[14]1 , 
        \P_Out[23]1 , \P_Out[10]1 , \P_Out[8]1 , \L_Out[9]1 , \R_Out[26]1 , 
        \R_Out[15]1 , \P_Out[22]1 , \P_Out[11]1 , \P_Out[5]1 , \R_Out[0]1 , 
        \R_Out[1]1 , \L_Out[22]1 , \L_Out[11]1 , \L_Out[4]1 , \R_Out[18]1 , 
        \R_Out[31] , \P_Out[4]1 , \L_Out[5]1 , \R_Out[19]1 , \L_Out[23]1 , 
        \L_Out[10]1 ;
    assign P_Out[31] = \P_Out[31] ;
    assign P_Out[30] = \P_Out[30]1 ;
    assign P_Out[29] = \P_Out[29]1 ;
    assign P_Out[28] = \P_Out[28]1 ;
    assign P_Out[27] = \P_Out[27]1 ;
    assign P_Out[26] = \P_Out[26]1 ;
    assign P_Out[25] = \P_Out[25]1 ;
    assign P_Out[24] = \P_Out[24]1 ;
    assign P_Out[23] = \P_Out[23]1 ;
    assign P_Out[22] = \P_Out[22]1 ;
    assign P_Out[21] = \P_Out[21]1 ;
    assign P_Out[20] = \P_Out[20]1 ;
    assign P_Out[19] = \P_Out[19]1 ;
    assign P_Out[18] = \P_Out[18]1 ;
    assign P_Out[17] = \P_Out[17]1 ;
    assign P_Out[16] = \P_Out[16]1 ;
    assign P_Out[15] = \P_Out[15]1 ;
    assign P_Out[14] = \P_Out[14]1 ;
    assign P_Out[13] = \P_Out[13]1 ;
    assign P_Out[12] = \P_Out[12]1 ;
    assign P_Out[11] = \P_Out[11]1 ;
    assign P_Out[10] = \P_Out[10]1 ;
    assign P_Out[9] = \P_Out[9]1 ;
    assign P_Out[8] = \P_Out[8]1 ;
    assign P_Out[7] = \P_Out[7]1 ;
    assign P_Out[6] = \P_Out[6]1 ;
    assign P_Out[5] = \P_Out[5]1 ;
    assign P_Out[4] = \P_Out[4]1 ;
    assign P_Out[3] = \P_Out[3]1 ;
    assign P_Out[2] = \P_Out[2]1 ;
    assign P_Out[1] = \P_Out[1]1 ;
    assign P_Out[0] = \P_Out[0]1 ;
    assign L_Out[31] = \L_Out[31] ;
    assign L_Out[30] = \L_Out[30]1 ;
    assign L_Out[29] = \L_Out[29]1 ;
    assign L_Out[28] = \L_Out[28]1 ;
    assign L_Out[27] = \L_Out[27]1 ;
    assign L_Out[26] = \L_Out[26]1 ;
    assign L_Out[25] = \L_Out[25]1 ;
    assign L_Out[24] = \L_Out[24]1 ;
    assign L_Out[23] = \L_Out[23]1 ;
    assign L_Out[22] = \L_Out[22]1 ;
    assign L_Out[21] = \L_Out[21]1 ;
    assign L_Out[20] = \L_Out[20]1 ;
    assign L_Out[19] = \L_Out[19]1 ;
    assign L_Out[18] = \L_Out[18]1 ;
    assign L_Out[17] = \L_Out[17]1 ;
    assign L_Out[16] = \L_Out[16]1 ;
    assign L_Out[15] = \L_Out[15]1 ;
    assign L_Out[14] = \L_Out[14]1 ;
    assign L_Out[13] = \L_Out[13]1 ;
    assign L_Out[12] = \L_Out[12]1 ;
    assign L_Out[11] = \L_Out[11]1 ;
    assign L_Out[10] = \L_Out[10]1 ;
    assign L_Out[9] = \L_Out[9]1 ;
    assign L_Out[8] = \L_Out[8]1 ;
    assign L_Out[7] = \L_Out[7]1 ;
    assign L_Out[6] = \L_Out[6]1 ;
    assign L_Out[5] = \L_Out[5]1 ;
    assign L_Out[4] = \L_Out[4]1 ;
    assign L_Out[3] = \L_Out[3]1 ;
    assign L_Out[2] = \L_Out[2]1 ;
    assign L_Out[1] = \L_Out[1]1 ;
    assign L_Out[0] = \L_Out[0]1 ;
    assign R_Out[31] = \R_Out[31] ;
    assign R_Out[30] = \R_Out[30]1 ;
    assign R_Out[29] = \R_Out[29]1 ;
    assign R_Out[28] = \R_Out[28]1 ;
    assign R_Out[27] = \R_Out[27]1 ;
    assign R_Out[26] = \R_Out[26]1 ;
    assign R_Out[25] = \R_Out[25]1 ;
    assign R_Out[24] = \R_Out[24]1 ;
    assign R_Out[23] = \R_Out[23]1 ;
    assign R_Out[22] = \R_Out[22]1 ;
    assign R_Out[21] = \R_Out[21]1 ;
    assign R_Out[20] = \R_Out[20]1 ;
    assign R_Out[19] = \R_Out[19]1 ;
    assign R_Out[18] = \R_Out[18]1 ;
    assign R_Out[17] = \R_Out[17]1 ;
    assign R_Out[16] = \R_Out[16]1 ;
    assign R_Out[15] = \R_Out[15]1 ;
    assign R_Out[14] = \R_Out[14]1 ;
    assign R_Out[13] = \R_Out[13]1 ;
    assign R_Out[12] = \R_Out[12]1 ;
    assign R_Out[11] = \R_Out[11]1 ;
    assign R_Out[10] = \R_Out[10]1 ;
    assign R_Out[9] = \R_Out[9]1 ;
    assign R_Out[8] = \R_Out[8]1 ;
    assign R_Out[7] = \R_Out[7]1 ;
    assign R_Out[6] = \R_Out[6]1 ;
    assign R_Out[5] = \R_Out[5]1 ;
    assign R_Out[4] = \R_Out[4]1 ;
    assign R_Out[3] = \R_Out[3]1 ;
    assign R_Out[2] = \R_Out[2]1 ;
    assign R_Out[1] = \R_Out[1]1 ;
    assign R_Out[0] = \R_Out[0]1 ;
    VMW_AO22 U54 ( .A(R_In[26]), .B(n417), .C(L_In[26]), .D(L_WR), .Z(n431) );
    VMW_AND3 U73 ( .A(n92), .B(Enable), .C(n90), .Z(L_WR) );
    VMW_BUFIZ U113 ( .A(P_In[3]), .E(L_WR), .Z(\L_Out[3]1 ) );
    VMW_BUFIZ U134 ( .A(P_In[22]), .E(R_WR), .Z(\R_Out[22]1 ) );
    VMW_AO22 U68 ( .A(R_In[13]), .B(n417), .C(L_In[13]), .D(L_WR), .Z(n426) );
    VMW_BUFIZ U96 ( .A(n421), .E(P_WR), .Z(\P_Out[17]1 ) );
    VMW_BUFIZ U108 ( .A(P_In[12]), .E(R_WR), .Z(\R_Out[12]1 ) );
    VMW_BUFIZ U141 ( .A(n444), .E(P_WR), .Z(\P_Out[3]1 ) );
    VMW_BUFIZ U166 ( .A(P_In[4]), .E(R_WR), .Z(\R_Out[4]1 ) );
    VMW_PULLDOWN U35 ( .Z(n451) );
    VMW_AO22 U41 ( .A(R_In[9]), .B(n417), .C(L_In[9]), .D(L_WR), .Z(n429) );
    VMW_AO22 U46 ( .A(R_In[4]), .B(n417), .C(L_In[4]), .D(L_WR), .Z(n433) );
    VMW_AO22 U61 ( .A(R_In[1]), .B(n417), .C(L_In[1]), .D(L_WR), .Z(n443) );
    VMW_BUFIZ U84 ( .A(P_In[24]), .E(L_WR), .Z(\L_Out[24]1 ) );
    VMW_BUFIZ U148 ( .A(P_In[13]), .E(R_WR), .Z(\R_Out[13]1 ) );
    VMW_BUFIZ U153 ( .A(n449), .E(P_WR), .Z(\P_Out[16]1 ) );
    VMW_BUFIZ U101 ( .A(n424), .E(P_WR), .Z(\P_Out[20]1 ) );
    VMW_BUFIZ U126 ( .A(n434), .E(P_WR), .Z(\P_Out[27]1 ) );
    VMW_AO22 U48 ( .A(R_In[31]), .B(n417), .C(L_In[31]), .D(L_WR), .Z(n440) );
    VMW_AO22 U66 ( .A(R_In[15]), .B(n417), .C(L_In[15]), .D(L_WR), .Z(n432) );
    VMW_BUFIZ U106 ( .A(P_In[28]), .E(R_WR), .Z(\R_Out[28]1 ) );
    VMW_BUFIZ U121 ( .A(n432), .E(P_WR), .Z(\P_Out[15]1 ) );
    VMW_BUFIZ U83 ( .A(P_In[15]), .E(L_WR), .Z(\L_Out[15]1 ) );
    VMW_BUFIZ U168 ( .A(P_In[9]), .E(R_WR), .Z(\R_Out[9]1 ) );
    VMW_BUFIZ U98 ( .A(P_In[16]), .E(R_WR), .Z(\R_Out[16]1 ) );
    VMW_BUFIZ U128 ( .A(n436), .E(P_WR), .Z(\P_Out[14]1 ) );
    VMW_BUFIZ U154 ( .A(P_In[24]), .E(R_WR), .Z(\R_Out[24]1 ) );
    VMW_AO22 U53 ( .A(R_In[27]), .B(n417), .C(L_In[27]), .D(L_WR), .Z(n434) );
    VMW_BUFIZ U91 ( .A(n420), .E(P_WR), .Z(\P_Out[6]1 ) );
    VMW_BUFIZ U146 ( .A(P_In[9]), .E(L_WR), .Z(\L_Out[9]1 ) );
    VMW_BUFIZ U161 ( .A(P_In[25]), .E(L_WR), .Z(\L_Out[25]1 ) );
    VMW_AND3 U74 ( .A(n98), .B(n100), .C(Enable), .Z(R_WR) );
    VMW_BUFIZ U114 ( .A(P_In[23]), .E(R_WR), .Z(\R_Out[23]1 ) );
    VMW_BUFIZ U133 ( .A(P_In[2]), .E(L_WR), .Z(\L_Out[2]1 ) );
    VMW_BUFIZ U99 ( .A(n422), .E(P_WR), .Z(\P_Out[29]1 ) );
    VMW_BUFIZ U155 ( .A(P_In[17]), .E(R_WR), .Z(\R_Out[17]1 ) );
    VMW_OR2 U40 ( .A(L_WR), .B(R_WR), .Z(P_WR) );
    VMW_BUFIZ U82 ( .A(P_In[26]), .E(L_WR), .Z(\L_Out[26]1 ) );
    VMW_BUFIZ U169 ( .A(P_In[23]), .E(L_WR), .Z(\L_Out[23]1 ) );
    VMW_AO22 U47 ( .A(R_In[3]), .B(n417), .C(L_In[3]), .D(L_WR), .Z(n444) );
    VMW_AO22 U49 ( .A(R_In[30]), .B(n417), .C(L_In[30]), .D(L_WR), .Z(n418) );
    VMW_AO22 U52 ( .A(R_In[28]), .B(n417), .C(L_In[28]), .D(L_WR), .Z(n441) );
    VMW_AO22 U67 ( .A(R_In[14]), .B(n417), .C(L_In[14]), .D(L_WR), .Z(n436) );
    VMW_BUFIZ U107 ( .A(P_In[21]), .E(R_WR), .Z(\R_Out[21]1 ) );
    VMW_BUFIZ U120 ( .A(n431), .E(P_WR), .Z(\P_Out[26]1 ) );
    VMW_INV U75 ( .A(L_WR), .Z(n417) );
    VMW_BUFIZ U115 ( .A(P_In[10]), .E(R_WR), .Z(\R_Out[10]1 ) );
    VMW_BUFIZ U132 ( .A(n439), .E(P_WR), .Z(\P_Out[8]1 ) );
    VMW_BUFIZ U90 ( .A(n419), .E(P_WR), .Z(\P_Out[24]1 ) );
    VMW_BUFIZ U129 ( .A(n437), .E(P_WR), .Z(\P_Out[5]1 ) );
    VMW_BUFIZ U147 ( .A(P_In[20]), .E(R_WR), .Z(\R_Out[20]1 ) );
    VMW_BUFIZ U160 ( .A(P_In[28]), .E(L_WR), .Z(\L_Out[28]1 ) );
    VMW_AO22 U55 ( .A(R_In[25]), .B(n417), .C(L_In[25]), .D(L_WR), .Z(n448) );
    VMW_AO22 U69 ( .A(R_In[12]), .B(n417), .C(L_In[12]), .D(L_WR), .Z(n446) );
    VMW_BUFIZ U109 ( .A(n426), .E(P_WR), .Z(\P_Out[13]1 ) );
    VMW_AO22 U72 ( .A(R_In[0]), .B(n417), .C(L_In[0]), .D(L_WR), .Z(n430) );
    VMW_BUFIZ U97 ( .A(P_In[25]), .E(R_WR), .Z(\R_Out[25]1 ) );
    VMW_BUFIZ U140 ( .A(n443), .E(P_WR), .Z(\P_Out[1]1 ) );
    VMW_BUFIZ U167 ( .A(P_In[19]), .E(L_WR), .Z(\L_Out[19]1 ) );
    VMW_BUFIZ U112 ( .A(n429), .E(P_WR), .Z(\P_Out[9]1 ) );
    VMW_BUFIZ U135 ( .A(P_In[11]), .E(R_WR), .Z(\R_Out[11]1 ) );
    VMW_AO22 U60 ( .A(R_In[20]), .B(n417), .C(L_In[20]), .D(L_WR), .Z(n424) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_1 gt_48_1 ( .A(L_In), .B(R_In), .LEQ(n452), 
        .TC(n452), .LT_LE(n100) );
    VMW_BUFIZ U100 ( .A(n423), .E(P_WR), .Z(\P_Out[22]1 ) );
    VMW_BUFIZ U127 ( .A(n435), .E(P_WR), .Z(\P_Out[23]1 ) );
    VMW_BUFIZ U85 ( .A(P_In[17]), .E(L_WR), .Z(\L_Out[17]1 ) );
    VMW_BUFIZ U149 ( .A(n446), .E(P_WR), .Z(\P_Out[12]1 ) );
    VMW_BUFIZ U152 ( .A(n448), .E(P_WR), .Z(\P_Out[25]1 ) );
    VMW_PULLUP U36 ( .Z(n450) );
    VMW_PULLDOWN U37 ( .Z(n452) );
    VMW_PULLDOWN U39 ( .Z(n454) );
    VMW_AO22 U57 ( .A(R_In[23]), .B(n417), .C(L_In[23]), .D(L_WR), .Z(n435) );
    VMW_BUFIZ U137 ( .A(n441), .E(P_WR), .Z(\P_Out[28]1 ) );
    VMW_AO22 U70 ( .A(R_In[11]), .B(n417), .C(L_In[11]), .D(L_WR), .Z(n428) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_2 gt_48 ( .A(P_In), .B(R_In), .LEQ(n453), 
        .TC(n453), .LT_LE(n98) );
    VMW_BUFIZ U110 ( .A(n427), .E(P_WR), .Z(\P_Out[18]1 ) );
    VMW_BUFIZ U159 ( .A(P_In[12]), .E(L_WR), .Z(\L_Out[12]1 ) );
    VMW_AO22 U42 ( .A(R_In[8]), .B(n417), .C(L_In[8]), .D(L_WR), .Z(n439) );
    VMW_AO22 U45 ( .A(R_In[5]), .B(n417), .C(L_In[5]), .D(L_WR), .Z(n437) );
    VMW_BUFIZ U79 ( .A(P_In[11]), .E(L_WR), .Z(\L_Out[11]1 ) );
    VMW_BUFIZ U95 ( .A(P_In[5]), .E(L_WR), .Z(\L_Out[5]1 ) );
    VMW_BUFIZ U119 ( .A(P_In[14]), .E(R_WR), .Z(\R_Out[14]1 ) );
    VMW_BUFIZ U142 ( .A(P_In[0]), .E(L_WR), .Z(\L_Out[0]1 ) );
    VMW_BUFIZ U165 ( .A(P_In[14]), .E(L_WR), .Z(\L_Out[14]1 ) );
    VMW_BUFIZ U87 ( .A(P_In[13]), .E(L_WR), .Z(\L_Out[13]1 ) );
    VMW_BUFIZ U150 ( .A(n447), .E(P_WR), .Z(\P_Out[7]1 ) );
    VMW_BUFIZ U125 ( .A(P_In[15]), .E(R_WR), .Z(\R_Out[15]1 ) );
    VMW_AO22 U62 ( .A(R_In[19]), .B(n417), .C(L_In[19]), .D(L_WR), .Z(n442) );
    VMW_AO22 U65 ( .A(R_In[16]), .B(n417), .C(L_In[16]), .D(L_WR), .Z(n449) );
    VMW_BUFIZ U102 ( .A(n425), .E(P_WR), .Z(\P_Out[2]1 ) );
    VMW_BUFIZ U105 ( .A(P_In[31]), .E(R_WR), .Z(\R_Out[31] ) );
    VMW_BUFIZ U80 ( .A(P_In[5]), .E(R_WR), .Z(\R_Out[5]1 ) );
    VMW_BUFIZ U122 ( .A(n433), .E(P_WR), .Z(\P_Out[4]1 ) );
    VMW_BUFIZ U157 ( .A(P_In[31]), .E(L_WR), .Z(\L_Out[31] ) );
    VMW_BUFIZ U170 ( .A(P_In[10]), .E(L_WR), .Z(\L_Out[10]1 ) );
    VMW_AO22 U50 ( .A(R_In[2]), .B(n417), .C(L_In[2]), .D(L_WR), .Z(n425) );
    VMW_AO22 U59 ( .A(R_In[21]), .B(n417), .C(L_In[21]), .D(L_WR), .Z(n445) );
    VMW_BUFIZ U139 ( .A(P_In[18]), .E(R_WR), .Z(\R_Out[18]1 ) );
    VMW_BUFIZ U77 ( .A(P_In[18]), .E(L_WR), .Z(\L_Out[18]1 ) );
    VMW_BUFIZ U89 ( .A(n418), .E(P_WR), .Z(\P_Out[30]1 ) );
    VMW_BUFIZ U92 ( .A(P_In[30]), .E(L_WR), .Z(\L_Out[30]1 ) );
    VMW_BUFIZ U145 ( .A(n445), .E(P_WR), .Z(\P_Out[21]1 ) );
    VMW_BUFIZ U162 ( .A(P_In[16]), .E(L_WR), .Z(\L_Out[16]1 ) );
    VMW_BUFIZ U117 ( .A(n430), .E(P_WR), .Z(\P_Out[0]1 ) );
    VMW_AO22 U58 ( .A(R_In[22]), .B(n417), .C(L_In[22]), .D(L_WR), .Z(n423) );
    VMW_BUFIZ U130 ( .A(P_In[6]), .E(L_WR), .Z(\L_Out[6]1 ) );
    VMW_BUFIZ U138 ( .A(n442), .E(P_WR), .Z(\P_Out[19]1 ) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_3 gt_47 ( .A(P_In), .B(L_In), .LEQ(n454), 
        .TC(n454), .LT_LE(n90) );
    VMW_BUFIZ U156 ( .A(P_In[2]), .E(R_WR), .Z(\R_Out[2]1 ) );
    VMW_BUFIZ U171 ( .A(P_In[0]), .E(R_WR), .Z(\R_Out[0]1 ) );
    VMW_PULLDOWN U38 ( .Z(n453) );
    VMW_AO22 U43 ( .A(R_In[7]), .B(n417), .C(L_In[7]), .D(L_WR), .Z(n447) );
    VMW_AO22 U64 ( .A(R_In[17]), .B(n417), .C(L_In[17]), .D(L_WR), .Z(n421) );
    VMW_BUFIZ U81 ( .A(P_In[1]), .E(R_WR), .Z(\R_Out[1]1 ) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_0 gte_47 ( .A(R_In), .B(L_In), .LEQ(n450), 
        .TC(n451), .LT_LE(n92) );
    VMW_BUFIZ U104 ( .A(P_In[1]), .E(L_WR), .Z(\L_Out[1]1 ) );
    VMW_AO22 U51 ( .A(R_In[29]), .B(n417), .C(L_In[29]), .D(L_WR), .Z(n422) );
    VMW_BUFIZ U76 ( .A(P_In[22]), .E(L_WR), .Z(\L_Out[22]1 ) );
    VMW_BUFIZ U116 ( .A(P_In[19]), .E(R_WR), .Z(\R_Out[19]1 ) );
    VMW_BUFIZ U123 ( .A(P_In[7]), .E(L_WR), .Z(\L_Out[7]1 ) );
    VMW_BUFIZ U88 ( .A(P_In[3]), .E(R_WR), .Z(\R_Out[3]1 ) );
    VMW_BUFIZ U93 ( .A(P_In[29]), .E(L_WR), .Z(\L_Out[29]1 ) );
    VMW_BUFIZ U131 ( .A(n438), .E(P_WR), .Z(\P_Out[10]1 ) );
    VMW_BUFIZ U143 ( .A(P_In[30]), .E(R_WR), .Z(\R_Out[30]1 ) );
    VMW_BUFIZ U144 ( .A(P_In[29]), .E(R_WR), .Z(\R_Out[29]1 ) );
    VMW_BUFIZ U163 ( .A(P_In[6]), .E(R_WR), .Z(\R_Out[6]1 ) );
    VMW_BUFIZ U158 ( .A(P_In[21]), .E(L_WR), .Z(\L_Out[21]1 ) );
    VMW_BUFIZ U164 ( .A(P_In[27]), .E(L_WR), .Z(\L_Out[27]1 ) );
    VMW_AO22 U44 ( .A(R_In[6]), .B(n417), .C(L_In[6]), .D(L_WR), .Z(n420) );
    VMW_AO22 U56 ( .A(R_In[24]), .B(n417), .C(L_In[24]), .D(L_WR), .Z(n419) );
    VMW_BUFIZ U94 ( .A(P_In[20]), .E(L_WR), .Z(\L_Out[20]1 ) );
    VMW_BUFIZ U136 ( .A(n440), .E(P_WR), .Z(\P_Out[31] ) );
    VMW_AO22 U71 ( .A(R_In[10]), .B(n417), .C(L_In[10]), .D(L_WR), .Z(n438) );
    VMW_BUFIZ U111 ( .A(n428), .E(P_WR), .Z(\P_Out[11]1 ) );
    VMW_BUFIZ U124 ( .A(P_In[26]), .E(R_WR), .Z(\R_Out[26]1 ) );
    VMW_AO22 U63 ( .A(R_In[18]), .B(n417), .C(L_In[18]), .D(L_WR), .Z(n427) );
    VMW_BUFIZ U78 ( .A(P_In[8]), .E(R_WR), .Z(\R_Out[8]1 ) );
    VMW_BUFIZ U86 ( .A(P_In[7]), .E(R_WR), .Z(\R_Out[7]1 ) );
    VMW_BUFIZ U103 ( .A(P_In[8]), .E(L_WR), .Z(\L_Out[8]1 ) );
    VMW_BUFIZ U118 ( .A(P_In[27]), .E(R_WR), .Z(\R_Out[27]1 ) );
    VMW_BUFIZ U151 ( .A(P_In[4]), .E(L_WR), .Z(\L_Out[4]1 ) );
endmodule


module BHeap_CtrlReg_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, In, 
    Out, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR, In;
output Out, Enable;
    wire n77, Out70;
    assign Enable = Out;
    VMW_NOR2 U12 ( .A(n77), .B(Reset), .Z(Out70) );
    VMW_INV U13 ( .A(In), .Z(n77) );
    VMW_FD Out_reg ( .D(Out70), .CP(Clk), .Q(Out) );
endmodule


module BHeap_Control_CWIDTH4_IDWIDTH1_WIDTH32_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, Go, Done );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR, Done;
output ScanEnable, Go;
    wire n379, \Count[0] , n362, n406, n345, n387, n339, n395, n357, n370, 
        n389, n377, n350, n392, n401, n380, n342, n365, \Count[2] , n359, n356, 
        n393, n376, n351, \ScanReg[15] , \ScanReg[26] , \ScanReg[2] , n388, 
        \ScanReg[18] , n358, n343, n364, n400, \ScanReg[11] , \ScanReg[6] , 
        \ScanReg[22] , n381, n344, \ScanReg[20] , \ScanReg[13] , \ScanReg[4] , 
        n386, n407, n363, n378, \ScanReg[29] , \ScanReg[30] , \ScanReg[17] , 
        \ScanReg[24] , \ScanReg[0] , n371, \ScanReg[9] , n338, n394, 
        \ScanReg[16] , \ScanReg[25] , Go259, \ScanReg[1] , n346, \ScanReg[8] , 
        n361, \ScanReg[7] , n405, n384, \ScanReg[5] , n396, \ScanReg[21] , 
        \ScanReg[12] , n373, n354, n368, \ScanReg[28] , \ScanReg[31] , n348, 
        \ScanReg[19] , n374, n353, n391, \ScanReg[10] , n383, \ScanReg[23] , 
        n402, n341, n366, \ScanReg[14] , \ScanReg[27] , n398, \ScanReg[3] , 
        n390, n375, n352, n349, \Count[3] , n399, n360, n340, n367, n403, n382, 
        n404, n385, n347, \Count[1] , n369, n355, n372, n397;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U68 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_AND2 U73 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_OAI211 U96 ( .A(n344), .B(n341), .C(n345), .D(n346), .Z(n405) );
    VMW_AND2 U113 ( .A(\ScanReg[21] ), .B(n349), .Z(n385) );
    VMW_AND2 U134 ( .A(n358), .B(n361), .Z(n360) );
    VMW_FD \Count_reg[0]  ( .D(n407), .CP(Clk), .Q(\Count[0] ) );
    VMW_AND2 U108 ( .A(\ScanReg[20] ), .B(n349), .Z(n391) );
    VMW_MUX2I U141 ( .A(n352), .B(DataIn[0]), .S(n354), .Z(n366) );
    VMW_BUFIZ U166 ( .A(n371), .E(n376), .Z(\arr[19] ) );
    VMW_BUFIZ U183 ( .A(n389), .E(n376), .Z(\arr[30] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AND2 U66 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U84 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_NAND3 U148 ( .A(n353), .B(n363), .C(n360), .Z(n346) );
    VMW_XNOR2 U153 ( .A(Addr[0]), .B(ScanId), .Z(n356) );
    VMW_BUFIZ U174 ( .A(n380), .E(n376), .Z(\arr[25] ) );
    VMW_BUFIZ U191 ( .A(n397), .E(n376), .Z(\arr[26] ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U101 ( .A(\ScanReg[18] ), .B(n349), .Z(n399) );
    VMW_AND2 U106 ( .A(\ScanReg[17] ), .B(n349), .Z(n394) );
    VMW_AND2 U121 ( .A(\ScanReg[4] ), .B(n349), .Z(n377) );
    VMW_AND2 U126 ( .A(\ScanReg[19] ), .B(n349), .Z(n371) );
    VMW_AND2 U74 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U83 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_BUFIZ U168 ( .A(n373), .E(n376), .Z(\arr[23] ) );
    VMW_AND2 U91 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_AND2 U98 ( .A(\ScanReg[8] ), .B(n349), .Z(n403) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_XOR2 U128 ( .A(Addr[0]), .B(Id), .Z(n349) );
    VMW_MUX2I U154 ( .A(n362), .B(n364), .S(\Count[3] ), .Z(n348) );
    VMW_BUFIZ U173 ( .A(n379), .E(n376), .Z(\arr[14] ) );
    VMW_BUFIZ U184 ( .A(n390), .E(n376), .Z(\arr[29] ) );
    VMW_BUFIZ U196 ( .A(n402), .E(n376), .Z(\arr[1] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_OR2 U146 ( .A(Done), .B(n365), .Z(n363) );
    VMW_INV U161 ( .A(\Count[2] ), .Z(n361) );
    VMW_AND2 U114 ( .A(\ScanReg[31] ), .B(n349), .Z(n384) );
    VMW_AND2 U133 ( .A(n359), .B(n352), .Z(n358) );
    VMW_AND2 U99 ( .A(\ScanReg[11] ), .B(n349), .Z(n401) );
    VMW_BUFIZ U197 ( .A(n403), .E(n376), .Z(\arr[8] ) );
    VMW_FD \Count_reg[2]  ( .D(n405), .CP(Clk), .Q(\Count[2] ) );
    VMW_OR2 U155 ( .A(Reset), .B(n366), .Z(n367) );
    VMW_BUFIZ U172 ( .A(n378), .E(n376), .Z(\arr[27] ) );
    VMW_AND2 U67 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U82 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_BUFIZ U169 ( .A(n374), .E(n376), .Z(\arr[10] ) );
    VMW_AND2 U107 ( .A(\ScanReg[24] ), .B(n349), .Z(n393) );
    VMW_AND2 U120 ( .A(\ScanReg[27] ), .B(n349), .Z(n378) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_AND2 U69 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U75 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AND2 U115 ( .A(\ScanReg[12] ), .B(n349), .Z(n383) );
    VMW_NAND2 U132 ( .A(n357), .B(n354), .Z(n341) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U90 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AND2 U109 ( .A(\ScanReg[29] ), .B(n349), .Z(n390) );
    VMW_NOR2 U129 ( .A(Reset), .B(n354), .Z(n353) );
    VMW_OR2 U147 ( .A(n358), .B(n365), .Z(n369) );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_INV U160 ( .A(Reset), .Z(n357) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_BUFIZ U185 ( .A(n391), .E(n376), .Z(\arr[20] ) );
    VMW_BUFIZ U182 ( .A(n388), .E(n376), .Z(\arr[13] ) );
    VMW_AND2 U72 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_OAI21 U97 ( .A(n347), .B(n341), .C(n348), .Z(n404) );
    VMW_OAI21 U140 ( .A(n360), .B(n365), .C(n363), .Z(n364) );
    VMW_BUFIZ U167 ( .A(n372), .E(n376), .Z(\arr[0] ) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD Go_reg ( .D(Go259), .CP(Clk), .Q(Go) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_AND2 U85 ( .A(WR), .B(DataIn[9]), .Z(ScanOut[9]) );
    VMW_AND2 U100 ( .A(\ScanReg[22] ), .B(n349), .Z(n400) );
    VMW_AND2 U112 ( .A(\ScanReg[28] ), .B(n349), .Z(n386) );
    VMW_AO22 U135 ( .A(\Count[3] ), .B(n350), .C(\ScanReg[3] ), .D(n349), .Z(
        n392) );
    VMW_OR4 U127 ( .A(n352), .B(\Count[2] ), .C(\Count[3] ), .D(\Count[1] ), 
        .Z(n351) );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_AO21 U149 ( .A(n363), .B(n369), .C(n361), .Z(n345) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_AO21 U152 ( .A(n363), .B(n370), .C(n359), .Z(n342) );
    VMW_BUFIZ U175 ( .A(n381), .E(n376), .Z(\arr[16] ) );
    VMW_NAND2 U62 ( .A(n338), .B(n339), .Z(Go259) );
    VMW_AND2 U70 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_AO22 U137 ( .A(\Count[1] ), .B(n350), .C(\ScanReg[1] ), .D(n349), .Z(
        n402) );
    VMW_BUFIZ U190 ( .A(n396), .E(n376), .Z(\arr[5] ) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AND2 U79 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_OAI211 U95 ( .A(n340), .B(n341), .C(n342), .D(n343), .Z(n406) );
    VMW_AND2 U110 ( .A(\ScanReg[30] ), .B(n349), .Z(n389) );
    VMW_INV U159 ( .A(DataIn[1]), .Z(n340) );
    VMW_AND2 U119 ( .A(\ScanReg[14] ), .B(n349), .Z(n379) );
    VMW_MUX2I U142 ( .A(n352), .B(n367), .S(n363), .Z(n407) );
    VMW_INV U165 ( .A(n355), .Z(ScanEnable) );
    VMW_BUFIZ U180 ( .A(n386), .E(n376), .Z(\arr[28] ) );
    VMW_BUFIZ U192 ( .A(n398), .E(n376), .Z(\arr[15] ) );
    VMW_AND2 U87 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_NAND2 U150 ( .A(\Count[0] ), .B(n353), .Z(n370) );
    VMW_BUFIZ U177 ( .A(n383), .E(n376), .Z(\arr[12] ) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO21 U125 ( .A(RD), .B(ScanEnable), .C(n350), .Z(n376) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U63 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U64 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U65 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U102 ( .A(\ScanReg[15] ), .B(n349), .Z(n398) );
    VMW_AND2 U105 ( .A(\ScanReg[7] ), .B(n349), .Z(n395) );
    VMW_BUFIZ U189 ( .A(n395), .E(n376), .Z(\arr[7] ) );
    VMW_AND2 U77 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AND2 U80 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U122 ( .A(\ScanReg[9] ), .B(n349), .Z(n375) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_AND2 U89 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_AND3 U139 ( .A(n360), .B(n363), .C(n353), .Z(n362) );
    VMW_INV U157 ( .A(DataIn[3]), .Z(n347) );
    VMW_BUFIZ U170 ( .A(n375), .E(n376), .Z(\arr[9] ) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_BUFIZ U195 ( .A(n401), .E(n376), .Z(\arr[11] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_BUFIZ U187 ( .A(n393), .E(n376), .Z(\arr[24] ) );
    VMW_AND2 U92 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_NAND3 U145 ( .A(n368), .B(n357), .C(n354), .Z(n338) );
    VMW_INV U162 ( .A(\Count[0] ), .Z(n352) );
    VMW_BUFIZ U179 ( .A(n385), .E(n376), .Z(\arr[21] ) );
    VMW_AND2 U117 ( .A(\ScanReg[16] ), .B(n349), .Z(n381) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AND2 U81 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_AND2 U130 ( .A(WR), .B(n350), .Z(n354) );
    VMW_AO22 U138 ( .A(\Count[0] ), .B(n350), .C(\ScanReg[0] ), .D(n349), .Z(
        n372) );
    VMW_BUFIZ U194 ( .A(n400), .E(n376), .Z(\arr[22] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_INV U156 ( .A(n349), .Z(n350) );
    VMW_BUFIZ U171 ( .A(n377), .E(n376), .Z(\arr[4] ) );
    VMW_AND2 U104 ( .A(\ScanReg[5] ), .B(n349), .Z(n396) );
    VMW_AND2 U71 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U76 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AND2 U116 ( .A(\ScanReg[6] ), .B(n349), .Z(n382) );
    VMW_AND2 U123 ( .A(\ScanReg[10] ), .B(n349), .Z(n374) );
    VMW_FD \Count_reg[3]  ( .D(n404), .CP(Clk), .Q(\Count[3] ) );
    VMW_AND2 U88 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_AND2 U93 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_OAI21 U131 ( .A(RD), .B(WR), .C(n356), .Z(n355) );
    VMW_BUFIZ U178 ( .A(n384), .E(n376), .Z(\arr[31] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_OR4 U143 ( .A(DataIn[0]), .B(DataIn[1]), .C(DataIn[2]), .D(DataIn[3]), 
        .Z(n368) );
    VMW_NAND3 U144 ( .A(n351), .B(n353), .C(Done), .Z(n339) );
    VMW_INV U163 ( .A(\Count[1] ), .Z(n359) );
    VMW_BUFIZ U181 ( .A(n387), .E(n376), .Z(\arr[2] ) );
    VMW_BUFIZ U186 ( .A(n392), .E(n376), .Z(\arr[3] ) );
    VMW_INV U158 ( .A(DataIn[2]), .Z(n344) );
    VMW_INV U164 ( .A(n353), .Z(n365) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(\Count[2] ), .B(n350), .C(\ScanReg[2] ), .D(n349), .Z(
        n387) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AND2 U111 ( .A(\ScanReg[13] ), .B(n349), .Z(n388) );
    VMW_AND2 U124 ( .A(\ScanReg[23] ), .B(n349), .Z(n373) );
    VMW_AND2 U78 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_AND2 U86 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U103 ( .A(\ScanReg[26] ), .B(n349), .Z(n397) );
    VMW_BUFIZ U188 ( .A(n394), .E(n376), .Z(\arr[17] ) );
    VMW_FD \Count_reg[1]  ( .D(n406), .CP(Clk), .Q(\Count[1] ) );
    VMW_AND2 U118 ( .A(\ScanReg[25] ), .B(n349), .Z(n380) );
    VMW_NAND3 U151 ( .A(n353), .B(n363), .C(n358), .Z(n343) );
    VMW_BUFIZ U176 ( .A(n382), .E(n376), .Z(\arr[6] ) );
    VMW_BUFIZ U193 ( .A(n399), .E(n376), .Z(\arr[18] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \wRegInTop_3_7[11] , \wRegOut_4_3[16] , \wRegInBot_6_51[8] , 
        \wRegOut_7_84[29] , \wRegOut_7_84[30] , \ScanLink213[0] , 
        \wRegInTop_7_104[29] , \wRegOut_7_116[6] , \wRegInTop_7_104[30] , 
        \wRegInTop_7_127[18] , \wRegInTop_7_20[4] , \ScanLink173[5] , 
        \ScanLink0[13] , \wRegInTop_1_0[15] , \ScanLink24[18] , 
        \ScanLink50[8] , \ScanLink51[31] , \ScanLink72[19] , 
        \wRegInTop_6_61[17] , \ScanLink51[28] , \wRegOut_6_5[6] , 
        \wRegInTop_6_14[27] , \wRegInTop_6_42[26] , \wRegInTop_7_121[9] , 
        \wRegOut_7_124[20] , \wRegInBot_6_22[25] , \wRegInTop_7_39[26] , 
        \wRegInTop_6_37[16] , \wRegOut_7_107[11] , \wRegOut_6_4[12] , 
        \wRegInBot_6_57[15] , \wRegInBot_6_14[20] , \wRegInTop_6_22[22] , 
        \wRegInBot_6_37[11] , \wRegInBot_6_42[21] , \wRegInTop_6_57[12] , 
        \wRegEnTop_7_6[0] , \ScanLink219[19] , \wRegInTop_7_59[22] , 
        \wRegOut_7_112[25] , \wRegInBot_5_5[11] , \wRegInTop_5_19[16] , 
        \wRegInBot_5_19[11] , \wRegOut_6_6[5] , \wRegInBot_6_61[10] , 
        \ScanLink89[18] , \wRegInTop_7_94[26] , \wRegInTop_7_81[12] , 
        \wRegOut_6_27[19] , \wRegInTop_7_0[9] , \wRegOut_6_52[29] , 
        \wRegOut_7_29[29] , \wRegOut_7_115[5] , \wRegOut_6_10[9] , 
        \wRegOut_7_29[30] , \ScanLink210[3] , \wRegInTop_1_0[26] , 
        \wRegInTop_6_22[11] , \wRegInBot_6_42[12] , \wRegOut_6_52[30] , 
        \wRegInTop_7_23[7] , \ScanLink170[6] , \wRegInTop_7_59[11] , 
        \wRegOut_7_112[16] , \wRegInBot_6_28[3] , \wRegInBot_6_37[22] , 
        \wRegInTop_6_57[21] , \wRegInBot_6_61[23] , \wRegOut_3_1[3] , 
        \wRegInBot_6_14[13] , \wRegInTop_3_7[22] , \wRegInTop_4_15[2] , 
        \wRegOut_5_1[7] , \wRegInTop_6_14[14] , \wRegOut_7_124[13] , 
        \wRegOut_6_4[21] , \wRegInTop_6_37[25] , \wRegInTop_6_61[24] , 
        \wRegInBot_6_57[26] , \wRegInBot_6_22[16] , \wRegInTop_6_42[15] , 
        \wRegOut_7_107[22] , \wRegInTop_7_39[15] , \wRegInTop_7_96[6] , 
        \ScanLink29[3] , \wRegOut_7_56[8] , \ScanLink1[19] , \ScanLink0[20] , 
        \wRegInBot_3_2[31] , \wRegInBot_3_2[28] , \wRegOut_4_3[25] , 
        \wRegOut_7_99[1] , \wRegInTop_5_0[31] , \ScanLink117[1] , 
        \wRegInTop_7_44[0] , \wRegInTop_5_0[28] , \ScanLink114[2] , 
        \wRegInTop_7_47[3] , \wRegOut_1_0[0] , \wRegEnBot_2_0[0] , 
        \wRegOut_3_2[0] , \wRegInTop_4_4[8] , \wRegInBot_5_5[22] , 
        \wRegInTop_5_19[25] , \ScanLink127[28] , \ScanLink152[18] , 
        \ScanLink171[30] , \wRegOut_7_48[4] , \wRegInTop_7_81[21] , 
        \wRegInTop_7_95[5] , \ScanLink171[29] , \wRegInBot_2_0[7] , 
        \wRegOut_3_0[20] , \ScanLink19[22] , \wRegInTop_4_4[27] , 
        \wRegOut_5_2[4] , \wRegInBot_5_19[22] , \ScanLink127[31] , 
        \ScanLink104[19] , \wRegInTop_7_94[15] , \wRegOut_7_110[8] , 
        \ScanLink84[0] , \ScanLink212[26] , \wRegInBot_6_57[6] , 
        \wRegOut_6_15[4] , \ScanLink244[27] , \wRegOut_7_34[2] , 
        \wRegInTop_7_47[30] , \wRegInTop_7_64[18] , \ScanLink194[10] , 
        \ScanLink231[17] , \ScanLink251[13] , \ScanLink181[24] , 
        \ScanLink224[23] , \ScanLink9[6] , \wRegOut_4_8[30] , 
        \wRegOut_4_8[29] , \wRegOut_5_21[17] , \ScanLink56[6] , 
        \wRegOut_6_3[8] , \ScanLink79[26] , \wRegInTop_7_11[28] , 
        \wRegInTop_6_49[19] , \wRegInTop_7_47[29] , \wRegInTop_7_11[31] , 
        \wRegInTop_7_32[19] , \ScanLink207[12] , \wRegInTop_7_127[7] , 
        \wRegInTop_6_3[23] , \ScanLink208[1] , \wRegOut_5_17[12] , 
        \wRegInBot_6_6[30] , \wRegInTop_7_5[4] , \wRegInTop_5_12[29] , 
        \ScanLink55[5] , \wRegInBot_6_6[29] , \ScanLink168[4] , 
        \wRegOut_6_39[12] , \wRegOut_7_14[13] , \wRegOut_7_37[22] , 
        \wRegOut_7_61[23] , \wRegInTop_7_124[4] , \wRegOut_7_42[12] , 
        \wRegInTop_6_19[0] , \wRegOut_6_59[16] , \wRegInTop_7_6[7] , 
        \wRegOut_7_22[16] , \ScanLink97[13] , \wRegInTop_7_38[6] , 
        \wRegOut_7_57[26] , \wRegOut_7_74[17] , \wRegInBot_6_54[5] , 
        \wRegInBot_4_0[3] , \wRegInTop_4_1[5] , \wRegInTop_5_12[30] , 
        \wRegOut_6_16[7] , \wRegOut_7_37[1] , \wRegOut_5_17[21] , 
        \wRegInBot_5_18[8] , \wRegInTop_5_31[18] , \ScanLink82[27] , 
        \ScanLink87[3] , \ScanLink139[10] , \wRegInTop_7_25[9] , 
        \ScanLink159[14] , \ScanLink176[8] , \wRegOut_7_82[0] , 
        \ScanLink32[2] , \wRegOut_5_20[2] , \wRegOut_5_7[9] , 
        \wRegOut_5_21[24] , \wRegInTop_7_90[8] , \ScanLink4[22] , 
        \ScanLink4[11] , \wRegInTop_2_1[1] , \wRegInTop_6_3[10] , 
        \wRegInTop_2_2[2] , \wRegInBot_2_3[4] , \wRegOut_3_0[13] , 
        \wRegInBot_6_29[30] , \ScanLink181[17] , \ScanLink224[10] , 
        \wRegInTop_4_2[6] , \ScanLink19[11] , \wRegInTop_4_4[14] , 
        \ScanLink79[15] , \wRegInBot_6_29[29] , \wRegInBot_6_33[2] , 
        \wRegOut_7_50[6] , \ScanLink251[20] , \ScanLink207[21] , 
        \wRegInTop_6_63[8] , \ScanLink212[15] , \wRegOut_7_119[29] , 
        \ScanLink194[23] , \ScanLink231[24] , \ScanLink31[1] , 
        \wRegOut_5_7[19] , \ScanLink82[14] , \wRegInBot_6_30[1] , 
        \ScanLink159[27] , \ScanLink244[14] , \wRegOut_7_119[30] , 
        \wRegOut_7_53[5] , \wRegInBot_5_24[18] , \ScanLink97[20] , 
        \ScanLink139[23] , \wRegEnTop_7_12[0] , \wRegOut_7_57[15] , 
        \wRegOut_5_23[1] , \wRegOut_7_22[25] , \wRegOut_6_59[25] , 
        \wRegOut_7_74[24] , \wRegInBot_4_3[0] , \wRegOut_7_81[3] , 
        \wRegOut_7_61[10] , \wRegInBot_2_2[25] , \wRegOut_5_3[31] , 
        \wRegInTop_5_31[9] , \wRegOut_6_39[21] , \wRegOut_7_14[20] , 
        \wRegOut_7_37[11] , \wRegOut_7_42[21] , \wRegOut_5_3[28] , 
        \ScanLink128[26] , \wRegInBot_2_2[16] , \wRegOut_3_4[22] , 
        \ScanLink15[7] , \wRegOut_4_9[0] , \ScanLink86[25] , 
        \wRegInBot_5_20[30] , \wRegInBot_6_14[7] , \ScanLink93[11] , 
        \wRegInTop_7_8[22] , \wRegOut_6_56[5] , \wRegOut_7_77[3] , 
        \wRegInBot_5_20[29] , \ScanLink148[22] , \wRegEnTop_6_17[0] , 
        \wRegOut_6_28[24] , \wRegInTop_6_59[2] , \wRegOut_7_26[14] , 
        \wRegOut_7_53[24] , \wRegInTop_7_78[4] , \wRegOut_6_48[20] , 
        \wRegOut_7_10[11] , \wRegOut_7_70[15] , \wRegOut_7_65[21] , 
        \wRegOut_7_33[20] , \wRegOut_7_46[10] , \ScanLink16[4] , 
        \wRegOut_5_13[10] , \wRegOut_5_30[21] , \ScanLink128[6] , 
        \wRegOut_5_25[15] , \wRegInTop_6_7[21] , \wRegOut_6_48[9] , 
        \ScanLink248[3] , \wRegInBot_6_58[31] , \ScanLink255[11] , 
        \ScanLink185[26] , \ScanLink220[21] , \wRegInTop_4_0[25] , 
        \wRegInBot_6_58[28] , \ScanLink135[9] , \wRegInTop_7_66[8] , 
        \ScanLink203[10] , \wRegInTop_5_16[18] , \wRegInBot_5_21[1] , 
        \ScanLink68[10] , \wRegInBot_6_17[4] , \ScanLink216[24] , 
        \ScanLink240[25] , \wRegOut_6_48[13] , \wRegOut_6_55[6] , 
        \wRegOut_7_10[22] , \ScanLink190[12] , \wRegOut_7_74[0] , 
        \ScanLink235[15] , \wRegOut_7_65[12] , \wRegOut_7_46[23] , 
        \wRegOut_7_33[13] , \ScanLink180[8] , \wRegOut_7_53[17] , 
        \wRegInTop_7_100[2] , \ScanLink71[3] , \wRegOut_6_28[17] , 
        \wRegOut_7_26[27] , \wRegOut_7_70[26] , \wRegInTop_6_20[9] , 
        \ScanLink93[22] , \wRegInTop_7_8[11] , \ScanLink86[16] , 
        \ScanLink128[15] , \ScanLink148[11] , \wRegOut_7_13[7] , 
        \wRegOut_6_32[1] , \wRegOut_3_4[11] , \wRegInTop_4_0[16] , 
        \wRegInBot_6_9[8] , \ScanLink216[17] , \ScanLink68[23] , 
        \wRegInTop_7_15[19] , \ScanLink185[15] , \ScanLink190[21] , 
        \ScanLink235[26] , \ScanLink240[16] , \ScanLink220[12] , 
        \wRegInBot_5_1[13] , \wRegInTop_5_4[19] , \wRegOut_5_13[23] , 
        \wRegOut_5_25[26] , \wRegOut_6_31[2] , \wRegOut_7_10[4] , 
        \wRegInTop_7_36[31] , \ScanLink231[8] , \ScanLink255[22] , 
        \wRegInTop_6_38[18] , \wRegInTop_7_36[28] , \wRegInTop_7_60[29] , 
        \ScanLink203[23] , \wRegInTop_7_43[18] , \wRegInTop_7_60[30] , 
        \wRegInTop_6_7[12] , \wRegInBot_5_22[2] , \wRegOut_5_30[12] , 
        \wRegInTop_7_103[1] , \wRegInBot_6_2[18] , \ScanLink72[0] , 
        \wRegInTop_6_42[3] , \ScanLink130[4] , \wRegInTop_7_63[5] , 
        \wRegInBot_5_8[4] , \wRegInBot_6_12[9] , \wRegInTop_5_9[2] , 
        \ScanLink250[1] , \wRegInTop_3_3[13] , \ScanLink13[9] , 
        \wRegInTop_4_13[24] , \wRegInTop_7_85[10] , \wRegInTop_5_13[1] , 
        \ScanLink100[31] , \ScanLink123[19] , \ScanLink156[29] , 
        \wRegInBot_4_13[23] , \ScanLink100[28] , \ScanLink156[30] , 
        \wRegInTop_7_90[24] , \ScanLink175[18] , \wRegOut_5_8[17] , 
        \wRegInTop_5_10[2] , \wRegInBot_6_10[22] , \wRegInTop_6_26[20] , 
        \wRegInBot_6_33[13] , \wRegInTop_7_28[10] , \wRegInBot_6_46[23] , 
        \wRegInTop_6_53[10] , \wRegOut_7_116[27] , \wRegOut_6_0[10] , 
        \wRegInTop_6_10[25] , \wRegInBot_6_26[27] , \wRegInTop_6_46[24] , 
        \wRegOut_7_120[22] , \wRegInTop_6_33[14] , \wRegInTop_7_48[14] , 
        \wRegOut_7_103[13] , \wRegInBot_6_53[17] , \wRegInBot_3_6[19] , 
        \wRegInTop_6_41[0] , \ScanLink133[7] , \wRegInTop_7_60[6] , 
        \ScanLink253[2] , \wRegOut_4_7[14] , \wRegInTop_4_13[17] , 
        \wRegInBot_4_13[10] , \wRegInBot_6_9[14] , \wRegOut_6_53[8] , 
        \ScanLink186[6] , \wRegOut_5_8[24] , \wRegEnBot_6_25[0] , 
        \wRegInTop_7_85[23] , \wRegInTop_7_90[17] , \wRegOut_6_23[28] , 
        \wRegInTop_6_26[7] , \wRegOut_6_29[0] , \wRegOut_6_56[18] , 
        \ScanLink154[0] , \wRegOut_7_58[28] , \wRegInTop_3_3[20] , 
        \wRegOut_4_7[27] , \wRegInBot_5_1[20] , \wRegOut_7_58[31] , 
        \wRegOut_6_23[31] , \wRegOut_7_15[9] , \ScanLink234[5] , 
        \wRegOut_7_80[18] , \wRegInTop_7_100[18] , \wRegInTop_7_123[30] , 
        \wRegInBot_6_9[27] , \wRegInTop_6_25[4] , \wRegInTop_7_123[29] , 
        \ScanLink157[3] , \wRegInTop_7_118[0] , \wRegInBot_4_4[16] , 
        \ScanLink20[30] , \ScanLink69[1] , \wRegInTop_6_10[16] , 
        \ScanLink237[6] , \wRegOut_7_120[11] , \ScanLink20[29] , 
        \wRegOut_6_0[23] , \ScanLink76[28] , \wRegInTop_6_33[27] , 
        \wRegInBot_6_53[24] , \wRegInTop_7_48[27] , \wRegOut_5_12[30] , 
        \ScanLink55[19] , \wRegInTop_6_46[17] , \wRegOut_7_103[20] , 
        \ScanLink185[5] , \wRegOut_5_31[18] , \wRegInTop_6_6[18] , 
        \wRegInBot_6_10[11] , \ScanLink76[31] , \wRegInBot_6_26[14] , 
        \wRegInTop_6_26[13] , \wRegInBot_6_46[10] , \wRegOut_7_116[14] , 
        \wRegInBot_6_33[20] , \wRegInTop_6_53[23] , \wRegInTop_7_28[23] , 
        \ScanLink193[1] , \wRegOut_5_12[29] , \wRegInBot_6_3[12] , 
        \wRegOut_7_3[7] , \ScanLink69[30] , \ScanLink69[29] , 
        \wRegInBot_6_39[15] , \wRegInTop_7_74[17] , \wRegInTop_6_33[0] , 
        \wRegInTop_6_59[16] , \wRegInTop_7_22[16] , \wRegInTop_7_12[6] , 
        \wRegInTop_7_57[26] , \wRegInTop_6_39[12] , \ScanLink141[7] , 
        \wRegInTop_7_37[22] , \ScanLink202[29] , \wRegOut_7_124[4] , 
        \ScanLink254[31] , \wRegInBot_6_59[11] , \wRegInTop_7_42[12] , 
        \ScanLink202[30] , \ScanLink221[18] , \wRegOut_7_109[15] , 
        \wRegOut_5_2[11] , \wRegInTop_5_17[12] , \wRegInBot_5_21[10] , 
        \wRegOut_6_21[8] , \wRegInTop_7_14[13] , \wRegInTop_7_61[23] , 
        \ScanLink221[2] , \ScanLink254[28] , \ScanLink92[31] , 
        \ScanLink92[28] , \wRegInTop_6_30[3] , \wRegInTop_7_11[5] , 
        \ScanLink142[4] , \wRegEnTop_7_107[0] , \wRegInBot_5_17[15] , 
        \wRegInBot_6_60[9] , \wRegInTop_5_21[17] , \ScanLink222[1] , 
        \wRegOut_7_127[7] , \wRegOut_7_47[29] , \wRegInBot_1_0[24] , 
        \wRegInBot_3_0[8] , \wRegOut_3_5[31] , \ScanLink61[9] , 
        \wRegInTop_6_6[8] , \wRegOut_6_49[19] , \wRegOut_7_0[4] , 
        \wRegOut_7_11[31] , \wRegOut_7_11[28] , \wRegOut_7_32[19] , 
        \ScanLink190[2] , \wRegOut_7_47[30] , \wRegOut_7_64[18] , 
        \wRegInTop_7_110[8] , \wRegInTop_6_39[21] , \wRegOut_7_5[15] , 
        \wRegInBot_6_59[22] , \wRegInTop_7_42[21] , \wRegOut_7_109[26] , 
        \ScanLink125[3] , \wRegOut_3_5[28] , \wRegInTop_6_57[4] , 
        \wRegInTop_7_14[20] , \wRegInTop_7_37[11] , \wRegInTop_7_76[2] , 
        \wRegInTop_7_61[10] , \wRegInBot_4_4[25] , \wRegOut_4_7[6] , 
        \wRegInBot_6_3[21] , \wRegInBot_6_39[26] , \wRegInTop_7_22[25] , 
        \wRegInTop_7_57[15] , \ScanLink191[18] , \wRegInTop_7_74[24] , 
        \ScanLink245[6] , \wRegEnTop_7_38[0] , \wRegInTop_6_59[25] , 
        \ScanLink18[2] , \wRegOut_4_4[5] , \wRegEnTop_5_4[0] , 
        \wRegEnBot_6_57[0] , \wRegOut_6_58[3] , \wRegOut_7_79[5] , 
        \wRegOut_5_2[22] , \wRegInTop_5_2[9] , \wRegInBot_6_19[2] , 
        \wRegInTop_6_49[8] , \wRegOut_7_5[26] , \wRegInBot_5_17[26] , 
        \wRegInTop_5_21[24] , \wRegInBot_5_21[23] , \wRegInTop_6_54[7] , 
        \ScanLink126[0] , \wRegInTop_7_75[1] , \wRegInTop_7_9[31] , 
        \ScanLink149[28] , \ScanLink21[23] , \wRegInTop_5_17[21] , 
        \wRegInTop_7_9[28] , \wRegInBot_6_2[3] , \ScanLink149[31] , 
        \wRegOut_7_67[9] , \ScanLink246[5] , \wRegOut_6_1[29] , 
        \wRegInBot_1_0[17] , \wRegOut_2_1[27] , \ScanLink5[28] , 
        \wRegInBot_3_7[20] , \ScanLink17[26] , \ScanLink54[13] , 
        \wRegInTop_6_3[5] , \wRegInTop_6_28[1] , \ScanLink209[16] , 
        \wRegOut_6_1[30] , \ScanLink77[22] , \wRegInBot_4_15[0] , 
        \ScanLink34[17] , \ScanLink62[16] , \wRegInTop_7_29[30] , 
        \wRegInTop_6_52[30] , \ScanLink41[27] , \wRegInTop_6_27[19] , 
        \wRegInTop_7_115[5] , \wRegInTop_7_29[29] , \ScanLink64[4] , 
        \wRegInTop_6_52[29] , \wRegOut_7_5[9] , \wRegInTop_7_14[8] , 
        \ScanLink188[0] , \wRegInTop_7_122[23] , \ScanLink147[9] , 
        \wRegOut_7_81[12] , \wRegOut_5_19[16] , \wRegInTop_7_101[12] , 
        \wRegInBot_5_29[9] , \wRegOut_6_27[6] , \wRegOut_7_94[26] , 
        \wRegInTop_7_114[26] , \ScanLink5[31] , \wRegInTop_3_2[19] , 
        \wRegInTop_5_5[20] , \wRegOut_6_22[22] , \wRegOut_6_57[12] , 
        \wRegOut_7_59[22] , \wRegOut_6_42[26] , \wRegInTop_6_0[6] , 
        \wRegInBot_6_1[0] , \wRegOut_6_14[27] , \wRegOut_6_37[16] , 
        \wRegOut_7_39[26] , \wRegOut_7_121[9] , \wRegOut_6_61[17] , 
        \wRegEnTop_7_96[0] , \wRegOut_6_24[5] , \ScanLink101[11] , 
        \ScanLink174[21] , \ScanLink157[10] , \ScanLink67[7] , 
        \ScanLink122[20] , \ScanLink159[5] , \ScanLink142[24] , 
        \wRegInTop_7_116[6] , \ScanLink99[17] , \wRegInTop_7_2[24] , 
        \ScanLink137[14] , \wRegInTop_7_84[30] , \ScanLink114[25] , 
        \ScanLink161[15] , \wRegInTop_7_84[29] , \wRegOut_7_94[15] , 
        \ScanLink239[0] , \wRegInTop_7_114[15] , \wRegInBot_3_6[6] , 
        \wRegInTop_3_7[0] , \wRegInBot_3_7[13] , \wRegOut_5_19[25] , 
        \wRegInTop_7_122[10] , \wRegOut_6_43[2] , \wRegOut_7_81[21] , 
        \wRegOut_7_62[4] , \wRegInTop_7_101[21] , \ScanLink62[25] , 
        \ScanLink243[8] , \wRegInBot_6_11[28] , \ScanLink17[15] , 
        \wRegInBot_6_47[30] , \wRegOut_4_1[8] , \ScanLink34[24] , 
        \ScanLink41[14] , \wRegInBot_6_11[31] , \wRegInBot_6_32[19] , 
        \wRegOut_5_12[0] , \ScanLink54[20] , \wRegInBot_6_47[29] , 
        \ScanLink209[25] , \wRegOut_7_121[31] , \wRegOut_2_1[14] , 
        \wRegInTop_3_4[3] , \ScanLink21[10] , \wRegInBot_5_6[2] , 
        \wRegOut_7_102[19] , \wRegInTop_5_7[4] , \ScanLink77[11] , 
        \wRegOut_7_121[28] , \ScanLink114[16] , \ScanLink137[27] , 
        \ScanLink142[17] , \wRegInBot_3_5[5] , \ScanLink99[24] , 
        \wRegInTop_7_2[17] , \wRegInBot_4_12[30] , \wRegInBot_4_12[29] , 
        \wRegInTop_5_4[7] , \wRegInBot_5_5[1] , \ScanLink101[22] , 
        \ScanLink161[26] , \ScanLink174[12] , \wRegOut_5_11[3] , 
        \ScanLink122[13] , \ScanLink157[23] , \wRegInBot_5_0[19] , 
        \wRegInTop_5_5[13] , \wRegOut_6_37[25] , \wRegOut_6_14[14] , 
        \wRegOut_6_42[15] , \wRegInTop_6_52[9] , \wRegOut_7_39[15] , 
        \wRegOut_6_61[24] , \wRegInBot_3_3[22] , \wRegInTop_3_6[31] , 
        \ScanLink27[5] , \wRegOut_6_22[11] , \wRegOut_6_40[1] , 
        \wRegOut_7_59[11] , \wRegOut_7_61[7] , \wRegOut_6_57[21] , 
        \ScanLink146[26] , \wRegOut_4_14[3] , \ScanLink133[16] , 
        \wRegInTop_5_1[22] , \wRegInBot_5_18[31] , \wRegInBot_5_18[28] , 
        \ScanLink88[21] , \ScanLink110[27] , \wRegInTop_7_6[26] , 
        \ScanLink165[17] , \wRegOut_7_97[7] , \ScanLink170[23] , 
        \ScanLink105[13] , \ScanLink153[12] , \wRegOut_6_46[24] , 
        \ScanLink119[7] , \ScanLink126[22] , \wRegInBot_5_4[31] , 
        \wRegInBot_5_4[28] , \wRegOut_6_10[25] , \wRegInBot_6_26[5] , 
        \wRegOut_6_33[14] , \wRegOut_7_48[14] , \wRegOut_7_45[1] , 
        \wRegOut_6_26[20] , \ScanLink104[8] , \wRegOut_6_53[10] , 
        \wRegOut_7_28[10] , \wRegInTop_7_98[0] , \wRegInTop_6_9[25] , 
        \wRegInTop_7_57[9] , \wRegInBot_6_25[6] , \wRegOut_7_90[24] , 
        \wRegInTop_7_110[24] , \wRegOut_7_46[2] , \wRegInTop_3_6[28] , 
        \ScanLink39[9] , \wRegOut_7_85[10] , \wRegInTop_7_126[21] , 
        \ScanLink13[24] , \wRegOut_4_13[24] , \wRegInTop_7_105[10] , 
        \ScanLink24[6] , \ScanLink30[15] , \ScanLink66[14] , 
        \wRegInBot_6_15[19] , \wRegInBot_6_38[9] , \wRegInBot_6_60[29] , 
        \wRegInBot_6_36[31] , \wRegInBot_6_43[18] , \wRegOut_7_94[4] , 
        \wRegInBot_6_60[30] , \ScanLink45[25] , \wRegInBot_6_36[28] , 
        \ScanLink25[21] , \ScanLink218[20] , \wRegOut_7_106[28] , 
        \ScanLink50[11] , \wRegInTop_7_49[5] , \ScanLink73[20] , 
        \wRegOut_7_106[31] , \wRegOut_7_125[19] , \wRegInBot_6_42[1] , 
        \wRegOut_7_21[5] , \ScanLink200[9] , \wRegInTop_2_2[27] , 
        \wRegInTop_2_2[14] , \wRegInBot_3_3[11] , \ScanLink13[17] , 
        \ScanLink25[12] , \wRegInTop_5_1[11] , \wRegOut_6_26[13] , 
        \ScanLink91[7] , \wRegOut_7_28[23] , \wRegOut_6_33[27] , 
        \wRegOut_6_53[23] , \wRegOut_7_48[27] , \ScanLink40[2] , 
        \wRegInBot_5_10[0] , \ScanLink43[1] , \wRegInBot_5_13[3] , 
        \wRegOut_6_10[16] , \wRegOut_6_46[17] , \ScanLink88[12] , 
        \ScanLink105[20] , \ScanLink170[10] , \ScanLink126[11] , 
        \ScanLink153[21] , \wRegOut_7_118[0] , \ScanLink110[14] , 
        \ScanLink133[25] , \wRegEnTop_7_60[0] , \ScanLink146[15] , 
        \wRegInTop_7_80[18] , \wRegInTop_7_6[15] , \ScanLink165[24] , 
        \ScanLink50[22] , \wRegOut_6_5[18] , \ScanLink66[27] , 
        \ScanLink73[13] , \wRegInTop_7_58[31] , \wRegOut_4_13[17] , 
        \ScanLink30[26] , \ScanLink45[16] , \wRegInTop_6_23[31] , 
        \wRegInTop_6_56[18] , \ScanLink218[13] , \wRegInTop_7_58[28] , 
        \wRegOut_6_8[3] , \wRegInTop_6_23[28] , \ScanLink92[4] , 
        \wRegInTop_7_126[12] , \wRegInBot_6_41[2] , \wRegOut_7_85[23] , 
        \wRegOut_7_22[6] , \wRegInTop_7_105[23] , \wRegOut_5_6[13] , 
        \wRegInBot_5_13[17] , \wRegInTop_5_21[3] , \wRegInTop_6_9[16] , 
        \wRegInTop_6_11[8] , \wRegOut_7_90[17] , \wRegInTop_7_110[17] , 
        \wRegOut_7_1[17] , \wRegOut_7_91[9] , \wRegInTop_7_83[1] , 
        \wRegInTop_5_25[15] , \wRegInBot_5_30[26] , \wRegOut_6_62[9] , 
        \wRegOut_3_1[19] , \wRegInBot_4_0[14] , \wRegInTop_5_13[10] , 
        \wRegInBot_5_25[12] , \wRegInTop_5_30[21] , \ScanLink102[6] , 
        \ScanLink138[29] , \ScanLink138[30] , \wRegInTop_7_51[7] , 
        \wRegInBot_6_23[8] , \wRegInBot_6_28[23] , \wRegInTop_6_48[20] , 
        \wRegInTop_7_33[20] , \wRegInTop_7_46[10] , \ScanLink22[8] , 
        \wRegOut_5_30[8] , \wRegInBot_6_7[10] , \wRegInTop_6_28[24] , 
        \wRegInBot_6_48[27] , \wRegInTop_7_10[11] , \wRegInTop_7_26[14] , 
        \wRegInTop_7_65[21] , \ScanLink195[29] , \wRegInTop_7_70[15] , 
        \wRegInTop_7_52[4] , \ScanLink195[30] , \wRegInTop_7_53[24] , 
        \wRegOut_7_118[23] , \ScanLink101[5] , \wRegOut_4_9[10] , 
        \wRegInTop_5_22[0] , \wRegInTop_5_30[12] , \wRegInTop_7_80[2] , 
        \ScanLink97[9] , \wRegOut_7_103[1] , \wRegOut_5_6[20] , 
        \wRegInTop_5_13[23] , \wRegInBot_5_25[21] , \ScanLink58[0] , 
        \ScanLink96[19] , \ScanLink206[7] , \wRegInBot_5_13[24] , 
        \wRegInTop_5_25[26] , \wRegInBot_5_30[15] , \wRegInTop_6_14[5] , 
        \wRegInTop_7_35[3] , \wRegOut_6_38[18] , \wRegOut_7_36[28] , 
        \ScanLink166[2] , \wRegOut_7_43[18] , \wRegOut_7_60[30] , 
        \wRegOut_0_0[6] , \wRegInBot_0_0[30] , \ScanLink4[3] , 
        \wRegInBot_6_59[0] , \wRegOut_7_36[31] , \wRegOut_7_15[19] , 
        \wRegOut_7_60[29] , \wRegInBot_0_0[29] , \wRegOut_7_1[24] , 
        \wRegInBot_0_0[20] , \wRegOut_1_0[9] , \wRegOut_2_1[5] , 
        \ScanLink7[0] , \wRegInTop_6_2[29] , \wRegInTop_3_2[10] , 
        \wRegInBot_4_0[27] , \ScanLink18[31] , \ScanLink18[28] , 
        \wRegOut_4_9[23] , \wRegInTop_6_2[30] , \wRegOut_6_18[1] , 
        \wRegOut_7_39[7] , \wRegInBot_6_7[23] , \ScanLink89[5] , 
        \wRegOut_5_16[18] , \wRegInTop_7_70[26] , \wRegInBot_6_48[14] , 
        \wRegOut_7_24[8] , \ScanLink205[4] , \wRegInTop_6_17[6] , 
        \wRegInTop_6_28[17] , \wRegInTop_7_53[17] , \wRegOut_7_100[2] , 
        \wRegOut_7_118[10] , \wRegInTop_6_48[13] , \wRegInTop_7_8[1] , 
        \wRegInTop_7_26[27] , \ScanLink165[1] , \wRegInTop_7_46[23] , 
        \ScanLink206[18] , \ScanLink225[30] , \wRegInBot_6_28[10] , 
        \wRegInTop_7_10[22] , \wRegInTop_7_33[13] , \wRegInTop_7_36[0] , 
        \wRegInTop_7_65[12] , \ScanLink250[19] , \ScanLink225[29] , 
        \wRegOut_4_6[17] , \wRegInBot_6_8[17] , \wRegOut_7_81[31] , 
        \wRegOut_7_81[28] , \wRegInTop_7_101[31] , \wRegInTop_7_122[19] , 
        \ScanLink243[1] , \wRegInTop_7_101[28] , \ScanLink21[19] , 
        \ScanLink54[29] , \wRegInBot_6_27[24] , \wRegInTop_6_47[27] , 
        \wRegInTop_6_51[3] , \ScanLink123[4] , \wRegInTop_7_70[5] , 
        \wRegInTop_6_32[17] , \wRegInTop_7_49[17] , \wRegOut_5_12[9] , 
        \wRegOut_7_102[10] , \wRegOut_6_1[13] , \wRegInBot_6_52[14] , 
        \ScanLink5[21] , \ScanLink5[12] , \wRegOut_2_2[6] , \wRegInTop_3_7[9] , 
        \ScanLink54[30] , \ScanLink77[18] , \wRegInTop_6_11[26] , 
        \wRegOut_7_121[21] , \wRegOut_4_1[1] , \wRegInBot_6_11[21] , 
        \wRegInTop_6_27[23] , \wRegInBot_6_32[10] , \wRegInTop_7_29[13] , 
        \wRegInBot_6_47[20] , \wRegInTop_6_52[13] , \wRegOut_7_117[24] , 
        \wRegEnTop_3_1[0] , \wRegInBot_4_12[20] , \wRegInBot_5_5[8] , 
        \wRegInTop_7_91[27] , \wRegOut_5_9[14] , \wRegInTop_7_84[13] , 
        \wRegOut_4_2[2] , \wRegInTop_4_12[27] , \wRegInBot_5_0[10] , 
        \wRegOut_6_40[8] , \ScanLink240[2] , \wRegInTop_3_2[23] , 
        \wRegInBot_4_15[9] , \wRegInBot_6_11[12] , \wRegOut_6_22[18] , 
        \wRegOut_6_57[31] , \wRegOut_7_59[18] , \wRegInTop_6_52[0] , 
        \wRegOut_6_57[28] , \ScanLink120[7] , \wRegInTop_7_73[6] , 
        \wRegInTop_6_27[10] , \wRegInBot_6_47[13] , \wRegOut_7_117[17] , 
        \wRegInBot_5_29[0] , \wRegOut_6_1[20] , \wRegInTop_6_32[24] , 
        \wRegInBot_6_32[23] , \wRegInTop_6_52[20] , \wRegOut_7_5[0] , 
        \wRegInTop_7_29[20] , \wRegEnBot_6_7[0] , \wRegInTop_6_11[15] , 
        \wRegInBot_6_27[17] , \wRegInTop_6_28[8] , \wRegInTop_6_47[14] , 
        \wRegInBot_6_52[27] , \wRegInTop_7_49[24] , \wRegOut_7_102[23] , 
        \ScanLink195[6] , \wRegEnBot_6_36[0] , \ScanLink227[5] , 
        \wRegOut_7_121[12] , \wRegInTop_7_108[3] , \wRegOut_7_122[3] , 
        \wRegInBot_3_7[30] , \ScanLink79[2] , \wRegInBot_3_7[29] , 
        \wRegOut_4_6[24] , \wRegInBot_6_8[24] , \wRegInTop_6_35[7] , 
        \wRegInTop_7_14[1] , \ScanLink188[9] , \ScanLink147[0] , 
        \wRegInTop_5_5[30] , \wRegInTop_5_5[29] , \wRegOut_7_121[0] , 
        \wRegEnTop_7_59[0] , \ScanLink224[6] , \wRegInBot_2_3[26] , 
        \wRegInBot_3_0[1] , \wRegInTop_3_1[7] , \wRegOut_3_5[21] , 
        \wRegInTop_4_1[26] , \wRegInTop_4_12[14] , \wRegInBot_5_0[23] , 
        \wRegInTop_6_36[4] , \ScanLink144[3] , \wRegInTop_7_17[2] , 
        \wRegOut_7_6[3] , \wRegOut_7_18[5] , \wRegInTop_7_84[20] , 
        \ScanLink239[9] , \wRegInBot_4_12[13] , \wRegOut_6_39[3] , 
        \ScanLink174[28] , \wRegOut_5_9[27] , \wRegInBot_6_1[9] , 
        \ScanLink101[18] , \ScanLink122[30] , \ScanLink157[19] , 
        \ScanLink174[31] , \wRegInTop_7_91[14] , \ScanLink69[13] , 
        \ScanLink122[29] , \ScanLink196[5] , \ScanLink241[26] , 
        \wRegOut_6_45[5] , \ScanLink191[11] , \wRegOut_7_64[3] , 
        \ScanLink234[16] , \wRegInTop_6_39[31] , \wRegInTop_6_39[28] , 
        \ScanLink217[27] , \wRegInTop_7_14[30] , \wRegInTop_7_37[18] , 
        \wRegInTop_7_42[28] , \ScanLink202[13] , \wRegInTop_7_14[29] , 
        \wRegInTop_7_42[31] , \wRegInTop_7_61[19] , \ScanLink254[12] , 
        \ScanLink184[25] , \ScanLink221[22] , \wRegInBot_5_0[5] , 
        \wRegInTop_6_6[22] , \wRegInTop_5_1[3] , \wRegOut_5_14[7] , 
        \wRegOut_5_24[16] , \wRegOut_5_31[22] , \ScanLink138[5] , 
        \wRegInBot_6_3[28] , \wRegOut_5_12[13] , \wRegInBot_6_3[31] , 
        \wRegInTop_3_2[4] , \wRegInTop_5_2[0] , \wRegInBot_5_3[6] , 
        \wRegOut_5_17[4] , \wRegOut_6_49[23] , \wRegOut_7_32[23] , 
        \wRegOut_7_11[12] , \wRegOut_7_47[13] , \wRegOut_7_64[22] , 
        \wRegInBot_3_3[2] , \wRegOut_7_71[16] , \wRegInTop_5_17[31] , 
        \wRegOut_6_29[27] , \wRegInTop_6_49[1] , \wRegOut_7_27[17] , 
        \wRegOut_7_52[27] , \wRegInTop_7_68[7] , \wRegInTop_5_17[28] , 
        \ScanLink149[21] , \ScanLink92[12] , \wRegOut_6_46[6] , 
        \wRegInTop_7_9[21] , \wRegOut_7_67[0] , \wRegInBot_2_3[15] , 
        \wRegOut_3_5[12] , \wRegInBot_4_13[7] , \wRegInTop_5_18[3] , 
        \ScanLink87[26] , \wRegOut_5_31[11] , \ScanLink126[9] , 
        \ScanLink129[25] , \wRegInTop_7_75[8] , \wRegOut_5_12[20] , 
        \ScanLink62[3] , \wRegInTop_7_113[2] , \wRegOut_5_24[25] , 
        \wRegInBot_6_4[4] , \wRegInTop_6_6[11] , \wRegInTop_6_5[2] , 
        \ScanLink193[8] , \wRegInBot_6_59[18] , \ScanLink202[20] , 
        \ScanLink184[16] , \ScanLink221[11] , \wRegInTop_4_1[15] , 
        \wRegEnTop_4_10[0] , \wRegOut_6_21[1] , \wRegInBot_6_63[3] , 
        \ScanLink254[21] , \ScanLink69[20] , \wRegInTop_6_33[9] , 
        \ScanLink191[22] , \ScanLink217[14] , \ScanLink234[25] , 
        \ScanLink241[15] , \ScanLink87[15] , \wRegInBot_6_60[0] , 
        \ScanLink222[8] , \wRegInBot_4_10[4] , \wRegOut_5_2[18] , 
        \wRegInBot_5_21[19] , \wRegOut_6_22[2] , \ScanLink129[16] , 
        \ScanLink92[21] , \ScanLink149[12] , \wRegInTop_7_9[12] , 
        \wRegOut_7_52[14] , \wRegOut_7_71[25] , \wRegInTop_7_110[1] , 
        \ScanLink61[0] , \wRegInBot_5_31[2] , \wRegOut_6_29[14] , 
        \wRegInBot_6_7[7] , \wRegOut_7_27[24] , \wRegOut_5_6[30] , 
        \wRegOut_5_6[29] , \wRegInTop_6_6[1] , \wRegOut_6_49[10] , 
        \wRegOut_7_47[20] , \wRegOut_7_11[21] , \wRegOut_7_32[10] , 
        \wRegOut_7_64[11] , \ScanLink83[24] , \ScanLink158[17] , 
        \wRegInBot_5_25[31] , \wRegInBot_5_25[28] , \ScanLink58[9] , 
        \ScanLink97[0] , \wRegOut_7_103[8] , \ScanLink138[13] , 
        \ScanLink96[10] , \wRegInBot_6_44[6] , \wRegOut_7_27[2] , 
        \wRegOut_6_58[15] , \wRegOut_7_23[15] , \wRegOut_7_75[14] , 
        \wRegInBot_0_0[13] , \ScanLink7[9] , \ScanLink45[6] , 
        \wRegInBot_5_15[4] , \wRegInTop_7_28[5] , \wRegOut_7_56[25] , 
        \wRegOut_6_38[11] , \wRegOut_7_36[21] , \wRegOut_7_43[11] , 
        \wRegOut_5_16[11] , \wRegInBot_6_59[9] , \wRegOut_7_15[10] , 
        \ScanLink178[7] , \wRegOut_7_60[20] , \wRegOut_3_1[23] , 
        \ScanLink46[5] , \wRegInBot_5_16[7] , \wRegInTop_6_2[20] , 
        \wRegOut_6_18[8] , \ScanLink218[2] , \wRegOut_5_20[14] , 
        \wRegInBot_6_28[19] , \wRegInTop_7_8[8] , \wRegInTop_7_36[9] , 
        \ScanLink165[8] , \ScanLink206[11] , \ScanLink180[27] , 
        \ScanLink225[20] , \ScanLink250[10] , \ScanLink18[21] , 
        \ScanLink78[25] , \wRegInBot_6_47[5] , \wRegInTop_4_5[24] , 
        \wRegEnTop_5_15[0] , \ScanLink245[24] , \wRegOut_7_24[1] , 
        \ScanLink195[13] , \ScanLink230[14] , \wRegOut_7_118[19] , 
        \ScanLink21[2] , \ScanLink94[3] , \ScanLink213[25] , 
        \wRegOut_6_38[22] , \wRegOut_7_15[23] , \wRegOut_7_36[12] , 
        \wRegOut_7_43[22] , \wRegInTop_7_83[8] , \wRegOut_7_60[13] , 
        \wRegOut_7_56[16] , \wRegOut_7_75[27] , \wRegOut_7_91[0] , 
        \wRegOut_7_23[26] , \ScanLink1[23] , \ScanLink1[10] , 
        \wRegOut_3_1[10] , \ScanLink18[12] , \wRegOut_4_12[4] , 
        \wRegOut_5_9[6] , \wRegInTop_5_30[28] , \wRegOut_6_58[26] , 
        \ScanLink138[20] , \wRegInTop_5_13[19] , \wRegInTop_5_30[31] , 
        \ScanLink96[23] , \ScanLink83[17] , \wRegInBot_6_20[2] , 
        \wRegOut_6_62[0] , \wRegOut_7_43[6] , \ScanLink158[24] , 
        \ScanLink195[20] , \ScanLink230[27] , \wRegInTop_4_5[17] , 
        \ScanLink213[16] , \ScanLink245[17] , \wRegInTop_6_48[30] , 
        \wRegInTop_6_48[29] , \ScanLink206[22] , \wRegInTop_7_33[29] , 
        \wRegInTop_7_46[19] , \wRegInTop_7_65[31] , \ScanLink180[14] , 
        \ScanLink225[13] , \ScanLink22[1] , \wRegOut_4_11[7] , 
        \wRegOut_5_20[27] , \wRegInTop_5_22[9] , \ScanLink78[16] , 
        \wRegInTop_7_10[18] , \wRegInBot_6_23[1] , \wRegOut_6_61[3] , 
        \wRegInTop_7_33[30] , \wRegOut_7_40[5] , \ScanLink250[23] , 
        \wRegInTop_7_65[28] , \wRegInTop_6_2[13] , \wRegInBot_6_7[19] , 
        \wRegOut_5_30[1] , \wRegOut_4_9[19] , \wRegOut_5_16[22] , 
        \wRegInTop_5_1[18] , \wRegOut_7_92[3] , \wRegInBot_5_4[12] , 
        \wRegInTop_6_12[2] , \wRegInBot_6_42[8] , \ScanLink160[5] , 
        \wRegInTop_7_33[4] , \ScanLink200[0] , \ScanLink1[7] , \ScanLink2[4] , 
        \wRegInTop_5_18[15] , \wRegInTop_7_80[11] , \wRegOut_7_105[6] , 
        \wRegInBot_5_18[12] , \ScanLink105[29] , \wRegInTop_1_1[16] , 
        \ScanLink43[8] , \ScanLink105[30] , \ScanLink153[31] , 
        \wRegInTop_7_95[25] , \ScanLink170[19] , \ScanLink126[18] , 
        \ScanLink153[28] , \wRegOut_7_118[9] , \wRegInBot_5_10[9] , 
        \wRegInBot_6_15[23] , \wRegInTop_6_23[21] , \wRegInBot_6_36[12] , 
        \wRegInBot_6_60[13] , \wRegInBot_6_43[22] , \wRegInTop_6_56[11] , 
        \wRegInTop_7_58[21] , \wRegOut_7_113[26] , \wRegInTop_6_43[25] , 
        \wRegOut_6_5[11] , \wRegInBot_6_23[26] , \wRegInTop_6_36[15] , 
        \wRegInTop_7_38[25] , \wRegInBot_6_56[16] , \wRegOut_7_106[12] , 
        \wRegInTop_6_60[14] , \wRegInBot_3_3[18] , \wRegInTop_3_6[12] , 
        \wRegInTop_6_15[24] , \wRegOut_7_125[23] , \wRegInTop_6_11[1] , 
        \ScanLink163[6] , \wRegInTop_7_30[7] , \wRegOut_7_106[5] , 
        \wRegOut_4_2[15] , \wRegInTop_5_18[26] , \wRegInBot_5_18[21] , 
        \ScanLink88[28] , \ScanLink203[3] , \wRegInTop_5_27[4] , 
        \wRegInTop_7_95[16] , \ScanLink88[31] , \wRegInTop_7_85[6] , 
        \wRegOut_7_58[7] , \wRegInTop_7_80[22] , \wRegInTop_1_1[25] , 
        \wRegInTop_3_6[21] , \wRegOut_4_2[26] , \wRegInBot_4_8[2] , 
        \wRegInTop_4_9[4] , \wRegInBot_5_4[21] , \wRegOut_5_28[3] , 
        \wRegOut_6_26[30] , \wRegOut_6_26[29] , \ScanLink104[1] , 
        \wRegOut_6_53[19] , \wRegOut_7_28[19] , \wRegInTop_7_98[9] , 
        \wRegInTop_7_57[0] , \wRegEnBot_5_27[0] , \wRegOut_7_45[8] , 
        \ScanLink107[2] , \wRegInTop_7_54[3] , \wRegInTop_7_126[28] , 
        \wRegOut_7_85[19] , \wRegInTop_7_105[19] , \wRegOut_7_89[2] , 
        \wRegInTop_7_126[31] , \ScanLink25[31] , \ScanLink25[28] , 
        \ScanLink39[0] , \wRegOut_6_5[22] , \wRegInTop_6_36[26] , 
        \wRegInBot_6_56[25] , \wRegOut_7_106[21] , \ScanLink50[18] , 
        \wRegInTop_6_43[16] , \wRegInTop_7_38[16] , \ScanLink73[30] , 
        \wRegInTop_7_86[5] , \wRegInTop_6_15[17] , \wRegInBot_6_23[15] , 
        \wRegOut_7_125[10] , \wRegInTop_5_24[7] , \ScanLink73[29] , 
        \wRegInTop_6_60[27] , \wRegInBot_6_15[10] , \wRegInBot_6_38[0] , 
        \wRegInBot_6_60[20] , \wRegInTop_2_1[8] , \wRegInTop_4_13[5] , 
        \wRegOut_5_7[0] , \wRegInTop_6_23[12] , \wRegInBot_6_43[11] , 
        \wRegInTop_7_58[12] , \ScanLink218[30] , \wRegOut_7_113[15] , 
        \wRegInBot_6_36[21] , \wRegInTop_6_56[22] , \ScanLink218[29] , 
        \wRegInTop_7_90[1] , \wRegInTop_6_3[19] , \wRegInTop_2_3[17] , 
        \wRegOut_3_7[4] , \wRegEnBot_4_5[0] , \wRegOut_5_17[28] , 
        \wRegInBot_4_1[17] , \ScanLink19[18] , \wRegOut_4_8[13] , 
        \wRegOut_7_82[9] , \wRegOut_5_17[31] , \wRegInBot_6_6[13] , 
        \wRegInTop_6_29[27] , \wRegInBot_6_49[24] , \wRegInTop_7_27[17] , 
        \wRegInTop_7_42[7] , \wRegInTop_7_52[27] , \wRegOut_7_119[20] , 
        \wRegInTop_6_63[1] , \ScanLink111[6] , \wRegInTop_7_71[16] , 
        \wRegInTop_7_11[12] , \ScanLink207[31] , \ScanLink224[19] , 
        \wRegInTop_5_12[13] , \wRegInBot_6_29[20] , \wRegInTop_6_49[23] , 
        \wRegInTop_7_64[22] , \ScanLink251[29] , \wRegInTop_7_32[23] , 
        \ScanLink207[28] , \wRegInTop_7_47[13] , \ScanLink251[30] , 
        \ScanLink97[29] , \wRegOut_3_0[30] , \wRegOut_3_0[29] , 
        \wRegOut_3_4[7] , \wRegInBot_4_3[9] , \wRegInTop_4_10[6] , 
        \wRegOut_5_4[3] , \wRegOut_5_7[10] , \wRegInBot_5_12[14] , 
        \wRegInTop_5_24[16] , \wRegInBot_5_24[11] , \wRegInTop_5_31[22] , 
        \ScanLink97[30] , \ScanLink112[5] , \wRegInBot_5_31[25] , 
        \wRegInTop_6_60[2] , \wRegInTop_7_41[4] , \wRegInBot_6_30[8] , 
        \wRegOut_6_39[31] , \wRegOut_7_42[31] , \wRegOut_7_61[19] , 
        \ScanLink31[8] , \wRegInTop_5_31[0] , \wRegOut_7_14[29] , 
        \wRegOut_6_39[28] , \wRegOut_7_14[30] , \wRegOut_7_42[28] , 
        \wRegInTop_7_93[2] , \wRegOut_7_37[18] , \wRegOut_5_23[8] , 
        \wRegOut_7_0[14] , \wRegInTop_7_64[11] , \wRegInBot_4_1[24] , 
        \wRegInTop_6_49[10] , \wRegInTop_7_11[21] , \wRegInTop_7_47[20] , 
        \ScanLink175[2] , \wRegOut_4_8[20] , \ScanLink84[9] , 
        \wRegInTop_6_29[14] , \wRegInBot_6_29[13] , \wRegInBot_6_49[17] , 
        \wRegInTop_7_26[3] , \wRegInTop_7_32[10] , \wRegInTop_7_52[14] , 
        \wRegOut_7_119[13] , \wRegOut_7_110[1] , \wRegInTop_7_27[24] , 
        \ScanLink194[19] , \wRegInTop_7_71[25] , \ScanLink215[7] , 
        \wRegOut_6_3[1] , \wRegInBot_6_6[20] , \wRegInTop_6_19[9] , 
        \ScanLink99[6] , \wRegOut_7_0[27] , \wRegOut_7_29[4] , 
        \ScanLink208[8] , \ScanLink0[30] , \wRegInTop_2_3[24] , 
        \wRegOut_5_7[23] , \wRegInTop_5_24[25] , \wRegOut_6_0[2] , 
        \wRegInBot_6_49[3] , \wRegInBot_5_31[16] , \wRegInTop_7_25[0] , 
        \ScanLink176[1] , \wRegInTop_5_12[20] , \wRegInBot_5_12[27] , 
        \wRegInBot_5_18[1] , \wRegInTop_5_31[11] , \wRegOut_7_37[8] , 
        \ScanLink216[4] , \wRegOut_7_113[2] , \wRegInBot_3_2[21] , 
        \ScanLink12[27] , \ScanLink24[22] , \ScanLink48[3] , 
        \wRegInBot_5_24[22] , \ScanLink139[19] , \wRegOut_6_4[31] , 
        \ScanLink72[23] , \ScanLink31[16] , \ScanLink51[12] , 
        \wRegOut_6_4[28] , \wRegInTop_7_59[6] , \wRegInTop_7_59[18] , 
        \ScanLink34[5] , \ScanLink44[26] , \wRegInTop_6_22[18] , 
        \wRegOut_5_26[5] , \wRegInTop_6_57[28] , \ScanLink219[23] , 
        \wRegInBot_4_6[4] , \wRegInTop_4_7[2] , \ScanLink67[17] , 
        \wRegInTop_6_57[31] , \wRegOut_7_84[7] , \wRegOut_7_84[13] , 
        \wRegOut_4_12[27] , \wRegInTop_5_29[2] , \wRegInTop_7_104[13] , 
        \wRegInTop_6_8[26] , \ScanLink117[8] , \wRegInTop_7_44[9] , 
        \wRegInTop_7_127[22] , \wRegInBot_6_35[5] , \wRegOut_7_91[27] , 
        \wRegInTop_7_111[27] , \wRegOut_7_29[13] , \wRegOut_7_56[1] , 
        \wRegOut_7_99[8] , \ScanLink0[29] , \wRegOut_6_27[23] , 
        \wRegOut_6_52[13] , \wRegInTop_7_88[3] , \wRegInTop_1_0[4] , 
        \wRegInBot_1_1[2] , \wRegOut_3_2[9] , \wRegInTop_4_4[1] , 
        \wRegInTop_5_0[21] , \wRegOut_6_11[26] , \wRegInBot_6_36[6] , 
        \wRegOut_7_55[2] , \ScanLink89[22] , \wRegOut_6_32[17] , 
        \wRegOut_6_47[27] , \ScanLink109[4] , \ScanLink127[21] , 
        \ScanLink152[11] , \wRegOut_7_49[17] , \ScanLink171[20] , 
        \ScanLink104[10] , \wRegInTop_7_7[25] , \ScanLink164[14] , 
        \wRegInTop_7_81[28] , \wRegOut_7_87[4] , \wRegInBot_3_2[12] , 
        \wRegInTop_3_7[18] , \wRegInBot_4_5[7] , \ScanLink37[6] , 
        \ScanLink111[24] , \ScanLink147[25] , \wRegInTop_7_81[31] , 
        \wRegOut_5_25[6] , \ScanLink132[15] , \wRegOut_4_12[14] , 
        \wRegInTop_6_8[15] , \wRegInBot_6_51[1] , \wRegOut_7_91[14] , 
        \wRegInTop_7_111[14] , \wRegOut_7_84[20] , \wRegOut_6_13[3] , 
        \wRegInTop_7_104[20] , \ScanLink213[9] , \ScanLink12[14] , 
        \ScanLink31[25] , \ScanLink44[15] , \ScanLink82[7] , \wRegOut_7_32[5] , 
        \wRegInBot_6_37[18] , \wRegInTop_7_127[11] , \wRegInTop_7_3[3] , 
        \wRegInBot_6_14[30] , \ScanLink219[10] , \ScanLink67[24] , 
        \wRegInBot_6_42[28] , \wRegInBot_6_14[29] , \wRegInBot_6_61[19] , 
        \ScanLink24[11] , \ScanLink50[1] , \ScanLink51[21] , \ScanLink72[10] , 
        \wRegInBot_6_42[31] , \wRegInTop_7_121[0] , \wRegOut_7_124[29] , 
        \wRegEnTop_7_73[0] , \wRegOut_7_107[18] , \wRegOut_7_124[30] , 
        \ScanLink111[17] , \ScanLink127[12] , \wRegInTop_7_0[0] , 
        \wRegInTop_7_7[16] , \ScanLink164[27] , \ScanLink132[26] , 
        \ScanLink147[16] , \wRegOut_7_108[3] , \wRegInTop_7_122[3] , 
        \wRegInBot_1_1[27] , \wRegOut_2_0[24] , \wRegInBot_4_13[19] , 
        \wRegInTop_5_0[12] , \wRegInBot_5_19[18] , \ScanLink53[2] , 
        \ScanLink152[22] , \ScanLink104[23] , \wRegOut_6_11[15] , 
        \ScanLink89[11] , \ScanLink171[13] , \wRegOut_6_32[24] , 
        \wRegOut_6_47[14] , \wRegOut_7_49[24] , \wRegInBot_5_5[18] , 
        \ScanLink81[4] , \wRegOut_6_27[10] , \wRegOut_7_29[20] , 
        \wRegOut_6_52[20] , \wRegInBot_5_27[6] , \wRegOut_6_10[0] , 
        \wRegInBot_6_52[2] , \wRegOut_6_29[9] , \ScanLink98[14] , 
        \wRegInTop_7_3[27] , \wRegOut_7_31[6] , \ScanLink160[16] , 
        \ScanLink115[26] , \ScanLink229[3] , \wRegInTop_7_106[5] , 
        \ScanLink77[4] , \ScanLink143[27] , \ScanLink123[23] , 
        \ScanLink136[17] , \ScanLink149[6] , \ScanLink156[13] , 
        \ScanLink175[22] , \wEnable_1[0] , \wRegInBot_5_1[30] , 
        \wRegInTop_5_4[23] , \wRegOut_6_15[24] , \ScanLink100[12] , 
        \wRegOut_6_60[14] , \wRegOut_6_34[6] , \wRegOut_7_15[0] , 
        \wRegEnTop_6_8[0] , \wRegOut_6_23[21] , \wRegOut_6_36[15] , 
        \wRegOut_6_43[25] , \wRegOut_7_38[25] , \wRegOut_6_56[11] , 
        \ScanLink154[9] , \wRegOut_7_58[21] , \wRegInTop_3_3[30] , 
        \wRegInTop_3_3[29] , \wRegInBot_5_1[29] , \wRegEnTop_7_85[0] , 
        \wRegInTop_7_118[9] , \ScanLink69[8] , \wRegOut_7_8[5] , 
        \wRegOut_7_16[3] , \wRegOut_7_95[25] , \wRegInTop_7_115[25] , 
        \wRegInBot_3_6[23] , \wRegOut_6_37[5] , \wRegOut_7_80[11] , 
        \ScanLink16[25] , \ScanLink35[14] , \wRegOut_5_18[15] , 
        \wRegInTop_7_100[11] , \wRegInBot_6_46[19] , \ScanLink198[3] , 
        \wRegInTop_7_123[20] , \ScanLink40[24] , \wRegInBot_5_24[5] , 
        \wRegInTop_7_105[6] , \ScanLink74[7] , \wRegInBot_6_33[29] , 
        \ScanLink20[20] , \ScanLink63[15] , \wRegInBot_6_10[18] , 
        \ScanLink76[21] , \wRegInBot_6_33[30] , \wRegOut_7_103[30] , 
        \wRegOut_7_120[18] , \wRegOut_7_103[29] , \wRegOut_2_0[17] , 
        \ScanLink55[10] , \wRegInTop_6_38[2] , \wRegInTop_7_19[4] , 
        \ScanLink208[15] , \wRegOut_6_23[12] , \wRegOut_7_58[12] , 
        \wRegOut_6_56[22] , \ScanLink4[18] , \wRegInBot_6_12[0] , 
        \wRegOut_6_50[2] , \wRegOut_7_71[4] , \ScanLink250[8] , 
        \wRegInTop_5_4[10] , \wRegOut_6_15[17] , \wRegOut_6_36[26] , 
        \wRegOut_6_60[27] , \wRegOut_6_43[16] , \ScanLink123[10] , 
        \wRegOut_7_38[16] , \ScanLink156[20] , \wRegInBot_1_1[14] , 
        \ScanLink10[3] , \ScanLink13[0] , \wRegInTop_5_13[8] , 
        \ScanLink98[27] , \ScanLink100[21] , \ScanLink115[15] , 
        \ScanLink175[11] , \wRegInTop_7_85[19] , \wRegInTop_7_3[14] , 
        \ScanLink55[23] , \ScanLink76[12] , \ScanLink136[24] , 
        \ScanLink160[25] , \ScanLink143[14] , \ScanLink208[26] , 
        \wRegInTop_2_2[10] , \wRegOut_3_4[18] , \wRegInBot_3_6[10] , 
        \ScanLink16[16] , \ScanLink20[13] , \wRegOut_6_0[19] , 
        \ScanLink35[27] , \ScanLink40[17] , \wRegInTop_7_28[19] , 
        \wRegInTop_6_53[19] , \ScanLink63[26] , \wRegInTop_6_26[29] , 
        \wRegOut_5_18[26] , \wRegInBot_6_11[3] , \wRegInTop_6_26[30] , 
        \wRegOut_6_53[1] , \wRegOut_7_80[22] , \wRegInTop_7_100[22] , 
        \wRegInBot_4_5[15] , \wRegOut_5_3[12] , \wRegInBot_5_16[16] , 
        \wRegInTop_5_20[14] , \wRegInBot_5_21[8] , \wRegInTop_6_41[9] , 
        \wRegOut_7_72[7] , \wRegInTop_7_123[13] , \wRegOut_7_95[16] , 
        \wRegInTop_7_115[16] , \wRegOut_7_4[16] , \ScanLink180[1] , 
        \wRegOut_6_32[8] , \wRegInTop_5_16[11] , \wRegInTop_7_8[18] , 
        \ScanLink232[2] , \wRegInBot_5_20[13] , \wRegInTop_6_20[0] , 
        \ScanLink148[18] , \ScanLink152[7] , \wRegInTop_7_15[10] , 
        \wRegInBot_4_0[10] , \wRegInBot_4_5[26] , \wRegOut_4_9[9] , 
        \wRegOut_5_3[21] , \wRegInTop_5_16[22] , \wRegInBot_6_2[11] , 
        \wRegInTop_6_8[7] , \wRegInBot_6_9[1] , \wRegInTop_6_38[11] , 
        \wRegInTop_7_36[21] , \wRegInTop_7_60[20] , \ScanLink231[1] , 
        \wRegInBot_6_58[12] , \wRegInTop_7_43[11] , \wRegOut_7_108[16] , 
        \wRegInTop_6_23[3] , \wRegInBot_6_38[16] , \wRegInTop_6_58[15] , 
        \wRegInTop_7_23[15] , \ScanLink190[31] , \wRegInTop_7_56[25] , 
        \ScanLink151[4] , \ScanLink190[28] , \wRegInTop_7_75[14] , 
        \wRegEnTop_7_114[0] , \ScanLink72[9] , \wRegInTop_7_103[8] , 
        \ScanLink93[18] , \ScanLink183[2] , \wRegInTop_5_20[27] , 
        \wRegInBot_5_20[20] , \wRegInTop_6_44[4] , \ScanLink136[3] , 
        \wRegInTop_7_65[2] , \wRegInBot_5_16[25] , \wRegOut_5_13[19] , 
        \wRegInTop_5_15[6] , \wRegOut_6_48[30] , \wRegOut_6_48[29] , 
        \wRegOut_7_10[18] , \wRegOut_7_33[30] , \wRegOut_7_65[28] , 
        \wRegOut_7_4[25] , \wRegOut_7_33[29] , \wRegOut_7_46[19] , 
        \wRegOut_7_65[31] , \wRegInTop_6_7[31] , \wRegInTop_6_7[28] , 
        \wRegEnBot_6_44[0] , \wRegOut_6_48[0] , \wRegOut_7_69[6] , 
        \wRegInTop_5_16[5] , \wRegOut_5_30[31] , \wRegOut_5_19[2] , 
        \wRegOut_5_30[28] , \wRegInBot_6_2[22] , \wRegInBot_6_38[25] , 
        \wRegInTop_7_23[26] , \wRegInTop_7_56[16] , \ScanLink68[19] , 
        \wRegInTop_6_58[26] , \wRegInTop_7_75[27] , \wRegInTop_7_60[13] , 
        \wRegOut_7_74[9] , \ScanLink255[5] , \ScanLink255[18] , 
        \ScanLink220[28] , \wRegOut_4_9[14] , \wRegInTop_5_22[4] , 
        \wRegInTop_6_38[22] , \wRegInTop_7_15[23] , \wRegInTop_6_47[7] , 
        \wRegInBot_6_58[21] , \wRegInTop_7_43[22] , \wRegOut_7_108[25] , 
        \ScanLink135[0] , \ScanLink203[19] , \ScanLink220[31] , 
        \wRegInTop_7_36[12] , \wRegInTop_7_66[1] , \wRegInTop_7_80[6] , 
        \wRegInBot_6_7[14] , \wRegInTop_6_28[20] , \wRegInBot_6_48[23] , 
        \wRegInTop_7_26[10] , \wRegInTop_7_52[0] , \wRegInTop_7_53[20] , 
        \wRegOut_7_118[27] , \ScanLink101[1] , \wRegInTop_7_10[15] , 
        \ScanLink180[19] , \wRegInTop_7_70[11] , \wRegInTop_5_13[14] , 
        \wRegInBot_6_28[27] , \wRegInTop_6_48[24] , \wRegOut_7_40[8] , 
        \wRegInTop_7_65[25] , \wRegInTop_7_33[24] , \wRegInTop_7_46[14] , 
        \ScanLink7[4] , \wRegInBot_4_0[23] , \wRegOut_4_12[9] , 
        \wRegOut_5_6[17] , \wRegInBot_5_13[13] , \wRegEnBot_5_22[0] , 
        \wRegInTop_5_25[11] , \wRegInBot_5_25[16] , \wRegInTop_5_30[25] , 
        \wRegInBot_5_30[22] , \ScanLink102[2] , \wRegInTop_7_51[3] , 
        \ScanLink158[29] , \ScanLink158[30] , \wRegInTop_5_21[7] , 
        \wRegInTop_7_83[5] , \wRegOut_7_1[13] , \wRegInTop_7_65[16] , 
        \wRegInTop_4_5[30] , \wRegInTop_4_5[29] , \ScanLink78[31] , 
        \ScanLink78[28] , \wRegInTop_7_10[26] , \wRegInTop_6_17[2] , 
        \wRegInTop_6_48[17] , \wRegInTop_7_8[5] , \ScanLink165[5] , 
        \wRegInTop_7_46[27] , \wRegInBot_6_28[14] , \wRegInBot_6_48[10] , 
        \wRegInTop_7_33[17] , \wRegInTop_7_36[4] , \wRegInTop_7_53[13] , 
        \wRegOut_7_100[6] , \wRegInTop_6_28[13] , \ScanLink245[30] , 
        \wRegOut_7_118[14] , \wRegEnTop_6_59[0] , \wRegInTop_7_26[23] , 
        \wRegInTop_7_70[22] , \ScanLink213[28] , \wRegOut_4_9[27] , 
        \wRegInBot_6_47[8] , \ScanLink205[0] , \ScanLink245[29] , 
        \ScanLink213[31] , \ScanLink230[19] , \ScanLink46[8] , 
        \wRegInBot_6_7[27] , \wRegOut_5_20[19] , \ScanLink89[1] , 
        \wRegOut_6_18[5] , \wRegOut_6_58[18] , \wRegOut_7_1[20] , 
        \wRegOut_7_23[18] , \wRegOut_7_39[3] , \wRegInTop_7_28[8] , 
        \wRegOut_7_56[28] , \wRegOut_7_56[31] , \wRegOut_7_75[19] , 
        \ScanLink4[7] , \wRegInBot_6_59[4] , \wRegInTop_2_2[23] , 
        \wRegOut_5_6[24] , \wRegInBot_5_15[9] , \wRegInTop_5_25[22] , 
        \ScanLink83[30] , \wRegInBot_5_30[11] , \wRegInTop_6_14[1] , 
        \ScanLink83[29] , \wRegInTop_7_35[7] , \ScanLink166[6] , 
        \wRegInTop_5_13[27] , \wRegInBot_5_13[20] , \wRegInTop_5_30[16] , 
        \ScanLink206[3] , \wRegOut_7_103[5] , \wRegInBot_5_25[25] , 
        \ScanLink58[4] , \ScanLink0[17] , \ScanEnable[0] , \wRegOut_1_0[4] , 
        \wRegInBot_1_0[20] , \ScanLink2[9] , \wRegInTop_1_1[31] , 
        \ScanLink25[25] , \ScanLink73[24] , \wRegInBot_6_56[31] , 
        \ScanLink30[11] , \ScanLink50[15] , \wRegInBot_6_23[18] , 
        \wRegInBot_6_56[28] , \wRegInTop_7_49[1] , \wRegInTop_7_86[8] , 
        \wRegOut_7_113[18] , \wRegInTop_1_1[28] , \ScanLink13[20] , 
        \ScanLink24[2] , \ScanLink45[21] , \ScanLink218[24] , 
        \wRegInBot_3_3[26] , \ScanLink66[10] , \wRegOut_7_85[14] , 
        \wRegOut_7_94[0] , \wRegInBot_3_3[15] , \wRegInTop_4_9[9] , 
        \wRegOut_4_13[20] , \wRegInTop_7_105[14] , \wRegInTop_6_9[21] , 
        \wRegInTop_7_110[20] , \wRegInTop_7_126[25] , \wRegInBot_6_25[2] , 
        \wRegOut_7_90[20] , \wRegOut_6_26[24] , \wRegOut_6_53[14] , 
        \wRegOut_7_28[14] , \wRegOut_7_46[6] , \wRegInTop_7_98[4] , 
        \wRegInBot_6_26[1] , \ScanLink27[1] , \wRegInTop_5_1[26] , 
        \wRegOut_6_10[21] , \wRegOut_7_45[5] , \wRegInTop_5_27[9] , 
        \ScanLink88[25] , \wRegOut_6_33[10] , \wRegOut_6_46[20] , 
        \ScanLink119[3] , \ScanLink153[16] , \wRegOut_7_48[10] , 
        \ScanLink126[26] , \ScanLink170[27] , \ScanLink105[17] , 
        \ScanLink110[23] , \wRegInTop_7_6[22] , \ScanLink165[13] , 
        \wRegOut_7_97[3] , \ScanLink146[22] , \wRegOut_4_13[13] , 
        \wRegOut_4_14[7] , \wRegInTop_6_9[12] , \ScanLink133[12] , 
        \wRegInTop_7_110[13] , \wRegInBot_6_41[6] , \wRegOut_7_90[13] , 
        \wRegOut_7_85[27] , \wRegInTop_7_105[27] , \ScanLink13[13] , 
        \wRegOut_4_2[18] , \ScanLink30[22] , \ScanLink45[12] , 
        \wRegOut_6_8[7] , \wRegOut_7_22[2] , \wRegOut_7_106[8] , 
        \ScanLink92[0] , \wRegInTop_7_126[16] , \ScanLink218[17] , 
        \ScanLink66[23] , \ScanLink25[16] , \ScanLink40[6] , 
        \wRegInBot_5_10[4] , \ScanLink73[17] , \wRegInTop_6_43[31] , 
        \wRegInTop_6_60[19] , \wRegInTop_7_38[31] , \wRegInTop_6_15[29] , 
        \wRegInTop_6_43[28] , \ScanLink50[26] , \wRegInTop_7_38[28] , 
        \wRegInTop_6_15[30] , \wRegInTop_6_36[18] , \ScanLink43[5] , 
        \wRegInBot_5_13[7] , \wRegInTop_5_18[18] , \ScanLink110[10] , 
        \ScanLink126[15] , \ScanLink133[21] , \wRegInTop_7_6[11] , 
        \ScanLink165[20] , \ScanLink146[11] , \ScanLink153[25] , 
        \wRegInTop_7_95[31] , \wRegOut_7_118[4] , \ScanLink105[24] , 
        \wRegInTop_7_95[28] , \wRegOut_2_1[23] , \wRegInTop_4_12[19] , 
        \wRegInTop_5_1[15] , \wRegOut_6_10[12] , \ScanLink88[16] , 
        \ScanLink170[14] , \wRegOut_6_33[23] , \wRegOut_6_46[13] , 
        \wRegInTop_7_33[9] , \wRegOut_7_48[23] , \wRegEnTop_5_10[0] , 
        \wRegOut_6_26[17] , \ScanLink160[8] , \ScanLink91[3] , 
        \wRegOut_7_28[27] , \wRegInBot_6_42[5] , \wRegOut_6_53[27] , 
        \wRegOut_7_21[1] , \ScanLink99[13] , \wRegInTop_7_2[20] , 
        \ScanLink161[11] , \wRegEnTop_4_15[0] , \wRegInTop_6_0[2] , 
        \wRegInBot_6_1[4] , \ScanLink67[3] , \ScanLink114[21] , 
        \ScanLink239[4] , \ScanLink142[20] , \wRegOut_7_18[8] , 
        \wRegInTop_7_116[2] , \ScanLink137[10] , \ScanLink157[14] , 
        \ScanLink101[15] , \ScanLink122[24] , \ScanLink159[1] , 
        \ScanLink174[25] , \ScanLink196[8] , \wRegOut_6_61[13] , 
        \wRegInTop_7_91[19] , \wRegInTop_5_5[24] , \wRegOut_6_14[23] , 
        \wRegOut_6_24[1] , \wRegOut_6_22[26] , \wRegOut_6_37[12] , 
        \wRegOut_6_42[22] , \wRegOut_7_39[22] , \wRegOut_6_57[16] , 
        \wRegOut_7_59[26] , \wRegInTop_6_36[9] , \wRegInBot_3_7[24] , 
        \wRegOut_4_6[29] , \wRegOut_6_27[2] , \wRegOut_7_94[22] , 
        \wRegInTop_7_114[22] , \ScanLink227[8] , \wRegOut_7_81[16] , 
        \ScanLink17[22] , \wRegOut_4_6[30] , \wRegOut_5_19[12] , 
        \wRegInTop_7_101[16] , \wRegInBot_6_8[30] , \wRegInTop_7_122[27] , 
        \wRegInBot_4_15[4] , \ScanLink34[13] , \wRegInBot_6_8[29] , 
        \ScanLink188[4] , \wRegInTop_7_115[1] , \ScanLink41[23] , 
        \ScanLink64[0] , \ScanLink21[27] , \ScanLink62[12] , 
        \wRegInBot_6_2[7] , \wRegInTop_6_11[18] , \wRegInTop_6_32[30] , 
        \ScanLink77[26] , \wRegInTop_7_49[30] , \wRegInTop_6_32[29] , 
        \wRegInTop_7_49[29] , \wRegInBot_1_0[13] , \wRegOut_2_1[10] , 
        \ScanLink54[17] , \wRegInTop_6_3[1] , \wRegInTop_6_28[5] , 
        \wRegInTop_6_47[19] , \ScanLink209[12] , \wRegOut_6_22[15] , 
        \wRegOut_7_59[15] , \wRegOut_6_57[25] , \wRegOut_2_1[8] , 
        \wRegInTop_3_4[7] , \wRegInTop_5_4[3] , \wRegInTop_5_5[17] , 
        \wRegOut_6_14[10] , \wRegOut_6_40[5] , \wRegOut_7_61[3] , 
        \wRegOut_6_37[21] , \wRegOut_6_61[20] , \wRegOut_6_42[11] , 
        \wRegInBot_5_5[5] , \wRegOut_5_11[7] , \ScanLink122[17] , 
        \wRegOut_7_39[11] , \ScanLink101[26] , \ScanLink157[27] , 
        \ScanLink174[16] , \wRegOut_5_9[19] , \ScanLink114[12] , 
        \wRegInBot_3_5[1] , \ScanLink99[20] , \wRegInTop_7_2[13] , 
        \wRegInBot_5_6[6] , \ScanLink137[23] , \ScanLink161[22] , 
        \ScanLink142[13] , \wRegInTop_5_7[0] , \ScanLink77[15] , 
        \wRegInBot_6_27[30] , \ScanLink54[24] , \ScanLink209[21] , 
        \wRegInBot_6_27[29] , \wRegInBot_3_6[2] , \wRegInTop_3_7[4] , 
        \ScanLink21[14] , \wRegOut_5_12[4] , \wRegInBot_6_52[19] , 
        \ScanLink34[20] , \ScanLink41[10] , \ScanLink62[21] , 
        \wRegOut_7_117[29] , \ScanLink17[11] , \wRegOut_7_117[30] , 
        \wRegInBot_3_7[17] , \wRegOut_5_19[21] , \wRegOut_6_43[6] , 
        \wRegOut_7_81[25] , \wRegInTop_7_101[25] , \wRegInBot_4_10[9] , 
        \ScanLink123[9] , \wRegOut_7_62[0] , \wRegInTop_7_122[14] , 
        \wRegInTop_7_70[8] , \wRegOut_7_71[31] , \wRegOut_7_94[11] , 
        \wRegInTop_7_114[11] , \wRegEnBot_6_2[0] , \wRegOut_6_29[19] , 
        \wRegOut_7_52[19] , \wRegEnBot_6_33[0] , \wRegOut_7_0[0] , 
        \wRegOut_7_27[29] , \wRegOut_7_5[11] , \wRegOut_7_27[30] , 
        \wRegOut_7_71[28] , \wRegInBot_1_1[19] , \wRegInBot_2_3[18] , 
        \wRegInBot_5_17[11] , \wRegInTop_5_21[13] , \ScanLink190[6] , 
        \wRegOut_7_127[3] , \wRegInTop_3_2[9] , \wRegInTop_4_1[18] , 
        \wRegInBot_4_4[12] , \wRegOut_5_2[15] , \wRegInTop_5_17[16] , 
        \ScanLink87[18] , \ScanLink222[5] , \wRegInBot_5_21[14] , 
        \wRegInTop_6_30[7] , \wRegInTop_7_11[1] , \ScanLink142[0] , 
        \wRegInTop_7_14[17] , \wRegInTop_6_39[16] , \wRegInTop_7_37[26] , 
        \wRegInTop_7_61[27] , \ScanLink221[6] , \wRegOut_7_124[0] , 
        \wRegInBot_6_39[11] , \wRegInBot_6_59[15] , \wRegInTop_7_42[16] , 
        \wRegOut_7_109[11] , \wRegInTop_6_59[12] , \wRegInTop_7_22[12] , 
        \ScanLink217[19] , \ScanLink234[31] , \ScanLink18[6] , 
        \wRegInTop_5_17[25] , \wRegOut_5_24[31] , \wRegOut_5_24[28] , 
        \wRegInBot_6_3[16] , \wRegInTop_6_33[4] , \wRegInTop_7_12[2] , 
        \wRegInTop_7_57[22] , \ScanLink141[3] , \wRegInTop_7_74[13] , 
        \ScanLink234[28] , \ScanLink241[18] , \wRegInBot_6_4[9] , 
        \wRegOut_7_3[3] , \ScanLink193[5] , \wRegInBot_5_21[27] , 
        \ScanLink246[1] , \wRegOut_5_2[26] , \wRegInTop_5_21[20] , 
        \wRegInTop_6_54[3] , \ScanLink126[4] , \ScanLink129[28] , 
        \wRegInTop_7_75[5] , \wRegOut_5_17[9] , \wRegInBot_5_17[22] , 
        \wRegInBot_6_19[6] , \ScanLink129[31] , \wRegOut_7_5[22] , 
        \wRegInTop_3_3[17] , \wRegEnTop_3_4[0] , \wRegOut_4_4[1] , 
        \wRegInBot_5_0[8] , \wRegOut_6_58[7] , \wRegOut_7_79[1] , 
        \wRegInBot_4_4[21] , \wRegOut_4_7[2] , \wRegInBot_6_3[25] , 
        \ScanLink138[8] , \wRegInBot_6_39[22] , \wRegInTop_7_22[21] , 
        \wRegInTop_7_57[11] , \wRegOut_6_45[8] , \wRegInTop_6_59[21] , 
        \wRegInTop_7_74[20] , \ScanLink245[2] , \ScanLink184[28] , 
        \wRegInTop_7_61[14] , \wRegOut_4_7[10] , \wRegInBot_6_9[10] , 
        \wRegInTop_6_39[25] , \wRegInTop_7_14[24] , \wRegInTop_6_57[0] , 
        \wRegInBot_6_59[26] , \wRegInTop_7_42[25] , \wRegOut_7_109[22] , 
        \ScanLink125[7] , \ScanLink184[31] , \wRegInTop_7_37[15] , 
        \wRegInTop_7_76[6] , \ScanLink253[6] , \wRegInBot_6_26[23] , 
        \wRegInTop_6_41[4] , \ScanLink133[3] , \wRegInTop_6_46[20] , 
        \wRegInTop_7_60[2] , \wRegInTop_6_33[10] , \wRegInBot_6_53[13] , 
        \wRegInTop_7_48[10] , \wRegOut_7_103[17] , \wRegOut_2_0[30] , 
        \wRegOut_2_0[29] , \ScanLink4[26] , \ScanLink4[15] , 
        \wRegInTop_4_13[20] , \wRegInBot_4_13[27] , \wRegOut_5_8[13] , 
        \wRegInTop_5_10[6] , \wRegOut_6_0[14] , \wRegInTop_6_10[21] , 
        \wRegInBot_6_10[26] , \wRegOut_7_120[26] , \wRegInTop_6_26[24] , 
        \wRegInBot_6_33[17] , \wRegInTop_7_28[14] , \wRegInBot_6_46[27] , 
        \wRegInTop_6_53[14] , \wRegOut_7_116[23] , \wRegInTop_7_90[20] , 
        \wRegEnBot_6_41[0] , \ScanLink136[29] , \ScanLink143[19] , 
        \ScanLink160[31] , \wRegInTop_7_85[14] , \ScanLink136[30] , 
        \wRegInBot_5_1[17] , \wRegInBot_5_8[0] , \wRegInTop_5_13[5] , 
        \ScanLink115[18] , \wRegInTop_7_3[19] , \ScanLink160[28] , 
        \wRegInTop_5_9[6] , \wRegOut_7_71[9] , \ScanLink250[5] , 
        \wRegInTop_3_3[24] , \ScanLink16[31] , \ScanLink16[28] , 
        \wRegInTop_6_42[7] , \ScanLink130[0] , \wRegInTop_7_63[1] , 
        \ScanLink35[19] , \ScanLink40[30] , \ScanLink63[18] , 
        \wRegInBot_6_10[15] , \wRegInBot_6_46[14] , \wRegOut_7_116[10] , 
        \ScanLink40[29] , \wRegInBot_5_24[8] , \wRegInTop_6_26[17] , 
        \wRegInBot_6_33[24] , \wRegInTop_7_28[27] , \wRegOut_6_0[27] , 
        \wRegInTop_6_33[23] , \wRegInTop_6_53[27] , \wRegInBot_6_53[20] , 
        \wRegInTop_6_10[12] , \wRegInBot_6_26[10] , \wRegInTop_6_46[13] , 
        \wRegInTop_7_48[23] , \wRegOut_7_103[24] , \wRegInTop_7_19[9] , 
        \ScanLink185[1] , \ScanLink208[18] , \wRegOut_6_37[8] , 
        \wRegOut_7_95[28] , \wRegInTop_7_115[28] , \wRegOut_7_120[15] , 
        \wRegOut_7_95[31] , \ScanLink237[2] , \wRegInTop_7_115[31] , 
        \wRegInTop_7_118[4] , \wRegOut_4_7[23] , \ScanLink69[5] , 
        \wRegOut_7_8[8] , \wRegInBot_6_9[23] , \wRegInTop_6_25[0] , 
        \ScanLink157[7] , \wRegOut_5_18[18] , \wRegOut_6_15[30] , 
        \wRegOut_6_36[18] , \wRegOut_6_43[28] , \wRegOut_7_38[28] , 
        \wRegOut_6_15[29] , \wRegOut_6_43[31] , \wRegOut_6_60[19] , 
        \wRegOut_7_38[31] , \ScanLink234[1] , \wRegEnTop_7_111[0] , 
        \wRegInBot_5_1[24] , \ScanLink154[4] , \wRegOut_3_4[26] , 
        \wRegInTop_4_0[21] , \wRegInTop_4_13[13] , \ScanLink77[9] , 
        \wRegInTop_6_26[3] , \wRegInTop_7_106[8] , \wRegOut_6_29[4] , 
        \ScanLink98[19] , \wRegInTop_7_85[27] , \wRegInBot_4_13[14] , 
        \wRegOut_5_8[20] , \ScanLink68[14] , \wRegInBot_6_17[0] , 
        \ScanLink186[2] , \wRegInTop_7_90[13] , \wRegInBot_6_38[31] , 
        \ScanLink240[21] , \wRegOut_6_55[2] , \ScanLink190[16] , 
        \wRegOut_7_74[4] , \ScanLink255[8] , \ScanLink235[11] , 
        \wRegInBot_6_38[28] , \ScanLink185[22] , \ScanLink203[14] , 
        \ScanLink216[20] , \wRegOut_7_108[28] , \wRegOut_7_108[31] , 
        \ScanLink255[15] , \ScanLink220[25] , \ScanLink15[3] , \ScanLink16[0] , 
        \wRegInTop_6_7[25] , \ScanLink248[7] , \wRegOut_5_13[14] , 
        \wRegOut_5_25[11] , \wRegOut_5_30[25] , \ScanLink128[2] , 
        \wRegInTop_5_16[8] , \wRegOut_6_48[24] , \wRegOut_7_33[24] , 
        \wRegOut_7_46[14] , \wRegOut_7_4[31] , \wRegOut_7_10[15] , 
        \wRegOut_7_65[25] , \wRegOut_7_26[10] , \wRegOut_7_70[11] , 
        \wRegInBot_2_0[3] , \wRegInTop_2_2[6] , \wRegInBot_2_2[21] , 
        \wRegInBot_6_14[3] , \wRegOut_6_28[20] , \wRegInTop_6_59[6] , 
        \wRegOut_7_4[28] , \wRegOut_7_53[20] , \wRegInTop_7_78[0] , 
        \ScanLink93[15] , \ScanLink148[26] , \wRegInTop_7_8[26] , 
        \wRegOut_6_56[1] , \wRegOut_7_77[7] , \wRegInBot_2_2[12] , 
        \wRegOut_3_4[15] , \wRegInBot_4_5[18] , \wRegOut_4_9[4] , 
        \ScanLink86[21] , \wRegOut_5_13[27] , \wRegInBot_5_16[31] , 
        \wRegInBot_5_16[28] , \ScanLink128[22] , \wRegInBot_5_22[6] , 
        \wRegOut_5_30[16] , \wRegInTop_6_44[9] , \wRegInTop_7_103[5] , 
        \ScanLink72[4] , \wRegOut_5_25[22] , \wRegInTop_6_7[16] , 
        \ScanLink185[11] , \ScanLink203[27] , \wEnable_4[0] , 
        \ScanLink220[16] , \wRegInTop_4_0[12] , \ScanLink68[27] , 
        \wRegOut_6_31[6] , \wRegOut_7_10[0] , \ScanLink255[26] , 
        \wRegInTop_6_58[18] , \wRegInTop_7_23[18] , \wRegInTop_7_56[31] , 
        \ScanLink190[25] , \ScanLink235[22] , \wRegInTop_7_75[19] , 
        \ScanLink240[12] , \wRegInTop_7_56[28] , \ScanLink216[13] , 
        \ScanLink86[12] , \ScanLink151[9] , \wRegOut_7_13[3] , 
        \wRegInTop_2_3[30] , \wRegInTop_2_3[29] , \wRegInTop_5_20[19] , 
        \wRegOut_6_32[5] , \ScanLink128[11] , \wRegEnTop_7_80[0] , 
        \wRegInBot_5_21[5] , \ScanLink93[26] , \ScanLink148[15] , 
        \wRegInTop_7_8[15] , \wRegOut_7_53[13] , \wRegOut_7_70[22] , 
        \wRegInTop_7_100[6] , \wRegInTop_5_24[31] , \ScanLink71[7] , 
        \wRegOut_6_28[13] , \wRegOut_6_48[17] , \wRegOut_7_26[23] , 
        \wRegOut_7_46[27] , \wRegOut_7_10[26] , \wRegOut_7_33[17] , 
        \wRegOut_7_65[16] , \wRegInTop_5_24[28] , \ScanLink82[23] , 
        \ScanLink159[10] , \ScanLink87[7] , \ScanLink9[2] , \ScanLink97[17] , 
        \ScanLink139[14] , \wRegInBot_6_54[1] , \wRegOut_6_16[3] , 
        \wRegOut_7_37[5] , \ScanLink216[9] , \wRegInBot_2_3[0] , 
        \wRegOut_3_0[24] , \wRegInBot_4_1[30] , \wRegOut_5_17[16] , 
        \ScanLink55[1] , \wRegInTop_6_19[4] , \wRegOut_6_59[12] , 
        \wRegOut_7_22[12] , \wRegOut_7_74[13] , \wRegInTop_7_6[3] , 
        \wRegOut_6_39[16] , \wRegOut_7_37[26] , \wRegInTop_7_38[2] , 
        \wRegOut_7_57[22] , \wRegInTop_7_124[0] , \wRegOut_7_42[16] , 
        \wRegEnTop_7_76[0] , \wRegInTop_7_5[0] , \wRegOut_7_14[17] , 
        \wRegOut_7_61[27] , \ScanLink168[0] , \wRegOut_5_21[13] , 
        \ScanLink56[2] , \wRegInTop_6_3[27] , \wRegOut_7_29[9] , 
        \ScanLink208[5] , \wRegInTop_7_127[3] , \ScanLink207[16] , 
        \ScanLink79[22] , \wRegEnBot_6_19[0] , \ScanLink251[17] , 
        \ScanLink181[20] , \ScanLink224[27] , \wRegInBot_4_1[29] , 
        \ScanLink19[26] , \wRegInBot_6_57[2] , \wRegInTop_7_71[28] , 
        \wRegInTop_4_4[23] , \wRegOut_6_15[0] , \wRegInTop_7_27[30] , 
        \ScanLink244[23] , \wRegOut_7_34[6] , \ScanLink231[13] , 
        \ScanLink194[14] , \ScanLink84[4] , \wRegInTop_6_29[19] , 
        \wRegInTop_7_52[19] , \wRegInTop_7_71[31] , \wRegInTop_7_27[29] , 
        \ScanLink212[22] , \wRegOut_6_39[25] , \wRegOut_7_37[15] , 
        \wRegOut_7_42[25] , \wRegOut_7_61[14] , \wRegOut_3_0[17] , 
        \wRegInTop_4_2[2] , \wRegOut_7_14[24] , \wRegOut_7_74[20] , 
        \wRegInBot_4_3[4] , \wRegOut_7_81[7] , \ScanLink19[15] , 
        \ScanLink31[5] , \wRegOut_7_57[11] , \wRegInBot_5_12[19] , 
        \wRegOut_5_23[5] , \wRegOut_6_59[21] , \wRegOut_7_0[19] , 
        \wRegOut_7_22[21] , \ScanLink97[24] , \ScanLink112[8] , 
        \ScanLink139[27] , \wRegInTop_7_41[9] , \wRegInBot_5_31[31] , 
        \wRegInBot_6_30[5] , \wRegInBot_5_31[28] , \ScanLink82[10] , 
        \wRegOut_7_53[1] , \wRegInBot_6_49[30] , \ScanLink159[23] , 
        \ScanLink194[27] , \ScanLink231[20] , \wRegInTop_4_4[10] , 
        \wRegInBot_6_49[29] , \ScanLink212[11] , \ScanLink244[10] , 
        \ScanLink79[11] , \ScanLink181[13] , \ScanLink207[25] , 
        \ScanLink224[14] , \wRegInBot_6_33[6] , \wRegOut_7_50[2] , 
        \ScanLink251[24] , \wRegInTop_2_1[5] , \wRegInTop_4_13[8] , 
        \wRegInTop_6_3[14] , \wRegOut_3_7[9] , \wRegInTop_4_1[1] , 
        \ScanLink32[6] , \wRegOut_5_20[6] , \wRegOut_5_21[20] , 
        \wRegOut_5_17[25] , \wRegOut_7_82[4] , \wRegInBot_4_0[7] , 
        \wRegInBot_5_5[15] , \wRegOut_6_11[18] , \wRegOut_6_32[29] , 
        \wRegOut_6_47[19] , \wRegOut_7_49[29] , \wRegInTop_7_23[3] , 
        \ScanLink170[2] , \wRegOut_6_32[30] , \wRegOut_7_49[30] , 
        \ScanLink210[7] , \wRegInTop_1_0[11] , \wRegInTop_1_0[9] , 
        \wRegInTop_5_19[12] , \ScanLink81[9] , \wRegOut_7_115[1] , 
        \wRegInTop_7_81[16] , \wRegInBot_5_19[15] , \wRegOut_6_6[1] , 
        \wRegInTop_7_94[22] , \ScanLink12[19] , \ScanLink67[29] , 
        \wRegInBot_6_14[24] , \ScanLink31[31] , \wRegInBot_6_61[14] , 
        \ScanLink31[28] , \ScanLink44[18] , \ScanLink67[30] , 
        \wRegInBot_6_37[15] , \wRegInBot_6_42[25] , \wRegInTop_6_57[16] , 
        \wRegInTop_7_59[26] , \wRegOut_7_112[21] , \wRegOut_6_4[16] , 
        \wRegOut_6_5[2] , \wRegInTop_6_22[26] , \wRegInBot_6_22[21] , 
        \wRegInTop_6_42[22] , \wRegInTop_6_37[12] , \wRegInTop_7_39[22] , 
        \wRegOut_7_107[15] , \wRegInTop_6_14[23] , \wRegInBot_6_57[11] , 
        \wRegInTop_6_61[13] , \wRegOut_7_124[24] , \ScanLink0[24] , 
        \wRegOut_3_2[4] , \wRegInTop_3_7[15] , \wRegInTop_6_8[18] , 
        \wRegOut_7_91[19] , \wRegInTop_7_111[19] , \wRegOut_4_3[12] , 
        \wRegInTop_7_20[0] , \ScanLink173[1] , \wRegOut_7_32[8] , 
        \ScanLink213[4] , \wRegOut_7_116[2] , \wRegOut_4_12[19] , 
        \wRegOut_5_2[0] , \wRegInTop_5_19[21] , \wRegInBot_5_19[26] , 
        \ScanLink109[9] , \wRegInTop_7_94[11] , \wRegInTop_7_95[1] , 
        \ScanLink111[30] , \wRegInTop_7_7[31] , \ScanLink147[28] , 
        \ScanLink132[18] , \wRegInTop_7_7[28] , \ScanLink147[31] , 
        \ScanLink164[19] , \wRegEnBot_4_0[0] , \ScanLink111[29] , 
        \wRegInTop_7_81[25] , \wRegOut_7_87[9] , \wRegOut_7_48[0] , 
        \wRegOut_4_3[21] , \wRegInBot_5_5[26] , \ScanLink114[6] , 
        \ScanLink117[5] , \wRegInTop_7_44[4] , \wRegInTop_7_47[7] , 
        \wRegInBot_6_35[8] , \wRegInTop_1_0[22] , \wRegInTop_3_7[26] , 
        \wRegOut_7_99[5] , \ScanLink29[7] , \wRegInTop_4_15[6] , 
        \wRegOut_5_1[3] , \wRegOut_6_4[25] , \wRegInTop_6_37[21] , 
        \wRegInBot_6_22[12] , \wRegInTop_6_42[11] , \wRegInBot_6_57[22] , 
        \wRegOut_7_107[26] , \wRegInTop_7_39[11] , \wRegInTop_7_96[2] , 
        \wRegInTop_6_14[10] , \wRegOut_7_124[17] , \wRegInBot_6_14[17] , 
        \wRegInBot_6_28[7] , \wRegInTop_6_61[20] , \wRegInBot_6_61[27] , 
        \wRegInBot_1_1[23] , \wRegInBot_2_2[31] , \wRegInBot_2_2[28] , 
        \wRegOut_3_1[7] , \wRegInBot_4_6[9] , \wRegInTop_4_0[31] , 
        \wRegInBot_4_5[22] , \wRegInBot_4_5[11] , \ScanLink34[8] , 
        \wRegOut_5_26[8] , \wRegInTop_6_22[15] , \wRegInBot_6_42[16] , 
        \wRegInTop_7_59[15] , \wRegOut_7_112[12] , \wRegInBot_6_37[26] , 
        \wRegInBot_6_2[15] , \wRegEnBot_6_20[0] , \wRegInTop_6_57[25] , 
        \ScanLink183[6] , \wRegInTop_6_8[3] , \wRegInBot_6_9[5] , 
        \wRegInTop_7_75[10] , \wRegInTop_6_23[7] , \wRegInBot_6_38[12] , 
        \wRegInTop_6_58[11] , \wRegInTop_7_23[11] , \wRegInTop_7_56[21] , 
        \wRegInTop_6_38[15] , \ScanLink151[0] , \wRegInTop_7_36[25] , 
        \wRegInBot_6_58[16] , \wRegInTop_7_43[15] , \wRegOut_7_108[12] , 
        \ScanLink185[18] , \wRegOut_5_3[16] , \wRegInTop_5_16[15] , 
        \wRegInBot_5_20[17] , \wRegOut_7_10[9] , \wRegInTop_7_15[14] , 
        \ScanLink231[5] , \wRegInTop_7_60[24] , \wRegInTop_6_20[4] , 
        \ScanLink152[3] , \wRegInBot_5_16[12] , \wRegInTop_5_20[10] , 
        \ScanLink128[18] , \ScanLink232[6] , \wRegInTop_6_38[26] , 
        \wRegOut_7_4[12] , \ScanLink180[5] , \wRegInTop_6_47[3] , 
        \wRegInBot_6_58[25] , \wRegInTop_7_43[26] , \wRegOut_7_108[21] , 
        \ScanLink135[4] , \wRegInTop_7_15[27] , \wRegInTop_7_36[16] , 
        \wRegInTop_7_60[17] , \wRegInTop_7_66[5] , \wRegInBot_6_17[9] , 
        \wRegInTop_7_75[23] , \wRegInTop_4_0[28] , \ScanLink216[30] , 
        \ScanLink235[18] , \ScanLink240[28] , \ScanLink255[1] , 
        \ScanLink16[9] , \wRegInTop_5_16[1] , \wRegOut_5_19[6] , 
        \wRegInBot_6_38[21] , \wRegInTop_7_23[22] , \wRegInTop_7_56[12] , 
        \ScanLink240[31] , \wRegInTop_6_58[22] , \wRegInBot_6_2[26] , 
        \ScanLink216[29] , \wRegOut_6_48[4] , \wRegOut_7_69[2] , 
        \wRegOut_5_3[25] , \wRegInTop_5_15[2] , \wRegOut_5_25[18] , 
        \ScanLink86[28] , \wRegOut_6_28[30] , \wRegOut_7_53[30] , 
        \wRegOut_7_70[18] , \wRegOut_6_28[29] , \wRegOut_7_4[21] , 
        \wRegOut_7_26[19] , \wRegOut_7_53[29] , \wRegInTop_7_78[9] , 
        \wRegInBot_5_16[21] , \ScanLink86[31] , \ScanLink20[24] , 
        \wRegInTop_5_16[26] , \wRegInTop_5_20[23] , \wRegInBot_5_20[24] , 
        \wRegInTop_6_44[0] , \ScanLink136[7] , \wRegInTop_7_65[6] , 
        \wRegOut_6_56[8] , \wRegInBot_1_1[10] , \wRegOut_2_0[20] , 
        \wRegInBot_3_6[27] , \ScanLink16[21] , \ScanLink55[14] , 
        \wRegInBot_6_26[19] , \wRegInTop_6_38[6] , \wRegInBot_6_53[29] , 
        \wRegInTop_7_19[0] , \ScanLink185[8] , \ScanLink208[11] , 
        \ScanLink76[25] , \wRegInBot_6_53[30] , \ScanLink35[10] , 
        \ScanLink63[11] , \ScanLink40[20] , \wRegInBot_5_24[1] , 
        \wRegInTop_7_105[2] , \wRegOut_7_116[19] , \ScanLink74[3] , 
        \wRegInTop_6_25[9] , \wRegInTop_7_123[24] , \ScanLink198[7] , 
        \wRegOut_7_80[15] , \wRegOut_5_18[11] , \wRegInTop_7_100[15] , 
        \wRegOut_6_37[1] , \wRegOut_7_16[7] , \wRegOut_7_95[21] , 
        \wRegInTop_7_115[21] , \wRegOut_7_8[1] , \ScanLink10[7] , 
        \wRegInBot_3_6[14] , \wRegInTop_5_4[27] , \wRegOut_6_23[25] , 
        \wRegOut_6_56[15] , \wRegOut_7_58[25] , \wRegOut_6_43[21] , 
        \wRegOut_5_8[30] , \wRegOut_5_8[29] , \wRegOut_6_15[20] , 
        \wRegOut_6_36[11] , \wRegOut_7_38[21] , \wRegOut_6_60[10] , 
        \wRegOut_6_34[2] , \wRegOut_7_15[4] , \ScanLink234[8] , 
        \ScanLink175[26] , \ScanLink100[16] , \ScanLink156[17] , 
        \wRegOut_5_18[22] , \wRegInBot_5_27[2] , \ScanLink123[27] , 
        \ScanLink149[2] , \wRegInTop_7_106[1] , \wRegInBot_6_9[19] , 
        \ScanLink77[0] , \ScanLink143[23] , \ScanLink98[10] , 
        \wRegInTop_7_3[23] , \ScanLink136[13] , \ScanLink115[22] , 
        \ScanLink160[12] , \ScanLink229[7] , \wRegOut_7_95[12] , 
        \wRegInTop_7_115[12] , \wRegInBot_6_11[7] , \wRegInTop_7_123[17] , 
        \wRegOut_6_53[5] , \wRegOut_7_80[26] , \wRegOut_7_72[3] , 
        \wRegInTop_7_100[26] , \ScanLink16[12] , \wRegOut_4_7[19] , 
        \ScanLink63[22] , \ScanLink35[23] , \ScanLink40[13] , \ScanLink55[27] , 
        \wRegInTop_6_46[29] , \ScanLink208[22] , \wRegInTop_6_10[31] , 
        \wRegEnTop_6_12[0] , \wRegInTop_6_33[19] , \wRegOut_2_0[13] , 
        \ScanLink13[4] , \ScanLink20[17] , \wRegInTop_7_48[19] , 
        \wRegInTop_4_13[30] , \wRegInTop_6_10[28] , \ScanLink76[16] , 
        \wRegInTop_6_46[30] , \ScanLink136[20] , \wRegInTop_4_13[29] , 
        \ScanLink115[11] , \ScanLink143[10] , \ScanLink98[23] , 
        \wRegInTop_7_3[10] , \ScanLink100[25] , \ScanLink160[21] , 
        \ScanLink123[14] , \ScanLink175[15] , \wRegInTop_7_90[29] , 
        \ScanLink156[24] , \wRegInTop_7_90[30] , \wRegInTop_5_4[14] , 
        \wRegOut_6_36[22] , \wRegInTop_7_63[8] , \wRegInBot_6_12[4] , 
        \wRegOut_6_15[13] , \wRegOut_6_43[12] , \ScanLink130[9] , 
        \wRegOut_7_38[12] , \wRegOut_6_60[23] , \wRegInTop_4_4[5] , 
        \ScanLink37[2] , \wRegInBot_5_8[9] , \wRegInTop_5_19[31] , 
        \wRegOut_6_23[16] , \wRegOut_6_50[6] , \wRegOut_7_58[16] , 
        \wRegOut_7_71[0] , \wRegOut_6_56[26] , \ScanLink147[21] , 
        \wRegInTop_5_19[28] , \wRegOut_5_25[2] , \ScanLink132[11] , 
        \wRegInTop_7_7[21] , \ScanLink164[10] , \wRegInBot_4_5[3] , 
        \wRegOut_7_87[0] , \wRegInTop_5_0[25] , \wRegOut_5_2[9] , 
        \ScanLink89[26] , \ScanLink111[20] , \wRegOut_7_48[9] , 
        \ScanLink171[24] , \ScanLink104[14] , \ScanLink109[0] , 
        \ScanLink152[15] , \wRegInTop_7_94[18] , \wRegInTop_7_95[8] , 
        \wRegOut_6_47[23] , \ScanLink127[25] , \wRegInTop_6_8[22] , 
        \wRegOut_6_11[22] , \wRegOut_6_32[13] , \wRegInBot_6_36[2] , 
        \wRegOut_7_49[13] , \wRegOut_6_27[27] , \wRegOut_6_52[17] , 
        \wRegOut_7_29[17] , \wRegOut_7_55[6] , \wRegInTop_7_88[7] , 
        \wRegInTop_7_111[23] , \wRegInBot_6_35[1] , \wRegOut_7_91[23] , 
        \wRegOut_7_56[5] , \wRegOut_0_0[2] , \wRegInTop_1_0[18] , 
        \wRegInTop_1_0[0] , \wRegInBot_1_1[6] , \wRegInBot_3_2[25] , 
        \wRegOut_4_3[31] , \wRegOut_4_3[28] , \wRegOut_7_84[17] , 
        \wRegInTop_7_127[26] , \ScanLink12[23] , \wRegOut_4_12[23] , 
        \wRegInTop_7_104[17] , \wRegInTop_5_29[6] , \wRegInBot_4_6[0] , 
        \wRegInTop_4_7[6] , \ScanLink67[13] , \wRegOut_7_84[3] , 
        \ScanLink24[26] , \ScanLink31[12] , \ScanLink34[1] , \ScanLink44[22] , 
        \wRegOut_5_26[1] , \wRegEnTop_7_17[0] , \wRegInTop_6_37[28] , 
        \ScanLink219[27] , \wRegInTop_5_0[16] , \ScanLink51[16] , 
        \wRegInTop_6_42[18] , \wRegInTop_6_61[30] , \wRegInTop_7_59[2] , 
        \wRegInTop_7_39[18] , \ScanLink72[27] , \wRegInTop_6_14[19] , 
        \wRegInTop_6_37[31] , \wRegInTop_6_61[29] , \wRegOut_6_10[4] , 
        \wRegInBot_6_52[6] , \ScanLink81[0] , \wRegOut_6_27[14] , 
        \wRegOut_7_31[2] , \wRegOut_7_115[8] , \wRegOut_7_29[24] , 
        \wRegOut_6_32[20] , \wRegOut_6_52[24] , \wRegOut_7_49[20] , 
        \wRegOut_6_6[8] , \wRegOut_6_11[11] , \wRegOut_6_47[10] , 
        \ScanLink89[15] , \ScanLink104[27] , \ScanLink171[17] , 
        \ScanLink127[16] , \wRegOut_7_108[7] , \wRegInTop_7_122[7] , 
        \ScanLink24[15] , \ScanLink50[5] , \ScanLink51[25] , \ScanLink53[6] , 
        \ScanLink152[26] , \ScanLink111[13] , \wRegInTop_7_0[4] , 
        \ScanLink132[22] , \ScanLink147[12] , \wRegInTop_7_7[12] , 
        \ScanLink164[23] , \wRegInTop_7_121[4] , \wRegInBot_6_22[28] , 
        \wRegInBot_6_57[18] , \ScanLink67[20] , \ScanLink72[14] , 
        \wRegInBot_6_22[31] , \wRegInTop_2_3[20] , \wRegInTop_2_3[13] , 
        \wRegInBot_2_3[9] , \wRegInBot_3_2[16] , \ScanLink12[10] , 
        \wRegOut_7_112[31] , \wRegOut_4_12[10] , \ScanLink31[21] , 
        \ScanLink44[11] , \wRegInTop_7_3[7] , \ScanLink219[14] , 
        \wRegOut_7_112[28] , \wRegOut_6_13[7] , \ScanLink82[3] , 
        \wRegInBot_6_51[5] , \wRegInTop_7_127[15] , \wRegOut_7_84[24] , 
        \wRegInTop_7_104[24] , \wRegOut_7_32[1] , \wRegOut_3_4[3] , 
        \wRegInTop_6_8[11] , \wRegInTop_7_111[10] , \wRegInTop_7_20[9] , 
        \ScanLink173[8] , \wRegOut_7_91[10] , \wRegOut_7_74[29] , 
        \wRegOut_6_59[31] , \wRegOut_7_22[31] , \wRegOut_6_59[28] , 
        \wRegOut_7_22[28] , \wRegOut_7_57[18] , \wRegOut_7_74[30] , 
        \wRegOut_7_0[10] , \wRegInTop_7_93[6] , \wRegInTop_4_10[2] , 
        \wRegOut_5_4[7] , \wRegOut_5_7[14] , \wRegInBot_5_12[10] , 
        \wRegInTop_5_31[4] , \wRegInTop_5_24[12] , \wRegInBot_5_31[21] , 
        \ScanLink82[19] , \wRegOut_7_53[8] , \wRegOut_3_7[0] , 
        \wRegInTop_4_1[8] , \wRegInBot_4_1[13] , \wRegInTop_5_12[17] , 
        \wRegInBot_5_24[15] , \wRegInTop_5_31[26] , \ScanLink112[1] , 
        \wRegInTop_6_60[6] , \wRegInTop_7_41[0] , \wRegInBot_6_29[24] , 
        \wRegInTop_6_49[27] , \wRegInTop_7_32[27] , \wRegInTop_7_47[17] , 
        \wRegInTop_4_4[19] , \wRegEnBot_5_31[0] , \ScanLink79[18] , 
        \wRegInTop_7_11[16] , \wRegInTop_7_64[26] , \wRegInTop_7_71[12] , 
        \ScanLink231[29] , \ScanLink244[19] , \wRegInTop_7_27[13] , 
        \wRegInTop_7_42[3] , \wRegInTop_7_52[23] , \ScanLink212[18] , 
        \ScanLink231[30] , \wRegInBot_6_6[17] , \wRegInTop_6_29[23] , 
        \wRegInBot_6_49[20] , \wRegInTop_6_63[5] , \wRegOut_7_119[24] , 
        \ScanLink111[2] , \wRegOut_4_8[17] , \wRegInTop_4_13[1] , 
        \wRegOut_5_7[4] , \wRegOut_5_21[30] , \wRegInBot_5_18[5] , 
        \wRegOut_5_21[29] , \wRegInTop_5_31[15] , \wRegInTop_7_90[5] , 
        \wRegOut_7_113[6] , \wRegOut_5_7[27] , \wRegInTop_5_12[24] , 
        \ScanLink48[7] , \wRegInBot_5_24[26] , \wRegInBot_6_54[8] , 
        \ScanLink216[0] , \wRegInBot_5_12[23] , \ScanLink55[8] , 
        \wRegInTop_5_24[21] , \ScanLink159[19] , \wRegInBot_5_31[12] , 
        \wRegOut_6_0[6] , \wRegInTop_7_25[4] , \ScanLink176[5] , 
        \wRegInTop_7_124[9] , \wRegInBot_6_49[7] , \wRegOut_7_0[23] , 
        \wRegEnTop_7_3[0] , \ScanLink1[27] , \ScanLink1[14] , \ScanLink1[3] , 
        \wRegInTop_3_6[16] , \wRegInBot_4_1[20] , \wRegOut_4_8[24] , 
        \wRegOut_6_3[5] , \wRegOut_7_29[0] , \wRegInBot_6_6[24] , 
        \ScanLink99[2] , \wRegInTop_7_5[9] , \ScanLink168[9] , 
        \wRegOut_6_15[9] , \wRegInTop_7_71[21] , \ScanLink215[3] , 
        \wRegInTop_6_29[10] , \wRegInBot_6_49[13] , \wRegInTop_7_52[10] , 
        \wRegOut_7_110[5] , \wRegOut_7_119[17] , \wRegInBot_6_29[17] , 
        \wRegInTop_6_49[14] , \wRegInTop_7_27[20] , \wRegInTop_7_47[24] , 
        \ScanLink175[6] , \ScanLink181[30] , \wRegInTop_7_11[25] , 
        \wRegInTop_7_26[7] , \wRegInTop_7_32[14] , \ScanLink181[29] , 
        \wRegInTop_7_64[15] , \wRegOut_4_2[11] , \ScanLink203[7] , 
        \ScanLink92[9] , \wRegOut_7_106[1] , \wRegInTop_6_11[5] , 
        \ScanLink163[2] , \wRegInTop_6_60[10] , \wRegInTop_7_30[3] , 
        \ScanLink2[0] , \wRegInTop_1_1[12] , \wRegOut_6_5[15] , 
        \wRegInTop_6_15[20] , \wRegInBot_6_23[22] , \wRegInTop_6_43[21] , 
        \wRegOut_7_125[27] , \wRegInTop_6_36[11] , \wRegInTop_7_38[21] , 
        \wRegOut_7_106[16] , \wRegInBot_6_15[27] , \wRegInTop_6_23[25] , 
        \wRegInBot_6_36[16] , \wRegInBot_6_56[12] , \wRegInBot_6_43[26] , 
        \wRegInTop_6_56[15] , \wRegInTop_7_58[25] , \wRegOut_7_113[22] , 
        \wRegInBot_5_18[16] , \wRegInBot_6_60[17] , \wRegInBot_5_4[16] , 
        \wRegInTop_5_18[11] , \ScanLink110[19] , \ScanLink133[31] , 
        \wRegInTop_7_80[15] , \wRegInTop_7_95[21] , \wRegInTop_7_6[18] , 
        \ScanLink133[28] , \ScanLink165[29] , \ScanLink146[18] , 
        \ScanLink165[30] , \wRegOut_7_105[2] , \wRegOut_7_21[8] , 
        \ScanLink200[4] , \wRegInTop_1_1[21] , \ScanLink13[30] , 
        \ScanLink30[18] , \wRegInTop_6_12[6] , \ScanLink160[1] , 
        \wRegInTop_7_33[0] , \wRegInTop_7_58[16] , \wRegOut_7_113[11] , 
        \ScanLink13[29] , \ScanLink45[28] , \wRegInTop_6_23[16] , 
        \wRegInBot_6_43[15] , \wRegInBot_6_36[25] , \wRegInTop_6_56[26] , 
        \wRegInBot_6_60[24] , \ScanLink45[31] , \ScanLink66[19] , 
        \wRegInBot_6_38[4] , \wRegInTop_3_6[25] , \wRegInTop_5_24[3] , 
        \wRegInTop_6_15[13] , \wRegInBot_6_15[14] , \wRegOut_7_94[9] , 
        \wRegOut_7_125[14] , \wRegOut_6_5[26] , \wRegInTop_6_36[22] , 
        \wRegInTop_6_60[23] , \wRegInTop_6_9[31] , \wRegInBot_6_23[11] , 
        \wRegInTop_6_43[12] , \wRegInBot_6_56[21] , \wRegOut_7_106[25] , 
        \wRegInTop_7_38[12] , \wRegInTop_7_49[8] , \wRegInTop_7_86[1] , 
        \wRegOut_7_90[30] , \wRegInTop_7_110[30] , \wRegOut_4_2[22] , 
        \wRegOut_4_13[29] , \ScanLink39[4] , \wRegInTop_6_9[28] , 
        \wRegOut_7_89[6] , \wRegOut_7_90[29] , \wRegInTop_7_110[29] , 
        \wRegInBot_4_8[6] , \wRegInTop_4_9[0] , \wRegOut_4_13[30] , 
        \wRegInBot_6_26[8] , \ScanLink107[6] , \wRegInTop_7_54[7] , 
        \wRegOut_6_46[30] , \wRegOut_6_10[28] , \wRegOut_5_28[7] , 
        \wRegOut_6_10[31] , \wRegOut_6_33[19] , \wRegOut_6_46[29] , 
        \wRegEnTop_6_38[0] , \wRegOut_7_48[19] , \ScanLink104[5] , 
        \wRegInTop_7_57[4] , \wRegOut_3_1[27] , \ScanLink18[25] , 
        \wRegInTop_4_5[20] , \ScanLink27[8] , \wRegInBot_5_4[25] , 
        \wRegInTop_5_18[22] , \wRegOut_7_58[3] , \wRegInTop_7_80[26] , 
        \wRegInBot_5_18[25] , \wRegInTop_7_85[2] , \wRegInTop_5_27[0] , 
        \wRegInTop_7_95[12] , \ScanLink94[7] , \wRegInBot_6_48[19] , 
        \ScanLink213[21] , \wRegInBot_6_47[1] , \ScanLink78[21] , 
        \wRegOut_7_24[5] , \ScanLink195[17] , \ScanLink245[20] , 
        \ScanLink230[10] , \ScanLink180[23] , \ScanLink205[9] , 
        \ScanLink225[24] , \ScanLink250[14] , \ScanLink46[1] , 
        \wRegInBot_5_16[3] , \ScanLink206[15] , \wRegOut_5_16[15] , 
        \wRegOut_5_20[10] , \ScanLink89[8] , \wRegEnTop_7_65[0] , 
        \wRegInTop_6_2[24] , \ScanLink218[6] , \ScanLink178[3] , 
        \wRegInBot_0_0[26] , \wRegInBot_0_0[24] , \ScanLink45[2] , 
        \wRegInBot_5_15[0] , \wRegOut_7_15[14] , \wRegOut_7_60[24] , 
        \wRegOut_6_38[15] , \wRegOut_7_36[25] , \wRegOut_7_43[15] , 
        \wRegOut_6_58[11] , \wRegOut_7_23[11] , \wRegOut_7_1[29] , 
        \wRegInBot_0_0[17] , \wRegInTop_2_2[19] , \wRegOut_3_1[14] , 
        \wRegInBot_4_0[19] , \ScanLink22[5] , \wRegOut_4_11[3] , 
        \wRegInBot_5_13[30] , \wRegInBot_5_30[18] , \ScanLink96[14] , 
        \wRegOut_7_1[30] , \wRegInTop_7_28[1] , \wRegOut_7_56[21] , 
        \wRegOut_7_75[10] , \ScanLink97[4] , \wRegInBot_6_44[2] , 
        \wRegOut_7_27[6] , \ScanLink138[17] , \ScanLink158[13] , 
        \wRegInTop_6_14[8] , \wRegInBot_5_13[29] , \ScanLink83[20] , 
        \wRegOut_5_16[26] , \wRegOut_7_92[7] , \wRegOut_5_30[5] , 
        \wRegOut_5_20[23] , \wRegInTop_6_2[17] , \ScanLink78[12] , 
        \ScanLink180[10] , \ScanLink225[17] , \ScanLink18[16] , 
        \wRegInTop_4_5[13] , \wRegInBot_6_23[5] , \wRegOut_6_61[7] , 
        \wRegOut_7_40[1] , \ScanLink250[27] , \wRegInTop_7_26[19] , 
        \ScanLink206[26] , \ScanLink213[12] , \wRegInTop_6_28[29] , 
        \ScanLink101[8] , \wRegInTop_7_52[9] , \wRegInTop_7_53[29] , 
        \ScanLink195[24] , \wRegInTop_7_70[18] , \ScanLink230[23] , 
        \wRegOut_5_9[2] , \wRegInTop_5_25[18] , \wRegInTop_6_28[30] , 
        \wRegInTop_7_53[30] , \ScanLink158[20] , \ScanLink245[13] , 
        \ScanLink83[13] , \wRegInBot_6_20[6] , \wRegOut_7_43[2] , 
        \wRegOut_6_62[4] , \ScanLink96[27] , \ScanLink21[6] , 
        \ScanLink138[24] , \wRegOut_7_56[12] , \wRegOut_4_12[0] , 
        \wRegOut_7_23[22] , \ScanLink1[25] , \ScanLink1[16] , 
        \wRegInBot_1_0[30] , \wRegOut_2_1[19] , \wRegInBot_2_3[22] , 
        \wRegInTop_5_21[30] , \wRegInTop_5_21[29] , \wRegOut_6_38[26] , 
        \wRegOut_6_58[22] , \wRegOut_7_15[27] , \wRegOut_7_60[17] , 
        \wRegOut_7_75[23] , \wRegOut_7_91[4] , \wRegOut_7_36[16] , 
        \wRegOut_7_43[26] , \ScanLink129[21] , \wRegInBot_2_3[11] , 
        \wRegInBot_3_0[5] , \wRegInTop_3_1[3] , \wRegInTop_3_2[0] , 
        \wRegInTop_5_18[7] , \ScanLink87[22] , \ScanLink92[16] , 
        \wRegOut_6_29[23] , \wRegOut_6_46[2] , \wRegInTop_7_9[25] , 
        \wRegInTop_6_49[5] , \ScanLink149[25] , \wRegOut_7_67[4] , 
        \ScanLink246[8] , \wRegOut_7_27[13] , \wRegOut_7_52[23] , 
        \wRegInTop_7_68[3] , \wRegInBot_3_3[6] , \wRegOut_7_71[12] , 
        \wRegOut_4_4[8] , \wRegInTop_5_2[4] , \wRegInBot_5_3[2] , 
        \wRegOut_7_11[16] , \wRegOut_5_17[0] , \wRegOut_6_49[27] , 
        \wRegOut_7_64[26] , \wRegOut_7_32[27] , \wRegOut_7_47[17] , 
        \wRegOut_5_12[17] , \wRegOut_3_5[25] , \wRegInBot_5_0[1] , 
        \wRegOut_5_14[3] , \wRegOut_5_31[26] , \ScanLink138[1] , 
        \wRegOut_5_24[12] , \wRegInTop_6_6[26] , \wRegInTop_5_1[7] , 
        \wRegOut_7_79[8] , \ScanLink184[21] , \ScanLink221[26] , 
        \ScanLink254[16] , \wRegInTop_4_1[22] , \wRegInBot_4_4[31] , 
        \wRegInBot_4_4[28] , \wRegInTop_6_57[9] , \ScanLink202[17] , 
        \wRegInTop_7_57[18] , \wRegInBot_4_10[0] , \ScanLink69[17] , 
        \wRegInTop_6_59[28] , \wRegInTop_7_22[28] , \wRegInTop_7_74[30] , 
        \ScanLink217[23] , \wRegInTop_7_74[29] , \ScanLink241[22] , 
        \wRegInTop_6_6[5] , \wRegInBot_6_7[3] , \wRegOut_6_45[1] , 
        \wRegInTop_7_22[31] , \wRegInTop_6_59[31] , \wRegOut_7_11[25] , 
        \ScanLink191[15] , \wRegOut_7_64[15] , \wRegOut_7_64[7] , 
        \ScanLink234[12] , \wRegOut_7_47[24] , \wRegOut_6_49[14] , 
        \wRegOut_7_32[14] , \wRegInBot_5_17[18] , \ScanLink61[4] , 
        \wRegInBot_5_31[6] , \wRegOut_7_52[10] , \wRegInTop_7_110[5] , 
        \wRegOut_6_29[10] , \ScanLink92[25] , \wRegOut_7_0[9] , 
        \wRegOut_7_5[18] , \wRegOut_7_27[20] , \wRegOut_7_71[21] , 
        \ScanLink129[12] , \wRegInTop_7_9[16] , \wRegInTop_7_11[8] , 
        \ScanLink142[9] , \ScanLink149[16] , \wRegOut_6_22[6] , 
        \ScanLink87[11] , \wRegInBot_6_60[4] , \wRegOut_3_5[16] , 
        \wRegInTop_4_1[11] , \wRegInBot_6_39[18] , \ScanLink217[10] , 
        \ScanLink69[24] , \ScanLink184[12] , \ScanLink191[26] , 
        \ScanLink221[15] , \ScanLink234[21] , \ScanLink241[11] , 
        \wRegInBot_4_13[3] , \wRegOut_5_12[24] , \wRegOut_5_24[21] , 
        \wRegInBot_6_4[0] , \wRegOut_6_21[5] , \wRegInBot_6_63[7] , 
        \ScanLink254[25] , \ScanLink202[24] , \wRegEnTop_7_93[0] , 
        \wRegOut_7_124[9] , \wRegOut_7_109[18] , \wRegInTop_6_5[6] , 
        \wRegInTop_6_6[15] , \wRegOut_5_31[15] , \wRegInTop_7_113[6] , 
        \wRegInBot_5_0[14] , \ScanLink62[7] , \wRegOut_6_14[19] , 
        \wRegEnTop_6_60[0] , \wRegOut_6_37[31] , \wRegOut_6_37[28] , 
        \wRegOut_6_61[29] , \wRegOut_6_42[18] , \wRegInTop_6_52[4] , 
        \ScanLink120[3] , \wRegOut_6_61[30] , \wRegInTop_7_73[2] , 
        \wRegOut_7_39[18] , \wRegOut_2_1[1] , \ScanLink5[16] , 
        \ScanLink240[6] , \wRegOut_2_2[2] , \wRegInBot_3_5[8] , 
        \wRegOut_4_2[6] , \wRegInTop_4_12[23] , \wRegInTop_7_84[17] , 
        \ScanLink99[30] , \ScanLink99[29] , \wRegOut_4_1[5] , \ScanLink17[18] , 
        \wRegInBot_4_12[24] , \wRegOut_5_9[10] , \wRegInTop_7_91[23] , 
        \wRegEnTop_5_1[0] , \ScanLink34[29] , \ScanLink41[19] , 
        \wRegInTop_7_29[17] , \ScanLink62[31] , \wRegInBot_6_32[14] , 
        \wRegInBot_6_47[24] , \wRegInTop_6_52[17] , \ScanLink62[28] , 
        \wRegInBot_6_11[25] , \wRegInTop_6_27[27] , \wRegOut_7_117[20] , 
        \wRegEnBot_6_52[0] , \ScanLink34[30] , \ScanLink5[25] , 
        \wRegInTop_3_2[14] , \wRegInTop_5_7[9] , \wRegInTop_6_11[22] , 
        \ScanLink209[31] , \wRegOut_6_1[17] , \wRegInBot_6_27[20] , 
        \wRegInTop_6_47[23] , \ScanLink209[28] , \wRegOut_7_121[25] , 
        \wRegInTop_6_32[13] , \wRegInBot_6_52[10] , \wRegInTop_7_49[13] , 
        \wRegOut_7_102[14] , \wRegOut_4_6[13] , \wRegOut_5_19[28] , 
        \wRegInTop_6_51[7] , \ScanLink123[0] , \wRegInTop_7_70[1] , 
        \wRegOut_7_94[18] , \wRegInTop_7_114[18] , \wRegInTop_4_12[10] , 
        \wRegInBot_4_12[17] , \wRegOut_5_9[23] , \wRegOut_5_19[31] , 
        \wRegOut_7_62[9] , \ScanLink243[5] , \wRegInBot_6_8[13] , 
        \ScanLink159[8] , \ScanLink196[1] , \wRegEnTop_5_29[0] , 
        \wRegInTop_7_2[29] , \wRegInTop_7_91[10] , \ScanLink142[30] , 
        \ScanLink161[18] , \wRegOut_6_39[7] , \ScanLink114[28] , 
        \wRegOut_7_18[1] , \wRegInTop_7_84[24] , \wRegInTop_6_36[0] , 
        \ScanLink114[31] , \wRegInTop_7_2[30] , \wRegOut_7_6[7] , 
        \ScanLink142[29] , \ScanLink137[19] , \ScanLink144[7] , 
        \wRegInTop_7_17[6] , \wRegInTop_3_2[27] , \wRegOut_4_6[20] , 
        \wRegInBot_5_0[27] , \wRegOut_6_24[8] , \ScanLink224[2] , 
        \wRegOut_7_121[4] , \wRegInBot_5_29[4] , \wRegInBot_6_8[20] , 
        \wRegInTop_6_35[3] , \wRegInTop_7_14[5] , \wRegEnTop_7_102[0] , 
        \ScanLink147[4] , \wRegInTop_7_108[7] , \wRegOut_7_122[7] , 
        \wRegInTop_6_11[11] , \ScanLink79[6] , \ScanLink227[1] , 
        \wRegInBot_1_0[29] , \wRegOut_6_1[24] , \wRegInTop_6_32[20] , 
        \wRegOut_7_121[16] , \wRegInBot_6_52[23] , \ScanLink64[9] , 
        \wRegInTop_6_3[8] , \wRegInTop_6_47[10] , \wRegInTop_7_49[20] , 
        \wRegOut_7_102[27] , \ScanLink195[2] , \wRegInTop_6_27[14] , 
        \wRegInBot_6_27[13] , \wRegInBot_6_47[17] , \wRegOut_7_117[13] , 
        \wRegInBot_6_32[27] , \wRegInTop_7_115[8] , \wRegInTop_6_52[24] , 
        \wRegInTop_7_29[24] , \wRegOut_6_10[19] , \wRegInBot_6_11[16] , 
        \wRegOut_7_5[4] , \wRegOut_6_33[31] , \wRegInTop_6_12[4] , 
        \wRegOut_6_46[18] , \wRegInTop_7_33[2] , \wRegOut_7_48[31] , 
        \ScanLink91[8] , \wRegOut_6_33[28] , \ScanLink160[3] , 
        \wRegOut_7_48[28] , \ScanLink200[6] , \wRegOut_7_105[0] , 
        \ScanLink1[1] , \ScanLink2[2] , \wRegInBot_5_4[14] , 
        \wRegInTop_5_18[13] , \wRegInBot_5_18[14] , \wRegInTop_7_80[17] , 
        \wRegInTop_7_95[23] , \wRegInTop_1_1[10] , \ScanLink13[18] , 
        \ScanLink30[30] , \ScanLink30[29] , \wRegOut_7_113[20] , 
        \ScanLink45[19] , \ScanLink66[31] , \wRegInTop_6_23[27] , 
        \wRegInBot_6_43[24] , \wRegInTop_7_58[27] , \wRegInBot_6_36[14] , 
        \wRegInTop_6_56[17] , \wRegInBot_6_60[15] , \ScanLink66[28] , 
        \wRegEnBot_6_12[0] , \wRegInBot_6_15[25] , \wRegInTop_6_15[22] , 
        \wRegOut_7_125[25] , \wRegInTop_3_6[14] , \wRegOut_6_5[17] , 
        \wRegInTop_6_36[13] , \wRegInTop_6_60[12] , \wRegInBot_6_56[10] , 
        \wRegInTop_6_11[7] , \wRegInBot_6_23[20] , \wRegInTop_6_43[23] , 
        \wRegOut_7_106[14] , \wRegInTop_7_38[23] , \wRegInTop_7_30[1] , 
        \ScanLink163[0] , \wRegOut_4_2[13] , \wRegOut_4_13[18] , 
        \wRegInTop_6_9[19] , \wRegInTop_7_110[18] , \wRegOut_7_90[18] , 
        \wRegOut_7_22[9] , \wRegInBot_5_4[27] , \wRegInTop_5_18[20] , 
        \wRegInBot_5_18[27] , \ScanLink119[8] , \ScanLink203[5] , 
        \wRegInTop_7_85[0] , \wRegOut_7_106[3] , \wRegInTop_5_27[2] , 
        \ScanLink110[28] , \wRegOut_7_58[1] , \wRegInTop_7_80[24] , 
        \wRegInTop_7_95[10] , \wRegOut_7_97[8] , \ScanLink104[7] , 
        \ScanLink110[31] , \ScanLink133[19] , \wRegInTop_7_6[29] , 
        \ScanLink146[30] , \ScanLink165[18] , \wRegInTop_7_6[30] , 
        \ScanLink146[29] , \wRegInTop_7_57[6] , \wRegInTop_1_1[23] , 
        \wRegInTop_3_6[27] , \wRegOut_4_2[20] , \wRegInBot_4_8[4] , 
        \wRegInTop_4_9[2] , \wRegOut_5_28[5] , \ScanLink107[4] , 
        \wRegInTop_7_54[5] , \ScanLink24[9] , \ScanLink39[6] , 
        \wRegInTop_5_24[1] , \wRegInBot_6_25[9] , \wRegOut_7_89[4] , 
        \wRegInTop_6_60[21] , \wRegOut_6_5[24] , \wRegInTop_6_15[11] , 
        \wRegInBot_6_23[13] , \wRegInTop_6_43[10] , \wRegOut_7_125[16] , 
        \wRegInTop_6_36[20] , \wRegInTop_7_38[10] , \wRegInTop_7_86[3] , 
        \wRegInBot_6_56[23] , \wRegOut_7_106[27] , \wRegInBot_6_36[27] , 
        \wRegInTop_6_56[24] , \wRegInBot_6_15[16] , \wRegInTop_6_23[14] , 
        \wRegInBot_6_43[17] , \wRegInTop_7_58[14] , \wRegOut_7_113[13] , 
        \wRegInTop_2_2[31] , \wRegInTop_5_25[30] , \wRegInTop_5_25[29] , 
        \wRegInBot_6_38[6] , \wRegInBot_6_60[26] , \ScanLink158[11] , 
        \ScanLink83[22] , \wRegInTop_2_2[28] , \ScanLink96[16] , 
        \wRegOut_7_27[4] , \ScanLink206[8] , \wRegInBot_6_44[0] , 
        \ScanLink97[6] , \ScanLink138[15] , \wRegOut_7_23[13] , 
        \wRegInTop_7_28[3] , \wRegOut_7_56[23] , \wRegInBot_0_0[15] , 
        \wRegOut_3_1[25] , \ScanLink45[0] , \wRegOut_6_38[17] , 
        \wRegOut_6_58[13] , \wRegOut_7_15[16] , \wRegOut_7_60[26] , 
        \wRegOut_7_75[12] , \ScanLink46[3] , \wRegInBot_5_15[2] , 
        \wRegOut_7_36[27] , \wRegOut_7_43[17] , \wRegOut_5_16[17] , 
        \ScanLink178[1] , \wRegInBot_5_16[1] , \wRegOut_5_20[12] , 
        \wRegInTop_6_2[26] , \wRegOut_7_39[8] , \ScanLink218[4] , 
        \ScanLink180[21] , \ScanLink225[26] , \wRegInBot_4_0[31] , 
        \wRegInBot_4_0[28] , \ScanLink78[23] , \wRegInTop_6_17[9] , 
        \ScanLink206[17] , \ScanLink250[16] , \ScanLink18[27] , 
        \wRegInTop_4_5[22] , \ScanLink94[5] , \wRegInTop_7_26[28] , 
        \wRegInTop_7_53[18] , \wRegInTop_7_70[30] , \ScanLink213[23] , 
        \wRegInTop_6_28[18] , \wRegOut_7_24[7] , \wRegInTop_7_26[31] , 
        \ScanLink230[12] , \ScanLink195[15] , \ScanLink21[4] , 
        \wRegOut_6_38[24] , \wRegInBot_6_47[3] , \wRegInTop_7_70[29] , 
        \wRegOut_7_15[25] , \ScanLink245[22] , \wRegOut_7_36[14] , 
        \wRegOut_7_60[15] , \wRegOut_7_23[20] , \wRegOut_7_43[24] , 
        \wRegOut_6_58[20] , \wRegInTop_1_0[30] , \wRegInTop_1_0[29] , 
        \wRegInBot_1_0[18] , \wRegOut_2_1[3] , \wRegInBot_2_3[20] , 
        \wRegInBot_3_0[7] , \wRegOut_3_1[16] , \ScanLink18[14] , 
        \wRegInTop_4_5[11] , \wRegOut_4_12[2] , \wRegOut_7_1[18] , 
        \wRegOut_5_9[0] , \ScanLink96[25] , \wRegOut_7_56[10] , 
        \wRegOut_7_75[21] , \wRegOut_7_91[6] , \wRegInBot_5_13[18] , 
        \wRegInBot_5_30[30] , \wRegInBot_5_30[29] , \ScanLink102[9] , 
        \ScanLink138[26] , \wRegInTop_7_51[8] , \ScanLink158[22] , 
        \ScanLink83[11] , \wRegOut_6_62[6] , \wRegOut_7_43[0] , 
        \wRegInBot_6_20[4] , \wRegInBot_6_48[28] , \ScanLink213[10] , 
        \wRegInBot_6_23[7] , \wRegInBot_6_48[31] , \wRegOut_6_61[5] , 
        \ScanLink195[26] , \ScanLink230[21] , \ScanLink245[11] , 
        \wRegOut_7_40[3] , \ScanLink180[12] , \ScanLink250[25] , 
        \ScanLink225[15] , \wRegOut_3_5[27] , \wRegInTop_4_1[20] , 
        \ScanLink22[7] , \wRegOut_4_11[1] , \wRegOut_5_16[24] , 
        \wRegOut_5_20[21] , \ScanLink78[10] , \ScanLink206[24] , 
        \wRegInTop_6_2[15] , \wRegOut_7_92[5] , \wRegOut_5_30[7] , 
        \wRegEnTop_6_20[0] , \wRegInBot_6_39[29] , \ScanLink217[21] , 
        \ScanLink69[15] , \wRegInBot_6_39[30] , \wRegOut_6_45[3] , 
        \ScanLink191[17] , \wRegOut_7_64[5] , \ScanLink234[10] , 
        \ScanLink245[9] , \ScanLink184[23] , \ScanLink241[20] , 
        \ScanLink221[24] , \wRegInBot_5_0[3] , \wRegInTop_5_1[5] , 
        \wRegOut_5_14[1] , \wRegOut_5_24[10] , \wRegEnTop_7_25[0] , 
        \ScanLink202[15] , \wRegOut_7_109[30] , \ScanLink254[14] , 
        \wRegOut_7_109[29] , \wRegOut_5_12[15] , \wRegInTop_6_6[24] , 
        \wRegInTop_3_1[1] , \wRegOut_4_7[9] , \wRegInTop_3_2[2] , 
        \wRegInBot_3_3[4] , \wRegInTop_5_2[6] , \wRegOut_5_31[24] , 
        \ScanLink138[3] , \wRegInBot_5_3[0] , \wRegOut_7_64[24] , 
        \wRegOut_5_17[2] , \wRegOut_7_11[14] , \wRegOut_6_29[21] , 
        \wRegOut_6_49[25] , \wRegOut_7_47[15] , \wRegInTop_6_49[7] , 
        \wRegOut_7_32[25] , \wRegOut_7_52[21] , \wRegInTop_7_68[1] , 
        \wRegOut_7_5[29] , \wRegOut_7_27[11] , \wRegOut_7_71[10] , 
        \wRegInBot_5_17[30] , \ScanLink92[14] , \wRegOut_6_46[0] , 
        \wRegOut_7_5[30] , \wRegOut_7_67[6] , \wRegInTop_7_9[27] , 
        \ScanLink149[27] , \wRegInBot_5_17[29] , \wRegInTop_6_54[8] , 
        \ScanLink129[23] , \wRegInTop_5_18[5] , \ScanLink87[20] , 
        \wRegInBot_2_3[13] , \wRegOut_3_5[14] , \wRegInBot_4_4[19] , 
        \wRegInBot_4_13[1] , \wRegOut_5_12[26] , \ScanLink62[5] , 
        \wRegOut_7_3[8] , \wRegOut_5_31[17] , \wRegOut_5_24[23] , 
        \wRegInBot_6_4[2] , \wRegInTop_6_5[4] , \wRegInTop_7_113[4] , 
        \wRegEnTop_5_31[0] , \wRegInTop_6_6[17] , \wRegOut_6_21[7] , 
        \ScanLink254[27] , \wRegInBot_6_63[5] , \ScanLink184[10] , 
        \ScanLink221[17] , \wRegInTop_4_1[13] , \wRegInTop_7_12[9] , 
        \ScanLink202[26] , \wRegInTop_5_21[18] , \ScanLink69[26] , 
        \wRegInTop_6_59[19] , \ScanLink141[8] , \wRegInTop_7_57[29] , 
        \wRegInTop_7_22[19] , \ScanLink217[12] , \wRegInTop_7_57[30] , 
        \wRegInTop_7_74[18] , \ScanLink241[13] , \ScanLink191[24] , 
        \ScanLink234[23] , \ScanLink129[10] , \wRegOut_7_127[8] , 
        \wRegInTop_3_2[16] , \wRegOut_4_6[11] , \wRegInBot_4_10[2] , 
        \ScanLink61[6] , \wRegOut_6_22[4] , \ScanLink87[13] , \ScanLink92[27] , 
        \wRegInBot_6_60[6] , \wRegInTop_7_9[14] , \ScanLink149[14] , 
        \wRegOut_7_27[22] , \wRegInBot_5_31[4] , \wRegOut_7_52[12] , 
        \wRegInTop_7_110[7] , \wRegInTop_6_6[7] , \wRegOut_6_29[12] , 
        \wRegOut_6_49[16] , \wRegOut_7_11[27] , \wRegOut_7_71[23] , 
        \wRegOut_7_64[17] , \wRegInBot_6_7[1] , \wRegOut_7_32[16] , 
        \wRegOut_7_47[26] , \ScanLink243[7] , \wRegInBot_6_8[11] , 
        \wRegInTop_6_51[5] , \ScanLink123[2] , \wRegInTop_7_70[3] , 
        \wRegInTop_6_11[20] , \wRegOut_7_121[27] , \wRegInTop_6_32[11] , 
        \wRegInBot_1_1[21] , \wRegOut_2_0[22] , \wRegOut_2_1[31] , 
        \ScanLink5[14] , \wRegOut_2_2[0] , \wRegInBot_3_6[9] , 
        \wRegOut_4_1[7] , \wRegOut_6_1[15] , \wRegInTop_6_27[25] , 
        \wRegInBot_6_27[22] , \wRegInTop_6_47[21] , \wRegInBot_6_52[12] , 
        \wRegInTop_7_49[11] , \wRegOut_7_102[16] , \wRegInBot_6_47[26] , 
        \wRegOut_7_117[22] , \wRegInBot_6_32[16] , \wRegInTop_6_52[15] , 
        \wRegInTop_7_29[15] , \wRegInBot_4_12[26] , \wRegInTop_5_4[8] , 
        \wRegInBot_6_11[27] , \wRegOut_5_9[12] , \wRegInTop_7_91[21] , 
        \wRegEnBot_3_0[0] , \wRegOut_4_2[4] , \wRegInTop_7_2[18] , 
        \wRegInTop_4_12[21] , \ScanLink114[19] , \ScanLink161[29] , 
        \wRegInTop_7_84[15] , \ScanLink137[31] , \ScanLink137[28] , 
        \ScanLink142[18] , \ScanLink161[30] , \wRegOut_7_61[8] , 
        \ScanLink240[4] , \wRegInTop_3_2[25] , \ScanLink17[30] , 
        \wRegInBot_5_0[16] , \ScanLink41[28] , \wRegInTop_6_52[6] , 
        \wRegInTop_7_73[0] , \ScanLink120[1] , \wRegInBot_6_32[25] , 
        \wRegInTop_7_29[26] , \wRegInTop_6_52[26] , \wRegOut_7_5[6] , 
        \ScanLink17[29] , \ScanLink34[18] , \wRegInBot_6_47[15] , 
        \ScanLink41[31] , \wRegInTop_6_27[16] , \wRegOut_7_117[11] , 
        \ScanLink62[19] , \wRegInBot_6_11[14] , \wRegOut_6_1[26] , 
        \wRegEnTop_6_6[0] , \wRegInTop_6_11[13] , \ScanLink195[0] , 
        \ScanLink209[19] , \wRegOut_7_121[14] , \wRegInBot_6_27[11] , 
        \wRegInTop_6_47[12] , \wRegInTop_6_32[22] , \wRegInTop_7_49[22] , 
        \wRegOut_7_102[25] , \wRegInBot_6_52[21] , \wRegOut_4_6[22] , 
        \wRegOut_5_19[19] , \wRegInBot_5_29[6] , \ScanLink79[4] , 
        \wRegOut_7_94[30] , \wRegInTop_7_114[30] , \wRegOut_6_27[9] , 
        \ScanLink227[3] , \wRegInTop_7_108[5] , \wRegOut_7_122[5] , 
        \wRegOut_7_94[29] , \wRegInTop_7_114[29] , \wRegInBot_6_8[22] , 
        \wRegInTop_6_35[1] , \wRegInTop_7_14[7] , \ScanLink147[6] , 
        \wRegOut_6_14[31] , \wRegOut_6_14[28] , \wRegOut_6_42[30] , 
        \ScanLink224[0] , \wRegOut_6_61[18] , \wRegOut_7_39[30] , 
        \wRegInTop_6_36[2] , \wRegOut_6_37[19] , \wRegOut_6_42[29] , 
        \ScanLink144[5] , \wRegOut_7_39[29] , \wRegOut_7_121[6] , 
        \wRegInTop_7_17[4] , \wRegOut_2_1[28] , \ScanLink5[27] , 
        \wRegInBot_5_0[25] , \wRegInBot_2_2[19] , \wRegInTop_4_12[12] , 
        \wRegInTop_7_84[26] , \wRegInBot_4_12[15] , \wRegInTop_6_0[9] , 
        \ScanLink67[8] , \ScanLink99[18] , \wRegOut_6_39[5] , 
        \wRegOut_7_18[3] , \wRegOut_7_6[5] , \wRegInTop_7_116[9] , 
        \ScanLink196[3] , \wRegInTop_7_91[12] , \wRegOut_5_9[21] , 
        \ScanLink86[19] , \wRegOut_6_28[18] , \wRegOut_7_4[10] , 
        \wRegOut_7_26[31] , \wRegOut_7_26[28] , \wRegOut_7_70[29] , 
        \wRegOut_7_53[18] , \wRegOut_7_70[30] , \ScanLink180[7] , 
        \wRegOut_7_13[8] , \ScanLink232[4] , \ScanLink15[8] , 
        \wRegInTop_4_0[19] , \wRegInBot_4_5[13] , \wRegOut_5_3[14] , 
        \wRegInTop_5_16[17] , \wRegInBot_5_16[10] , \wRegInTop_5_20[12] , 
        \wRegInBot_5_20[15] , \wRegInTop_6_20[6] , \ScanLink152[1] , 
        \wRegInTop_6_38[17] , \wRegInBot_6_58[14] , \wRegInTop_7_43[17] , 
        \wRegOut_7_108[10] , \wRegInTop_7_15[16] , \wRegInTop_7_36[27] , 
        \wRegInTop_7_60[26] , \ScanLink231[7] , \wRegInTop_6_23[5] , 
        \wRegInTop_7_75[12] , \ScanLink235[29] , \ScanLink240[19] , 
        \wRegInTop_7_56[23] , \wRegOut_5_3[27] , \wRegInTop_5_16[24] , 
        \wRegInBot_5_20[26] , \wRegOut_5_25[30] , \wRegInBot_6_2[17] , 
        \wRegInTop_6_8[1] , \ScanLink151[2] , \wRegInBot_6_9[7] , 
        \wRegInBot_6_38[10] , \wRegInTop_7_23[13] , \wRegInTop_6_58[13] , 
        \ScanLink216[18] , \ScanLink235[30] , \wRegOut_5_25[29] , 
        \ScanLink183[4] , \wRegInBot_5_16[23] , \wRegInBot_6_14[8] , 
        \ScanLink128[30] , \wRegInTop_5_20[21] , \wRegInTop_6_44[2] , 
        \ScanLink128[29] , \wRegInTop_7_65[4] , \ScanLink136[5] , 
        \wRegInBot_4_5[20] , \wRegInTop_5_15[0] , \wRegInTop_5_16[3] , 
        \wRegInBot_6_2[24] , \wRegOut_6_48[6] , \wRegOut_7_4[23] , 
        \wRegOut_7_69[0] , \ScanLink128[9] , \wRegOut_5_19[4] , 
        \wRegInBot_6_38[23] , \wRegOut_6_55[9] , \wRegInTop_7_75[21] , 
        \ScanLink255[3] , \wRegInTop_7_23[20] , \wRegInTop_6_38[24] , 
        \wRegInTop_6_47[1] , \wRegInTop_6_58[20] , \ScanLink135[6] , 
        \wRegInTop_7_56[10] , \ScanLink185[30] , \wRegInTop_7_36[14] , 
        \wRegInTop_7_66[7] , \wRegInBot_6_58[27] , \wRegInTop_7_43[24] , 
        \ScanLink185[29] , \wRegOut_7_108[23] , \wRegInTop_4_13[18] , 
        \wRegInBot_5_27[0] , \ScanLink77[2] , \wRegInTop_7_15[25] , 
        \wRegInTop_7_60[15] , \ScanLink136[11] , \ScanLink115[20] , 
        \ScanLink143[21] , \wRegInTop_7_106[3] , \ScanLink229[5] , 
        \wRegInTop_5_4[25] , \ScanLink98[12] , \wRegOut_6_36[13] , 
        \ScanLink100[14] , \wRegInTop_7_3[21] , \ScanLink160[10] , 
        \ScanLink123[25] , \ScanLink149[0] , \ScanLink175[24] , 
        \wRegInTop_7_90[18] , \ScanLink156[15] , \ScanLink186[9] , 
        \wRegOut_6_15[22] , \wRegOut_6_43[23] , \wRegOut_7_38[23] , 
        \wRegOut_6_34[0] , \wRegOut_6_60[12] , \wRegOut_7_15[6] , 
        \wRegInBot_3_6[25] , \wRegOut_4_7[31] , \wRegEnBot_6_9[0] , 
        \wRegOut_6_23[27] , \wRegInTop_6_26[8] , \wRegEnBot_6_38[0] , 
        \wRegOut_7_58[27] , \wRegInBot_6_9[28] , \wRegOut_6_37[3] , 
        \wRegOut_6_56[17] , \wRegOut_7_8[3] , \wRegOut_7_16[5] , 
        \ScanLink237[9] , \wRegOut_7_95[23] , \wRegInTop_7_115[23] , 
        \ScanLink198[5] , \wRegOut_4_7[28] , \wRegOut_5_18[13] , 
        \wRegInTop_7_123[26] , \wRegInBot_6_9[31] , \wRegOut_7_80[17] , 
        \wRegInTop_7_100[17] , \ScanLink16[23] , \ScanLink63[13] , 
        \ScanLink35[12] , \ScanLink40[22] , \ScanLink74[1] , 
        \wRegEnTop_7_57[0] , \ScanLink55[16] , \wRegInBot_5_24[3] , 
        \wRegInTop_6_38[4] , \wRegInTop_6_46[18] , \wRegInTop_7_105[0] , 
        \wRegInTop_7_19[2] , \ScanLink208[13] , \wRegInTop_6_33[28] , 
        \wRegInBot_1_1[12] , \wRegOut_2_0[11] , \ScanLink20[26] , 
        \wRegInTop_6_10[19] , \ScanLink76[27] , \wRegInTop_7_48[28] , 
        \wRegInTop_6_33[31] , \wRegOut_6_50[4] , \wRegInTop_7_48[31] , 
        \wRegOut_7_71[2] , \ScanLink10[5] , \ScanLink13[6] , 
        \wRegInTop_5_4[16] , \wRegInBot_6_12[6] , \wRegOut_6_23[14] , 
        \wRegOut_6_56[24] , \wRegOut_7_58[14] , \wRegOut_6_43[10] , 
        \wRegOut_5_8[18] , \wRegOut_6_15[11] , \wRegOut_6_36[20] , 
        \wRegOut_7_38[10] , \wRegOut_6_60[21] , \ScanLink175[17] , 
        \ScanLink100[27] , \ScanLink156[26] , \ScanLink98[21] , 
        \ScanLink123[16] , \ScanLink136[22] , \ScanLink143[12] , 
        \ScanLink115[13] , \wRegInTop_7_3[12] , \ScanLink160[23] , 
        \ScanLink20[15] , \wRegInBot_6_53[18] , \wRegInBot_3_6[16] , 
        \ScanLink16[10] , \ScanLink55[25] , \wRegInBot_6_26[28] , 
        \ScanLink208[20] , \ScanLink76[14] , \wRegInBot_6_26[31] , 
        \ScanLink35[21] , \ScanLink63[20] , \wRegOut_7_116[31] , 
        \ScanLink40[11] , \wRegOut_7_116[28] , \wRegOut_7_80[24] , 
        \wRegInTop_7_123[15] , \ScanLink24[24] , \wRegOut_5_18[20] , 
        \wRegOut_6_53[7] , \wRegOut_7_72[1] , \wRegInTop_7_100[24] , 
        \ScanLink51[14] , \wRegInBot_6_11[5] , \ScanLink133[8] , 
        \wRegOut_7_95[10] , \wRegInTop_7_115[10] , \wRegInTop_7_59[0] , 
        \wRegInTop_7_60[9] , \wRegInTop_7_96[9] , \wRegInBot_6_22[19] , 
        \wRegInBot_6_57[29] , \wRegOut_5_1[8] , \ScanLink72[25] , 
        \ScanLink67[11] , \wRegInBot_6_57[30] , \ScanLink12[21] , 
        \wRegInBot_4_6[2] , \wRegInTop_4_7[4] , \wRegOut_7_84[1] , 
        \ScanLink44[20] , \wRegOut_5_26[3] , \wRegInBot_3_2[27] , 
        \wRegOut_4_12[21] , \ScanLink31[10] , \ScanLink34[3] , 
        \ScanLink219[25] , \wRegOut_7_112[19] , \wRegInTop_5_29[4] , 
        \wRegInTop_7_127[24] , \wRegOut_7_84[15] , \wRegInTop_7_104[15] , 
        \wRegInTop_4_4[7] , \wRegInBot_4_5[1] , \wRegInTop_5_0[27] , 
        \wRegInTop_6_8[20] , \wRegOut_7_56[7] , \wRegOut_6_27[25] , 
        \wRegInBot_6_35[3] , \wRegInTop_7_111[21] , \wRegInTop_7_88[5] , 
        \wRegOut_7_91[21] , \wRegOut_6_32[11] , \wRegOut_6_52[15] , 
        \wRegOut_7_29[15] , \wRegOut_7_49[11] , \ScanLink37[0] , 
        \wRegEnBot_5_29[0] , \wRegOut_6_11[20] , \wRegOut_6_47[21] , 
        \ScanLink89[24] , \wRegInBot_6_36[0] , \wRegOut_7_55[4] , 
        \ScanLink104[16] , \ScanLink171[26] , \ScanLink109[2] , 
        \ScanLink127[27] , \ScanLink152[17] , \wRegOut_5_25[0] , 
        \ScanLink132[13] , \ScanLink147[23] , \ScanLink111[22] , 
        \wRegOut_7_87[2] , \wRegInTop_7_7[23] , \wRegInTop_6_8[13] , 
        \ScanLink164[12] , \wRegOut_7_91[12] , \wRegInTop_7_111[12] , 
        \wRegOut_0_0[9] , \wRegOut_0_0[0] , \wRegInTop_1_0[2] , 
        \wRegInBot_3_2[14] , \ScanLink82[1] , \wRegInTop_7_127[17] , 
        \wRegOut_7_84[26] , \wRegOut_7_116[9] , \ScanLink12[12] , 
        \wRegOut_4_3[19] , \wRegOut_4_12[12] , \wRegOut_7_32[3] , 
        \wRegOut_6_13[5] , \wRegInBot_6_51[7] , \wRegInTop_7_104[26] , 
        \ScanLink24[17] , \ScanLink31[23] , \ScanLink67[22] , \ScanLink44[13] , 
        \ScanLink50[7] , \wRegInTop_6_37[19] , \wRegInTop_7_3[5] , 
        \ScanLink219[16] , \wRegInTop_6_14[31] , \wRegEnTop_6_52[0] , 
        \wRegInTop_5_19[19] , \ScanLink51[27] , \wRegOut_6_5[9] , 
        \wRegInTop_7_121[6] , \wRegInTop_6_42[29] , \ScanLink72[16] , 
        \wRegInTop_6_14[28] , \wRegInTop_7_39[29] , \wRegInTop_6_42[30] , 
        \wRegInTop_6_61[18] , \wRegInTop_7_0[6] , \ScanLink132[20] , 
        \ScanLink147[10] , \wRegInTop_7_39[30] , \wRegInTop_7_7[10] , 
        \ScanLink89[17] , \ScanLink111[11] , \ScanLink164[21] , 
        \ScanLink171[15] , \ScanLink104[25] , \ScanLink152[24] , 
        \wRegInTop_7_94[29] , \wRegInBot_1_1[4] , \ScanLink53[4] , 
        \ScanLink127[14] , \wRegInTop_7_94[30] , \wRegOut_7_108[5] , 
        \wRegInTop_7_122[5] , \wRegInBot_2_0[8] , \wRegInTop_4_13[3] , 
        \wRegInTop_5_0[14] , \wRegOut_6_47[12] , \wRegOut_6_10[6] , 
        \wRegOut_6_11[13] , \wRegOut_6_32[22] , \wRegInTop_7_23[8] , 
        \ScanLink170[9] , \wRegOut_7_49[22] , \wRegOut_7_31[0] , 
        \ScanLink81[2] , \wRegInBot_6_52[4] , \wRegOut_6_27[16] , 
        \wRegOut_6_52[26] , \wRegOut_7_29[26] , \wRegEnBot_6_60[0] , 
        \wRegInTop_2_3[11] , \wRegOut_3_7[2] , \wRegOut_4_8[15] , 
        \wRegOut_5_7[6] , \wRegInBot_6_6[15] , \wRegInTop_7_90[7] , 
        \wRegInBot_4_1[11] , \wRegEnTop_4_4[0] , \wRegInTop_6_29[21] , 
        \ScanLink111[0] , \wRegInBot_6_49[22] , \wRegInTop_7_71[10] , 
        \wRegInTop_6_63[7] , \wRegInTop_7_42[1] , \wRegOut_7_119[26] , 
        \wRegInTop_7_52[21] , \wRegInBot_6_29[26] , \wRegInTop_6_49[25] , 
        \wRegInTop_7_27[11] , \wRegInTop_7_47[15] , \wRegInTop_7_11[14] , 
        \wRegInTop_7_32[25] , \wRegOut_7_50[9] , \ScanLink181[18] , 
        \wRegInTop_7_64[24] , \wRegInTop_5_31[24] , \ScanLink112[3] , 
        \wRegInTop_6_60[4] , \wRegInTop_7_41[2] , \wRegOut_3_4[1] , 
        \wRegInTop_4_10[0] , \wRegOut_5_7[16] , \wRegInTop_5_12[15] , 
        \wRegInBot_5_24[17] , \ScanLink159[31] , \wRegInBot_5_12[12] , 
        \wRegInTop_5_24[10] , \ScanLink159[28] , \wRegInTop_5_31[6] , 
        \wRegInBot_5_31[23] , \wRegInTop_7_93[4] , \wRegOut_5_4[5] , 
        \wRegInBot_4_1[22] , \wRegInTop_4_2[9] , \ScanLink79[30] , 
        \wRegInTop_6_49[16] , \wRegOut_7_0[12] , \wRegInTop_7_26[5] , 
        \wRegInTop_7_32[16] , \ScanLink175[4] , \ScanLink79[29] , 
        \wRegInBot_6_29[15] , \wRegInTop_7_47[26] , \wRegInTop_4_4[31] , 
        \wRegInBot_6_57[9] , \wRegInTop_7_11[27] , \wRegInTop_7_64[17] , 
        \ScanLink212[30] , \ScanLink215[1] , \ScanLink231[18] , 
        \wRegInTop_4_4[28] , \wRegInTop_7_27[22] , \wRegInTop_7_71[23] , 
        \ScanLink244[28] , \ScanLink212[29] , \wRegOut_7_119[15] , 
        \wRegOut_4_8[26] , \wRegInBot_6_6[26] , \wRegInTop_6_29[12] , 
        \wRegInBot_6_49[11] , \wRegInTop_7_52[12] , \wRegOut_7_110[7] , 
        \ScanLink244[31] , \wRegOut_5_21[18] , \ScanLink56[9] , 
        \wRegOut_7_29[2] , \ScanLink99[0] , \wRegOut_6_3[7] , 
        \wRegOut_7_57[30] , \wRegOut_7_74[18] , \wRegInTop_7_127[8] , 
        \wRegInBot_1_1[31] , \wRegInBot_1_1[28] , \wRegOut_2_0[18] , 
        \ScanLink4[17] , \wRegInTop_2_3[22] , \wRegOut_5_7[25] , 
        \wRegInBot_5_12[21] , \wRegOut_6_0[4] , \wRegOut_6_59[19] , 
        \wRegOut_7_22[19] , \wRegInTop_7_38[9] , \wRegOut_7_57[29] , 
        \wRegOut_7_0[21] , \wRegInTop_7_6[8] , \wRegInBot_6_49[5] , 
        \wRegInTop_5_24[23] , \wRegInBot_5_31[10] , \ScanLink82[28] , 
        \wRegInTop_7_25[6] , \ScanLink176[7] , \ScanLink82[31] , 
        \ScanLink9[9] , \wRegInTop_5_12[26] , \ScanLink48[5] , 
        \wRegInBot_5_18[7] , \wRegInBot_5_24[24] , \wRegInTop_5_31[17] , 
        \wRegOut_7_113[4] , \wRegOut_6_16[8] , \ScanLink216[2] , 
        \wRegInTop_5_9[4] , \wRegEnBot_5_10[0] , \wRegOut_6_36[29] , 
        \wRegInTop_6_42[5] , \wRegOut_6_60[31] , \wRegInTop_7_63[3] , 
        \wRegOut_6_43[19] , \ScanLink130[2] , \wRegOut_7_38[19] , 
        \wRegOut_6_15[18] , \wRegOut_6_36[30] , \wRegOut_6_60[28] , 
        \ScanLink250[7] , \wRegInBot_5_1[15] , \ScanLink4[24] , 
        \wRegInTop_3_3[15] , \ScanLink16[19] , \wRegInTop_4_13[22] , 
        \wRegInBot_5_8[2] , \wRegInTop_5_13[7] , \ScanLink98[31] , 
        \ScanLink98[28] , \wRegInTop_7_85[16] , \wRegInBot_4_13[25] , 
        \ScanLink35[31] , \wRegOut_5_8[11] , \wRegInTop_7_90[22] , 
        \ScanLink35[28] , \wRegInTop_5_10[4] , \ScanLink63[29] , 
        \wRegInBot_6_10[24] , \ScanLink40[18] , \ScanLink63[30] , 
        \wRegInTop_6_26[26] , \wRegInBot_6_46[25] , \wRegOut_7_116[21] , 
        \wRegInBot_6_33[15] , \wRegOut_6_0[16] , \wRegInTop_6_33[12] , 
        \wRegInTop_6_53[16] , \wRegInTop_7_28[16] , \wRegInTop_6_10[23] , 
        \wRegInBot_6_26[21] , \wRegInTop_6_46[22] , \wRegInBot_6_53[11] , 
        \wRegInTop_7_48[12] , \wRegOut_7_103[15] , \ScanLink208[29] , 
        \wRegInTop_6_41[6] , \ScanLink133[1] , \ScanLink208[30] , 
        \wRegOut_7_120[24] , \wRegOut_7_95[19] , \wRegInTop_7_115[19] , 
        \wRegInTop_7_60[0] , \wRegOut_4_7[12] , \wRegOut_5_18[30] , 
        \wRegInBot_6_9[12] , \ScanLink253[4] , \wRegInTop_4_13[11] , 
        \wRegInBot_4_13[16] , \wRegOut_5_18[29] , \wRegOut_7_72[8] , 
        \wRegInTop_7_90[11] , \wRegOut_5_8[22] , \wRegInBot_5_27[9] , 
        \ScanLink115[30] , \ScanLink136[18] , \ScanLink149[9] , 
        \ScanLink186[0] , \wRegInTop_7_3[31] , \ScanLink143[28] , 
        \wRegInTop_7_85[25] , \wRegInBot_5_1[26] , \wRegOut_6_29[6] , 
        \ScanLink115[29] , \wRegInTop_7_3[28] , \ScanLink143[31] , 
        \ScanLink160[19] , \wRegInTop_3_3[26] , \wRegOut_4_7[21] , 
        \wRegInBot_6_9[21] , \wRegInTop_6_25[2] , \wRegInTop_6_26[1] , 
        \ScanLink154[6] , \wRegOut_6_34[9] , \ScanLink234[3] , 
        \ScanLink157[5] , \ScanLink237[0] , \wRegOut_6_0[25] , \ScanLink69[7] , 
        \wRegInBot_6_26[12] , \wRegInTop_6_46[11] , \ScanLink185[3] , 
        \wRegInTop_7_118[6] , \wRegInTop_6_33[21] , \wRegInTop_7_48[21] , 
        \wRegOut_7_103[26] , \wRegInTop_6_10[10] , \wRegInBot_6_53[22] , 
        \wRegOut_7_120[17] , \wRegInBot_2_2[23] , \wRegOut_4_9[6] , 
        \wRegInBot_6_10[17] , \ScanLink74[8] , \wRegInBot_6_33[26] , 
        \wRegInTop_7_28[25] , \wRegEnTop_7_98[0] , \wRegInTop_6_26[15] , 
        \wRegInBot_6_46[16] , \wRegInTop_6_53[25] , \wRegInTop_7_105[9] , 
        \wRegOut_7_116[12] , \ScanLink86[23] , \wRegInBot_2_2[10] , 
        \wRegOut_3_4[24] , \ScanLink15[1] , \wRegInTop_5_15[9] , 
        \wRegInTop_5_20[31] , \wRegInTop_5_20[28] , \ScanLink128[20] , 
        \wRegInBot_6_14[1] , \ScanLink93[17] , \wRegOut_6_56[3] , 
        \ScanLink148[24] , \wRegOut_7_77[5] , \wRegInTop_7_8[24] , 
        \wRegOut_6_28[22] , \wRegInTop_6_59[4] , \wRegOut_7_53[22] , 
        \wRegOut_7_70[13] , \wRegInTop_7_78[2] , \wRegOut_7_26[12] , 
        \wRegEnTop_7_36[0] , \ScanLink16[2] , \wRegOut_5_13[16] , 
        \wRegOut_5_30[27] , \wRegOut_6_48[26] , \wRegOut_7_46[16] , 
        \ScanLink128[0] , \wRegOut_7_10[17] , \wRegOut_7_33[26] , 
        \wRegOut_7_65[27] , \wRegInTop_6_7[27] , \wRegOut_7_69[9] , 
        \ScanLink248[5] , \wCtrlOut_1[0] , \wRegInBot_4_5[30] , 
        \wRegOut_5_25[13] , \ScanLink203[16] , \wRegInTop_6_47[8] , 
        \ScanLink185[20] , \ScanLink220[27] , \wRegInTop_4_0[23] , 
        \wRegInBot_4_5[29] , \ScanLink68[16] , \wRegEnBot_6_59[0] , 
        \ScanLink255[17] , \wRegInTop_7_23[30] , \wRegInBot_6_17[2] , 
        \wRegOut_6_55[0] , \wRegInTop_6_58[30] , \ScanLink190[14] , 
        \wRegOut_7_74[6] , \ScanLink235[13] , \wRegInTop_7_75[28] , 
        \wRegInTop_6_58[29] , \wRegInTop_7_23[29] , \ScanLink240[23] , 
        \wRegInTop_7_75[31] , \ScanLink216[22] , \wRegInBot_5_21[7] , 
        \ScanLink71[5] , \wRegOut_6_48[15] , \wRegInTop_7_56[19] , 
        \wRegOut_7_10[24] , \wRegOut_7_33[15] , \wRegOut_7_46[25] , 
        \wRegOut_7_26[21] , \wRegOut_7_65[14] , \wRegOut_7_70[20] , 
        \wRegOut_7_4[19] , \wRegEnTop_5_22[0] , \wRegOut_6_28[11] , 
        \wRegOut_7_53[11] , \wRegInTop_7_100[4] , \ScanLink93[24] , 
        \wRegInTop_7_8[17] , \ScanLink148[17] , \ScanLink152[8] , 
        \wRegOut_6_32[7] , \wRegOut_3_0[26] , \wRegOut_3_4[17] , 
        \wRegInTop_4_0[10] , \wRegInBot_5_16[19] , \ScanLink86[10] , 
        \wRegOut_7_13[1] , \ScanLink68[25] , \ScanLink128[13] , 
        \ScanLink240[10] , \ScanLink190[27] , \ScanLink235[20] , 
        \wRegInTop_6_8[8] , \wRegOut_6_31[4] , \wRegInBot_6_38[19] , 
        \ScanLink203[25] , \ScanLink216[11] , \wRegOut_7_108[19] , 
        \wRegOut_7_10[2] , \ScanLink255[24] , \ScanLink185[13] , 
        \ScanLink220[14] , \ScanLink19[24] , \wRegOut_5_13[25] , 
        \wRegInBot_5_22[4] , \wRegOut_5_25[20] , \wRegInTop_6_7[14] , 
        \wRegEnTop_7_109[0] , \wRegOut_5_30[14] , \ScanLink72[6] , 
        \wRegInTop_7_103[7] , \wRegOut_6_15[2] , \wRegOut_7_34[4] , 
        \ScanLink194[16] , \ScanLink215[8] , \ScanLink231[11] , 
        \wRegInTop_4_4[21] , \ScanLink84[6] , \wRegInBot_6_57[0] , 
        \ScanLink244[21] , \wRegInBot_6_49[18] , \ScanLink212[20] , 
        \ScanLink181[22] , \ScanLink207[14] , \ScanLink224[25] , 
        \wRegOut_5_17[14] , \wRegOut_5_21[11] , \ScanLink56[0] , 
        \wRegInTop_6_3[25] , \ScanLink79[20] , \ScanLink208[7] , 
        \ScanLink251[15] , \ScanLink99[9] , \wRegInTop_7_5[2] , 
        \ScanLink168[2] , \wRegInTop_7_127[1] , \ScanLink55[3] , 
        \wRegOut_6_39[14] , \wRegOut_7_0[31] , \wRegOut_7_14[15] , 
        \wRegOut_7_37[24] , \wRegOut_7_42[14] , \wRegOut_7_61[25] , 
        \wRegInTop_7_124[2] , \wRegOut_7_74[11] , \wRegInTop_7_38[0] , 
        \wRegOut_7_57[20] , \wRegInBot_2_0[1] , \wRegInTop_2_1[7] , 
        \ScanLink9[0] , \wRegOut_6_16[1] , \wRegInTop_6_19[6] , 
        \ScanLink87[5] , \wRegOut_6_59[10] , \wRegOut_7_0[28] , 
        \wRegOut_7_22[10] , \wRegInTop_7_6[1] , \ScanLink139[16] , 
        \wRegOut_7_37[7] , \ScanLink97[15] , \wRegInBot_4_0[5] , 
        \ScanLink32[4] , \wRegInBot_5_12[31] , \wRegInBot_5_12[28] , 
        \wRegInBot_6_54[3] , \ScanLink82[21] , \wRegOut_5_20[4] , 
        \wRegInBot_5_31[19] , \ScanLink159[12] , \wRegInTop_4_1[3] , 
        \wRegOut_7_82[6] , \wRegOut_5_17[27] , \wRegInTop_6_3[16] , 
        \wRegInTop_2_2[4] , \wRegInTop_2_3[18] , \wRegOut_3_0[15] , 
        \wRegInBot_4_1[18] , \wRegOut_5_21[22] , \wRegInBot_6_33[4] , 
        \wRegOut_7_50[0] , \ScanLink207[27] , \ScanLink181[11] , 
        \ScanLink224[16] , \ScanLink251[26] , \ScanLink19[17] , 
        \ScanLink79[13] , \wRegInTop_7_52[31] , \wRegInTop_4_4[12] , 
        \wRegInTop_6_29[31] , \wRegInTop_7_71[19] , \ScanLink244[12] , 
        \wRegInTop_7_52[28] , \ScanLink194[25] , \ScanLink231[22] , 
        \wRegInTop_5_24[19] , \ScanLink82[12] , \wRegInTop_6_29[28] , 
        \wRegInTop_7_42[8] , \ScanLink111[9] , \wRegInTop_7_27[18] , 
        \ScanLink212[13] , \wRegInBot_6_30[7] , \wRegOut_7_53[3] , 
        \ScanLink159[21] , \wRegOut_3_4[8] , \ScanLink97[26] , 
        \ScanLink139[25] , \wRegInTop_4_2[0] , \wRegInBot_4_3[6] , 
        \wRegOut_7_74[22] , \wRegOut_7_81[5] , \ScanLink31[7] , 
        \wRegEnTop_6_33[0] , \wRegOut_7_22[23] , \wRegOut_5_23[7] , 
        \wRegOut_6_39[27] , \wRegOut_6_59[23] , \wRegOut_7_37[17] , 
        \wRegOut_7_57[13] , \wRegOut_7_42[27] , \wRegInBot_2_3[2] , 
        \wRegInTop_4_10[9] , \wRegOut_7_14[26] , \wRegOut_4_3[10] , 
        \ScanLink82[8] , \wRegOut_7_61[16] , \wRegOut_7_116[0] , 
        \ScanLink213[6] , \ScanLink0[15] , \wRegInTop_1_0[13] , 
        \wRegInTop_3_7[17] , \wRegInTop_7_20[2] , \ScanLink173[3] , 
        \wRegOut_6_4[14] , \wRegInTop_6_37[10] , \wRegInBot_6_57[13] , 
        \wRegOut_6_5[0] , \wRegInTop_6_42[20] , \wRegOut_7_107[17] , 
        \wRegInTop_6_14[21] , \wRegInBot_6_22[23] , \wRegInTop_7_39[20] , 
        \wRegInBot_6_14[26] , \wRegInTop_6_61[11] , \wRegOut_7_124[26] , 
        \wRegInBot_6_61[16] , \wRegInTop_5_19[10] , \wRegInBot_5_19[17] , 
        \wRegInTop_6_22[24] , \wRegInBot_6_42[27] , \wRegInTop_7_59[24] , 
        \wRegOut_7_112[23] , \wRegInBot_6_37[17] , \wRegInTop_6_57[14] , 
        \wRegOut_6_6[3] , \wRegInTop_7_94[20] , \ScanLink132[29] , 
        \ScanLink147[19] , \ScanLink164[31] , \ScanLink111[18] , 
        \wRegInTop_7_7[19] , \ScanLink164[28] , \wRegInTop_7_81[14] , 
        \ScanLink132[30] , \wRegOut_7_31[9] , \ScanLink210[5] , 
        \wRegInTop_1_0[20] , \wRegInBot_5_5[17] , \wRegInTop_7_23[1] , 
        \wRegOut_7_115[3] , \ScanLink170[0] , \wRegOut_3_1[5] , 
        \ScanLink44[30] , \wRegInBot_6_14[15] , \ScanLink67[18] , 
        \wRegOut_7_84[8] , \ScanLink12[31] , \ScanLink12[28] , 
        \ScanLink44[29] , \wRegInBot_6_28[5] , \wRegInBot_6_61[25] , 
        \wRegInBot_6_37[24] , \wRegInBot_6_42[14] , \wRegInTop_6_57[27] , 
        \wRegInTop_4_15[4] , \ScanLink31[19] , \wRegOut_7_112[10] , 
        \wRegOut_6_4[27] , \wRegInTop_6_22[17] , \wRegInTop_7_59[17] , 
        \wRegInBot_6_22[10] , \wRegInTop_6_42[13] , \wRegInTop_7_59[9] , 
        \wRegInTop_6_37[23] , \wRegInTop_7_39[13] , \wRegInTop_7_96[0] , 
        \wRegInBot_6_57[20] , \wRegOut_7_107[24] , \wRegInTop_6_61[22] , 
        \wRegOut_5_1[1] , \wRegInTop_6_14[12] , \wRegOut_7_99[7] , 
        \wRegOut_7_124[15] , \ScanLink0[26] , \wRegInTop_3_7[24] , 
        \wRegInTop_6_8[29] , \wRegInTop_7_111[28] , \wRegOut_7_91[28] , 
        \wRegOut_4_3[23] , \wRegOut_4_12[31] , \ScanLink29[5] , 
        \wRegInTop_6_8[30] , \wRegInTop_7_111[31] , \ScanLink117[7] , 
        \wRegInTop_7_44[6] , \wRegOut_7_91[31] , \wRegOut_4_12[28] , 
        \wRegInBot_5_5[24] , \wRegOut_6_11[30] , \wRegOut_6_11[29] , 
        \wRegOut_6_32[18] , \wRegOut_6_47[28] , \wRegOut_7_49[18] , 
        \wRegInBot_6_36[9] , \wRegOut_6_47[31] , \wRegEnTop_2_1[0] , 
        \wRegOut_3_2[6] , \wRegInBot_4_5[8] , \wRegEnBot_4_15[0] , 
        \ScanLink114[4] , \wRegInTop_7_47[5] , \ScanLink37[9] , 
        \wRegOut_5_25[9] , \wRegInTop_7_81[27] , \wRegInTop_5_19[23] , 
        \wRegOut_7_48[2] , \wRegInBot_5_19[24] , \wRegInTop_2_2[21] , 
        \wRegInTop_2_2[12] , \wRegOut_5_2[2] , \wRegInTop_7_94[13] , 
        \wRegOut_5_6[15] , \wRegInTop_5_21[5] , \wRegOut_6_58[30] , 
        \wRegOut_6_58[29] , \wRegOut_7_1[11] , \wRegOut_7_23[29] , 
        \wRegInTop_7_95[3] , \wRegOut_7_23[30] , \wRegOut_7_56[19] , 
        \wRegOut_7_75[31] , \wRegOut_7_75[28] , \wRegInTop_5_25[13] , 
        \wRegInTop_7_83[7] , \wRegInBot_5_30[20] , \ScanLink83[18] , 
        \wRegOut_7_43[9] , \wRegOut_5_9[9] , \wRegInTop_5_13[16] , 
        \wRegInBot_5_13[11] , \wRegInTop_5_30[27] , \ScanLink102[0] , 
        \wRegInTop_7_51[1] , \wRegInBot_4_0[12] , \wRegInBot_5_25[14] , 
        \ScanLink78[19] , \wRegInTop_7_65[27] , \wRegInTop_4_5[18] , 
        \wRegInBot_6_28[25] , \wRegInTop_6_48[26] , \wRegInTop_7_10[17] , 
        \wRegInTop_7_46[16] , \wRegInBot_6_48[21] , \wRegInTop_7_33[26] , 
        \wRegInTop_7_52[2] , \wRegOut_7_118[25] , \wRegOut_4_9[16] , 
        \wRegInTop_6_28[22] , \ScanLink101[3] , \wRegInTop_7_53[22] , 
        \wRegInTop_7_26[12] , \wRegInTop_7_70[13] , \ScanLink213[19] , 
        \ScanLink230[31] , \ScanLink230[28] , \ScanLink245[18] , 
        \wRegOut_4_11[8] , \wRegInTop_5_13[25] , \wRegOut_5_20[31] , 
        \wRegOut_5_20[28] , \wRegInBot_6_7[16] , \wRegInTop_7_80[4] , 
        \wRegInTop_5_22[6] , \ScanLink206[1] , \wRegInBot_6_44[9] , 
        \wRegOut_5_6[26] , \wRegInBot_5_13[22] , \wRegInTop_5_25[20] , 
        \wRegInBot_5_25[27] , \ScanLink58[6] , \wRegInTop_5_30[14] , 
        \wRegInBot_5_30[13] , \wRegInTop_7_35[5] , \wRegOut_7_103[7] , 
        \wRegInTop_6_14[3] , \ScanLink158[18] , \ScanLink166[4] , 
        \wRegEnTop_7_123[0] , \wRegOut_0_0[4] , \ScanLink1[8] , \ScanLink4[5] , 
        \ScanLink7[6] , \ScanLink45[9] , \wRegInBot_6_59[6] , 
        \wRegInBot_5_16[8] , \ScanLink89[3] , \wRegOut_7_1[22] , 
        \wRegOut_6_18[7] , \wRegOut_7_39[1] , \wRegInBot_3_3[24] , 
        \wRegInBot_4_0[21] , \wRegOut_4_9[25] , \wRegInBot_6_7[25] , 
        \ScanLink178[8] , \wRegInTop_6_28[11] , \wRegInBot_6_48[12] , 
        \wRegInTop_7_26[21] , \wRegInTop_7_53[11] , \wRegOut_7_118[16] , 
        \wRegOut_7_100[4] , \wRegInTop_7_10[24] , \ScanLink180[28] , 
        \wRegInTop_7_70[20] , \ScanLink205[2] , \wRegOut_4_2[29] , 
        \ScanLink27[3] , \wRegInTop_5_18[29] , \wRegInTop_6_17[0] , 
        \wRegInBot_6_28[16] , \wRegInTop_6_48[15] , \wRegInTop_7_65[14] , 
        \wRegInTop_7_33[15] , \ScanLink165[7] , \ScanLink180[31] , 
        \wRegInTop_7_36[6] , \ScanLink110[21] , \wRegInTop_7_8[7] , 
        \wRegInTop_7_46[25] , \wRegOut_7_97[1] , \wRegInTop_7_6[20] , 
        \wRegOut_7_58[8] , \ScanLink165[11] , \wRegOut_4_13[22] , 
        \wRegOut_4_14[5] , \wRegInTop_5_1[24] , \wRegInTop_5_18[30] , 
        \ScanLink133[10] , \wRegOut_6_10[23] , \ScanLink88[27] , 
        \ScanLink105[15] , \ScanLink119[1] , \ScanLink126[24] , 
        \ScanLink146[20] , \wRegInTop_7_85[9] , \ScanLink153[14] , 
        \ScanLink170[25] , \wRegInTop_7_95[19] , \wRegInBot_6_26[3] , 
        \wRegOut_7_45[7] , \wRegOut_6_33[12] , \wRegOut_6_46[22] , 
        \wRegOut_7_48[12] , \wRegInTop_6_9[23] , \wRegOut_6_26[26] , 
        \wRegInTop_7_98[6] , \wRegOut_6_53[16] , \wRegOut_7_28[16] , 
        \wRegOut_7_46[4] , \wRegInBot_6_25[0] , \wRegInTop_7_110[22] , 
        \wRegOut_7_85[16] , \wRegOut_7_90[22] , \wRegInTop_7_105[16] , 
        \ScanLink13[22] , \wRegOut_4_2[30] , \wRegInTop_7_126[27] , 
        \ScanLink24[0] , \ScanLink45[23] , \ScanLink218[26] , \ScanLink30[13] , 
        \ScanLink66[12] , \wRegOut_7_94[2] , \ScanLink25[27] , 
        \ScanLink50[17] , \wRegInTop_5_24[8] , \ScanLink73[26] , 
        \wRegInTop_6_60[28] , \wRegInTop_6_15[18] , \wRegInTop_6_36[30] , 
        \wRegInTop_6_43[19] , \wRegInTop_6_60[31] , \wRegInTop_7_49[3] , 
        \wRegInTop_6_36[29] , \wRegInTop_7_38[19] , \wRegInTop_5_1[17] , 
        \wRegOut_6_10[10] , \wRegOut_6_26[15] , \ScanLink91[1] , 
        \wRegOut_6_53[25] , \wRegOut_7_28[25] , \wRegInBot_6_42[7] , 
        \wRegOut_7_21[3] , \wRegOut_7_105[9] , \ScanLink43[7] , 
        \wRegOut_6_33[21] , \wRegOut_6_46[11] , \wRegEnTop_7_8[0] , 
        \ScanLink153[27] , \wRegOut_7_48[21] , \wRegInBot_5_13[5] , 
        \wRegEnTop_6_41[0] , \ScanLink126[17] , \wRegOut_7_118[6] , 
        \ScanLink88[14] , \ScanLink170[16] , \ScanLink105[26] , 
        \ScanLink110[12] , \wRegInTop_7_6[13] , \ScanLink165[22] , 
        \ScanLink133[23] , \ScanLink146[13] , \wRegOut_1_0[6] , 
        \wRegInBot_1_0[22] , \wRegInTop_1_1[19] , \ScanLink13[11] , 
        \ScanLink25[14] , \ScanLink40[4] , \ScanLink73[15] , 
        \wRegInBot_6_23[30] , \ScanLink30[20] , \wRegInBot_5_10[6] , 
        \wRegInBot_6_56[19] , \ScanLink50[24] , \wRegInBot_6_23[29] , 
        \wRegOut_7_113[29] , \ScanLink45[10] , \ScanLink218[15] , 
        \wRegOut_7_113[30] , \wRegInBot_3_3[17] , \ScanLink66[21] , 
        \wRegOut_7_22[0] , \wRegOut_7_85[25] , \wRegOut_4_13[11] , 
        \ScanLink54[15] , \wRegOut_6_8[5] , \ScanLink92[2] , 
        \wRegInBot_6_41[4] , \wRegInTop_7_105[25] , \wRegInTop_7_126[14] , 
        \wRegInTop_6_9[10] , \wRegInTop_7_30[8] , \ScanLink163[9] , 
        \ScanLink77[24] , \wRegOut_7_90[11] , \wRegInTop_7_110[11] , 
        \wRegInTop_6_28[7] , \wRegInBot_6_52[31] , \ScanLink195[9] , 
        \ScanLink209[10] , \wRegInBot_6_2[5] , \wRegInTop_6_3[3] , 
        \wRegInBot_6_27[18] , \wRegInBot_6_52[28] , \wRegInBot_1_0[11] , 
        \wRegOut_2_1[21] , \wRegInBot_3_7[26] , \ScanLink17[20] , 
        \ScanLink21[25] , \wRegInBot_4_15[6] , \ScanLink34[11] , 
        \ScanLink41[21] , \ScanLink64[2] , \wRegOut_7_117[18] , 
        \ScanLink62[10] , \wRegInTop_7_115[3] , \wRegOut_5_19[10] , 
        \wRegOut_7_81[14] , \wRegInTop_7_101[14] , \wRegOut_6_22[24] , 
        \wRegOut_6_27[0] , \wRegInTop_6_35[8] , \ScanLink188[6] , 
        \wRegInTop_7_122[25] , \wRegOut_7_59[24] , \wRegOut_7_94[20] , 
        \wRegInTop_7_114[20] , \wRegOut_6_57[14] , \wRegInBot_3_6[0] , 
        \wRegInBot_3_7[15] , \wRegInTop_5_5[26] , \wRegOut_6_14[21] , 
        \wRegOut_6_24[3] , \wRegOut_6_37[10] , \wRegOut_6_61[11] , 
        \ScanLink224[9] , \wRegOut_6_42[20] , \wRegOut_5_9[31] , 
        \wRegInTop_6_0[0] , \ScanLink122[26] , \ScanLink159[3] , 
        \wRegOut_7_39[20] , \ScanLink157[16] , \wRegOut_5_9[28] , 
        \wRegInBot_6_1[6] , \ScanLink101[17] , \ScanLink174[27] , 
        \ScanLink67[1] , \ScanLink99[11] , \ScanLink114[23] , \ScanLink239[6] , 
        \wRegInTop_7_2[22] , \ScanLink161[13] , \ScanLink137[12] , 
        \wRegEnTop_7_44[0] , \ScanLink142[22] , \wRegInTop_7_116[0] , 
        \wRegOut_7_62[2] , \wRegOut_7_81[27] , \wRegOut_7_94[13] , 
        \wRegInTop_7_114[13] , \ScanLink17[13] , \wRegOut_4_6[18] , 
        \ScanLink34[22] , \wRegOut_5_19[23] , \wRegOut_6_43[4] , 
        \wRegInTop_7_101[27] , \wRegInBot_6_8[18] , \wRegInTop_7_122[16] , 
        \ScanLink41[12] , \wRegInTop_3_7[6] , \ScanLink21[16] , 
        \wRegInBot_5_6[4] , \wRegInTop_5_7[2] , \ScanLink62[23] , 
        \wRegInTop_6_11[29] , \wRegInTop_6_11[30] , \ScanLink77[17] , 
        \wRegInTop_6_47[31] , \wRegInTop_6_32[18] , \wRegOut_5_12[6] , 
        \wRegInTop_7_49[18] , \wRegOut_2_1[12] , \wRegOut_2_2[9] , 
        \wRegInTop_3_4[5] , \wRegInBot_3_5[3] , \ScanLink54[26] , 
        \wRegInTop_6_47[28] , \ScanLink209[23] , \ScanLink99[22] , 
        \wRegInTop_7_2[11] , \ScanLink161[20] , \wRegInTop_4_12[31] , 
        \wRegInTop_4_12[28] , \ScanLink114[10] , \ScanLink137[21] , 
        \ScanLink142[11] , \wRegInTop_5_4[1] , \wRegOut_5_11[5] , 
        \ScanLink157[25] , \ScanLink122[15] , \wRegInTop_7_91[31] , 
        \wRegInBot_5_5[7] , \ScanLink101[24] , \ScanLink174[14] , 
        \wRegInTop_5_5[15] , \wRegOut_6_14[12] , \wRegOut_6_61[22] , 
        \wRegInTop_7_91[28] , \wRegOut_6_22[17] , \wRegOut_6_37[23] , 
        \wRegOut_6_42[13] , \ScanLink120[8] , \wRegOut_7_39[13] , 
        \wRegInTop_7_73[9] , \wRegOut_6_57[27] , \wRegOut_7_59[17] , 
        \wRegOut_6_40[7] , \wRegOut_7_61[1] , \wRegInBot_4_4[10] , 
        \wRegInBot_4_13[8] , \wRegOut_7_3[1] , \ScanLink193[7] , 
        \wRegInBot_6_3[14] , \wRegInTop_6_33[6] , \wRegInBot_6_39[13] , 
        \wRegInTop_7_12[0] , \wRegInTop_7_57[20] , \ScanLink141[1] , 
        \wRegInTop_7_22[10] , \wRegInTop_6_59[10] , \ScanLink184[19] , 
        \wRegInTop_7_61[25] , \wRegInTop_7_74[11] , \ScanLink221[4] , 
        \wRegOut_5_2[17] , \wRegInTop_5_17[14] , \wRegInTop_6_39[14] , 
        \wRegInTop_7_14[15] , \wRegInBot_6_59[17] , \wRegInTop_7_42[14] , 
        \wRegOut_7_109[13] , \wRegInTop_7_37[24] , \wRegOut_7_124[2] , 
        \wRegInTop_5_21[11] , \wRegInBot_5_21[16] , \wRegInTop_6_30[5] , 
        \ScanLink142[2] , \wRegInTop_7_11[3] , \ScanLink129[19] , 
        \wRegOut_7_127[1] , \ScanLink222[7] , \wRegInBot_5_17[13] , 
        \ScanLink190[4] , \wRegInTop_2_2[9] , \wRegInBot_2_3[30] , 
        \wRegInTop_3_1[8] , \wRegInTop_4_1[30] , \wRegInTop_4_1[29] , 
        \wRegInBot_4_4[23] , \wRegInBot_6_7[8] , \wRegOut_7_0[2] , 
        \wRegOut_7_5[13] , \wRegInTop_7_14[26] , \wRegEnTop_6_19[0] , 
        \wRegInTop_6_39[27] , \wRegInTop_6_57[2] , \ScanLink125[5] , 
        \wRegInTop_7_61[16] , \wRegInTop_7_37[17] , \wRegInTop_7_76[4] , 
        \wRegInBot_6_39[20] , \wRegInBot_6_59[24] , \wRegInTop_7_42[27] , 
        \wRegOut_7_109[20] , \wRegInTop_6_59[23] , \wRegInTop_7_22[23] , 
        \ScanLink217[28] , \wRegInTop_7_57[13] , \ScanLink217[31] , 
        \ScanLink241[30] , \ScanLink234[19] , \ScanLink245[0] , 
        \wRegOut_4_7[0] , \wRegInTop_7_74[22] , \ScanLink241[29] , 
        \wRegOut_4_4[3] , \wRegEnBot_5_5[0] , \wRegOut_5_14[8] , 
        \wRegInBot_6_3[27] , \wRegOut_5_24[19] , \wRegOut_6_58[5] , 
        \wRegOut_7_79[3] , \wRegOut_6_29[28] , \wRegOut_7_52[28] , 
        \wRegInTop_7_68[8] , \wRegOut_7_5[20] , \wRegOut_7_27[18] , 
        \wRegOut_7_52[31] , \wRegOut_7_71[19] , \wRegInBot_5_3[9] , 
        \wRegInBot_6_19[4] , \wRegOut_6_29[31] , \wRegInTop_5_21[22] , 
        \wRegInTop_6_54[1] , \wRegInTop_7_75[7] , \ScanLink126[6] , 
        \wRegInBot_2_3[29] , \wRegOut_5_2[24] , \wRegInBot_5_17[20] , 
        \ScanLink87[30] , \wRegOut_3_4[5] , \ScanLink18[4] , 
        \wRegInTop_5_17[27] , \ScanLink87[29] , \wRegOut_6_46[9] , 
        \ScanLink246[3] , \wRegInBot_5_21[25] , \wRegOut_7_0[16] , 
        \wRegOut_7_81[8] , \wRegInTop_2_3[26] , \wRegInTop_2_3[15] , 
        \wRegInTop_4_10[4] , \wRegInTop_5_31[2] , \wRegOut_5_4[1] , 
        \wRegOut_5_7[12] , \wRegInTop_5_24[14] , \wRegInTop_7_93[0] , 
        \wRegInBot_5_31[27] , \wRegInTop_5_12[11] , \wRegInBot_5_12[16] , 
        \wRegInTop_5_31[20] , \ScanLink139[31] , \ScanLink112[7] , 
        \wRegInTop_6_60[0] , \wRegInTop_7_41[6] , \wRegOut_3_0[18] , 
        \wRegInBot_4_1[15] , \wRegInBot_5_24[13] , \ScanLink139[28] , 
        \wRegInTop_7_64[20] , \wRegOut_3_7[6] , \wRegInBot_4_0[8] , 
        \wRegOut_4_8[11] , \wRegEnBot_4_10[0] , \wRegInTop_6_29[25] , 
        \wRegInBot_6_29[22] , \wRegInBot_6_33[9] , \wRegInTop_7_11[10] , 
        \wRegInTop_6_49[21] , \wRegInTop_7_47[11] , \ScanLink111[4] , 
        \wRegInBot_6_49[26] , \wRegInTop_6_63[3] , \wRegInTop_7_32[21] , 
        \wRegInTop_7_42[5] , \wRegInTop_7_52[25] , \wRegOut_7_119[22] , 
        \wRegInTop_7_27[15] , \ScanLink194[31] , \ScanLink194[28] , 
        \wRegInTop_7_71[14] , \wRegInTop_4_13[7] , \ScanLink32[9] , 
        \wRegOut_5_20[9] , \wRegInBot_6_6[11] , \wRegInTop_7_90[3] , 
        \wRegOut_5_7[2] , \wRegInTop_5_12[22] , \ScanLink97[18] , 
        \ScanLink216[6] , \wRegOut_5_7[21] , \wRegInBot_5_12[25] , 
        \ScanLink48[1] , \ScanLink87[8] , \wRegInBot_5_18[3] , 
        \wRegInBot_5_24[20] , \wRegInTop_5_31[13] , \wRegOut_7_113[0] , 
        \wRegInTop_5_24[27] , \wRegInBot_5_31[14] , \wRegInTop_7_25[2] , 
        \ScanLink176[3] , \wRegOut_6_0[0] , \wRegOut_6_39[19] , 
        \wRegInBot_6_49[1] , \wRegOut_7_14[18] , \wRegOut_7_61[28] , 
        \wRegOut_7_37[30] , \wRegOut_7_42[19] , \wRegOut_7_61[31] , 
        \wRegOut_7_37[29] , \ScanLink0[18] , \wRegOut_3_1[8] , 
        \wRegInBot_3_2[23] , \wRegInTop_3_7[30] , \wRegInTop_3_7[29] , 
        \wRegInBot_4_1[26] , \ScanLink19[30] , \wRegOut_4_8[22] , 
        \wRegOut_5_17[19] , \wRegOut_6_3[3] , \ScanLink99[4] , 
        \wRegOut_7_0[25] , \wRegInTop_6_3[31] , \wRegInTop_6_3[28] , 
        \wRegOut_7_29[6] , \wRegInBot_6_6[22] , \wRegInTop_7_27[26] , 
        \wRegInTop_7_52[16] , \wRegOut_7_110[3] , \wRegOut_7_119[11] , 
        \ScanLink19[29] , \wRegInTop_6_29[16] , \wRegInBot_6_49[15] , 
        \wRegOut_7_34[9] , \ScanLink215[5] , \wRegInTop_7_11[23] , 
        \wRegInTop_7_71[27] , \ScanLink224[28] , \wRegInTop_4_4[3] , 
        \wRegInBot_4_5[5] , \wRegInBot_6_29[11] , \wRegInTop_6_49[12] , 
        \wRegInTop_7_64[13] , \ScanLink251[18] , \wRegInTop_7_26[1] , 
        \ScanLink175[0] , \ScanLink207[19] , \ScanLink224[31] , 
        \wRegInTop_7_32[12] , \wRegInTop_7_47[22] , \ScanLink111[26] , 
        \wRegOut_7_87[6] , \wRegInTop_7_7[27] , \wRegInTop_5_0[23] , 
        \ScanLink37[4] , \ScanLink164[16] , \wRegInBot_5_19[30] , 
        \wRegOut_5_25[4] , \ScanLink109[6] , \ScanLink132[17] , 
        \ScanLink147[27] , \ScanLink127[23] , \wRegInBot_5_19[29] , 
        \ScanLink104[12] , \ScanLink152[13] , \wRegOut_6_11[24] , 
        \ScanLink89[20] , \ScanLink171[22] , \wRegOut_6_32[15] , 
        \wRegInBot_6_36[4] , \wRegOut_7_55[0] , \wRegOut_6_47[25] , 
        \wRegOut_7_49[15] , \wRegInBot_5_5[30] , \ScanLink114[9] , 
        \wRegInTop_7_88[1] , \wRegInTop_7_47[8] , \wRegInBot_5_5[29] , 
        \wRegOut_6_27[21] , \wRegOut_6_52[11] , \wRegOut_7_29[11] , 
        \ScanLink29[8] , \wRegOut_4_12[25] , \wRegInTop_5_29[0] , 
        \wRegInTop_6_8[24] , \wRegOut_7_56[3] , \wRegInTop_7_111[25] , 
        \wRegInBot_6_35[7] , \wRegOut_7_91[25] , \wRegOut_7_84[11] , 
        \wRegInTop_7_104[11] , \ScanLink31[14] , \ScanLink34[7] , 
        \ScanLink44[24] , \wRegOut_5_26[7] , \wRegInTop_7_127[20] , 
        \wRegInBot_6_37[29] , \wRegEnTop_6_36[0] , \ScanLink219[21] , 
        \ScanLink67[15] , \wRegInBot_6_42[19] , \wRegInBot_6_61[31] , 
        \wRegInBot_6_14[18] , \wRegInBot_6_37[30] , \ScanLink12[25] , 
        \wRegInBot_4_6[6] , \wRegInTop_4_7[0] , \wRegOut_7_84[5] , 
        \wRegInBot_6_61[28] , \ScanLink24[20] , \wRegInTop_4_15[9] , 
        \wRegInBot_6_28[8] , \ScanLink51[10] , \ScanLink72[21] , 
        \wRegInTop_7_59[4] , \wRegOut_7_107[30] , \wRegOut_7_124[18] , 
        \wRegOut_7_107[29] , \wRegOut_6_10[2] , \ScanLink81[6] , 
        \wRegOut_6_27[12] , \wRegOut_6_52[22] , \wRegOut_7_29[22] , 
        \wRegOut_7_31[4] , \ScanLink210[8] , \wRegInTop_1_0[6] , 
        \wRegInTop_5_0[10] , \wRegOut_6_11[17] , \wRegInBot_6_52[0] , 
        \wRegOut_6_32[26] , \wRegOut_6_47[16] , \ScanLink152[20] , 
        \wRegOut_7_49[26] , \wRegInBot_1_1[25] , \wRegInBot_1_1[0] , 
        \ScanLink53[0] , \ScanLink127[10] , \wRegOut_7_108[1] , 
        \wRegInTop_7_122[1] , \wRegInBot_3_2[10] , \ScanLink12[16] , 
        \ScanLink24[13] , \ScanLink50[3] , \ScanLink72[12] , \ScanLink89[13] , 
        \ScanLink171[11] , \ScanLink104[21] , \ScanLink111[15] , 
        \wRegInTop_7_7[14] , \ScanLink164[25] , \wRegInTop_7_81[19] , 
        \wRegInTop_7_0[2] , \ScanLink132[24] , \ScanLink147[14] , 
        \ScanLink31[27] , \ScanLink51[23] , \wRegOut_6_4[19] , 
        \wRegInTop_7_121[2] , \ScanLink44[17] , \wRegInTop_6_22[29] , 
        \wRegInTop_7_59[29] , \wRegInTop_6_57[19] , \wRegInTop_7_3[1] , 
        \ScanLink219[12] , \ScanLink67[26] , \wRegInTop_6_22[30] , 
        \wRegInTop_7_59[30] , \wRegOut_7_32[7] , \wRegOut_7_84[22] , 
        \wRegOut_4_12[16] , \wRegOut_6_13[1] , \wRegInTop_7_104[22] , 
        \ScanLink55[12] , \wRegOut_6_0[31] , \wRegInTop_6_8[17] , 
        \ScanLink82[5] , \wRegInBot_6_51[3] , \wRegInTop_7_127[13] , 
        \wRegInTop_7_111[16] , \ScanLink76[23] , \wRegOut_7_91[16] , 
        \wRegInTop_6_38[0] , \wRegInTop_7_19[6] , \ScanLink208[17] , 
        \wRegOut_6_0[28] , \wRegInBot_1_1[16] , \wRegOut_2_0[26] , 
        \ScanLink4[30] , \wRegInBot_3_6[21] , \ScanLink16[27] , 
        \ScanLink20[22] , \ScanLink35[16] , \ScanLink40[26] , \ScanLink74[5] , 
        \wRegInTop_7_28[28] , \wRegInTop_6_53[28] , \wRegInBot_5_24[7] , 
        \wRegInTop_6_26[18] , \ScanLink63[17] , \wRegInTop_7_105[4] , 
        \wRegInTop_6_53[31] , \wRegInTop_7_28[31] , \wRegOut_5_18[17] , 
        \wRegOut_7_80[13] , \wRegInTop_7_100[13] , \wRegEnTop_5_27[0] , 
        \wRegOut_6_37[7] , \wRegOut_7_8[7] , \ScanLink157[8] , 
        \ScanLink198[1] , \wRegInTop_7_123[22] , \wRegOut_7_16[1] , 
        \wRegOut_6_23[23] , \wRegOut_7_58[23] , \wRegOut_7_95[27] , 
        \wRegInTop_7_115[27] , \wRegOut_6_56[13] , \ScanLink4[29] , 
        \ScanLink10[1] , \wRegInTop_3_3[18] , \wRegInTop_5_4[21] , 
        \wRegOut_6_15[26] , \wRegOut_6_34[4] , \wRegOut_6_36[17] , 
        \wRegOut_6_60[16] , \wRegOut_7_15[2] , \wRegOut_6_43[27] , 
        \wRegInBot_5_27[4] , \ScanLink77[6] , \ScanLink98[16] , 
        \ScanLink100[10] , \ScanLink123[21] , \wRegOut_7_38[27] , 
        \ScanLink149[4] , \ScanLink156[11] , \ScanLink115[24] , 
        \ScanLink175[20] , \wRegInTop_7_85[28] , \ScanLink229[1] , 
        \wRegInTop_7_3[25] , \ScanLink160[14] , \wRegInTop_7_85[31] , 
        \ScanLink136[15] , \ScanLink143[25] , \wRegInTop_7_106[7] , 
        \wRegInBot_3_6[12] , \wRegOut_7_72[5] , \wRegOut_7_80[20] , 
        \wRegOut_7_95[14] , \wRegInTop_7_115[14] , \ScanLink253[9] , 
        \ScanLink16[14] , \ScanLink35[25] , \wRegOut_5_18[24] , 
        \wRegOut_6_53[3] , \wRegInTop_7_100[20] , \wRegInBot_6_11[1] , 
        \wRegInBot_6_46[28] , \wRegInTop_7_123[11] , \ScanLink40[15] , 
        \wRegInBot_6_10[30] , \wRegInBot_6_33[18] , \wRegInTop_5_10[9] , 
        \wRegInBot_6_46[31] , \ScanLink63[24] , \wRegInBot_6_10[29] , 
        \ScanLink76[10] , \wRegOut_7_120[29] , \wRegEnTop_7_33[0] , 
        \ScanLink20[11] , \wRegOut_7_103[18] , \ScanLink13[2] , 
        \ScanLink55[21] , \ScanLink208[24] , \wRegOut_7_120[30] , 
        \ScanLink98[25] , \ScanLink115[17] , \wRegInTop_7_3[16] , 
        \ScanLink160[27] , \ScanLink136[26] , \ScanLink143[16] , 
        \ScanLink156[22] , \wRegInBot_4_13[31] , \wRegInBot_0_0[22] , 
        \wRegOut_2_0[15] , \wRegInBot_4_13[28] , \ScanLink123[12] , 
        \ScanLink175[13] , \wRegInBot_5_1[18] , \wRegInTop_5_4[12] , 
        \wRegOut_6_15[15] , \ScanLink100[23] , \wRegOut_6_60[25] , 
        \wCtrlOut_4[0] , \wRegInTop_5_9[9] , \wRegOut_6_23[10] , 
        \wRegOut_6_36[24] , \wRegInTop_6_42[8] , \wRegOut_6_43[14] , 
        \wRegOut_7_38[14] , \wRegOut_6_56[20] , \wRegOut_7_58[10] , 
        \wRegOut_7_71[6] , \wRegInBot_6_12[2] , \wRegOut_6_50[0] , 
        \ScanLink4[8] , \wRegOut_2_1[7] , \ScanLink5[10] , \wRegOut_3_4[30] , 
        \wRegOut_3_4[29] , \wRegInBot_4_5[17] , \wRegOut_5_13[31] , 
        \wRegOut_5_13[28] , \wRegInTop_6_7[19] , \ScanLink183[0] , 
        \wRegInBot_5_22[9] , \wRegOut_5_30[19] , \wRegInBot_6_2[13] , 
        \ScanLink68[31] , \wRegInTop_6_8[5] , \wRegInTop_6_23[1] , 
        \ScanLink151[6] , \wRegInTop_7_56[27] , \wRegInTop_7_23[17] , 
        \ScanLink68[28] , \wRegInBot_6_9[3] , \wRegInBot_6_38[14] , 
        \wRegInTop_6_58[17] , \wRegInTop_7_75[16] , \wRegOut_6_31[9] , 
        \ScanLink231[3] , \ScanLink255[29] , \wRegInTop_7_60[22] , 
        \ScanLink203[31] , \ScanLink220[19] , \wRegOut_5_3[10] , 
        \wRegInTop_5_16[13] , \wRegInTop_6_38[13] , \wRegInTop_7_15[12] , 
        \wRegInBot_6_58[10] , \wRegInTop_7_43[13] , \wRegOut_7_108[14] , 
        \ScanLink255[30] , \wRegInTop_7_36[23] , \ScanLink203[28] , 
        \wRegInTop_5_20[16] , \wRegInBot_5_20[11] , \wRegInTop_6_20[2] , 
        \ScanLink93[30] , \ScanLink93[29] , \ScanLink152[5] , \ScanLink232[0] , 
        \wRegInBot_5_16[14] , \ScanLink71[8] , \wRegOut_6_48[18] , 
        \wRegOut_7_10[29] , \wRegOut_7_46[31] , \wRegOut_7_65[19] , 
        \wRegOut_7_10[30] , \wRegOut_7_33[18] , \ScanLink180[3] , 
        \wRegOut_7_46[28] , \wRegOut_7_4[14] , \wRegInTop_7_15[21] , 
        \wRegInTop_7_100[9] , \wRegInBot_4_5[24] , \wRegInTop_6_47[5] , 
        \ScanLink135[2] , \wRegInTop_7_60[11] , \wRegInTop_7_36[10] , 
        \wRegInTop_7_66[3] , \wRegOut_5_3[23] , \wRegInTop_5_15[4] , 
        \wRegEnBot_5_15[0] , \wRegInTop_6_38[20] , \wRegInBot_6_58[23] , 
        \wRegInTop_7_43[20] , \wRegOut_7_108[27] , \wRegInTop_5_16[7] , 
        \wRegOut_5_19[0] , \wRegInBot_6_38[27] , \wRegInTop_6_58[24] , 
        \wRegInTop_7_23[24] , \wRegInTop_7_56[14] , \ScanLink190[19] , 
        \wRegInTop_7_75[25] , \ScanLink255[7] , \wRegInBot_6_2[20] , 
        \wRegOut_6_48[2] , \wRegOut_7_69[4] , \ScanLink248[8] , 
        \wRegInTop_6_59[9] , \wRegOut_7_4[27] , \wRegInBot_5_16[27] , 
        \wRegInTop_5_20[25] , \wRegInTop_6_44[6] , \wRegInTop_7_65[0] , 
        \ScanLink136[1] , \wRegInTop_5_5[18] , \wRegInTop_5_16[20] , 
        \wRegOut_7_77[8] , \wRegInBot_5_20[22] , \wRegInTop_7_8[29] , 
        \ScanLink148[30] , \wRegInTop_6_52[2] , \wRegInTop_7_8[30] , 
        \ScanLink148[29] , \wRegInTop_7_73[4] , \ScanLink120[5] , 
        \ScanLink240[0] , \wRegOut_2_2[4] , \wRegInTop_3_4[8] , 
        \wRegOut_4_2[0] , \wRegInBot_5_0[12] , \wRegInTop_7_84[11] , 
        \wRegInTop_4_12[25] , \wRegInBot_4_12[22] , \wRegOut_5_9[16] , 
        \ScanLink157[31] , \ScanLink174[19] , \wRegEnBot_5_0[0] , 
        \ScanLink101[29] , \wRegInTop_7_91[25] , \wRegOut_4_1[3] , 
        \wRegOut_5_11[8] , \ScanLink101[30] , \ScanLink122[18] , 
        \ScanLink157[28] , \wRegOut_6_1[11] , \wRegInBot_6_11[23] , 
        \wRegInTop_6_27[21] , \wRegInBot_6_47[22] , \wRegOut_7_117[26] , 
        \wRegInTop_6_32[15] , \wRegInBot_6_32[12] , \wRegInTop_6_52[11] , 
        \wRegInTop_7_29[11] , \wRegInBot_6_52[16] , \wRegInTop_6_11[24] , 
        \wRegInBot_6_27[26] , \wRegInTop_6_47[25] , \wRegInTop_7_49[15] , 
        \wRegOut_7_102[12] , \wRegOut_7_121[23] , \ScanLink5[23] , 
        \wRegInTop_3_2[12] , \wRegInBot_5_6[9] , \wRegInTop_6_51[1] , 
        \ScanLink123[6] , \wRegInTop_7_70[7] , \wRegInBot_3_7[18] , 
        \wRegInBot_6_8[15] , \wRegOut_6_43[9] , \wRegOut_4_6[15] , 
        \wRegInTop_4_12[16] , \wRegInBot_4_12[11] , \wRegOut_5_9[25] , 
        \wRegInTop_7_91[16] , \ScanLink243[3] , \wRegOut_6_39[1] , 
        \wRegOut_7_6[1] , \ScanLink196[7] , \wRegInTop_7_84[22] , 
        \wRegInBot_5_0[21] , \wRegOut_6_22[30] , \wRegOut_7_18[7] , 
        \wRegOut_7_59[30] , \wRegInBot_2_3[24] , \wRegInTop_3_2[21] , 
        \wRegOut_4_6[26] , \wRegInBot_6_8[26] , \wRegOut_6_22[29] , 
        \ScanLink144[1] , \wRegOut_7_59[29] , \wRegInTop_6_35[5] , 
        \wRegInTop_6_36[6] , \wRegOut_6_57[19] , \wRegInTop_7_17[0] , 
        \ScanLink224[4] , \wRegOut_7_121[2] , \wRegInTop_7_14[3] , 
        \ScanLink147[2] , \wRegOut_7_81[19] , \wRegInTop_7_122[28] , 
        \ScanLink227[7] , \wRegInTop_7_101[19] , \wRegInTop_7_122[31] , 
        \ScanLink21[31] , \ScanLink21[28] , \ScanLink54[18] , 
        \wRegInBot_5_29[2] , \ScanLink79[0] , \ScanLink77[30] , 
        \wRegInTop_6_47[16] , \ScanLink195[4] , \wRegInTop_7_108[1] , 
        \wRegOut_7_122[1] , \wRegInBot_6_27[15] , \wRegInBot_6_2[8] , 
        \wRegInTop_6_32[26] , \wRegOut_6_1[22] , \wRegInBot_6_52[25] , 
        \wRegInTop_7_49[26] , \wRegOut_7_102[21] , \wRegInTop_6_11[17] , 
        \ScanLink77[29] , \wRegOut_5_2[29] , \wRegInTop_5_18[1] , 
        \wRegInBot_6_11[10] , \wRegOut_7_121[10] , \wRegInTop_6_27[12] , 
        \wRegInBot_6_32[21] , \wRegInTop_7_29[22] , \wRegInBot_6_47[11] , 
        \wRegInTop_6_52[22] , \wRegOut_7_5[2] , \wRegOut_7_117[15] , 
        \ScanLink87[24] , \wRegInBot_2_3[17] , \wRegInBot_3_0[3] , 
        \wRegInTop_3_2[6] , \wRegInBot_3_3[0] , \ScanLink18[9] , 
        \wRegOut_5_2[30] , \ScanLink129[27] , \wRegInBot_5_21[28] , 
        \wRegInBot_5_21[31] , \wRegOut_6_46[4] , \ScanLink149[23] , 
        \wRegOut_7_67[2] , \ScanLink92[10] , \wRegInTop_7_9[23] , 
        \wRegOut_7_71[14] , \wRegInTop_5_2[2] , \wRegOut_5_17[6] , 
        \wRegOut_6_29[25] , \wRegInTop_6_49[3] , \wRegOut_7_52[25] , 
        \wRegInTop_7_68[5] , \wRegOut_7_27[15] , \wRegOut_6_49[21] , 
        \wRegOut_7_47[11] , \wRegOut_7_32[21] , \wRegInBot_5_3[4] , 
        \wRegInBot_6_19[9] , \wRegOut_7_64[20] , \wRegOut_5_12[11] , 
        \wRegOut_5_31[20] , \wRegOut_7_11[10] , \ScanLink138[7] , 
        \wRegInTop_3_1[5] , \wRegOut_3_5[23] , \wRegInBot_5_0[7] , 
        \wRegInTop_5_1[1] , \wRegOut_6_58[8] , \wRegOut_5_14[5] , 
        \wRegOut_5_24[14] , \wRegInTop_6_6[20] , \wRegInBot_6_59[29] , 
        \ScanLink125[8] , \ScanLink202[11] , \wRegInTop_7_76[9] , 
        \ScanLink184[27] , \ScanLink221[20] , \wRegInTop_4_1[24] , 
        \ScanLink69[11] , \wRegInBot_6_59[30] , \ScanLink254[10] , 
        \wRegOut_6_45[7] , \ScanLink191[13] , \wRegOut_7_64[1] , 
        \ScanLink234[14] , \ScanLink217[25] , \ScanLink241[24] , 
        \wRegInBot_4_10[6] , \ScanLink61[2] , \wRegInTop_6_6[3] , 
        \wRegInBot_6_7[5] , \wRegOut_6_49[12] , \wRegOut_7_32[12] , 
        \ScanLink190[9] , \wRegOut_7_47[22] , \wRegOut_7_11[23] , 
        \wRegOut_7_27[26] , \wRegOut_7_64[13] , \wRegOut_7_71[27] , 
        \wRegInBot_5_31[0] , \wRegInTop_5_17[19] , \ScanLink92[23] , 
        \wRegOut_6_29[16] , \wRegOut_7_52[16] , \wRegInTop_7_110[3] , 
        \wRegInTop_6_30[8] , \ScanLink149[10] , \wRegInTop_7_9[10] , 
        \wRegOut_6_22[0] , \wRegOut_3_1[21] , \wRegOut_3_5[10] , 
        \wRegInTop_4_1[17] , \ScanLink69[22] , \ScanLink87[17] , 
        \wRegInBot_6_60[2] , \ScanLink129[14] , \ScanLink241[17] , 
        \ScanLink191[20] , \ScanLink234[27] , \wRegOut_6_21[3] , 
        \wRegInTop_6_39[19] , \ScanLink217[16] , \wRegInTop_7_37[29] , 
        \wRegInTop_7_42[19] , \wRegInTop_7_61[31] , \ScanLink202[22] , 
        \wRegInBot_6_63[1] , \ScanLink184[14] , \wRegInTop_7_61[28] , 
        \ScanLink221[9] , \ScanLink254[23] , \ScanLink221[13] , 
        \wRegInTop_7_14[18] , \wRegInTop_7_37[30] , \ScanLink18[23] , 
        \wRegInBot_4_13[5] , \wRegOut_5_24[27] , \wRegInBot_6_4[6] , 
        \wRegInTop_6_5[0] , \wRegInTop_6_6[13] , \ScanLink62[1] , 
        \wRegOut_5_31[13] , \wRegEnTop_7_41[0] , \wRegInBot_6_3[19] , 
        \wRegInTop_7_113[0] , \wRegOut_5_12[22] , \wRegOut_7_24[3] , 
        \ScanLink195[11] , \ScanLink230[16] , \wRegInTop_4_5[26] , 
        \ScanLink94[1] , \wRegInBot_6_47[7] , \ScanLink245[26] , 
        \ScanLink213[27] , \ScanLink78[27] , \wRegInTop_6_48[18] , 
        \ScanLink206[13] , \wRegOut_7_100[9] , \wRegInTop_7_10[30] , 
        \wRegInTop_7_33[18] , \wRegInTop_7_46[28] , \ScanLink180[25] , 
        \ScanLink225[22] , \wRegOut_4_9[31] , \ScanLink46[7] , 
        \wRegInTop_6_2[22] , \wRegInTop_7_10[29] , \wRegInTop_7_46[31] , 
        \ScanLink250[12] , \wRegInTop_7_65[19] , \ScanLink218[0] , 
        \wRegInBot_5_16[5] , \wRegOut_5_20[16] , \wRegEnTop_6_44[0] , 
        \wRegInBot_6_7[28] , \ScanLink178[5] , \wRegOut_4_9[28] , 
        \wRegOut_5_16[13] , \wRegInBot_6_7[31] , \ScanLink45[4] , 
        \wRegOut_6_38[13] , \wRegInBot_5_15[6] , \wRegOut_7_36[23] , 
        \wRegOut_7_43[13] , \wRegOut_7_60[22] , \wRegOut_7_15[12] , 
        \wRegOut_7_23[17] , \wRegInTop_7_28[7] , \wRegOut_7_75[16] , 
        \wRegOut_7_56[27] , \wRegInBot_0_0[18] , \wRegInBot_0_0[11] , 
        \wRegOut_3_1[12] , \ScanLink22[3] , \wRegOut_4_11[5] , 
        \wRegInTop_5_13[31] , \wRegInTop_5_30[19] , \ScanLink97[2] , 
        \wRegOut_6_58[17] , \ScanLink138[11] , \wRegInTop_5_13[28] , 
        \wRegOut_7_27[0] , \wRegOut_5_30[3] , \ScanLink83[26] , 
        \ScanLink96[12] , \wRegInBot_6_44[4] , \ScanLink158[15] , 
        \wRegInTop_7_35[8] , \ScanLink166[9] , \wRegOut_5_16[20] , 
        \wRegOut_7_92[1] , \wRegOut_5_20[25] , \wRegInTop_6_2[11] , 
        \wRegInTop_7_80[9] , \ScanLink78[14] , \wRegInBot_6_23[3] , 
        \wRegInBot_6_28[28] , \ScanLink206[20] , \wRegOut_6_61[1] , 
        \wRegOut_7_40[7] , \ScanLink180[16] , \ScanLink250[21] , 
        \ScanLink225[11] , \wRegInBot_6_28[31] , \ScanLink18[10] , 
        \wRegOut_7_118[31] , \wRegInTop_4_5[15] , \ScanLink195[22] , 
        \ScanLink230[25] , \ScanLink245[15] , \ScanLink21[0] , 
        \wRegOut_5_6[18] , \wRegOut_6_62[2] , \ScanLink213[14] , 
        \wRegOut_7_118[28] , \wRegOut_5_9[4] , \wRegInBot_5_25[19] , 
        \ScanLink83[15] , \wRegOut_7_43[4] , \wRegInBot_6_20[0] , 
        \ScanLink138[22] , \ScanLink158[26] , \ScanLink96[21] , 
        \wRegOut_7_23[24] , \wRegOut_7_75[25] , \wRegOut_7_91[2] , 
        \wRegOut_4_12[6] , \wRegOut_6_58[24] , \ScanLink1[31] , 
        \ScanLink1[28] , \ScanLink1[21] , \ScanLink1[12] , \ScanLink1[5] , 
        \wRegInTop_3_6[10] , \wRegOut_4_2[17] , \wRegInTop_5_21[8] , 
        \wRegOut_6_38[20] , \wRegOut_7_36[10] , \wRegOut_7_56[14] , 
        \wRegOut_7_15[21] , \wRegOut_7_43[20] , \wRegOut_6_8[8] , 
        \wRegOut_7_60[11] , \wRegOut_7_85[31] , \wRegInTop_7_105[31] , 
        \wRegOut_7_106[7] , \wRegInTop_7_126[19] , \ScanLink203[1] , 
        \wRegOut_7_85[28] , \wRegInTop_7_105[28] , \wRegInTop_6_11[3] , 
        \wRegInBot_6_41[9] , \wRegInTop_7_30[5] , \ScanLink163[4] , 
        \wRegEnTop_7_126[0] , \ScanLink25[19] , \ScanLink40[9] , 
        \wRegInTop_6_36[17] , \wRegOut_6_5[13] , \wRegInBot_6_56[14] , 
        \wRegOut_7_106[10] , \ScanLink50[29] , \wRegInTop_6_43[27] , 
        \wRegInTop_6_15[26] , \wRegInBot_6_23[24] , \wRegInTop_7_38[27] , 
        \wRegOut_7_125[21] , \ScanLink2[6] , \wRegInTop_1_1[14] , 
        \ScanLink50[30] , \wRegInTop_6_60[16] , \ScanLink73[18] , 
        \wRegInBot_6_15[21] , \wRegInBot_6_60[11] , \wRegInBot_5_18[10] , 
        \wRegInTop_6_23[23] , \wRegInBot_6_43[20] , \wRegInTop_7_58[23] , 
        \wRegOut_7_113[24] , \ScanLink88[19] , \wRegInBot_6_36[10] , 
        \wRegInTop_6_56[13] , \ScanLink218[18] , \wRegInTop_7_95[27] , 
        \wRegInBot_5_13[8] , \wRegInTop_5_18[17] , \wRegOut_6_53[31] , 
        \wRegOut_7_28[31] , \wRegInTop_7_80[13] , \ScanLink200[2] , 
        \wRegInTop_1_1[27] , \wRegInBot_5_4[10] , \wRegInTop_6_12[0] , 
        \wRegOut_6_26[18] , \wRegOut_6_53[28] , \wRegOut_7_28[28] , 
        \wRegOut_7_105[4] , \wRegInTop_7_33[6] , \ScanLink160[7] , 
        \wRegInBot_3_3[30] , \wRegInTop_3_6[23] , \wRegInTop_5_24[5] , 
        \wRegOut_6_5[20] , \wRegInBot_6_15[12] , \wRegInTop_6_23[10] , 
        \wRegInBot_6_36[23] , \wRegInBot_6_38[2] , \wRegInBot_6_60[22] , 
        \wRegInBot_6_43[13] , \wRegInTop_6_56[20] , \wRegInTop_7_58[10] , 
        \wRegOut_7_113[17] , \wRegInBot_6_23[17] , \wRegInTop_6_43[14] , 
        \wRegInTop_6_36[24] , \wRegInTop_7_38[14] , \wRegInTop_7_86[7] , 
        \wRegOut_7_106[23] , \wRegInBot_6_56[27] , \wRegInTop_6_60[25] , 
        \wRegInTop_6_15[15] , \wRegOut_7_46[9] , \wRegOut_7_125[12] , 
        \wRegOut_7_89[0] , \ScanLink39[2] , \ScanLink107[0] , 
        \wRegInTop_7_54[1] , \wRegInBot_3_3[29] , \wRegOut_4_2[24] , 
        \wRegInBot_4_8[0] , \wRegInTop_5_1[29] , \wRegOut_5_28[1] , 
        \wRegEnTop_7_19[0] , \wRegInTop_4_9[6] , \wRegInTop_5_1[30] , 
        \wRegInBot_5_4[23] , \wRegOut_1_0[2] , \wRegOut_4_14[8] , 
        \ScanLink104[3] , \wRegInTop_7_57[2] , \wRegInTop_5_18[24] , 
        \wRegOut_7_58[5] , \wRegInTop_7_80[20] , \wRegInBot_5_18[23] , 
        \wRegInTop_5_27[6] , \ScanLink105[18] , \ScanLink126[30] , 
        \wRegInBot_5_31[9] , \ScanLink126[29] , \ScanLink170[28] , 
        \wRegInTop_7_95[14] , \wRegOut_7_0[6] , \ScanLink153[19] , 
        \wRegInTop_7_85[4] , \ScanLink170[31] , \wRegOut_7_5[17] , 
        \wRegEnTop_6_3[0] , \ScanLink190[0] , \wRegInBot_1_0[26] , 
        \wRegOut_2_1[25] , \wRegInBot_3_3[9] , \wRegOut_3_5[19] , 
        \wRegInBot_4_4[14] , \wRegOut_5_2[13] , \wRegOut_6_22[9] , 
        \ScanLink222[3] , \wRegInTop_5_17[10] , \wRegInBot_5_17[17] , 
        \wRegInTop_5_21[15] , \wRegInBot_5_21[12] , \wRegInTop_6_30[1] , 
        \ScanLink142[6] , \wRegOut_7_127[5] , \wRegInTop_7_11[7] , 
        \ScanLink149[19] , \wRegInTop_6_39[10] , \wRegInTop_7_9[19] , 
        \wRegInBot_6_59[13] , \wRegInTop_7_42[10] , \wRegOut_7_109[17] , 
        \wRegInTop_7_14[11] , \wRegInTop_7_37[20] , \wRegInTop_7_61[21] , 
        \ScanLink221[0] , \wRegOut_7_124[6] , \ScanLink18[0] , \ScanLink62[8] , 
        \wRegInTop_6_33[2] , \wRegInBot_6_63[8] , \ScanLink191[29] , 
        \wRegInTop_7_74[15] , \wRegInBot_6_39[17] , \wRegInTop_7_12[4] , 
        \ScanLink141[5] , \wRegInTop_7_57[24] , \wRegInTop_7_22[14] , 
        \wRegInTop_6_59[14] , \ScanLink191[30] , \wRegInBot_6_3[10] , 
        \wRegOut_7_3[5] , \wRegInTop_7_113[9] , \wRegInTop_6_5[9] , 
        \ScanLink193[3] , \wRegOut_4_4[7] , \wRegOut_5_2[20] , 
        \wRegInTop_5_17[23] , \wRegInBot_5_21[21] , \ScanLink246[7] , 
        \wRegInBot_5_17[24] , \wRegInTop_5_18[8] , \ScanLink92[19] , 
        \wRegInTop_5_21[26] , \wRegInTop_6_54[5] , \wRegInTop_7_75[3] , 
        \ScanLink126[2] , \wRegInBot_6_19[0] , \wRegOut_6_49[31] , 
        \wRegOut_6_49[28] , \wRegOut_7_47[18] , \wRegOut_7_64[30] , 
        \wRegOut_7_32[28] , \wRegOut_7_64[29] , \wRegOut_7_11[19] , 
        \wRegOut_7_32[31] , \wRegEnBot_3_5[0] , \wRegInTop_5_1[8] , 
        \wRegOut_6_58[1] , \wRegOut_7_5[24] , \wRegOut_7_79[7] , 
        \wRegOut_5_31[29] , \wRegInTop_6_6[30] , \wRegInTop_6_6[29] , 
        \wRegInBot_6_3[23] , \wRegInBot_4_4[27] , \wRegOut_4_7[4] , 
        \wRegOut_5_12[18] , \wRegOut_5_31[30] , \ScanLink69[18] , 
        \wRegInTop_6_39[23] , \wRegInBot_6_39[24] , \wRegOut_7_64[8] , 
        \wRegInTop_7_74[26] , \ScanLink245[4] , \wRegInTop_6_57[6] , 
        \wRegInTop_6_59[27] , \wRegInTop_7_22[27] , \ScanLink125[1] , 
        \wRegInTop_7_57[17] , \ScanLink221[30] , \wRegInTop_7_37[13] , 
        \ScanLink202[18] , \wRegInTop_7_76[0] , \wRegInBot_6_59[20] , 
        \wRegInTop_7_42[23] , \wRegOut_7_109[24] , \ScanLink221[29] , 
        \wRegInBot_4_12[18] , \ScanLink67[5] , \wRegInTop_7_14[22] , 
        \wRegInTop_7_61[12] , \ScanLink254[19] , \ScanLink99[15] , 
        \wRegOut_6_39[8] , \ScanLink114[27] , \wRegOut_7_6[8] , 
        \ScanLink137[16] , \ScanLink142[26] , \wRegInTop_7_116[4] , 
        \ScanLink239[2] , \ScanLink101[13] , \wRegInTop_7_2[26] , 
        \ScanLink161[17] , \ScanLink174[23] , \wRegInTop_5_5[22] , 
        \wRegInTop_6_0[4] , \ScanLink122[22] , \ScanLink159[7] , 
        \wRegInBot_6_1[2] , \ScanLink157[12] , \wRegOut_6_37[14] , 
        \wRegOut_6_14[25] , \wRegOut_6_42[24] , \wRegOut_7_39[24] , 
        \wRegOut_6_24[7] , \wRegOut_6_61[15] , \wRegInTop_3_2[31] , 
        \wRegInBot_5_0[31] , \wRegInBot_5_0[28] , \ScanLink144[8] , 
        \wRegOut_7_59[20] , \wRegOut_6_22[20] , \wRegInTop_7_17[9] , 
        \wRegOut_6_27[4] , \wRegOut_6_57[10] , \wRegInTop_3_2[28] , 
        \wRegOut_7_94[24] , \wRegInTop_7_114[24] , \wRegInBot_3_7[22] , 
        \wRegOut_5_19[14] , \ScanLink79[9] , \ScanLink188[2] , 
        \wRegInTop_7_108[8] , \wRegOut_7_122[8] , \wRegInTop_7_122[21] , 
        \wRegOut_7_81[10] , \wRegInTop_7_101[10] , \ScanLink17[24] , 
        \ScanLink62[14] , \wRegInBot_6_32[31] , \wRegInBot_6_11[19] , 
        \wRegInBot_4_15[2] , \ScanLink34[15] , \ScanLink41[25] , 
        \wRegInBot_6_32[28] , \ScanLink64[6] , \wRegInBot_6_47[18] , 
        \wRegInTop_7_115[7] , \ScanLink54[11] , \wRegInTop_6_28[3] , 
        \ScanLink209[14] , \wRegInBot_6_2[1] , \wRegInTop_6_3[7] , 
        \wRegInBot_1_0[15] , \wRegOut_2_1[16] , \ScanLink5[19] , 
        \ScanLink21[21] , \ScanLink77[20] , \wRegOut_7_102[28] , 
        \wRegOut_6_40[3] , \wRegOut_7_61[5] , \wRegOut_7_102[31] , 
        \wRegOut_7_121[19] , \ScanLink240[9] , \wRegInTop_3_4[1] , 
        \wRegInBot_3_5[7] , \wRegInTop_5_4[5] , \wRegInTop_5_5[11] , 
        \wRegOut_6_22[13] , \wRegOut_6_57[23] , \wRegOut_7_59[13] , 
        \wRegOut_6_42[17] , \wRegOut_6_14[16] , \wRegOut_6_37[27] , 
        \wRegOut_7_39[17] , \wRegOut_6_61[26] , \wRegInBot_5_5[3] , 
        \ScanLink101[20] , \ScanLink174[10] , \wRegOut_5_11[1] , 
        \ScanLink157[21] , \ScanLink122[11] , \wRegEnTop_7_20[0] , 
        \ScanLink137[25] , \ScanLink142[15] , \wRegOut_4_2[9] , 
        \ScanLink99[26] , \wRegInTop_7_2[15] , \ScanLink161[24] , 
        \wRegInTop_7_84[18] , \ScanLink21[12] , \ScanLink114[14] , 
        \wRegInBot_3_3[20] , \ScanLink13[26] , \wRegInBot_3_6[4] , 
        \ScanLink17[17] , \wRegInBot_5_6[0] , \wRegInTop_5_7[6] , 
        \wRegOut_5_12[2] , \wRegOut_6_1[18] , \ScanLink54[22] , 
        \ScanLink209[27] , \ScanLink77[13] , \wRegInTop_3_7[2] , 
        \wRegInTop_6_27[31] , \wRegInBot_3_7[11] , \ScanLink34[26] , 
        \ScanLink62[27] , \ScanLink41[16] , \wRegInTop_6_27[28] , 
        \wRegInTop_6_52[18] , \wRegInTop_7_29[18] , \wRegOut_7_81[23] , 
        \wRegInTop_7_122[12] , \ScanLink25[23] , \ScanLink50[13] , 
        \wRegOut_5_19[27] , \wRegOut_6_43[0] , \wRegOut_7_62[6] , 
        \wRegInTop_7_101[23] , \wRegInTop_6_51[8] , \wRegOut_7_94[17] , 
        \wRegInTop_7_114[17] , \wRegInTop_7_49[7] , \wRegOut_6_5[29] , 
        \ScanLink66[16] , \wRegOut_6_5[30] , \ScanLink73[22] , 
        \wRegInTop_6_56[30] , \wRegOut_7_94[6] , \ScanLink24[4] , 
        \ScanLink45[27] , \wRegInTop_6_56[29] , \ScanLink218[22] , 
        \wRegOut_4_13[26] , \ScanLink30[17] , \wRegInTop_6_23[19] , 
        \wRegInTop_7_58[19] , \ScanLink107[9] , \wRegInTop_7_54[8] , 
        \wRegOut_7_85[12] , \wRegInTop_7_126[23] , \wRegInTop_7_105[12] , 
        \wRegInTop_6_9[27] , \wRegOut_7_46[0] , \wRegOut_7_89[9] , 
        \wRegInTop_7_110[26] , \wRegInBot_6_25[4] , \wRegOut_7_90[26] , 
        \wRegOut_6_26[22] , \wRegInTop_7_98[2] , \wRegOut_6_53[12] , 
        \wRegOut_7_28[12] , \wRegInTop_2_2[16] , \wRegInBot_3_3[13] , 
        \wRegInTop_3_6[19] , \wRegInBot_4_8[9] , \wRegInTop_5_1[20] , 
        \wRegOut_5_28[8] , \wRegOut_6_33[16] , \wRegOut_7_48[16] , 
        \wRegOut_6_10[27] , \wRegOut_6_46[26] , \ScanLink27[7] , 
        \ScanLink88[23] , \wRegInBot_6_26[7] , \wRegOut_7_45[3] , 
        \ScanLink105[11] , \ScanLink170[21] , \wRegEnTop_6_25[0] , 
        \ScanLink119[5] , \ScanLink126[20] , \ScanLink153[10] , 
        \wRegOut_4_14[1] , \ScanLink133[14] , \wRegInTop_7_80[30] , 
        \wRegInTop_6_9[14] , \ScanLink110[25] , \ScanLink146[24] , 
        \wRegInTop_7_80[29] , \wRegOut_7_97[5] , \wRegInTop_7_6[24] , 
        \ScanLink165[15] , \wRegInTop_7_110[15] , \wRegOut_7_90[15] , 
        \wRegOut_6_8[1] , \ScanLink92[6] , \wRegInTop_7_126[10] , 
        \wRegOut_7_85[21] , \ScanLink13[15] , \wRegOut_4_13[15] , 
        \wRegOut_7_22[4] , \ScanLink203[8] , \wRegInTop_7_105[21] , 
        \wRegInBot_6_41[0] , \wRegInBot_6_43[30] , \wRegInBot_4_0[16] , 
        \ScanLink18[19] , \wRegOut_4_9[12] , \ScanLink25[10] , 
        \ScanLink30[24] , \ScanLink66[25] , \wRegInBot_6_15[28] , 
        \wRegInBot_6_60[18] , \wRegInBot_6_43[29] , \ScanLink40[0] , 
        \ScanLink45[14] , \wRegInBot_6_15[31] , \wRegInBot_6_36[19] , 
        \ScanLink218[11] , \wRegOut_7_106[19] , \wRegInTop_5_1[13] , 
        \wRegInBot_5_10[2] , \wRegOut_7_125[31] , \ScanLink43[3] , 
        \wRegInBot_5_18[19] , \ScanLink50[20] , \ScanLink73[11] , 
        \wRegOut_7_125[28] , \ScanLink88[10] , \ScanLink110[16] , 
        \ScanLink133[27] , \ScanLink146[17] , \wRegInTop_7_6[17] , 
        \ScanLink165[26] , \ScanLink170[12] , \ScanLink105[22] , 
        \ScanLink153[23] , \wRegInBot_5_13[1] , \ScanLink126[13] , 
        \wRegOut_7_118[2] , \wRegInTop_6_12[9] , \wRegOut_6_46[15] , 
        \wRegInBot_5_4[19] , \wRegOut_6_10[14] , \wRegOut_6_33[25] , 
        \wRegOut_7_48[25] , \wRegOut_7_21[7] , \wRegOut_5_16[30] , 
        \wRegInTop_5_22[2] , \wRegInTop_6_2[18] , \wRegOut_6_26[11] , 
        \ScanLink91[5] , \wRegInBot_6_42[3] , \wRegOut_6_53[21] , 
        \wRegOut_7_28[21] , \wRegInTop_7_80[0] , \wRegInBot_6_7[12] , 
        \wRegOut_7_92[8] , \wRegOut_5_16[29] , \wRegInTop_6_28[26] , 
        \ScanLink101[7] , \wRegInBot_6_48[25] , \wRegInTop_7_70[17] , 
        \wRegInTop_7_52[6] , \wRegInTop_7_53[26] , \wRegOut_7_118[21] , 
        \wRegInBot_6_28[21] , \wRegInTop_6_48[22] , \wRegInTop_7_26[16] , 
        \wRegInTop_7_46[12] , \ScanLink250[31] , \ScanLink206[29] , 
        \wRegOut_6_61[8] , \wRegInTop_7_33[22] , \ScanLink250[28] , 
        \wRegInTop_7_10[13] , \wRegInTop_7_65[23] , \ScanLink206[30] , 
        \ScanLink225[18] , \wRegInTop_5_30[23] , \ScanLink96[31] , 
        \ScanLink102[4] , \wRegInTop_7_51[5] , \ScanLink21[9] , 
        \wRegOut_5_6[11] , \wRegInTop_5_13[12] , \wRegInBot_5_25[10] , 
        \ScanLink96[28] , \wRegInBot_5_13[15] , \wRegInTop_5_21[1] , 
        \wRegInTop_5_25[17] , \wRegInBot_6_20[9] , \wRegInBot_5_30[24] , 
        \wRegOut_6_38[29] , \wRegOut_7_15[31] , \wRegOut_7_36[19] , 
        \wRegInTop_7_83[3] , \wRegOut_7_43[29] , \wRegOut_6_38[30] , 
        \wRegOut_7_15[28] , \wRegOut_7_43[30] , \wRegOut_7_60[18] , 
        \ScanLink7[2] , \wRegOut_3_1[31] , \wRegInTop_6_48[11] , 
        \wRegOut_7_1[15] , \wRegInTop_7_33[11] , \wRegInTop_7_36[2] , 
        \ScanLink165[3] , \wRegOut_3_1[28] , \wRegInTop_6_17[4] , 
        \wRegInBot_6_28[12] , \wRegInTop_7_8[3] , \wRegInTop_7_46[21] , 
        \wRegInBot_4_0[25] , \wRegOut_4_9[21] , \wRegInBot_6_7[21] , 
        \wRegInTop_6_28[15] , \ScanLink94[8] , \wRegInTop_7_10[20] , 
        \wRegInTop_7_26[25] , \wRegInTop_7_65[10] , \ScanLink195[18] , 
        \ScanLink205[6] , \wRegInTop_7_70[24] , \wRegEnTop_7_78[0] , 
        \wRegInBot_6_48[16] , \wRegInTop_7_53[15] , \wRegOut_7_100[0] , 
        \wRegOut_7_118[12] , \wRegOut_6_18[3] , \wRegOut_7_39[5] , 
        \ScanLink218[9] , \wRegEnBot_6_17[0] , \ScanLink89[7] , 
        \wRegOut_7_1[26] , \ScanLink0[11] , \ScanLink4[1] , 
        \wRegInTop_2_2[25] , \wRegOut_5_6[22] , \wRegInBot_5_13[26] , 
        \wRegInBot_6_59[2] , \wRegInTop_5_25[24] , \wRegInBot_5_30[17] , 
        \wRegInTop_6_14[7] , \wRegInTop_7_35[1] , \ScanLink166[0] , 
        \wRegInTop_5_0[19] , \wRegInTop_5_13[21] , \wRegInBot_5_25[23] , 
        \ScanLink58[2] , \wRegInTop_5_30[10] , \ScanLink138[18] , 
        \wRegOut_7_27[9] , \wRegOut_7_103[3] , \ScanLink206[5] , 
        \wRegInTop_7_23[5] , \ScanLink170[4] , \ScanLink210[1] , 
        \wRegOut_7_115[7] , \wRegInTop_1_0[17] , \wRegInBot_1_1[9] , 
        \wRegInBot_5_5[13] , \wRegInBot_6_52[9] , \wRegInTop_5_19[14] , 
        \ScanLink53[9] , \ScanLink152[29] , \wRegInTop_7_81[10] , 
        \ScanLink104[31] , \ScanLink127[19] , \wRegInBot_5_19[13] , 
        \wRegOut_6_6[7] , \ScanLink152[30] , \ScanLink171[18] , 
        \wRegOut_7_108[8] , \wRegInTop_7_122[8] , \wRegInTop_6_22[20] , 
        \ScanLink104[28] , \wRegInBot_6_42[23] , \wRegInTop_7_59[20] , 
        \wRegInTop_7_94[24] , \wRegOut_7_112[27] , \wRegInBot_6_37[13] , 
        \wRegInTop_6_57[10] , \wRegInTop_7_3[8] , \wRegInBot_6_61[12] , 
        \wRegInTop_3_7[13] , \wRegOut_6_4[10] , \wRegInTop_6_14[25] , 
        \wRegInBot_6_14[22] , \wRegInTop_6_37[14] , \wRegInTop_6_61[15] , 
        \wRegOut_7_124[22] , \wRegOut_6_5[4] , \wRegInBot_6_57[17] , 
        \wRegOut_7_107[13] , \wRegInBot_6_22[27] , \wRegInTop_6_42[24] , 
        \wRegInTop_7_39[24] , \wRegInTop_7_20[6] , \ScanLink173[7] , 
        \ScanLink0[22] , \wRegOut_3_2[2] , \wRegInBot_3_2[19] , 
        \wRegOut_6_13[8] , \ScanLink213[2] , \wRegOut_4_3[14] , 
        \wRegOut_5_2[6] , \wRegInBot_5_19[20] , \ScanLink89[30] , 
        \wRegInTop_7_95[7] , \wRegOut_7_116[4] , \ScanLink89[29] , 
        \wRegInTop_7_94[17] , \wRegInTop_7_81[23] , \wRegEnTop_4_1[0] , 
        \wRegOut_7_48[6] , \wRegInBot_5_5[20] , \wRegInTop_5_19[27] , 
        \wRegOut_6_27[31] , \wRegOut_6_27[28] , \ScanLink114[0] , 
        \wRegInTop_7_88[8] , \wRegOut_6_52[18] , \wRegOut_7_29[18] , 
        \wRegInTop_7_47[1] , \wRegInTop_3_7[20] , \wRegOut_4_3[27] , 
        \wRegInTop_5_29[9] , \wRegOut_7_55[9] , \wRegOut_7_84[18] , 
        \wRegInTop_7_127[30] , \ScanLink117[3] , \wRegInTop_7_44[2] , 
        \wRegInTop_7_104[18] , \wRegInTop_7_127[29] , \ScanLink29[1] , 
        \wRegOut_7_99[3] , \wRegInTop_1_0[24] , \ScanLink24[30] , 
        \wRegInTop_4_15[0] , \wRegInTop_6_61[26] , \wRegOut_5_1[5] , 
        \ScanLink72[28] , \wRegInTop_6_14[16] , \ScanLink24[29] , 
        \ScanLink51[19] , \ScanLink72[31] , \wRegInBot_6_22[14] , 
        \wRegInTop_6_42[17] , \wRegOut_7_124[11] , \wRegInTop_6_37[27] , 
        \wRegInTop_7_39[17] , \wRegInTop_7_96[4] , \wRegOut_7_107[20] , 
        \wRegOut_6_4[23] , \wRegInBot_6_14[11] , \wRegInTop_6_22[13] , 
        \wRegInBot_6_37[20] , \wRegInBot_6_57[24] , \wRegInBot_6_42[10] , 
        \wRegInTop_6_57[23] , \ScanLink219[28] , \wRegInTop_7_59[13] , 
        \wRegOut_7_112[14] , \wRegInBot_1_0[4] , \ScanLink2[24] , 
        \wRegInBot_2_0[5] , \wRegInTop_2_1[3] , \wRegInTop_2_2[0] , 
        \wRegOut_3_0[22] , \wRegOut_3_1[1] , \ScanLink219[31] , \ScanLink9[4] , 
        \wRegInTop_4_7[9] , \wRegInBot_6_61[21] , \wRegOut_5_7[31] , 
        \wRegInBot_6_28[1] , \ScanLink159[16] , \wRegOut_5_7[28] , 
        \ScanLink82[25] , \wRegInBot_5_24[30] , \wRegOut_6_16[5] , 
        \wRegOut_7_37[3] , \ScanLink97[11] , \ScanLink48[8] , 
        \wRegInBot_5_24[29] , \ScanLink87[1] , \wRegInBot_6_54[7] , 
        \ScanLink139[12] , \wRegOut_5_17[10] , \ScanLink55[7] , 
        \wRegInTop_6_19[2] , \wRegInTop_7_38[4] , \wRegOut_7_113[9] , 
        \wRegOut_7_57[24] , \wRegOut_6_39[10] , \wRegInBot_6_49[8] , 
        \wRegOut_6_59[14] , \wRegOut_7_22[14] , \wRegInTop_7_6[5] , 
        \wRegOut_7_61[21] , \wRegOut_7_74[15] , \wRegOut_7_14[11] , 
        \wRegOut_6_0[9] , \wRegEnTop_6_57[0] , \wRegOut_7_37[20] , 
        \wRegOut_7_42[10] , \wRegInTop_7_124[6] , \wRegOut_5_21[15] , 
        \ScanLink56[4] , \wRegInTop_7_5[6] , \ScanLink168[6] , 
        \wRegInTop_6_3[21] , \ScanLink208[3] , \wRegInTop_7_127[5] , 
        \ScanLink79[24] , \ScanLink181[26] , \ScanLink224[21] , 
        \ScanLink19[20] , \wRegInTop_4_4[25] , \ScanLink84[2] , 
        \wRegInBot_6_29[18] , \ScanLink175[9] , \ScanLink251[11] , 
        \ScanLink207[10] , \wRegInTop_7_26[8] , \ScanLink212[24] , 
        \wRegOut_6_15[6] , \wRegOut_7_34[0] , \ScanLink194[12] , 
        \wRegOut_7_119[18] , \ScanLink231[15] , \wRegInBot_6_57[4] , 
        \ScanLink244[25] , \wRegInBot_2_3[6] , \wRegOut_5_4[8] , 
        \wRegOut_7_14[22] , \wRegOut_3_0[11] , \wRegInTop_4_2[4] , 
        \wRegInBot_4_3[2] , \ScanLink31[3] , \wRegOut_6_39[23] , 
        \wRegOut_7_37[13] , \wRegOut_7_61[12] , \wRegInTop_7_93[9] , 
        \wRegOut_7_22[27] , \wRegOut_7_42[23] , \wRegOut_5_23[3] , 
        \wRegOut_6_59[27] , \wRegOut_7_57[17] , \wRegOut_7_74[26] , 
        \wRegOut_7_81[1] , \ScanLink19[13] , \wRegInTop_4_4[16] , 
        \wRegInTop_5_12[18] , \wRegInTop_5_31[30] , \ScanLink97[22] , 
        \wRegInTop_5_31[29] , \ScanLink82[16] , \wRegInTop_6_60[9] , 
        \ScanLink139[21] , \ScanLink159[25] , \wRegOut_7_53[7] , 
        \wRegInBot_6_30[3] , \ScanLink212[17] , \ScanLink79[17] , 
        \wRegInBot_6_33[0] , \wRegInTop_6_49[31] , \wRegOut_7_50[4] , 
        \ScanLink194[21] , \ScanLink244[16] , \ScanLink231[26] , 
        \ScanLink181[15] , \wRegInTop_7_64[29] , \ScanLink251[22] , 
        \ScanLink224[12] , \wRegInTop_7_32[31] , \wRegOut_5_21[26] , 
        \wRegInTop_6_49[28] , \wRegInTop_7_11[19] , \wRegInTop_7_47[18] , 
        \wRegInTop_7_64[30] , \wRegInTop_7_32[28] , \ScanLink207[23] , 
        \wRegInTop_6_3[12] , \ScanLink4[20] , \ScanLink4[13] , 
        \wRegInBot_2_2[27] , \wRegOut_3_4[20] , \wRegInTop_4_0[27] , 
        \wRegInBot_4_0[1] , \wRegInTop_4_1[7] , \wRegOut_4_8[18] , 
        \wRegOut_7_82[2] , \ScanLink32[0] , \wRegOut_5_17[23] , 
        \wRegOut_5_20[0] , \wRegOut_5_19[9] , \wRegInBot_6_6[18] , 
        \ScanLink216[26] , \ScanLink68[12] , \wRegInBot_6_17[6] , 
        \wRegOut_6_55[4] , \ScanLink190[10] , \wRegOut_7_74[2] , 
        \ScanLink235[17] , \wRegInTop_7_15[28] , \ScanLink185[24] , 
        \ScanLink220[23] , \ScanLink240[27] , \ScanLink15[5] , \ScanLink16[6] , 
        \wRegInTop_6_38[30] , \ScanLink255[13] , \wRegInTop_6_38[29] , 
        \wRegInTop_7_15[31] , \wRegInTop_7_43[30] , \wRegInTop_7_60[18] , 
        \ScanLink203[12] , \wRegInTop_7_36[19] , \wRegInTop_7_43[29] , 
        \wRegOut_5_13[12] , \wRegOut_5_25[17] , \wRegInTop_6_7[23] , 
        \ScanLink248[1] , \wRegOut_5_30[23] , \wRegInBot_6_2[30] , 
        \wRegInBot_6_2[29] , \ScanLink128[4] , \wRegOut_7_10[13] , 
        \wRegOut_7_65[23] , \wRegOut_4_9[2] , \wRegInTop_5_16[30] , 
        \wRegInTop_5_16[29] , \wRegOut_6_28[26] , \wRegOut_6_48[22] , 
        \wRegOut_7_46[12] , \wRegInTop_6_59[0] , \wRegOut_7_33[22] , 
        \wRegOut_7_53[26] , \wRegInTop_7_78[6] , \ScanLink93[13] , 
        \wRegOut_6_56[7] , \wRegOut_7_26[16] , \wRegOut_7_70[17] , 
        \wRegOut_7_77[1] , \wRegInTop_7_8[20] , \wRegInBot_6_14[5] , 
        \ScanLink128[24] , \ScanLink148[20] , \ScanLink136[8] , 
        \wRegInTop_7_65[9] , \ScanLink86[27] , \wRegInBot_2_2[14] , 
        \wRegOut_3_4[13] , \wRegOut_5_13[21] , \wRegInBot_5_22[0] , 
        \wRegOut_5_30[10] , \ScanLink72[2] , \wRegOut_5_25[24] , 
        \ScanLink183[9] , \wRegInTop_7_103[3] , \wRegInTop_6_7[10] , 
        \wRegOut_6_31[0] , \wRegOut_7_10[6] , \ScanLink255[20] , 
        \ScanLink185[17] , \ScanLink220[10] , \wRegInTop_4_0[14] , 
        \wRegInBot_6_58[19] , \ScanLink203[21] , \ScanLink68[21] , 
        \wRegInTop_6_23[8] , \ScanLink216[15] , \ScanLink240[14] , 
        \ScanLink128[17] , \ScanLink190[23] , \ScanLink235[24] , 
        \ScanLink10[8] , \wRegInTop_3_3[11] , \wRegOut_4_7[16] , 
        \wRegOut_5_3[19] , \wRegInBot_5_20[18] , \ScanLink86[14] , 
        \wRegOut_6_32[3] , \ScanLink232[9] , \ScanLink93[20] , 
        \wRegInTop_7_8[13] , \wRegOut_7_13[5] , \ScanLink148[13] , 
        \wRegInBot_5_21[3] , \ScanLink71[1] , \wRegOut_7_26[25] , 
        \wRegEnTop_7_52[0] , \wRegOut_6_28[15] , \wRegOut_7_53[15] , 
        \wRegInTop_7_100[0] , \wRegOut_6_48[11] , \wRegOut_7_10[20] , 
        \wRegOut_7_70[24] , \wRegOut_7_65[10] , \wRegOut_7_33[11] , 
        \wRegOut_7_46[21] , \wRegOut_7_80[29] , \wRegInTop_7_100[29] , 
        \wRegInBot_6_9[16] , \wRegInBot_6_11[8] , \ScanLink253[0] , 
        \wRegOut_7_80[30] , \wRegInTop_7_100[30] , \wRegInTop_7_123[18] , 
        \wRegInTop_6_41[2] , \ScanLink133[5] , \wRegInTop_7_60[4] , 
        \ScanLink55[31] , \wRegInTop_6_10[27] , \wRegOut_7_120[20] , 
        \ScanLink76[19] , \ScanLink20[18] , \wRegOut_6_0[12] , 
        \wRegInTop_6_33[16] , \wRegInBot_6_53[15] , \wRegInTop_4_13[26] , 
        \wRegInBot_4_13[21] , \wRegOut_5_8[15] , \wRegInTop_5_10[0] , 
        \ScanLink55[28] , \wRegInTop_6_46[26] , \wRegInTop_7_48[16] , 
        \wRegOut_7_103[11] , \wRegInTop_6_26[22] , \wRegInBot_6_26[25] , 
        \wRegInBot_6_46[21] , \wRegOut_7_116[25] , \wRegInBot_6_33[11] , 
        \wRegInTop_6_53[12] , \wRegInTop_7_28[12] , \wRegInBot_6_10[20] , 
        \wRegInTop_5_13[3] , \wRegInTop_7_90[26] , \wRegInTop_7_85[12] , 
        \wRegInTop_5_9[0] , \wRegOut_6_23[19] , \wRegOut_6_56[29] , 
        \wRegOut_7_58[19] , \wRegOut_6_50[9] , \wRegOut_6_56[30] , 
        \ScanLink250[3] , \wRegInTop_3_3[22] , \wRegInBot_5_1[11] , 
        \wRegInBot_5_8[6] , \wRegOut_6_0[21] , \wRegInTop_6_10[14] , 
        \wRegInBot_6_10[13] , \wRegInTop_6_26[11] , \wRegInBot_6_33[22] , 
        \wRegInTop_6_42[1] , \wRegInTop_7_63[7] , \ScanLink130[6] , 
        \wRegInTop_7_28[21] , \wRegInBot_6_46[12] , \wRegInTop_6_53[21] , 
        \wRegOut_7_116[16] , \wRegInBot_6_26[16] , \wRegInTop_6_38[9] , 
        \wRegInTop_6_46[15] , \ScanLink185[7] , \wRegOut_7_120[13] , 
        \wRegInTop_6_33[25] , \wRegInBot_6_53[26] , \wRegInTop_7_48[25] , 
        \wRegOut_7_103[22] , \wRegInBot_3_6[31] , \wRegInBot_3_6[28] , 
        \wRegOut_4_7[25] , \ScanLink69[3] , \wRegOut_7_16[8] , 
        \ScanLink237[4] , \wRegInTop_7_118[2] , \wRegInBot_6_9[25] , 
        \wRegInTop_6_25[6] , \ScanLink157[1] , \ScanLink198[8] , 
        \wRegInBot_5_1[22] , \wRegInTop_5_4[31] , \ScanLink234[7] , 
        \wRegInTop_5_4[28] , \wRegInTop_6_26[5] , \ScanLink154[2] , 
        \wRegInTop_4_13[15] , \wRegOut_6_29[2] , \wRegInTop_7_85[21] , 
        \wRegInBot_4_13[12] , \wRegOut_5_8[26] , \ScanLink100[19] , 
        \ScanLink123[28] , \ScanLink229[8] , \ScanLink156[18] , 
        \ScanLink186[4] , \ScanLink175[30] , \ScanLink123[31] , 
        \ScanLink175[29] , \wRegInTop_7_90[15] , \wRegInTop_4_15[11] , 
        \ScanLink113[29] , \wRegOut_7_68[0] , \wRegInBot_4_15[16] , 
        \wRegInTop_5_17[3] , \wRegOut_6_49[6] , \ScanLink113[30] , 
        \wRegInTop_7_5[28] , \ScanLink145[31] , \wRegInTop_7_83[25] , 
        \ScanLink166[19] , \ScanLink129[9] , \ScanLink130[18] , 
        \wRegInTop_7_5[31] , \ScanLink145[28] , \wRegInTop_7_96[11] , 
        \wRegInBot_5_7[26] , \wRegOut_5_18[4] , \wRegOut_6_54[9] , 
        \ScanLink254[3] , \wRegInTop_6_46[1] , \wRegInTop_7_67[7] , 
        \ScanLink134[6] , \wRegOut_7_9[26] , \ScanLink2[17] , 
        \wRegInTop_3_5[26] , \ScanLink14[8] , \wRegOut_4_1[21] , 
        \wRegInBot_6_15[8] , \wRegInTop_6_45[2] , \ScanLink137[5] , 
        \wRegInTop_7_64[4] , \wRegInBot_4_8[25] , \wRegInBot_6_16[17] , 
        \wRegInTop_6_20[15] , \wRegInBot_6_35[26] , \wRegInTop_6_55[25] , 
        \wRegInBot_6_40[16] , \wRegOut_7_110[12] , \wRegInBot_6_63[27] , 
        \wRegInTop_7_18[20] , \wRegInTop_7_78[24] , \wRegInTop_5_14[0] , 
        \wRegOut_6_6[25] , \wRegInTop_6_16[10] , \wRegInTop_6_63[20] , 
        \wRegOut_7_126[17] , \wRegInBot_6_20[12] , \wRegInTop_6_40[11] , 
        \wRegInTop_6_35[21] , \wRegInBot_6_55[22] , \wRegOut_7_105[26] , 
        \wRegOut_7_9[15] , \wRegInTop_1_1[2] , \wRegInTop_2_1[30] , 
        \wRegOut_3_2[17] , \ScanLink10[19] , \wRegInBot_4_8[16] , 
        \wRegInTop_4_15[22] , \wRegInBot_4_15[25] , \wRegInBot_5_7[15] , 
        \ScanLink230[7] , \wRegInBot_6_8[7] , \wRegInTop_6_9[1] , 
        \wRegOut_6_13[18] , \wRegOut_7_68[18] , \wRegOut_6_30[30] , 
        \ScanLink150[2] , \wRegInTop_6_22[5] , \wRegOut_6_45[19] , 
        \wRegOut_6_30[29] , \wRegInTop_7_96[22] , \wRegInTop_6_16[23] , 
        \ScanLink182[4] , \wRegInTop_7_83[16] , \wRegOut_7_126[24] , 
        \ScanLink33[28] , \wRegOut_6_6[16] , \wRegInTop_6_63[13] , 
        \wRegInTop_7_18[13] , \wRegOut_7_105[15] , \wRegInTop_6_20[26] , 
        \wRegInBot_6_20[21] , \wRegInTop_6_35[12] , \wRegInBot_6_55[11] , 
        \wRegInTop_6_40[22] , \ScanLink181[7] , \wRegInBot_6_40[25] , 
        \ScanLink46[18] , \wRegInTop_6_55[16] , \wRegOut_7_110[21] , 
        \ScanLink65[30] , \wRegInBot_6_35[15] , \ScanLink11[5] , 
        \wRegInTop_3_5[15] , \wRegOut_4_1[12] , \ScanLink33[31] , 
        \wRegInBot_6_63[14] , \wRegInTop_7_78[17] , \ScanLink65[29] , 
        \wRegInBot_6_16[24] , \ScanLink233[4] , \wRegOut_4_10[19] , 
        \wRegOut_7_12[8] , \wRegInTop_6_21[6] , \ScanLink153[1] , 
        \wRegOut_7_2[19] , \wRegOut_7_93[19] , \wRegInTop_7_113[19] , 
        \wRegInTop_5_9[13] , \wRegOut_6_18[14] , \wRegOut_7_16[24] , 
        \wRegOut_7_20[21] , \wRegOut_7_55[11] , \wRegOut_7_76[20] , 
        \wRegOut_7_63[14] , \wRegOut_7_35[15] , \wRegInBot_5_10[19] , 
        \ScanLink80[10] , \wRegOut_7_40[25] , \wRegOut_7_73[1] , 
        \wRegOut_6_52[7] , \ScanLink178[12] , \wRegInBot_6_10[5] , 
        \ScanLink95[24] , \wRegOut_6_51[4] , \ScanLink118[16] , 
        \ScanLink132[8] , \wRegInTop_7_61[9] , \wRegOut_7_70[2] , 
        \ScanLink253[24] , \ScanLink12[6] , \wRegInTop_4_6[10] , 
        \ScanLink38[24] , \ScanLink58[20] , \wRegInBot_6_13[6] , 
        \ScanLink183[13] , \ScanLink226[14] , \ScanLink205[25] , 
        \wRegOut_5_15[25] , \ScanLink196[27] , \ScanLink210[11] , 
        \ScanLink246[10] , \ScanLink233[20] , \wRegOut_5_23[20] , 
        \wRegInTop_6_1[14] , \wRegOut_7_98[15] , \wRegInTop_7_118[15] , 
        \wRegOut_6_36[3] , \ScanLink118[25] , \wRegOut_7_17[5] , 
        \ScanLink236[9] , \wRegInTop_7_88[29] , \wRegInTop_2_1[29] , 
        \ScanLink95[17] , \wRegOut_7_9[3] , \wRegInTop_7_88[30] , 
        \ScanLink9[31] , \wRegInTop_5_9[20] , \wRegInBot_5_25[3] , 
        \wRegInTop_5_26[31] , \wRegInTop_5_26[28] , \ScanLink199[5] , 
        \ScanLink75[1] , \ScanLink80[23] , \wRegOut_6_18[27] , 
        \ScanLink178[21] , \wRegOut_7_63[27] , \wRegOut_7_16[17] , 
        \wRegOut_7_40[16] , \wRegEnTop_7_56[0] , \wRegOut_7_35[26] , 
        \wRegInTop_7_104[0] , \wRegInTop_6_39[4] , \wRegInTop_7_18[2] , 
        \wRegOut_7_55[22] , \ScanLink9[28] , \wRegOut_7_20[12] , 
        \wRegOut_7_76[13] , \wRegOut_3_2[24] , \wRegInBot_4_3[29] , 
        \wRegInTop_4_6[23] , \ScanLink38[17] , \wRegOut_5_15[16] , 
        \wRegOut_5_23[13] , \wRegInBot_5_26[0] , \ScanLink76[2] , 
        \wRegInTop_6_1[27] , \wRegOut_7_98[26] , \ScanLink228[5] , 
        \wRegInTop_7_107[3] , \wRegInTop_7_118[26] , \ScanLink148[0] , 
        \ScanLink187[9] , \wRegInTop_7_25[29] , \ScanLink210[22] , 
        \wRegOut_6_35[0] , \wRegInTop_7_50[19] , \wRegInTop_7_73[31] , 
        \wRegOut_7_14[6] , \ScanLink196[14] , \ScanLink233[13] , 
        \wRegInTop_7_25[30] , \wRegInTop_7_73[28] , \ScanLink246[23] , 
        \wRegInBot_4_3[30] , \ScanLink58[13] , \wRegEnBot_6_39[0] , 
        \ScanLink183[20] , \ScanLink226[27] , \ScanLink253[17] , 
        \wRegOut_5_11[27] , \wRegOut_5_27[22] , \wRegEnBot_6_8[0] , 
        \wRegInTop_6_27[8] , \ScanLink205[16] , \wRegInTop_6_5[16] , 
        \wRegInTop_7_1[6] , \wRegOut_7_89[23] , \wRegInTop_7_109[23] , 
        \ScanLink52[4] , \wRegOut_7_109[5] , \wRegInTop_7_123[5] , 
        \wRegOut_1_1[22] , \wRegOut_1_1[11] , \wRegInBot_2_0[12] , 
        \wRegOut_3_6[15] , \wRegInTop_4_2[12] , \ScanLink171[9] , 
        \wRegInTop_7_54[28] , \ScanLink49[16] , \wRegInTop_7_22[8] , 
        \ScanLink214[13] , \wRegOut_6_11[6] , \wRegInTop_7_21[18] , 
        \wRegOut_7_30[0] , \wRegInTop_7_54[31] , \wRegInTop_7_77[19] , 
        \ScanLink242[12] , \ScanLink192[25] , \ScanLink237[22] , 
        \wRegInBot_4_7[18] , \ScanLink29[12] , \wRegInBot_6_53[4] , 
        \ScanLink187[11] , \ScanLink222[16] , \wRegInTop_5_22[19] , 
        \wRegOut_6_9[18] , \ScanLink80[2] , \ScanLink83[1] , \ScanLink91[26] , 
        \ScanLink169[24] , \ScanLink201[27] , \wRegOut_6_12[5] , 
        \ScanLink84[12] , \wRegOut_7_117[9] , \wRegOut_7_33[3] , 
        \wRegOut_3_6[26] , \ScanLink51[7] , \ScanLink109[20] , 
        \wRegInBot_6_50[7] , \wRegInTop_7_2[5] , \wRegOut_7_12[26] , 
        \wRegOut_7_31[17] , \wRegOut_7_67[16] , \wRegOut_7_44[27] , 
        \wRegOut_6_4[9] , \wRegEnTop_6_53[0] , \wRegOut_7_24[23] , 
        \wRegOut_7_51[13] , \wRegInTop_7_120[6] , \wRegOut_7_72[22] , 
        \wRegInTop_4_2[21] , \ScanLink29[21] , \ScanLink187[22] , 
        \ScanLink222[25] , \ScanLink201[14] , \wRegInTop_7_89[5] , 
        \ScanLink49[25] , \ScanLink214[20] , \wRegOut_5_11[14] , 
        \wRegInBot_6_19[19] , \wRegOut_7_54[4] , \ScanLink192[16] , 
        \ScanLink237[11] , \wRegInBot_6_37[0] , \ScanLink242[21] , 
        \wRegOut_7_89[10] , \wRegInTop_7_109[10] , \wRegInBot_2_0[21] , 
        \wRegInBot_4_4[1] , \ScanLink36[0] , \wRegOut_5_24[0] , 
        \wRegEnBot_5_28[0] , \ScanLink108[2] , \wRegOut_5_27[11] , 
        \wRegInTop_4_5[7] , \wRegOut_7_86[2] , \wRegInTop_4_6[4] , 
        \wRegInBot_4_7[2] , \wRegOut_5_0[8] , \wRegInBot_5_8[31] , 
        \wRegInTop_6_5[25] , \wRegInBot_5_8[28] , \wRegOut_7_6[28] , 
        \wRegOut_7_51[20] , \wRegInTop_7_97[9] , \wRegInTop_7_58[0] , 
        \wRegOut_7_24[10] , \wRegOut_7_6[31] , \wRegOut_7_72[11] , 
        \wRegOut_7_12[15] , \wRegOut_7_67[25] , \wRegOut_7_85[1] , 
        \ScanLink35[3] , \wRegOut_7_44[14] , \wRegInBot_5_14[31] , 
        \wRegOut_5_27[3] , \wRegOut_7_31[24] , \wRegInBot_5_14[28] , 
        \wRegInTop_5_28[4] , \ScanLink109[13] , \wRegOut_2_2[30] , 
        \ScanLink8[9] , \wRegInTop_3_1[24] , \ScanLink14[31] , 
        \ScanLink37[19] , \ScanLink42[29] , \wRegOut_6_2[27] , 
        \wRegInTop_6_12[12] , \ScanLink84[21] , \ScanLink91[15] , 
        \wRegInBot_6_34[3] , \wRegOut_7_57[7] , \ScanLink169[17] , 
        \wRegInTop_7_69[12] , \ScanLink229[29] , \wRegOut_7_122[15] , 
        \wRegInBot_6_24[10] , \wRegInTop_6_44[13] , \ScanLink229[30] , 
        \wRegInBot_6_51[20] , \wRegInTop_7_39[9] , \wRegInTop_6_31[23] , 
        \wRegInTop_7_7[8] , \wRegOut_7_101[24] , \wRegInBot_6_31[24] , 
        \wRegInTop_6_51[27] , \wRegOut_6_1[4] , \wRegInTop_6_24[17] , 
        \wRegOut_7_114[10] , \wRegInBot_6_44[14] , \ScanLink14[28] , 
        \ScanLink42[30] , \ScanLink61[18] , \wRegInBot_6_12[15] , 
        \wRegInBot_6_48[5] , \wRegOut_4_5[23] , \wRegOut_4_14[28] , 
        \wRegOut_4_14[31] , \wRegInTop_7_24[6] , \ScanLink177[7] , 
        \ScanLink49[5] , \wRegInBot_5_19[7] , \wRegOut_7_112[4] , 
        \wRegOut_6_17[8] , \wRegOut_7_97[31] , \wRegInTop_7_117[31] , 
        \ScanLink217[2] , \wRegOut_7_97[28] , \wRegInTop_7_117[28] , 
        \wRegOut_2_2[29] , \wRegInBot_5_3[24] , \wRegInTop_7_27[5] , 
        \ScanLink174[4] , \ScanLink6[26] , \wRegInTop_3_1[17] , 
        \wRegInTop_4_11[13] , \wRegInBot_4_11[14] , \wRegInTop_5_29[26] , 
        \wRegOut_6_17[30] , \wRegOut_6_17[29] , \ScanLink214[1] , 
        \wRegOut_6_34[18] , \wRegOut_6_41[31] , \wRegInBot_6_56[9] , 
        \wRegOut_7_19[19] , \wRegOut_6_62[19] , \wRegOut_6_41[28] , 
        \wRegOut_7_111[7] , \wRegInTop_7_92[13] , \wRegOut_7_28[2] , 
        \ScanLink57[9] , \wRegInBot_5_29[21] , \ScanLink98[0] , 
        \wRegInTop_7_87[27] , \wRegOut_6_2[7] , \ScanLink113[3] , 
        \wRegInTop_6_61[4] , \wRegInTop_7_126[8] , \wRegInTop_7_40[2] , 
        \wRegOut_3_5[1] , \wRegOut_4_5[10] , \wRegInTop_4_11[0] , 
        \wRegInTop_5_30[6] , \wRegInTop_6_24[24] , \wRegInBot_6_31[17] , 
        \wRegInBot_6_44[27] , \wRegInTop_6_51[14] , \wRegInTop_7_92[4] , 
        \wRegOut_7_114[23] , \ScanLink199[30] , \wRegOut_5_5[5] , 
        \ScanLink199[29] , \wRegInTop_6_12[21] , \wRegInBot_6_12[26] , 
        \wRegInTop_7_69[21] , \wRegOut_7_122[26] , \wRegInTop_4_3[9] , 
        \wRegOut_6_2[14] , \wRegInBot_6_51[13] , \wRegOut_7_101[17] , 
        \wRegInTop_6_31[10] , \ScanLink0[1] , \wRegOut_1_0[31] , 
        \wRegOut_1_0[28] , \wRegInBot_2_1[8] , \wRegInTop_4_11[20] , 
        \wRegInTop_4_12[3] , \wRegInBot_6_24[23] , \wRegInTop_6_44[20] , 
        \ScanLink162[28] , \wRegInTop_7_1[19] , \ScanLink117[18] , 
        \ScanLink134[30] , \wRegEnBot_6_61[0] , \wRegInTop_7_87[14] , 
        \ScanLink6[15] , \wRegOut_3_6[2] , \wRegOut_5_6[6] , 
        \wRegInTop_5_29[15] , \wRegInBot_5_29[12] , \ScanLink141[19] , 
        \ScanLink162[31] , \wRegInTop_7_91[7] , \ScanLink134[29] , 
        \wRegEnTop_4_5[0] , \wRegInBot_4_11[27] , \ScanLink110[0] , 
        \wRegInTop_7_92[20] , \wRegInTop_6_62[7] , \wRegInTop_7_43[1] , 
        \ScanLink25[9] , \wRegOut_5_0[26] , \wRegInBot_5_3[17] , 
        \wRegOut_7_51[9] , \wRegInBot_5_15[22] , \wRegInTop_7_98[15] , 
        \ScanLink108[19] , \ScanLink38[6] , \wRegInTop_5_23[20] , 
        \ScanLink106[4] , \wRegInTop_7_55[5] , \wRegInBot_5_23[27] , 
        \wRegInBot_5_9[22] , \wRegInTop_5_15[25] , \wRegInBot_6_24[9] , 
        \wRegOut_7_88[4] , \wRegInTop_5_25[1] , \wRegOut_7_7[22] , 
        \wRegInTop_7_87[3] , \wRegInBot_6_1[25] , \wRegInBot_6_39[6] , 
        \wRegInTop_5_26[2] , \ScanLink118[8] , \wRegInTop_7_84[0] , 
        \wRegInBot_4_6[21] , \wRegOut_6_8[21] , \ScanLink105[7] , 
        \wRegInTop_7_35[15] , \wRegOut_7_59[1] , \wRegOut_7_96[8] , 
        \wRegInTop_7_56[6] , \wRegInTop_7_40[25] , \ScanLink186[31] , 
        \wRegInTop_7_16[24] , \wRegInTop_4_8[2] , \wRegInBot_4_9[4] , 
        \wRegInTop_6_18[14] , \ScanLink186[28] , \wRegInTop_7_63[14] , 
        \wRegInBot_6_18[13] , \wRegInBot_5_9[11] , \wRegOut_5_29[5] , 
        \wRegInTop_7_76[20] , \wRegEnBot_6_13[0] , \wRegInTop_7_20[21] , 
        \wRegInTop_7_55[11] , \wRegOut_7_25[30] , \wRegOut_7_73[28] , 
        \ScanLink3[2] , \wRegInBot_2_1[18] , \wRegOut_5_0[15] , 
        \wRegInTop_5_15[16] , \wRegInBot_5_23[14] , \wRegInTop_6_10[7] , 
        \wRegOut_7_7[11] , \wRegOut_7_25[29] , \wRegInTop_7_31[1] , 
        \wRegOut_7_50[19] , \wRegOut_7_73[31] , \ScanLink162[0] , 
        \wRegInTop_4_3[18] , \wRegInBot_5_15[11] , \ScanLink85[18] , 
        \wRegOut_7_23[9] , \ScanLink202[5] , \wRegInTop_7_98[26] , 
        \wRegInTop_5_23[13] , \wRegInBot_6_18[20] , \wRegInTop_7_76[13] , 
        \wRegOut_7_107[3] , \ScanLink243[18] , \ScanLink236[28] , 
        \wRegInTop_7_32[2] , \ScanLink161[3] , \wRegInBot_4_6[12] , 
        \ScanLink28[18] , \wRegOut_6_8[12] , \wRegInTop_6_13[4] , 
        \wRegInTop_7_55[22] , \wRegInTop_7_20[12] , \ScanLink215[19] , 
        \ScanLink236[31] , \wRegInTop_6_18[27] , \ScanLink90[8] , 
        \wRegInTop_7_40[16] , \wRegInTop_7_35[26] , \wRegOut_7_104[0] , 
        \wRegInTop_7_63[27] , \ScanLink201[6] , \wRegOut_5_26[31] , 
        \wRegInTop_7_16[17] , \wRegOut_5_26[28] , \wRegInBot_6_1[16] , 
        \wRegOut_7_88[30] , \wRegInTop_7_108[30] , \wRegOut_7_88[29] , 
        \wRegInTop_7_108[29] , \wRegOut_2_3[23] , \wRegOut_2_3[10] , 
        \wRegInTop_5_7[17] , \wRegOut_6_16[10] , \wRegOut_6_35[21] , 
        \wRegOut_6_40[11] , \wRegOut_6_63[20] , \wRegOut_7_18[20] , 
        \wRegInBot_6_22[7] , \wRegOut_6_60[5] , \wRegOut_7_41[3] , 
        \wRegInBot_3_5[17] , \ScanLink15[11] , \ScanLink23[7] , 
        \wRegInBot_5_28[18] , \wRegOut_6_20[15] , \wRegOut_6_55[25] , 
        \wRegOut_7_78[24] , \ScanLink135[23] , \ScanLink140[13] , 
        \wRegEnTop_6_21[0] , \ScanLink103[26] , \ScanLink116[12] , 
        \wRegInTop_7_0[13] , \ScanLink163[22] , \ScanLink176[16] , 
        \wRegOut_7_93[5] , \wRegOut_4_10[1] , \wRegOut_5_31[7] , 
        \ScanLink120[17] , \ScanLink155[27] , \wRegOut_7_115[30] , 
        \ScanLink248[14] , \ScanLink20[4] , \ScanLink23[14] , 
        \wRegInTop_4_8[14] , \ScanLink36[20] , \ScanLink60[21] , 
        \ScanLink198[23] , \wRegOut_7_115[29] , \wRegOut_4_13[2] , 
        \ScanLink43[10] , \wRegInBot_6_50[19] , \wRegOut_4_15[11] , 
        \wRegOut_5_8[0] , \ScanLink56[24] , \ScanLink75[15] , 
        \wRegInBot_6_25[30] , \wRegInBot_6_25[29] , \wRegOut_7_90[6] , 
        \wRegOut_7_96[11] , \ScanLink228[10] , \wRegInTop_7_116[11] , 
        \ScanLink103[9] , \wRegInTop_7_50[8] , \wRegInTop_7_120[14] , 
        \wRegOut_6_63[6] , \wRegOut_7_42[0] , \wRegInTop_7_103[25] , 
        \wRegInTop_4_10[19] , \ScanLink47[3] , \wRegInBot_6_21[4] , 
        \wRegOut_7_83[25] , \ScanLink103[15] , \wRegInTop_7_93[19] , 
        \ScanLink120[24] , \ScanLink176[25] , \ScanLink135[10] , 
        \ScanLink155[14] , \ScanLink179[1] , \wRegInBot_5_17[1] , 
        \ScanLink140[20] , \ScanLink116[21] , \ScanLink219[4] , 
        \wRegInTop_7_0[20] , \ScanLink163[11] , \wRegOut_7_38[8] , 
        \wRegInTop_6_16[9] , \wRegOut_6_20[26] , \wRegOut_7_78[17] , 
        \wRegInBot_3_1[15] , \wRegInBot_3_5[24] , \wRegOut_4_4[30] , 
        \wRegInTop_5_7[24] , \ScanLink95[5] , \wRegOut_6_55[16] , 
        \wRegOut_6_35[12] , \wRegOut_6_40[22] , \wRegOut_6_16[23] , 
        \wRegOut_7_25[7] , \wRegInBot_6_46[3] , \wRegOut_6_63[13] , 
        \wRegOut_7_18[13] , \wRegInTop_7_120[27] , \ScanLink15[22] , 
        \wRegOut_4_4[29] , \ScanLink23[27] , \wRegOut_4_15[22] , 
        \ScanLink56[17] , \ScanLink96[6] , \wRegInBot_6_45[0] , 
        \wRegOut_7_26[4] , \wRegOut_7_83[16] , \wRegInTop_7_103[16] , 
        \ScanLink207[8] , \wRegOut_7_96[22] , \wRegInTop_7_116[22] , 
        \wRegInTop_6_45[19] , \wRegInTop_7_29[3] , \ScanLink60[12] , 
        \ScanLink75[26] , \wRegInTop_6_30[29] , \wRegInTop_6_13[18] , 
        \wRegInTop_6_30[30] , \wRegInTop_7_68[18] , \ScanLink228[23] , 
        \ScanLink198[10] , \ScanLink248[27] , \wRegOut_4_0[18] , 
        \wRegInTop_4_8[27] , \ScanLink36[13] , \ScanLink43[23] , 
        \ScanLink44[0] , \wRegInBot_5_14[2] , \wRegOut_4_11[13] , 
        \wRegOut_6_23[4] , \wRegInTop_7_107[27] , \wRegInTop_7_124[16] , 
        \wRegOut_7_126[8] , \wRegOut_5_29[26] , \wRegInBot_6_61[6] , 
        \wRegOut_7_87[27] , \wRegOut_7_92[13] , \wRegInTop_7_112[13] , 
        \wRegOut_0_0[16] , \ScanLink11[13] , \wRegInBot_4_11[2] , 
        \ScanLink27[16] , \ScanLink52[26] , \ScanLink60[6] , 
        \wRegInTop_6_17[30] , \wRegInTop_6_34[18] , \wRegInBot_5_30[4] , 
        \wRegInTop_6_41[28] , \wRegInTop_7_111[7] , \ScanLink71[17] , 
        \wRegInTop_6_17[29] , \wRegInTop_6_41[31] , \wRegInTop_7_19[19] , 
        \ScanLink189[15] , \wRegInTop_6_62[19] , \wRegInBot_4_12[1] , 
        \ScanLink32[22] , \ScanLink64[23] , \ScanLink239[26] , 
        \ScanLink47[12] , \wRegInBot_6_6[1] , \wRegInTop_6_7[7] , 
        \ScanLink63[5] , \ScanLink107[24] , \ScanLink172[14] , 
        \wRegInTop_7_97[28] , \wRegOut_7_2[8] , \ScanLink151[25] , 
        \wRegInTop_7_97[31] , \wRegInBot_3_2[4] , \ScanLink11[20] , 
        \wRegInTop_4_14[31] , \wRegInTop_6_4[4] , \ScanLink124[15] , 
        \wRegInTop_7_112[4] , \ScanLink144[11] , \ScanLink131[21] , 
        \wRegInTop_4_14[28] , \wRegInBot_6_5[2] , \ScanLink112[10] , 
        \wRegInTop_7_4[11] , \ScanLink167[20] , \wRegInBot_5_2[0] , 
        \wRegInTop_5_3[15] , \wRegEnTop_5_30[0] , \wRegOut_6_20[7] , 
        \wRegOut_6_24[17] , \wRegOut_6_51[27] , \wRegInBot_6_62[5] , 
        \ScanLink140[8] , \wRegInTop_7_13[9] , \wRegInTop_5_3[6] , 
        \wRegOut_6_12[12] , \wRegOut_6_31[23] , \wRegOut_6_44[13] , 
        \wRegOut_7_69[12] , \ScanLink239[15] , \ScanLink64[10] , 
        \ScanLink27[25] , \ScanLink32[11] , \ScanLink47[21] , 
        \wRegOut_5_16[2] , \ScanLink52[15] , \wRegInBot_6_21[18] , 
        \wRegOut_7_111[18] , \wRegInTop_6_48[7] , \wRegInTop_7_69[1] , 
        \ScanLink71[24] , \wRegInBot_6_54[28] , \wRegInTop_3_3[2] , 
        \ScanLink189[26] , \wRegOut_5_29[15] , \wRegOut_6_47[0] , 
        \wRegInBot_6_54[31] , \wRegOut_7_66[6] , \wRegOut_7_92[20] , 
        \wRegInTop_7_112[20] , \wRegOut_0_0[25] , \wRegInTop_3_0[1] , 
        \wRegInBot_3_1[26] , \wRegInTop_5_19[5] , \wRegInTop_6_55[8] , 
        \wRegInTop_7_124[25] , \wRegInBot_3_1[7] , \wRegOut_4_11[20] , 
        \wRegInTop_7_107[14] , \wRegInTop_5_0[5] , \wRegInTop_5_3[26] , 
        \wRegOut_6_31[10] , \wRegOut_7_87[14] , \wRegOut_6_44[20] , 
        \wRegOut_5_15[1] , \wRegOut_6_12[21] , \wRegOut_6_44[3] , 
        \wRegOut_7_65[5] , \wRegOut_7_69[21] , \ScanLink244[9] , 
        \wRegOut_6_24[24] , \wRegOut_6_51[14] , \ScanLink131[12] , 
        \ScanLink144[22] , \wRegEnTop_7_24[0] , \wRegInBot_5_1[3] , 
        \ScanLink112[23] , \ScanLink167[13] , \wRegInTop_7_4[22] , 
        \wRegOut_4_6[9] , \ScanLink107[17] , \ScanLink172[27] , 
        \wRegInBot_0_0[2] , \ScanLink0[8] , \wRegOut_2_0[3] , 
        \wRegInTop_2_0[23] , \ScanLink8[22] , \wRegInBot_4_2[23] , 
        \wRegInTop_4_7[30] , \ScanLink124[26] , \ScanLink139[3] , 
        \ScanLink151[16] , \wRegInTop_7_72[22] , \ScanLink211[31] , 
        \ScanLink225[0] , \ScanLink232[19] , \ScanLink247[29] , 
        \wRegInTop_4_7[29] , \wRegInTop_7_24[23] , \ScanLink211[28] , 
        \wRegInTop_7_51[13] , \ScanLink247[30] , \wRegOut_7_120[6] , 
        \ScanLink59[19] , \wRegInTop_6_37[2] , \wRegInTop_7_12[26] , 
        \wRegInTop_7_16[4] , \ScanLink145[5] , \wRegInTop_7_31[17] , 
        \wRegInTop_7_44[27] , \wRegOut_5_22[19] , \wRegOut_6_38[5] , 
        \wRegInTop_7_67[16] , \wRegOut_7_19[3] , \wRegInTop_6_1[9] , 
        \ScanLink66[8] , \wRegOut_7_7[5] , \wRegInBot_6_5[27] , 
        \ScanLink197[3] , \wRegInTop_7_117[9] , \wRegOut_7_4[6] , 
        \wRegOut_7_54[31] , \wRegOut_7_77[19] , \wRegInBot_5_27[25] , 
        \wRegEnTop_6_7[0] , \wRegOut_7_54[28] , \ScanLink194[0] , 
        \wRegOut_7_3[20] , \wRegOut_7_21[18] , \ScanLink78[4] , 
        \wRegInTop_2_0[10] , \wRegOut_2_3[0] , \wRegOut_5_4[24] , 
        \wRegInTop_5_11[27] , \wRegInBot_5_28[6] , \wRegOut_6_26[9] , 
        \wRegInTop_7_89[23] , \wRegInTop_7_109[5] , \wRegOut_7_123[5] , 
        \ScanLink226[3] , \wRegInBot_5_11[20] , \ScanLink81[29] , 
        \wRegInTop_5_5[8] , \wRegInTop_5_27[22] , \ScanLink81[30] , 
        \wRegInTop_6_34[1] , \ScanLink146[6] , \wRegInTop_7_15[7] , 
        \wRegInBot_6_5[14] , \wRegEnBot_3_1[0] , \wRegInBot_4_2[10] , 
        \wRegOut_4_3[4] , \wRegInTop_7_31[24] , \wRegInTop_7_44[14] , 
        \wRegOut_7_60[8] , \wRegInTop_7_67[25] , \ScanLink241[4] , 
        \wRegOut_5_4[17] , \wRegInTop_6_53[6] , \ScanLink121[1] , 
        \wRegInTop_7_12[15] , \ScanLink182[19] , \wRegInTop_7_72[11] , 
        \wRegInTop_7_51[20] , \wRegInTop_7_72[0] , \wRegInTop_7_24[10] , 
        \wRegInBot_5_11[13] , \ScanLink179[18] , \ScanLink242[7] , 
        \wRegInTop_5_27[11] , \wRegInBot_5_27[16] , \wRegInTop_6_50[5] , 
        \wRegInTop_7_71[3] , \ScanLink122[2] , \ScanLink8[11] , 
        \wRegInTop_5_11[14] , \wRegInTop_7_89[10] , \ScanLink5[5] , 
        \ScanLink6[6] , \wRegInBot_3_7[9] , \wRegOut_4_0[7] , 
        \wRegInTop_5_8[19] , \wRegOut_7_3[13] , \wRegInTop_4_10[10] , 
        \wRegInBot_5_17[8] , \wRegInBot_5_28[22] , \ScanLink88[3] , 
        \ScanLink116[31] , \ScanLink135[19] , \ScanLink140[29] , 
        \wRegOut_6_19[7] , \ScanLink116[28] , \wRegInTop_7_0[30] , 
        \wRegOut_7_38[1] , \ScanLink140[30] , \wRegInTop_7_86[24] , 
        \ScanLink163[18] , \ScanLink7[25] , \wRegInBot_4_10[17] , 
        \wRegInTop_7_0[29] , \wRegInTop_7_93[10] , \wRegInBot_5_2[27] , 
        \wRegInTop_5_28[25] , \ScanLink179[8] , \ScanLink204[2] , 
        \wRegOut_7_101[4] , \wRegInTop_3_0[27] , \ScanLink59[6] , 
        \wRegInTop_6_16[0] , \wRegInTop_7_37[6] , \wRegInBot_6_45[9] , 
        \wRegInTop_7_9[7] , \ScanLink164[7] , \ScanLink207[1] , 
        \wRegOut_4_4[20] , \wRegInTop_6_15[3] , \wRegInTop_7_34[5] , 
        \ScanLink167[4] , \wRegOut_7_102[7] , \wRegEnTop_7_122[0] , 
        \wRegInBot_6_13[16] , \ScanLink198[19] , \wRegOut_2_3[19] , 
        \ScanLink7[16] , \ScanLink44[9] , \wRegInTop_6_50[24] , 
        \wRegInBot_6_58[6] , \wRegOut_6_3[24] , \wRegInTop_6_25[14] , 
        \wRegInBot_6_30[27] , \wRegInBot_6_25[13] , \wRegInBot_6_45[17] , 
        \wRegOut_7_115[13] , \wRegInTop_6_45[10] , \wRegInBot_6_50[23] , 
        \wRegInTop_6_13[11] , \wRegInTop_6_30[20] , \wRegOut_7_100[27] , 
        \wRegInTop_7_68[11] , \wRegOut_7_123[16] , \wRegInTop_3_0[14] , 
        \ScanLink15[18] , \wRegOut_4_10[8] , \wRegInBot_4_10[24] , 
        \wRegInBot_5_2[14] , \wRegOut_6_16[19] , \wRegOut_6_35[28] , 
        \ScanLink100[3] , \wRegOut_6_40[18] , \wRegOut_7_18[30] , 
        \wRegOut_6_63[30] , \wRegInTop_7_53[2] , \wRegOut_6_63[29] , 
        \wRegOut_7_18[29] , \wRegOut_6_35[31] , \wRegInTop_5_28[16] , 
        \wRegInTop_7_93[23] , \wRegInTop_4_10[23] , \wRegInTop_5_23[6] , 
        \wRegInBot_5_28[11] , \wRegInTop_7_81[4] , \wRegInTop_5_20[5] , 
        \wRegOut_6_3[17] , \wRegInBot_6_50[10] , \wRegInTop_7_86[17] , 
        \wRegOut_7_100[14] , \wRegInTop_6_13[22] , \wRegInBot_6_25[20] , 
        \wRegInTop_6_30[13] , \wRegInTop_6_45[23] , \wRegInTop_7_68[22] , 
        \wRegOut_7_123[25] , \ScanLink228[19] , \wRegOut_4_4[13] , 
        \ScanLink36[30] , \ScanLink36[29] , \ScanLink60[28] , 
        \wRegInBot_6_13[25] , \wRegInTop_6_25[27] , \wRegInBot_6_45[24] , 
        \wRegInTop_7_82[7] , \wRegOut_7_115[20] , \ScanLink43[19] , 
        \wRegInTop_6_50[17] , \ScanLink60[31] , \wRegInBot_6_30[14] , 
        \wRegOut_7_42[9] , \wRegOut_4_15[18] , \wRegOut_5_8[9] , 
        \wRegOut_7_96[18] , \wRegInTop_7_116[18] , \ScanLink103[0] , 
        \wRegInTop_7_50[1] , \wRegInBot_5_9[18] , \wRegOut_7_73[21] , 
        \wRegOut_1_0[21] , \wRegOut_1_0[12] , \wRegInBot_2_1[11] , 
        \ScanLink41[4] , \wRegOut_7_7[18] , \wRegInBot_5_11[6] , 
        \wRegOut_7_25[20] , \wRegOut_7_50[10] , \ScanLink85[11] , 
        \wRegOut_7_13[25] , \wRegOut_7_30[14] , \wRegOut_7_45[24] , 
        \wRegOut_7_66[15] , \wRegOut_7_23[0] , \wRegOut_3_7[16] , 
        \ScanLink28[11] , \wRegInBot_5_15[18] , \ScanLink108[23] , 
        \wRegOut_6_9[5] , \ScanLink93[2] , \wRegInBot_6_40[4] , 
        \ScanLink90[25] , \wRegInTop_7_31[8] , \ScanLink162[9] , 
        \ScanLink168[27] , \ScanLink90[1] , \wRegOut_7_20[3] , 
        \ScanLink200[24] , \wRegOut_7_104[9] , \wRegInTop_4_3[11] , 
        \wRegInBot_6_18[29] , \wRegInBot_6_43[7] , \ScanLink186[12] , 
        \ScanLink193[26] , \ScanLink223[15] , \ScanLink236[21] , 
        \ScanLink243[11] , \ScanLink42[7] , \ScanLink48[15] , 
        \ScanLink215[10] , \wRegInBot_6_18[30] , \wRegEnTop_7_9[0] , 
        \wRegEnTop_6_40[0] , \wRegOut_7_119[6] , \wRegInBot_2_1[22] , 
        \wRegOut_5_10[24] , \wRegInBot_5_12[5] , \wRegOut_7_88[20] , 
        \wRegInTop_7_108[20] , \wRegInTop_5_23[30] , \wRegOut_5_26[21] , 
        \wRegInTop_6_4[15] , \wRegInBot_6_24[0] , \wRegOut_7_47[4] , 
        \ScanLink90[16] , \ScanLink168[14] , \ScanLink108[10] , 
        \ScanLink25[0] , \wRegInTop_5_23[29] , \ScanLink85[22] , 
        \wRegOut_7_45[17] , \ScanLink26[3] , \wRegOut_4_15[5] , 
        \wRegInTop_5_25[8] , \wRegOut_7_13[16] , \wRegOut_7_30[27] , 
        \wRegOut_7_66[26] , \wRegOut_7_95[2] , \wRegOut_7_73[12] , 
        \wRegOut_5_26[12] , \wRegInTop_6_4[26] , \wRegOut_7_25[13] , 
        \wRegInTop_7_48[3] , \wRegOut_7_50[23] , \wRegOut_7_59[8] , 
        \wRegOut_7_96[1] , \wRegInTop_2_0[19] , \wRegOut_2_3[9] , 
        \wRegInBot_3_4[3] , \wRegOut_3_7[25] , \wRegInTop_4_3[22] , 
        \wRegOut_5_10[17] , \ScanLink118[1] , \wRegInTop_7_84[9] , 
        \ScanLink48[26] , \wRegInBot_6_27[3] , \wRegInTop_7_20[31] , 
        \wRegOut_7_44[7] , \wRegOut_7_88[13] , \wRegInTop_7_108[13] , 
        \ScanLink193[15] , \ScanLink236[12] , \ScanLink243[22] , 
        \wRegInTop_7_76[29] , \ScanLink215[23] , \wRegInTop_7_20[28] , 
        \wRegInTop_7_55[18] , \wRegInBot_4_6[31] , \wRegInTop_7_76[30] , 
        \wRegInBot_4_6[28] , \ScanLink28[22] , \wRegOut_6_8[28] , 
        \ScanLink200[17] , \wRegInTop_7_99[6] , \wRegOut_6_8[31] , 
        \ScanLink186[21] , \ScanLink223[26] , \wRegOut_7_99[16] , 
        \wRegInTop_7_119[16] , \wRegInTop_3_5[5] , \wRegInTop_6_0[17] , 
        \wRegInBot_5_4[7] , \wRegInTop_5_5[1] , \wRegOut_5_10[5] , 
        \wRegOut_5_22[23] , \wRegOut_3_3[14] , \wRegInTop_4_7[13] , 
        \ScanLink39[27] , \wRegOut_5_14[26] , \ScanLink121[8] , 
        \wRegInTop_7_51[30] , \wRegInTop_7_72[18] , \ScanLink247[13] , 
        \ScanLink197[24] , \ScanLink232[23] , \wRegInTop_7_72[9] , 
        \ScanLink59[23] , \wRegInTop_7_24[19] , \wRegInTop_7_51[29] , 
        \ScanLink211[12] , \wRegOut_6_41[7] , \wRegOut_7_60[1] , 
        \ScanLink204[26] , \ScanLink252[27] , \wRegInBot_4_2[19] , 
        \ScanLink182[10] , \ScanLink227[17] , \ScanLink8[18] , 
        \wRegInTop_3_6[6] , \wRegInBot_3_7[0] , \wRegInTop_5_8[10] , 
        \wRegInTop_5_27[18] , \ScanLink81[13] , \ScanLink94[27] , 
        \ScanLink119[15] , \wRegOut_7_63[2] , \wRegInTop_7_89[19] , 
        \wRegOut_6_42[4] , \ScanLink179[11] , \wRegOut_7_34[16] , 
        \wRegOut_7_41[26] , \wRegOut_6_19[17] , \wRegOut_7_17[27] , 
        \wRegOut_7_62[17] , \wRegInTop_5_6[2] , \wRegOut_3_3[27] , 
        \wRegInBot_5_7[4] , \wRegOut_5_13[6] , \wRegOut_7_77[23] , 
        \ScanLink59[10] , \wRegOut_7_21[22] , \wRegOut_7_54[12] , 
        \ScanLink204[15] , \wRegInTop_4_7[20] , \ScanLink39[14] , 
        \wRegOut_6_25[3] , \ScanLink182[23] , \ScanLink227[24] , 
        \ScanLink252[14] , \ScanLink197[17] , \ScanLink232[10] , 
        \ScanLink211[21] , \ScanLink225[9] , \ScanLink247[20] , 
        \wRegOut_5_14[15] , \wRegInBot_6_0[6] , \wRegInTop_6_1[0] , 
        \ScanLink158[3] , \wRegOut_5_22[10] , \wRegInTop_6_0[24] , 
        \wRegOut_7_99[25] , \ScanLink238[6] , \wRegInTop_7_119[25] , 
        \ScanLink66[1] , \ScanLink11[30] , \ScanLink11[29] , \wRegOut_4_5[3] , 
        \wRegInBot_4_9[26] , \wRegInBot_4_14[6] , \ScanLink65[2] , 
        \wRegInTop_6_2[3] , \wRegOut_7_3[30] , \wRegEnTop_7_45[0] , 
        \wRegOut_7_77[10] , \wRegInTop_7_117[0] , \wRegInBot_6_3[5] , 
        \wRegInTop_6_29[7] , \wRegOut_7_3[29] , \wRegOut_7_54[21] , 
        \ScanLink194[9] , \wRegOut_7_21[11] , \wRegOut_7_41[15] , 
        \wRegInTop_5_8[23] , \wRegOut_7_34[25] , \wRegInTop_7_114[3] , 
        \wRegInBot_5_11[30] , \wRegInBot_5_11[29] , \wRegOut_6_19[24] , 
        \wRegOut_7_62[24] , \wRegOut_7_17[14] , \ScanLink81[20] , 
        \ScanLink179[22] , \ScanLink189[6] , \wRegOut_6_7[26] , 
        \wRegInBot_6_21[11] , \wRegOut_6_26[0] , \wRegInTop_6_34[8] , 
        \ScanLink119[26] , \ScanLink94[14] , \wRegInTop_6_41[12] , 
        \wRegInTop_7_69[8] , \wRegInTop_6_34[22] , \wRegInBot_6_54[21] , 
        \wRegOut_7_104[25] , \wRegInTop_6_62[23] , \wRegInTop_7_19[23] , 
        \wRegInBot_5_2[9] , \ScanLink47[31] , \ScanLink64[19] , 
        \wRegInTop_6_17[13] , \wRegOut_7_127[14] , \wRegInBot_6_17[14] , 
        \wRegInBot_6_18[4] , \wRegInBot_6_62[24] , \ScanLink32[18] , 
        \ScanLink47[28] , \wRegInBot_6_34[25] , \wRegInTop_6_54[26] , 
        \wRegInTop_7_79[27] , \wRegInTop_6_21[16] , \wRegOut_7_111[11] , 
        \wRegInTop_3_4[25] , \wRegOut_4_0[22] , \wRegOut_4_11[30] , 
        \wRegInBot_6_41[15] , \wRegInTop_6_55[1] , \ScanLink127[6] , 
        \wRegInTop_7_74[7] , \wRegOut_4_11[29] , \ScanLink19[4] , 
        \wRegOut_6_47[9] , \wRegOut_7_92[29] , \ScanLink247[3] , 
        \wRegInTop_7_112[29] , \wRegOut_1_1[6] , \ScanLink3[27] , 
        \wRegInBot_5_6[25] , \wRegOut_7_92[30] , \wRegInTop_7_112[30] , 
        \wRegInTop_3_0[8] , \wRegOut_4_6[0] , \wRegOut_6_12[31] , 
        \wRegEnTop_6_18[0] , \wRegOut_6_31[19] , \wRegInTop_6_56[2] , 
        \wRegInTop_7_77[4] , \ScanLink124[5] , \wRegOut_7_8[25] , 
        \wRegOut_7_69[31] , \wRegOut_6_12[28] , \wRegOut_6_44[29] , 
        \wRegOut_7_69[28] , \ScanLink244[0] , \wRegOut_6_44[30] , 
        \wRegInTop_7_97[12] , \wRegInBot_4_14[15] , \wRegInTop_3_4[16] , 
        \wRegInTop_4_14[12] , \wRegOut_5_15[8] , \wRegOut_7_78[3] , 
        \wRegEnBot_5_4[0] , \wRegOut_6_59[5] , \wRegInTop_7_82[26] , 
        \wRegInTop_6_31[5] , \wRegInTop_7_10[3] , \ScanLink143[2] , 
        \wRegOut_4_0[11] , \ScanLink223[7] , \wRegOut_7_126[1] , 
        \wRegInBot_6_17[27] , \wRegInBot_6_62[17] , \wRegInTop_7_79[14] , 
        \wRegInTop_6_21[25] , \ScanLink191[4] , \wRegInBot_6_41[26] , 
        \wRegOut_7_111[22] , \wRegInBot_4_9[15] , \wRegInBot_6_6[8] , 
        \wRegOut_6_7[15] , \wRegInBot_6_34[16] , \wRegInTop_6_54[15] , 
        \wRegOut_7_104[16] , \wRegInTop_6_17[20] , \wRegInBot_6_21[22] , 
        \wRegInTop_6_34[11] , \wRegInBot_6_54[12] , \wRegOut_7_1[2] , 
        \wRegInTop_6_41[21] , \wRegOut_7_127[27] , \wRegInTop_7_19[10] , 
        \wRegInTop_6_62[10] , \ScanLink131[28] , \ScanLink144[18] , 
        \ScanLink167[30] , \ScanLink192[7] , \wRegOut_0_0[12] , 
        \wRegOut_1_1[18] , \ScanLink3[14] , \wRegInBot_4_12[8] , 
        \wRegInTop_4_14[21] , \ScanLink131[31] , \wRegInTop_7_4[18] , 
        \ScanLink167[29] , \wRegInBot_4_14[26] , \ScanLink112[19] , 
        \wRegInTop_7_82[15] , \wRegOut_7_2[1] , \wRegInTop_7_97[21] , 
        \wRegInTop_6_32[6] , \ScanLink140[1] , \wRegInTop_7_13[0] , 
        \wRegEnTop_2_0[0] , \wRegInTop_2_0[7] , \wRegInTop_2_1[20] , 
        \wRegOut_5_5[27] , \wRegInBot_5_6[16] , \ScanLink220[4] , 
        \wRegInBot_5_10[23] , \wRegInTop_5_26[21] , \wRegInTop_6_24[2] , 
        \wRegOut_7_8[16] , \ScanLink156[5] , \wRegOut_7_125[2] , 
        \ScanLink178[31] , \wRegInTop_5_10[24] , \ScanLink178[28] , 
        \wRegInTop_7_88[20] , \ScanLink236[0] , \wRegInBot_5_26[26] , 
        \ScanLink68[7] , \wRegInTop_2_1[13] , \ScanLink9[21] , 
        \wRegOut_7_2[23] , \ScanLink184[3] , \wRegInTop_7_119[6] , 
        \ScanLink9[12] , \wRegInBot_4_3[20] , \wRegInTop_5_9[30] , 
        \wRegInTop_5_9[29] , \ScanLink75[8] , \wRegEnTop_7_99[0] , 
        \wRegInTop_7_104[9] , \wRegInBot_5_26[9] , \wRegInBot_6_4[24] , 
        \ScanLink187[0] , \ScanLink148[9] , \wRegOut_6_28[6] , 
        \wRegInTop_5_11[4] , \wRegInTop_6_27[1] , \wRegInTop_7_13[25] , 
        \ScanLink183[29] , \wRegInTop_7_66[15] , \wRegOut_6_35[9] , 
        \wRegInTop_7_25[20] , \ScanLink155[6] , \wRegInTop_7_30[14] , 
        \wRegInTop_7_45[24] , \ScanLink183[30] , \wRegInTop_7_50[10] , 
        \ScanLink235[3] , \wRegInTop_7_73[21] , \wRegOut_7_2[10] , 
        \wRegOut_7_20[28] , \wRegOut_7_55[18] , \wRegOut_7_76[30] , 
        \wRegInTop_5_10[17] , \wRegOut_7_20[31] , \wRegOut_7_76[29] , 
        \wRegInBot_5_26[15] , \wRegInTop_6_40[6] , \wRegInTop_7_61[0] , 
        \wRegInTop_7_88[13] , \ScanLink132[1] , \wRegInBot_2_2[2] , 
        \wRegInTop_2_3[4] , \wRegInBot_3_0[25] , \wRegInBot_3_0[16] , 
        \ScanLink10[10] , \wRegInBot_4_3[13] , \wRegInTop_4_6[19] , 
        \wRegOut_5_5[14] , \wRegInTop_5_26[12] , \wRegInBot_5_10[10] , 
        \ScanLink80[19] , \wRegOut_7_73[8] , \ScanLink252[4] , 
        \ScanLink131[2] , \wRegInTop_7_50[23] , \wRegInTop_5_8[4] , 
        \wRegEnBot_5_11[0] , \wRegInTop_6_43[5] , \wRegInTop_7_62[3] , 
        \ScanLink210[18] , \ScanLink233[30] , \wRegInTop_7_25[13] , 
        \wRegInTop_7_66[26] , \wRegInTop_7_73[12] , \ScanLink246[19] , 
        \ScanLink233[29] , \wRegInBot_5_9[2] , \ScanLink58[30] , 
        \ScanLink251[7] , \wRegInTop_7_13[16] , \ScanLink33[21] , 
        \wRegInTop_5_2[16] , \wRegInTop_5_12[7] , \wRegOut_5_23[29] , 
        \ScanLink58[29] , \wRegInTop_7_45[17] , \wRegInTop_7_30[27] , 
        \wRegOut_5_23[30] , \wRegInBot_6_4[17] , \wRegInTop_6_9[8] , 
        \wRegOut_6_13[11] , \wRegOut_7_68[11] , \wRegOut_6_45[10] , 
        \wRegInBot_5_23[4] , \ScanLink73[6] , \wRegOut_6_25[14] , 
        \wRegOut_6_30[20] , \wRegOut_6_50[24] , \wRegOut_6_30[4] , 
        \ScanLink113[13] , \wRegInTop_7_5[12] , \wRegOut_7_11[2] , 
        \ScanLink166[23] , \wRegEnTop_7_108[0] , \ScanLink130[22] , 
        \ScanLink145[12] , \ScanLink150[26] , \ScanLink106[27] , 
        \ScanLink125[16] , \wRegInTop_7_102[7] , \ScanLink173[17] , 
        \ScanLink46[11] , \wRegOut_7_110[28] , \wRegOut_7_110[31] , 
        \wRegOut_4_10[10] , \ScanLink26[15] , \ScanLink65[20] , 
        \ScanLink238[25] , \ScanLink70[14] , \wRegInBot_6_20[31] , 
        \wRegInBot_6_55[18] , \ScanLink188[16] , \wRegInBot_5_20[7] , 
        \ScanLink53[25] , \ScanLink70[5] , \wRegInBot_6_20[28] , 
        \wRegOut_5_28[25] , \ScanLink153[8] , \wRegInTop_7_101[4] , 
        \wRegOut_6_33[7] , \wRegOut_7_93[10] , \wRegInTop_7_106[24] , 
        \wRegInTop_7_113[10] , \ScanLink17[2] , \wRegInTop_4_15[18] , 
        \wRegEnTop_5_23[0] , \wRegOut_7_12[1] , \ScanLink106[14] , 
        \ScanLink125[25] , \ScanLink129[0] , \wRegOut_7_86[24] , 
        \wRegInTop_7_125[15] , \ScanLink150[15] , \wRegInTop_7_96[18] , 
        \ScanLink173[24] , \ScanLink113[20] , \wRegOut_7_68[9] , 
        \ScanLink130[11] , \wRegInTop_7_5[21] , \ScanLink166[10] , 
        \ScanLink249[5] , \wCtrlOut_0[0] , \wRegOut_4_8[6] , 
        \wRegInTop_5_2[25] , \wRegOut_6_13[22] , \wRegOut_6_25[27] , 
        \wRegInTop_6_46[8] , \ScanLink145[21] , \wRegOut_6_50[17] , 
        \wRegOut_6_54[0] , \wRegEnBot_6_58[0] , \wRegOut_7_68[22] , 
        \wRegOut_7_75[6] , \wRegInBot_6_16[2] , \wRegOut_6_30[13] , 
        \wRegOut_6_45[23] , \ScanLink10[23] , \ScanLink14[1] , 
        \wRegOut_4_1[31] , \wRegOut_4_1[28] , \wRegOut_4_10[23] , 
        \wRegInTop_7_106[17] , \wRegOut_7_86[17] , \ScanLink26[26] , 
        \wRegInTop_5_14[9] , \wRegOut_5_28[16] , \wRegInTop_7_125[26] , 
        \ScanLink70[27] , \wRegInBot_6_15[1] , \wRegOut_6_57[3] , 
        \wRegOut_7_76[5] , \wRegOut_7_93[23] , \wRegInTop_7_113[23] , 
        \wRegInTop_6_63[29] , \wRegInTop_7_18[29] , \ScanLink53[16] , 
        \wRegInTop_6_16[19] , \wRegInTop_6_35[31] , \ScanLink188[25] , 
        \wRegInTop_7_18[30] , \wRegInTop_6_40[18] , \wRegInTop_6_58[4] , 
        \wRegInTop_6_63[30] , \wRegInTop_7_79[2] , \wRegInTop_6_35[28] , 
        \wRegEnTop_7_37[0] , \ScanLink33[12] , \ScanLink46[22] , 
        \ScanLink65[13] , \ScanLink238[16] , \wRegInBot_3_4[14] , 
        \wRegOut_4_5[19] , \wRegOut_4_14[12] , \wRegInTop_7_102[26] , 
        \wRegOut_3_5[8] , \wRegInBot_6_31[7] , \wRegOut_7_52[3] , 
        \wRegOut_7_82[26] , \wRegInTop_7_69[28] , \wRegOut_7_97[12] , 
        \wRegInTop_7_121[17] , \wRegInTop_7_117[12] , \wRegInBot_4_2[6] , 
        \wRegInTop_6_12[28] , \wRegInTop_4_3[0] , \wRegOut_7_80[5] , 
        \ScanLink22[17] , \wRegOut_5_22[7] , \ScanLink74[16] , 
        \wRegInTop_6_44[30] , \ScanLink229[13] , \wRegInTop_7_69[31] , 
        \wRegInTop_4_9[17] , \ScanLink30[7] , \wRegInTop_6_12[31] , 
        \wRegEnTop_6_32[0] , \wRegInTop_6_31[19] , \ScanLink37[23] , 
        \ScanLink57[27] , \wRegInTop_6_44[29] , \wRegInTop_4_11[9] , 
        \ScanLink42[13] , \ScanLink249[17] , \ScanLink14[12] , 
        \wRegInTop_4_0[3] , \wRegInBot_4_1[5] , \ScanLink33[4] , 
        \ScanLink61[22] , \ScanLink199[20] , \wRegOut_5_21[4] , 
        \ScanLink121[14] , \ScanLink154[24] , \wRegInTop_7_92[30] , 
        \ScanLink177[15] , \wRegOut_7_83[6] , \wRegInTop_7_92[29] , 
        \ScanLink102[25] , \wRegInBot_2_1[1] , \wRegInTop_4_11[29] , 
        \ScanLink117[11] , \wRegInTop_7_1[10] , \ScanLink162[21] , 
        \wRegOut_2_2[20] , \wRegOut_2_2[13] , \wRegInTop_4_11[30] , 
        \ScanLink141[10] , \wRegOut_6_21[16] , \wRegOut_6_54[26] , 
        \ScanLink134[20] , \wRegOut_7_51[0] , \ScanLink8[0] , \ScanLink14[21] , 
        \wRegInTop_4_9[24] , \ScanLink37[10] , \wRegInTop_5_6[14] , 
        \wRegOut_6_17[13] , \wRegInBot_6_32[4] , \wRegOut_6_62[23] , 
        \wRegOut_7_19[23] , \wRegOut_7_79[27] , \wRegOut_6_41[12] , 
        \ScanLink110[9] , \wRegInTop_7_43[8] , \ScanLink42[20] , 
        \ScanLink54[3] , \wRegOut_6_34[22] , \wRegOut_7_114[19] , 
        \wRegInTop_7_125[2] , \ScanLink61[11] , \ScanLink199[13] , 
        \ScanLink249[24] , \ScanLink22[24] , \ScanLink57[14] , 
        \ScanLink74[25] , \wRegInBot_6_24[19] , \wRegInBot_6_51[30] , 
        \ScanLink229[20] , \wRegInTop_6_18[6] , \wRegInTop_7_39[0] , 
        \wRegOut_6_17[1] , \ScanLink86[5] , \wRegInBot_6_51[29] , 
        \wRegInTop_7_7[1] , \wRegOut_7_36[7] , \wRegInBot_3_4[27] , 
        \wRegInBot_6_55[3] , \wRegOut_7_97[21] , \wRegInTop_7_117[21] , 
        \wRegOut_4_14[21] , \wRegInTop_5_6[27] , \wRegOut_6_14[2] , 
        \wRegOut_7_35[4] , \wRegOut_7_82[15] , \wRegInTop_7_102[15] , 
        \ScanLink214[8] , \wRegInTop_7_121[24] , \wRegOut_6_17[20] , 
        \ScanLink85[6] , \wRegInBot_6_56[0] , \wRegOut_6_62[10] , 
        \wRegOut_7_19[10] , \wRegOut_6_34[11] , \wRegOut_6_21[25] , 
        \wRegOut_6_41[21] , \wRegOut_6_54[15] , \wRegOut_3_3[6] , 
        \wRegInTop_4_2[31] , \wRegInTop_4_2[28] , \ScanLink57[0] , 
        \wRegInBot_5_29[31] , \wRegOut_7_79[14] , \wRegInBot_5_29[28] , 
        \ScanLink117[22] , \ScanLink209[7] , \wRegInTop_7_1[23] , 
        \ScanLink162[12] , \ScanLink134[13] , \ScanLink98[9] , 
        \ScanLink102[16] , \ScanLink121[27] , \ScanLink141[23] , 
        \wRegInTop_7_126[1] , \wRegInTop_7_4[2] , \ScanLink154[17] , 
        \ScanLink169[2] , \wRegInTop_7_21[22] , \ScanLink177[26] , 
        \ScanLink214[29] , \ScanLink242[31] , \wRegInBot_6_19[10] , 
        \wRegInTop_7_54[12] , \ScanLink214[30] , \ScanLink237[18] , 
        \wRegInBot_6_37[9] , \wRegInTop_7_77[23] , \ScanLink242[28] , 
        \wRegInBot_4_4[8] , \wRegInBot_4_7[22] , \ScanLink29[31] , 
        \wRegInTop_7_17[27] , \ScanLink29[28] , \wRegInTop_6_19[17] , 
        \wRegInTop_7_62[17] , \ScanLink115[4] , \wRegInTop_7_34[16] , 
        \wRegInTop_7_46[5] , \wRegEnBot_4_14[0] , \wRegOut_6_9[22] , 
        \wRegInTop_7_41[26] , \ScanLink36[9] , \wRegOut_5_24[9] , 
        \wRegOut_5_27[18] , \wRegOut_7_49[2] , \wRegInBot_2_0[31] , 
        \wRegOut_3_0[5] , \wRegOut_5_3[2] , \wRegInTop_7_109[19] , 
        \wRegInBot_6_0[26] , \wRegOut_7_89[19] , \wRegOut_7_85[8] , 
        \wRegInTop_7_94[3] , \ScanLink28[5] , \wRegInTop_4_14[4] , 
        \wRegInBot_5_8[21] , \wRegInBot_6_29[5] , \wRegOut_7_6[21] , 
        \wRegOut_7_51[29] , \wRegInTop_7_58[9] , \wRegInTop_7_97[0] , 
        \wRegOut_7_24[19] , \wRegOut_7_51[30] , \wRegOut_7_72[18] , 
        \wRegOut_5_0[1] , \wRegInTop_5_14[26] , \wRegOut_7_98[7] , 
        \wRegInBot_5_22[24] , \ScanLink84[31] , \ScanLink116[7] , 
        \wRegInTop_7_45[6] , \wRegInBot_2_0[28] , \wRegInBot_5_14[21] , 
        \wRegInTop_5_22[23] , \wRegInTop_7_99[16] , \ScanLink84[28] , 
        \wRegOut_5_1[25] , \wRegOut_6_7[3] , \ScanLink3[19] , \wRegOut_2_0[7] , 
        \wRegInTop_2_0[27] , \wRegInBot_4_7[11] , \wRegInBot_6_0[15] , 
        \wRegInTop_6_19[24] , \wRegInTop_7_62[24] , \wRegInTop_7_17[14] , 
        \wRegOut_7_30[9] , \ScanLink211[5] , \wRegOut_5_1[16] , 
        \wRegInTop_5_22[10] , \wRegOut_6_9[11] , \ScanLink187[18] , 
        \wRegInBot_6_19[23] , \wRegInTop_7_21[11] , \wRegInTop_7_22[1] , 
        \wRegInTop_7_34[25] , \wRegInTop_7_41[15] , \wRegOut_7_114[3] , 
        \ScanLink171[0] , \wRegInTop_7_54[21] , \wRegInTop_7_77[10] , 
        \ScanLink83[8] , \ScanLink109[30] , \wRegOut_7_117[0] , 
        \wRegOut_5_4[20] , \wRegInBot_5_8[12] , \wRegInTop_5_14[15] , 
        \wRegInBot_5_14[12] , \ScanLink212[6] , \wRegInTop_7_99[25] , 
        \ScanLink109[29] , \wRegInBot_5_22[17] , \wRegInTop_7_21[2] , 
        \ScanLink172[3] , \wRegOut_6_4[0] , \wRegOut_7_6[12] , 
        \wRegInBot_5_11[24] , \wRegInTop_5_27[26] , \wRegInTop_6_34[5] , 
        \ScanLink146[2] , \wRegInTop_7_15[3] , \wRegInTop_5_11[23] , 
        \wRegInTop_7_89[27] , \ScanLink226[7] , \wRegInBot_5_27[21] , 
        \ScanLink94[19] , \ScanLink78[0] , \ScanLink8[26] , 
        \wRegInBot_5_28[2] , \wRegInBot_6_3[8] , \wRegOut_7_3[24] , 
        \ScanLink194[4] , \wRegInTop_7_109[1] , \wRegOut_7_123[1] , 
        \ScanLink8[15] , \wRegOut_4_0[3] , \wRegInBot_4_2[27] , 
        \wRegOut_5_14[18] , \wRegOut_6_19[30] , \wRegOut_6_19[29] , 
        \wRegOut_7_62[29] , \wRegOut_7_4[2] , \wRegOut_7_17[19] , 
        \wRegOut_7_34[31] , \wRegOut_7_62[30] , \wRegOut_7_41[18] , 
        \wRegOut_7_34[28] , \wRegInTop_6_0[30] , \wRegInBot_6_5[23] , 
        \ScanLink197[7] , \wRegOut_7_7[1] , \wRegOut_7_99[31] , 
        \wRegInTop_7_119[31] , \wRegInTop_6_0[29] , \wRegOut_6_38[1] , 
        \wRegOut_7_19[7] , \wRegOut_7_99[28] , \wRegInTop_7_119[28] , 
        \ScanLink39[19] , \wRegInTop_6_37[6] , \wRegInTop_7_12[22] , 
        \wRegInTop_7_67[12] , \ScanLink227[29] , \ScanLink252[19] , 
        \wRegInTop_7_16[0] , \wRegInTop_7_31[13] , \ScanLink145[1] , 
        \wRegInTop_7_24[27] , \wRegInTop_7_44[23] , \ScanLink204[18] , 
        \ScanLink227[30] , \wRegInTop_7_51[17] , \wRegInTop_7_72[26] , 
        \ScanLink225[4] , \wRegOut_7_120[2] , \wRegOut_7_3[17] , 
        \wRegInTop_2_0[14] , \wRegInBot_5_7[9] , \wRegInTop_5_11[10] , 
        \wRegInBot_5_27[12] , \wRegInTop_6_50[1] , \ScanLink119[18] , 
        \wRegInTop_7_71[7] , \wRegInTop_7_89[14] , \ScanLink122[6] , 
        \wRegOut_2_3[4] , \wRegOut_3_3[19] , \wRegOut_5_4[13] , 
        \wRegInTop_5_27[15] , \wRegOut_6_42[9] , \wRegInBot_5_11[17] , 
        \ScanLink242[3] , \wRegInTop_6_53[2] , \ScanLink121[5] , 
        \wRegInTop_7_51[24] , \wRegInTop_7_72[4] , \wRegInTop_7_12[11] , 
        \wRegInTop_7_24[14] , \ScanLink197[30] , \wRegInTop_7_67[21] , 
        \ScanLink197[29] , \wRegInTop_7_72[15] , \ScanLink241[0] , 
        \wRegInTop_3_5[8] , \wRegInBot_4_2[14] , \wRegOut_4_3[0] , 
        \wRegInTop_7_31[20] , \wRegInTop_7_44[10] , \wRegEnBot_5_1[0] , 
        \wRegInTop_5_3[11] , \wRegOut_5_10[8] , \wRegInBot_6_5[10] , 
        \wRegOut_6_12[16] , \wRegOut_7_69[16] , \wRegOut_6_44[17] , 
        \wRegOut_6_24[13] , \wRegOut_6_31[27] , \wRegOut_6_51[23] , 
        \ScanLink63[1] , \wRegInTop_6_4[0] , \wRegOut_6_20[3] , 
        \ScanLink112[14] , \wRegInBot_6_62[1] , \ScanLink220[9] , 
        \wRegInTop_7_4[15] , \ScanLink167[24] , \ScanLink144[15] , 
        \wRegInTop_7_82[18] , \wRegInBot_6_5[6] , \ScanLink131[25] , 
        \ScanLink151[21] , \wRegEnTop_7_40[0] , \ScanLink11[17] , 
        \wRegInBot_4_12[5] , \wRegInTop_7_112[0] , \ScanLink32[26] , 
        \wRegInTop_6_21[28] , \ScanLink107[20] , \ScanLink124[11] , 
        \ScanLink172[10] , \ScanLink191[9] , \ScanLink47[16] , 
        \wRegInBot_6_6[5] , \wRegInTop_6_7[3] , \wRegInTop_6_54[18] , 
        \wRegInTop_6_21[31] , \wRegInBot_4_9[18] , \ScanLink64[27] , 
        \wRegInTop_7_79[19] , \ScanLink239[22] , \wRegInBot_4_11[6] , 
        \ScanLink27[12] , \wRegOut_6_7[18] , \ScanLink71[13] , 
        \ScanLink189[11] , \ScanLink52[22] , \ScanLink60[2] , 
        \wRegInBot_5_30[0] , \wRegOut_5_29[22] , \wRegInTop_6_31[8] , 
        \wRegInTop_7_111[3] , \wRegOut_0_0[21] , \wRegInBot_3_1[11] , 
        \wRegOut_4_11[17] , \wRegOut_7_92[17] , \wRegInTop_7_112[17] , 
        \wRegOut_6_23[0] , \wRegInTop_7_107[23] , \wRegInBot_6_61[2] , 
        \wRegOut_7_87[23] , \wRegInTop_7_124[12] , \wRegInTop_3_0[5] , 
        \wRegInBot_3_1[3] , \ScanLink124[22] , \ScanLink139[7] , 
        \ScanLink151[12] , \wRegInBot_4_14[18] , \ScanLink107[13] , 
        \wRegInBot_3_1[22] , \wRegInTop_5_0[1] , \ScanLink172[23] , 
        \wRegInBot_5_1[7] , \ScanLink112[27] , \wRegOut_6_59[8] , 
        \ScanLink167[17] , \wRegInTop_5_3[22] , \wRegInBot_5_6[31] , 
        \wRegOut_5_15[5] , \ScanLink131[16] , \wRegInTop_7_4[26] , 
        \wRegOut_6_24[20] , \ScanLink144[26] , \wRegInBot_5_6[28] , 
        \wRegOut_6_51[10] , \ScanLink124[8] , \wRegInTop_7_77[9] , 
        \wRegOut_7_8[28] , \wRegOut_6_12[25] , \wRegOut_6_44[7] , 
        \wRegOut_7_8[31] , \wRegOut_7_65[1] , \wRegOut_7_69[25] , 
        \wRegOut_6_31[14] , \wRegInTop_5_19[1] , \wRegOut_6_44[24] , 
        \ScanLink19[9] , \wRegOut_4_11[24] , \wRegOut_5_29[11] , 
        \wRegOut_7_87[10] , \wRegInTop_7_107[10] , \wRegInTop_7_124[21] , 
        \ScanLink0[5] , \ScanLink3[6] , \ScanLink5[8] , \wRegOut_2_3[14] , 
        \wRegInTop_3_0[19] , \wRegInBot_3_2[0] , \wRegInTop_3_4[31] , 
        \wRegInTop_3_4[28] , \wRegOut_6_47[4] , \wRegOut_7_66[2] , 
        \ScanLink71[20] , \wRegOut_7_92[24] , \wRegInTop_7_112[24] , 
        \wRegInTop_3_3[6] , \ScanLink189[22] , \wRegOut_7_104[31] , 
        \ScanLink11[24] , \ScanLink27[21] , \ScanLink52[11] , 
        \wRegOut_7_127[19] , \wRegInTop_6_48[3] , \wRegInTop_7_69[5] , 
        \ScanLink32[15] , \ScanLink47[25] , \wRegOut_7_104[28] , 
        \wRegOut_5_16[6] , \wRegInBot_6_34[28] , \wRegInBot_6_41[18] , 
        \wRegInBot_6_62[30] , \wRegInBot_5_2[4] , \wRegInTop_5_3[2] , 
        \ScanLink239[11] , \ScanLink64[14] , \wRegInBot_6_17[19] , 
        \wRegInBot_6_34[31] , \wRegInBot_6_18[9] , \wRegInBot_3_5[13] , 
        \wRegOut_4_15[15] , \wRegInBot_6_62[29] , \wRegOut_6_63[2] , 
        \wRegInTop_7_103[21] , \wRegInBot_6_21[0] , \wRegOut_7_42[4] , 
        \wRegOut_7_83[21] , \wRegInTop_7_120[10] , \ScanLink15[15] , 
        \ScanLink20[0] , \ScanLink23[10] , \wRegOut_5_8[4] , 
        \wRegOut_7_96[15] , \wRegInTop_7_116[15] , \ScanLink75[11] , 
        \wRegOut_7_90[2] , \wRegOut_7_123[28] , \wRegOut_7_100[19] , 
        \ScanLink228[14] , \wRegOut_7_123[31] , \wRegOut_4_13[6] , 
        \wRegInTop_4_8[10] , \ScanLink36[24] , \ScanLink56[20] , 
        \ScanLink43[14] , \wRegInBot_6_13[31] , \wRegInBot_6_30[19] , 
        \wRegInBot_6_45[29] , \wRegInTop_5_20[8] , \ScanLink248[10] , 
        \wRegInBot_6_45[30] , \ScanLink23[3] , \wRegInBot_4_10[30] , 
        \ScanLink60[25] , \ScanLink198[27] , \wRegInBot_6_13[28] , 
        \wRegOut_4_10[5] , \wRegOut_5_31[3] , \wRegInBot_4_10[29] , 
        \ScanLink120[13] , \ScanLink155[23] , \wRegOut_6_20[11] , 
        \ScanLink103[22] , \ScanLink176[12] , \wRegOut_7_93[1] , 
        \ScanLink116[16] , \wRegInTop_7_0[17] , \ScanLink163[26] , 
        \wRegOut_6_55[21] , \ScanLink135[27] , \ScanLink140[17] , 
        \wRegInTop_7_81[9] , \wRegOut_6_60[1] , \wRegOut_7_41[7] , 
        \wRegInTop_4_8[23] , \wRegInBot_5_2[19] , \ScanLink36[17] , 
        \wRegInTop_5_7[13] , \wRegOut_6_16[14] , \wRegInBot_6_22[3] , 
        \wRegOut_6_63[24] , \wRegOut_7_18[24] , \wRegOut_7_78[20] , 
        \wRegOut_6_40[15] , \ScanLink43[27] , \ScanLink44[4] , 
        \wRegOut_6_35[25] , \wRegInTop_6_50[29] , \wRegInBot_5_14[6] , 
        \wRegInTop_6_25[19] , \ScanLink60[16] , \wRegInTop_6_50[30] , 
        \ScanLink198[14] , \ScanLink248[23] , \wRegOut_2_3[27] , 
        \ScanLink7[31] , \wRegInBot_3_5[20] , \ScanLink15[26] , 
        \ScanLink23[23] , \ScanLink56[13] , \wRegOut_6_3[30] , 
        \ScanLink75[22] , \ScanLink228[27] , \wRegInTop_7_29[7] , 
        \wRegOut_6_3[29] , \ScanLink96[2] , \wRegInBot_6_45[4] , 
        \wRegOut_7_26[0] , \wRegOut_7_96[26] , \wRegInTop_7_116[26] , 
        \wRegOut_4_15[26] , \wRegInTop_7_103[12] , \wRegInTop_5_7[20] , 
        \wRegOut_6_16[27] , \wRegOut_7_25[3] , \wRegInTop_7_34[8] , 
        \ScanLink167[9] , \wRegOut_7_83[12] , \wRegInTop_7_120[23] , 
        \ScanLink95[1] , \wRegInBot_6_46[7] , \wRegOut_7_18[17] , 
        \wRegOut_6_63[17] , \wRegOut_6_35[16] , \wRegOut_6_20[22] , 
        \wRegOut_6_40[26] , \wRegOut_7_101[9] , \wRegOut_6_55[12] , 
        \ScanLink7[28] , \wRegOut_7_78[13] , \wRegOut_3_7[31] , 
        \wRegOut_3_7[28] , \wRegInBot_4_6[25] , \wRegInTop_4_8[6] , 
        \wRegInBot_4_9[0] , \ScanLink47[7] , \ScanLink116[25] , 
        \wRegInTop_7_0[24] , \ScanLink163[15] , \wRegInTop_7_86[29] , 
        \ScanLink219[0] , \ScanLink135[14] , \wRegInBot_5_17[5] , 
        \wRegEnTop_6_45[0] , \wRegInTop_7_86[30] , \ScanLink140[24] , 
        \wRegInTop_5_28[31] , \wRegInTop_5_28[28] , \ScanLink120[20] , 
        \ScanLink179[5] , \ScanLink103[11] , \ScanLink155[10] , 
        \wRegOut_5_29[1] , \ScanLink176[21] , \wRegInBot_6_18[17] , 
        \wRegEnTop_7_18[0] , \wRegInTop_7_20[25] , \wRegInTop_7_55[15] , 
        \ScanLink193[18] , \wRegInTop_7_76[24] , \wRegInTop_6_18[10] , 
        \wRegInTop_7_16[20] , \wRegInTop_7_63[10] , \wRegOut_4_15[8] , 
        \wRegOut_6_8[25] , \ScanLink105[3] , \wRegInTop_7_35[11] , 
        \wRegInTop_7_56[2] , \wRegInTop_7_40[21] , \wRegOut_5_0[22] , 
        \ScanLink38[2] , \wRegInBot_5_9[26] , \wRegInTop_5_26[6] , 
        \wRegOut_7_59[5] , \wRegInBot_6_1[21] , \wRegInBot_6_39[2] , 
        \wRegInTop_7_84[4] , \wRegOut_7_7[26] , \wRegInTop_7_87[7] , 
        \wRegInTop_5_15[21] , \wRegInTop_5_25[5] , \ScanLink168[19] , 
        \wRegOut_7_47[9] , \wRegOut_7_88[0] , \wRegInBot_5_23[23] , 
        \wRegInBot_5_15[26] , \wRegInTop_5_23[24] , \ScanLink106[0] , 
        \wRegInTop_7_55[1] , \wRegInTop_7_98[11] , \wRegInBot_4_6[16] , 
        \wRegOut_5_10[30] , \wRegOut_5_10[29] , \wRegInBot_5_12[8] , 
        \wRegInBot_6_1[12] , \wRegInTop_6_4[18] , \wRegInTop_6_18[23] , 
        \wRegInTop_7_63[23] , \wRegInTop_7_16[13] , \ScanLink201[2] , 
        \wRegOut_5_0[11] , \ScanLink48[18] , \wRegOut_6_8[16] , 
        \ScanLink200[30] , \ScanLink223[18] , \wRegInTop_6_13[0] , 
        \wRegInTop_7_32[6] , \ScanLink161[7] , \wRegInTop_7_35[22] , 
        \wRegInTop_7_40[12] , \wRegOut_7_104[4] , \ScanLink200[29] , 
        \wRegInTop_7_55[26] , \wRegInTop_5_23[17] , \wRegInBot_6_18[24] , 
        \wRegInTop_7_20[16] , \wRegInTop_7_76[17] , \wRegOut_6_9[8] , 
        \wRegOut_7_107[7] , \wRegInBot_5_9[15] , \ScanLink41[9] , 
        \wRegInTop_5_15[12] , \wRegInBot_5_15[15] , \wRegInBot_6_40[9] , 
        \ScanLink202[1] , \wRegInTop_7_98[22] , \ScanLink90[28] , 
        \wRegEnTop_7_127[0] , \wRegInBot_5_23[10] , \wRegInTop_6_10[3] , 
        \wRegInTop_7_31[5] , \ScanLink90[31] , \ScanLink162[4] , 
        \wRegOut_7_7[15] , \ScanLink6[22] , \wRegInTop_4_11[17] , 
        \wRegInBot_5_29[25] , \ScanLink98[4] , \wRegOut_7_13[31] , 
        \wRegOut_7_13[28] , \wRegOut_7_45[30] , \wRegOut_7_66[18] , 
        \wRegOut_7_30[19] , \wRegOut_7_45[29] , \wRegOut_6_2[3] , 
        \wRegOut_7_28[6] , \wRegInBot_4_11[10] , \wRegInTop_7_87[23] , 
        \wRegInTop_7_92[17] , \wRegInBot_5_3[20] , \wRegInTop_5_29[22] , 
        \wRegOut_7_35[9] , \ScanLink214[5] , \wRegOut_7_111[3] , 
        \wRegOut_6_21[31] , \wRegOut_7_79[19] , \ScanLink6[11] , 
        \wRegInTop_3_1[20] , \ScanLink49[1] , \wRegOut_6_21[28] , 
        \wRegInTop_7_27[1] , \wRegOut_6_54[18] , \ScanLink174[0] , 
        \ScanLink217[6] , \wRegOut_4_5[27] , \wRegInBot_5_19[3] , 
        \ScanLink86[8] , \wRegOut_7_112[0] , \wRegInTop_7_24[2] , 
        \ScanLink177[3] , \wRegInTop_7_102[18] , \wRegInTop_7_121[29] , 
        \wRegInTop_7_121[30] , \ScanLink22[30] , \ScanLink22[29] , 
        \wRegInTop_4_9[30] , \wRegInBot_6_12[11] , \wRegOut_7_82[18] , 
        \wRegInBot_6_48[1] , \ScanLink249[29] , \wRegInTop_4_9[29] , 
        \wRegOut_6_1[0] , \wRegInTop_6_24[13] , \wRegInBot_6_31[20] , 
        \wRegInTop_6_51[23] , \ScanLink249[30] , \ScanLink57[19] , 
        \wRegInBot_6_44[10] , \wRegOut_7_114[14] , \wRegOut_6_2[23] , 
        \ScanLink74[31] , \wRegInBot_6_24[14] , \wRegInTop_6_44[17] , 
        \wRegInBot_6_51[24] , \wRegOut_7_101[20] , \ScanLink74[28] , 
        \wRegInTop_6_31[27] , \wRegInTop_7_69[16] , \wRegOut_7_122[11] , 
        \wRegInTop_6_12[16] , \wRegOut_3_6[6] , \wRegInBot_4_1[8] , 
        \wRegEnBot_4_11[0] , \wRegInBot_5_3[13] , \wRegInBot_6_32[9] , 
        \wRegInTop_5_6[19] , \ScanLink110[4] , \wRegInTop_6_62[3] , 
        \wRegInTop_7_43[5] , \wRegInBot_4_11[23] , \wRegInTop_4_11[24] , 
        \wRegInTop_4_12[7] , \ScanLink33[9] , \ScanLink102[28] , 
        \ScanLink154[30] , \ScanLink177[18] , \wRegInTop_7_92[24] , 
        \wRegOut_5_21[9] , \wRegInTop_5_29[11] , \ScanLink154[29] , 
        \wRegInBot_5_29[16] , \ScanLink102[31] , \ScanLink121[19] , 
        \wRegInTop_7_91[3] , \wRegOut_5_6[2] , \wRegInTop_7_87[10] , 
        \wRegOut_6_2[10] , \wRegOut_7_101[13] , \wRegInTop_6_31[14] , 
        \wRegInBot_6_51[17] , \wRegOut_0_0[31] , \wRegOut_0_0[28] , 
        \wRegInBot_1_0[9] , \wRegInBot_1_0[0] , \wRegOut_1_1[15] , 
        \wRegInTop_1_1[6] , \wRegInBot_2_0[16] , \wRegInTop_2_3[9] , 
        \wRegOut_3_5[5] , \wRegInBot_6_24[27] , \wRegInTop_6_44[24] , 
        \wRegInTop_7_69[25] , \wRegOut_7_122[22] , \wRegOut_7_80[8] , 
        \wRegInTop_4_11[4] , \wRegInTop_5_30[2] , \wRegInTop_6_12[25] , 
        \wRegInTop_3_1[13] , \wRegInBot_3_4[19] , \wRegOut_4_5[14] , 
        \wRegOut_5_5[1] , \wRegInBot_6_12[22] , \wRegInTop_6_24[20] , 
        \wRegInBot_6_31[13] , \wRegInBot_6_44[23] , \wRegInTop_6_51[10] , 
        \wRegInTop_7_92[0] , \wRegOut_7_114[27] , \ScanLink113[7] , 
        \wRegInTop_6_61[0] , \wRegInTop_7_40[6] , \ScanLink51[3] , 
        \wRegOut_7_72[26] , \ScanLink84[16] , \wRegInTop_7_2[1] , 
        \wRegOut_7_24[27] , \wRegOut_7_31[13] , \wRegOut_7_51[17] , 
        \wRegInTop_7_120[2] , \wRegOut_7_44[23] , \wRegOut_7_12[22] , 
        \wRegOut_7_33[7] , \wRegOut_7_67[12] , \wRegOut_3_6[11] , 
        \ScanLink29[16] , \wRegInTop_5_14[18] , \wRegOut_6_12[1] , 
        \ScanLink83[5] , \ScanLink109[24] , \wRegInTop_7_99[28] , 
        \wRegInBot_6_50[3] , \ScanLink169[20] , \wRegInTop_7_99[31] , 
        \ScanLink91[22] , \wRegOut_6_11[2] , \ScanLink80[6] , 
        \wRegInTop_7_41[18] , \wRegInTop_7_62[30] , \wRegInTop_6_19[30] , 
        \wRegInTop_6_19[29] , \wRegOut_7_30[4] , \wRegInTop_7_34[28] , 
        \wRegInTop_7_62[29] , \ScanLink201[23] , \ScanLink211[8] , 
        \wRegInTop_4_2[16] , \wRegInBot_6_53[0] , \wRegInTop_7_17[19] , 
        \wRegInTop_7_34[31] , \ScanLink187[15] , \ScanLink222[12] , 
        \ScanLink192[21] , \ScanLink242[16] , \ScanLink237[26] , 
        \ScanLink49[12] , \ScanLink214[17] , \ScanLink52[0] , 
        \wRegOut_7_109[1] , \wRegInTop_7_123[1] , \wRegInBot_6_0[18] , 
        \ScanLink2[20] , \wRegOut_1_1[26] , \wRegInBot_2_0[25] , 
        \ScanLink28[8] , \wRegOut_5_11[23] , \wRegOut_7_89[27] , 
        \wRegInTop_7_109[27] , \wRegOut_5_27[26] , \wRegInTop_6_5[12] , 
        \wRegInTop_7_1[2] , \wRegInBot_5_22[30] , \wRegInBot_5_22[29] , 
        \wRegInTop_5_28[0] , \ScanLink91[11] , \wRegInBot_6_34[7] , 
        \wRegOut_7_57[3] , \ScanLink169[13] , \ScanLink109[17] , 
        \wRegOut_3_0[8] , \wRegOut_5_1[31] , \wRegOut_5_1[28] , 
        \ScanLink84[25] , \ScanLink35[7] , \wRegEnTop_6_37[0] , 
        \wRegOut_7_44[10] , \wRegOut_5_27[7] , \wRegOut_7_31[20] , 
        \wRegInBot_4_4[5] , \wRegInTop_4_6[0] , \wRegInBot_4_7[6] , 
        \wRegInBot_6_29[8] , \wRegOut_7_12[11] , \wRegOut_7_67[21] , 
        \wRegOut_7_85[5] , \wRegInTop_4_14[9] , \wRegOut_7_72[15] , 
        \wRegOut_7_24[14] , \wRegOut_7_51[24] , \wRegInTop_7_58[4] , 
        \wRegInTop_4_5[3] , \wRegOut_7_86[6] , \ScanLink36[4] , 
        \wRegOut_5_24[4] , \wRegInTop_6_5[21] , \wRegOut_5_27[15] , 
        \wRegInBot_3_0[31] , \wRegOut_3_2[20] , \wRegOut_3_2[13] , 
        \ScanLink12[2] , \wRegOut_3_6[22] , \wRegInTop_4_2[25] , 
        \wRegOut_5_11[10] , \ScanLink108[6] , \ScanLink49[21] , 
        \wRegInBot_6_37[4] , \wRegOut_7_54[0] , \ScanLink192[12] , 
        \wRegOut_7_89[14] , \wRegInTop_7_109[14] , \ScanLink237[15] , 
        \ScanLink242[25] , \ScanLink214[24] , \ScanLink29[25] , 
        \ScanLink115[9] , \wRegInTop_7_46[8] , \ScanLink201[10] , 
        \wRegInTop_7_89[1] , \wRegOut_5_23[24] , \wRegInTop_6_1[10] , 
        \ScanLink187[26] , \ScanLink222[21] , \wRegOut_7_98[11] , 
        \wRegInTop_7_118[11] , \wRegInTop_4_6[14] , \ScanLink38[20] , 
        \wRegOut_5_15[21] , \wCtrlOut_5[0] , \wRegInTop_6_43[8] , 
        \ScanLink196[23] , \ScanLink246[14] , \ScanLink233[24] , 
        \wRegInTop_5_8[9] , \ScanLink58[24] , \ScanLink210[15] , 
        \wRegOut_6_51[0] , \wRegOut_7_70[6] , \ScanLink205[21] , 
        \ScanLink253[20] , \ScanLink11[1] , \wRegOut_5_5[19] , 
        \wRegInBot_5_26[18] , \wRegInBot_6_13[2] , \ScanLink183[17] , 
        \ScanLink226[10] , \ScanLink80[14] , \ScanLink95[20] , 
        \ScanLink118[12] , \ScanLink252[9] , \wRegOut_7_73[5] , 
        \wRegInTop_5_9[17] , \wRegInBot_6_10[1] , \wRegOut_6_52[3] , 
        \ScanLink178[16] , \wRegOut_7_35[11] , \wRegInTop_5_11[9] , 
        \wRegOut_7_40[21] , \wRegOut_6_18[10] , \wRegOut_7_16[20] , 
        \wRegOut_7_63[10] , \wRegEnTop_7_32[0] , \wRegOut_7_76[24] , 
        \ScanLink58[17] , \wRegOut_7_20[25] , \wRegOut_7_55[15] , 
        \wRegInTop_7_13[31] , \wRegInTop_7_30[19] , \wRegInTop_7_13[28] , 
        \wRegInTop_7_45[29] , \ScanLink205[12] , \wRegInTop_4_6[27] , 
        \ScanLink38[13] , \wRegOut_6_35[4] , \wRegInTop_7_45[30] , 
        \ScanLink183[24] , \ScanLink226[23] , \wRegInTop_7_66[18] , 
        \ScanLink253[13] , \wRegOut_7_14[2] , \ScanLink196[10] , 
        \ScanLink210[26] , \ScanLink233[17] , \ScanLink246[27] , 
        \wRegInBot_4_8[21] , \wRegInTop_5_9[24] , \wRegOut_5_15[12] , 
        \wRegInBot_6_4[30] , \wRegInBot_6_4[29] , \ScanLink148[4] , 
        \wRegOut_5_23[17] , \wRegInTop_6_1[23] , \wRegOut_7_98[22] , 
        \ScanLink228[1] , \wRegInTop_7_118[22] , \wRegInBot_5_25[7] , 
        \wRegInBot_5_26[4] , \ScanLink76[6] , \ScanLink75[5] , 
        \wRegInTop_6_39[0] , \wRegOut_7_76[17] , \wRegInTop_7_107[7] , 
        \wRegInTop_7_18[6] , \wRegOut_7_55[26] , \wRegOut_7_20[16] , 
        \wRegOut_7_40[12] , \wRegOut_7_35[22] , \wRegInTop_7_104[4] , 
        \wRegInTop_5_10[30] , \ScanLink80[27] , \wRegOut_6_18[23] , 
        \wRegOut_7_63[23] , \wRegOut_7_16[13] , \wRegOut_7_9[7] , 
        \ScanLink156[8] , \ScanLink178[25] , \ScanLink199[1] , 
        \wRegInTop_5_10[29] , \wRegEnTop_5_26[0] , \ScanLink95[13] , 
        \wRegOut_6_36[7] , \ScanLink118[21] , \wRegOut_7_17[1] , 
        \wRegOut_6_6[21] , \wRegInBot_6_20[16] , \wRegInTop_6_40[15] , 
        \wRegInTop_6_58[9] , \wRegInBot_6_55[26] , \ScanLink188[31] , 
        \wRegInTop_6_35[25] , \wRegOut_7_105[22] , \wRegInTop_5_14[4] , 
        \wRegInTop_7_18[24] , \ScanLink188[28] , \wRegInTop_6_16[14] , 
        \wRegInTop_6_63[24] , \wRegOut_7_126[13] , \wRegInBot_6_16[13] , 
        \wRegInTop_6_20[11] , \wRegInBot_6_35[22] , \wRegInTop_6_55[21] , 
        \wRegInBot_6_63[23] , \wRegInTop_7_78[20] , \wRegInBot_6_40[12] , 
        \wRegOut_7_110[16] , \wRegInTop_6_45[6] , \ScanLink137[1] , 
        \wRegInTop_7_64[0] , \wRegInBot_3_0[28] , \wRegInTop_3_5[22] , 
        \wRegOut_4_1[25] , \wRegOut_7_76[8] , \wRegInBot_5_7[22] , 
        \ScanLink2[13] , \wRegInTop_3_5[11] , \wRegInTop_4_15[15] , 
        \wRegInBot_4_15[12] , \wRegInTop_5_2[31] , \wRegInTop_5_2[28] , 
        \wRegEnBot_5_14[0] , \wRegInTop_6_46[5] , \wRegInTop_7_67[3] , 
        \ScanLink134[2] , \wRegOut_7_9[22] , \wRegOut_5_18[0] , 
        \ScanLink254[7] , \wRegInTop_5_17[7] , \wRegInTop_7_96[15] , 
        \ScanLink106[19] , \ScanLink125[31] , \wRegOut_6_49[2] , 
        \ScanLink125[28] , \ScanLink173[29] , \ScanLink150[18] , 
        \ScanLink173[30] , \wRegOut_7_68[4] , \ScanLink249[8] , 
        \wRegOut_5_28[31] , \wRegInTop_7_83[21] , \wRegOut_5_28[28] , 
        \wRegInTop_6_21[2] , \ScanLink153[5] , \wRegOut_4_1[16] , 
        \wRegOut_7_86[30] , \wRegInTop_7_106[30] , \wRegInTop_7_125[18] , 
        \wRegInBot_4_8[12] , \ScanLink26[18] , \wRegInBot_6_16[20] , 
        \wRegInBot_6_63[10] , \wRegInTop_7_78[13] , \wRegOut_7_86[29] , 
        \ScanLink233[0] , \wRegInTop_7_106[29] , \ScanLink238[28] , 
        \wRegInTop_6_20[22] , \ScanLink181[3] , \wRegInBot_6_35[11] , 
        \wRegInBot_6_40[21] , \wRegInTop_6_55[12] , \wRegOut_7_110[25] , 
        \ScanLink238[31] , \ScanLink53[28] , \wRegOut_6_6[12] , 
        \wRegInBot_6_55[15] , \wRegOut_7_105[11] , \ScanLink70[8] , 
        \wRegInBot_6_20[25] , \wRegInTop_6_35[16] , \ScanLink70[19] , 
        \wRegInTop_6_16[27] , \wRegInTop_6_40[26] , \wRegInTop_7_101[9] , 
        \wRegOut_7_126[20] , \wRegInTop_7_18[17] , \wRegInTop_4_15[26] , 
        \ScanLink53[31] , \wRegInTop_6_63[17] , \ScanLink182[0] , 
        \wRegInBot_4_15[21] , \wRegInTop_7_83[12] , \wRegInBot_5_23[9] , 
        \wRegInTop_7_96[26] , \wRegInBot_6_8[3] , \wRegInTop_6_9[5] , 
        \ScanLink150[6] , \wRegInTop_6_22[1] , \wRegOut_3_0[1] , 
        \ScanLink28[1] , \wRegOut_5_1[21] , \wRegInBot_5_7[11] , 
        \wRegOut_6_30[9] , \wRegOut_6_50[30] , \ScanLink230[3] , 
        \wRegInBot_5_14[25] , \wRegOut_6_25[19] , \wRegOut_6_50[29] , 
        \wRegOut_7_9[11] , \wRegInTop_7_99[12] , \wRegInTop_5_28[9] , 
        \wRegInTop_5_22[27] , \ScanLink116[3] , \wRegInTop_7_45[2] , 
        \wRegInBot_5_22[20] , \wRegInTop_4_14[0] , \wRegInBot_5_8[25] , 
        \wRegInTop_5_14[22] , \ScanLink91[18] , \wRegOut_7_98[3] , 
        \wRegOut_5_0[5] , \wRegOut_7_6[25] , \wRegInTop_7_97[4] , 
        \wRegOut_7_31[29] , \wRegOut_7_44[19] , \wRegOut_7_67[31] , 
        \wRegOut_7_67[28] , \wRegOut_3_3[2] , \wRegInTop_4_6[9] , 
        \wRegInBot_6_29[1] , \wRegOut_7_12[18] , \wRegOut_7_31[30] , 
        \wRegOut_5_3[6] , \wRegOut_5_11[19] , \wRegInBot_6_0[22] , 
        \wRegInTop_7_94[7] , \wRegOut_7_49[6] , \wRegOut_3_6[18] , 
        \wRegEnTop_4_0[0] , \wRegInBot_4_7[26] , \wRegInTop_6_5[31] , 
        \wRegInTop_6_5[28] , \wRegOut_6_9[26] , \ScanLink115[0] , 
        \wRegInTop_7_34[12] , \wRegInTop_7_46[1] , \ScanLink201[19] , 
        \wRegInTop_7_41[22] , \wRegInTop_7_89[8] , \ScanLink222[31] , 
        \wRegInTop_7_17[23] , \wRegOut_5_1[12] , \wRegInBot_5_8[16] , 
        \ScanLink49[31] , \wRegInTop_6_19[13] , \wRegInTop_7_62[13] , 
        \ScanLink222[28] , \wRegOut_7_54[9] , \ScanLink49[28] , 
        \wRegInBot_6_19[14] , \wRegInTop_7_77[27] , \wRegInTop_7_2[8] , 
        \wRegInTop_7_21[26] , \wRegInTop_7_54[16] , \wRegInTop_5_14[11] , 
        \wRegInBot_5_22[13] , \wRegOut_6_4[4] , \wRegOut_7_6[16] , 
        \wRegInTop_7_21[6] , \ScanLink169[30] , \ScanLink172[7] , 
        \ScanLink169[29] , \wRegInBot_5_14[16] , \wRegOut_6_12[8] , 
        \ScanLink212[2] , \wRegInTop_7_99[21] , \wRegInTop_5_22[14] , 
        \wRegOut_6_9[15] , \wRegInBot_6_19[27] , \ScanLink192[28] , 
        \wRegInTop_7_77[14] , \wRegOut_7_117[4] , \wRegInTop_7_21[15] , 
        \wRegInTop_7_22[5] , \ScanLink171[4] , \wRegInTop_7_54[25] , 
        \ScanLink192[31] , \wRegInTop_6_19[20] , \wRegInTop_7_34[21] , 
        \wRegInTop_7_41[11] , \wRegOut_7_114[7] , \wRegInTop_7_62[20] , 
        \wRegInBot_6_53[9] , \ScanLink211[1] , \wRegInBot_4_7[15] , 
        \ScanLink52[9] , \wRegInTop_7_17[10] , \ScanLink2[30] , 
        \ScanLink2[29] , \wRegInTop_2_0[3] , \wRegOut_2_2[17] , 
        \ScanLink6[18] , \wRegInTop_5_6[10] , \wRegInBot_6_0[11] , 
        \wRegOut_6_7[7] , \wRegOut_7_109[8] , \wRegInTop_7_123[8] , 
        \wRegOut_6_17[17] , \wRegOut_6_34[26] , \wRegOut_6_41[16] , 
        \wRegOut_6_62[27] , \wRegOut_7_19[27] , \wRegInBot_6_32[0] , 
        \wRegOut_7_51[4] , \wRegOut_6_21[12] , \wRegOut_6_54[22] , 
        \wRegOut_7_79[23] , \ScanLink134[24] , \ScanLink141[14] , 
        \wRegInBot_2_1[5] , \ScanLink117[15] , \wRegInTop_7_1[14] , 
        \ScanLink162[25] , \wRegOut_2_2[24] , \wRegInBot_2_2[6] , 
        \wRegInTop_2_3[0] , \wRegInTop_4_0[7] , \wRegInBot_4_1[1] , 
        \wRegInTop_7_87[19] , \ScanLink177[11] , \wRegOut_7_83[2] , 
        \ScanLink33[0] , \wRegInTop_5_29[18] , \ScanLink102[21] , 
        \wRegOut_5_21[0] , \wRegInTop_6_24[30] , \ScanLink121[10] , 
        \ScanLink154[20] , \ScanLink249[13] , \ScanLink14[16] , 
        \wRegOut_5_5[8] , \wRegInBot_3_4[10] , \wRegInBot_4_2[2] , 
        \ScanLink22[13] , \wRegInTop_4_9[13] , \ScanLink37[27] , 
        \ScanLink61[26] , \ScanLink199[24] , \wRegInTop_6_24[29] , 
        \ScanLink42[17] , \wRegInTop_6_51[19] , \wRegInTop_7_92[9] , 
        \wRegOut_5_22[3] , \wRegOut_6_2[19] , \ScanLink30[3] , 
        \ScanLink57[23] , \wRegInTop_4_3[4] , \wRegOut_7_80[1] , 
        \wRegOut_4_14[16] , \ScanLink74[12] , \wRegInTop_6_61[9] , 
        \wRegOut_7_97[16] , \ScanLink229[17] , \wRegInTop_7_117[16] , 
        \wRegInTop_7_102[22] , \wRegInTop_7_121[13] , \wRegOut_7_52[7] , 
        \wRegInBot_4_11[19] , \wRegInBot_6_31[3] , \wRegOut_7_82[22] , 
        \ScanLink102[12] , \wRegInBot_5_3[29] , \ScanLink57[4] , 
        \ScanLink121[23] , \ScanLink169[6] , \ScanLink177[22] , 
        \wRegInTop_7_4[6] , \ScanLink154[13] , \ScanLink134[17] , 
        \ScanLink117[26] , \ScanLink141[27] , \wRegInTop_7_126[5] , 
        \wRegInTop_7_1[27] , \ScanLink162[16] , \ScanLink209[3] , 
        \wRegInBot_3_0[21] , \wRegInBot_3_0[12] , \ScanLink8[4] , 
        \wRegInTop_3_1[30] , \wRegInBot_3_4[23] , \wRegInBot_5_3[30] , 
        \wRegOut_6_21[21] , \wRegOut_7_79[10] , \wRegInTop_7_27[8] , 
        \wRegInTop_5_6[23] , \ScanLink85[2] , \wRegOut_6_54[11] , 
        \ScanLink174[9] , \wRegOut_6_34[15] , \wRegOut_6_41[25] , 
        \wRegOut_6_14[6] , \wRegOut_7_35[0] , \wRegOut_6_17[24] , 
        \wRegInBot_6_56[4] , \wRegOut_7_19[14] , \wRegOut_6_62[14] , 
        \wRegInTop_7_121[20] , \wRegOut_4_14[25] , \wRegInTop_7_102[11] , 
        \wRegOut_7_36[3] , \wRegOut_7_82[11] , \wRegOut_6_17[5] , 
        \wRegInTop_3_1[29] , \ScanLink49[8] , \wRegInBot_6_55[7] , 
        \wRegOut_7_97[25] , \wRegInTop_7_117[25] , \ScanLink86[1] , 
        \ScanLink14[25] , \ScanLink22[20] , \ScanLink57[10] , 
        \wRegOut_7_112[9] , \wRegInTop_6_18[2] , \wRegInTop_7_39[4] , 
        \wRegOut_7_101[29] , \ScanLink61[15] , \ScanLink74[21] , 
        \wRegInTop_7_7[5] , \wRegInBot_6_12[18] , \ScanLink199[17] , 
        \wRegOut_7_101[30] , \ScanLink229[24] , \wRegOut_7_122[18] , 
        \wRegInBot_6_31[30] , \wRegInBot_6_48[8] , \ScanLink249[20] , 
        \wRegInTop_4_9[20] , \ScanLink37[14] , \ScanLink42[24] , 
        \ScanLink54[7] , \wRegEnTop_6_56[0] , \wRegOut_6_1[9] , 
        \wRegInBot_6_31[29] , \wRegInTop_7_125[6] , \wRegInBot_6_44[19] , 
        \wRegOut_4_10[14] , \wRegInTop_7_125[11] , \wRegOut_6_33[3] , 
        \wRegInTop_7_106[20] , \wRegOut_7_12[5] , \ScanLink233[9] , 
        \ScanLink10[27] , \ScanLink10[14] , \wRegInTop_3_5[18] , 
        \wRegOut_5_28[21] , \wRegOut_7_86[20] , \wRegOut_7_93[14] , 
        \wRegInTop_7_113[14] , \ScanLink26[11] , \wRegOut_7_126[30] , 
        \wRegInBot_5_20[3] , \ScanLink53[21] , \ScanLink70[1] , 
        \wRegEnTop_7_53[0] , \wRegOut_7_105[18] , \ScanLink70[10] , 
        \wRegInTop_7_101[0] , \wRegOut_7_126[29] , \wRegInBot_6_63[19] , 
        \ScanLink188[12] , \wRegInBot_4_15[31] , \wRegInBot_4_15[28] , 
        \ScanLink33[25] , \ScanLink65[24] , \wRegInBot_6_40[31] , 
        \ScanLink238[21] , \wRegInBot_6_16[29] , \ScanLink46[15] , 
        \wRegInBot_6_35[18] , \wRegInBot_6_40[28] , \wRegInBot_6_16[30] , 
        \ScanLink106[23] , \ScanLink173[13] , \wRegInTop_5_2[12] , 
        \wRegInBot_5_7[18] , \wRegInBot_5_23[0] , \ScanLink73[2] , 
        \ScanLink150[22] , \wRegOut_6_30[0] , \ScanLink113[17] , 
        \ScanLink125[12] , \wRegInTop_7_102[3] , \ScanLink130[26] , 
        \ScanLink145[16] , \ScanLink182[9] , \wRegInTop_7_5[16] , 
        \ScanLink166[27] , \wRegOut_7_11[6] , \wRegOut_6_25[10] , 
        \wRegOut_6_50[20] , \wRegOut_7_9[18] , \ScanLink65[17] , 
        \wRegOut_6_13[15] , \wRegInTop_6_22[8] , \wRegOut_6_45[14] , 
        \wRegOut_6_30[24] , \wRegOut_7_68[15] , \wRegInTop_6_55[31] , 
        \ScanLink238[12] , \ScanLink14[5] , \wRegInTop_7_78[29] , 
        \wRegOut_4_8[2] , \wRegInBot_4_8[31] , \ScanLink33[16] , 
        \ScanLink46[26] , \wRegInTop_6_55[28] , \wRegInTop_6_20[18] , 
        \wRegInTop_7_78[30] , \wRegInBot_4_8[28] , \ScanLink26[22] , 
        \ScanLink53[12] , \wRegInTop_6_58[0] , \wRegInTop_7_79[6] , 
        \wRegOut_6_6[28] , \wRegOut_5_28[12] , \wRegOut_6_6[31] , 
        \ScanLink70[23] , \ScanLink188[21] , \wRegInBot_6_15[5] , 
        \wRegOut_6_57[7] , \wRegOut_7_76[1] , \wRegOut_7_93[27] , 
        \wRegInTop_7_113[27] , \ScanLink137[8] , \wRegInTop_7_64[9] , 
        \wRegInTop_7_125[22] , \wRegOut_4_10[27] , \wRegInTop_5_2[21] , 
        \wRegOut_5_18[9] , \wRegOut_7_86[13] , \wRegInTop_7_106[13] , 
        \wRegOut_6_30[17] , \wRegOut_6_45[27] , \wRegOut_6_13[26] , 
        \wRegOut_6_54[4] , \wRegOut_7_68[26] , \wRegOut_7_75[2] , 
        \wRegInBot_6_16[6] , \wRegOut_6_25[23] , \wRegInTop_2_1[24] , 
        \ScanLink9[25] , \wRegOut_3_2[30] , \ScanLink17[6] , 
        \wRegOut_6_50[13] , \ScanLink130[15] , \wRegInTop_7_83[31] , 
        \wRegInTop_6_27[5] , \ScanLink106[10] , \ScanLink113[24] , 
        \ScanLink145[25] , \ScanLink249[1] , \wRegInTop_7_5[25] , 
        \ScanLink166[14] , \wRegInTop_7_83[28] , \ScanLink125[21] , 
        \ScanLink173[20] , \ScanLink129[4] , \ScanLink150[11] , 
        \wRegInTop_7_25[24] , \ScanLink196[19] , \wRegInTop_7_73[25] , 
        \ScanLink235[7] , \wRegInTop_7_50[14] , \wRegOut_3_2[29] , 
        \wRegInBot_4_3[24] , \wRegInTop_7_13[21] , \ScanLink155[2] , 
        \wRegInTop_7_30[10] , \wRegInTop_7_45[20] , \wRegInBot_6_4[20] , 
        \wRegOut_6_28[2] , \wRegInTop_7_66[11] , \ScanLink187[4] , 
        \ScanLink228[8] , \wRegInBot_5_26[22] , \wRegInTop_6_39[9] , 
        \ScanLink184[7] , \wRegOut_7_2[27] , \ScanLink68[3] , 
        \ScanLink118[31] , \wRegInTop_2_1[17] , \wRegInBot_4_3[17] , 
        \wRegOut_5_5[23] , \wRegInTop_5_10[20] , \ScanLink118[28] , 
        \wRegInTop_7_119[2] , \wRegOut_7_17[8] , \wRegInTop_7_88[24] , 
        \ScanLink236[4] , \wRegInBot_5_10[27] , \wRegInTop_5_8[0] , 
        \wRegInTop_5_12[3] , \wRegOut_5_15[31] , \wRegInTop_5_26[25] , 
        \wRegInTop_6_24[6] , \ScanLink156[1] , \ScanLink199[8] , 
        \wRegInBot_6_4[13] , \wRegOut_5_15[28] , \wRegOut_7_98[18] , 
        \wRegInTop_7_118[18] , \wRegInTop_6_1[19] , \wRegOut_6_51[9] , 
        \wRegInTop_7_30[23] , \wRegInTop_7_45[13] , \ScanLink253[30] , 
        \wRegInTop_7_66[22] , \ScanLink205[28] , \wRegInBot_5_9[6] , 
        \ScanLink251[3] , \ScanLink253[29] , \wRegOut_5_5[10] , 
        \ScanLink38[30] , \wRegInTop_7_13[12] , \ScanLink205[31] , 
        \ScanLink226[19] , \ScanLink38[29] , \ScanLink131[6] , 
        \wRegInTop_7_73[16] , \wRegInTop_7_62[7] , \wRegInTop_6_43[1] , 
        \wRegInTop_7_50[27] , \wRegInTop_7_25[17] , \wRegInBot_5_10[14] , 
        \wRegInBot_6_10[8] , \ScanLink252[0] , \wRegInTop_5_26[16] , 
        \wRegInBot_5_26[11] , \ScanLink95[30] , \wRegInTop_6_40[2] , 
        \wRegInTop_7_61[4] , \ScanLink132[5] , \ScanLink9[16] , 
        \wRegInTop_5_10[13] , \ScanLink95[29] , \wRegInTop_7_88[17] , 
        \ScanLink11[8] , \wRegOut_7_2[14] , \wRegInTop_4_14[16] , 
        \wRegInTop_5_0[8] , \wRegInTop_5_11[0] , \wRegOut_7_16[30] , 
        \wRegOut_7_16[29] , \wRegOut_7_35[18] , \wRegOut_7_40[28] , 
        \wRegOut_6_18[19] , \wRegOut_7_40[31] , \wRegOut_7_63[19] , 
        \wRegOut_7_78[7] , \wRegOut_6_59[1] , \wRegInTop_7_82[22] , 
        \wRegInTop_7_97[16] , \ScanLink3[23] , \wRegEnBot_3_4[0] , 
        \wRegOut_4_6[4] , \wRegInBot_4_14[11] , \wRegInBot_5_6[21] , 
        \wRegOut_6_24[29] , \wRegOut_7_65[8] , \wRegInTop_7_77[0] , 
        \ScanLink244[4] , \wRegOut_6_51[19] , \wRegInTop_6_56[6] , 
        \ScanLink124[1] , \wRegOut_7_8[21] , \wRegOut_6_24[30] , 
        \ScanLink3[10] , \wRegInBot_3_2[9] , \wRegInTop_3_4[21] , 
        \ScanLink19[0] , \wRegOut_5_29[18] , \wRegOut_4_0[26] , 
        \wRegInTop_5_19[8] , \ScanLink247[7] , \wRegInTop_7_107[19] , 
        \wRegOut_4_5[7] , \wRegInBot_4_9[22] , \ScanLink71[29] , 
        \wRegInBot_6_17[10] , \wRegInTop_6_21[12] , \wRegInBot_6_34[21] , 
        \wRegInTop_6_54[22] , \wRegInTop_6_55[5] , \ScanLink127[2] , 
        \wRegOut_7_87[19] , \wRegInTop_7_124[31] , \wRegInTop_7_74[3] , 
        \wRegInTop_7_124[28] , \wRegInBot_6_41[11] , \wRegOut_7_111[15] , 
        \ScanLink239[18] , \wRegInBot_6_18[0] , \wRegInBot_6_62[20] , 
        \wRegInTop_7_79[23] , \wRegInTop_7_19[27] , \ScanLink27[31] , 
        \wRegInTop_6_62[27] , \wRegOut_7_127[10] , \ScanLink27[28] , 
        \ScanLink52[18] , \wRegInTop_6_17[17] , \wRegOut_6_7[22] , 
        \ScanLink71[30] , \wRegInBot_6_21[15] , \wRegInTop_6_41[16] , 
        \wRegInBot_6_54[25] , \wRegInTop_6_34[26] , \wRegOut_7_104[21] , 
        \wRegOut_7_8[12] , \wRegOut_7_125[6] , \wRegInBot_4_14[22] , 
        \wRegInTop_5_3[18] , \wRegInBot_5_6[12] , \ScanLink220[0] , 
        \wRegInTop_6_32[2] , \wRegInBot_6_62[8] , \ScanLink140[5] , 
        \ScanLink63[8] , \wRegInTop_7_13[4] , \ScanLink107[30] , 
        \wRegOut_7_2[5] , \ScanLink151[28] , \wRegInTop_7_112[9] , 
        \ScanLink124[18] , \ScanLink107[29] , \ScanLink151[31] , 
        \ScanLink172[19] , \wRegInTop_7_97[25] , \wRegInBot_0_0[6] , 
        \wRegOut_1_1[2] , \wRegInBot_4_9[11] , \wRegInTop_4_14[25] , 
        \wRegInTop_6_4[9] , \wRegInTop_7_82[11] , \wRegInTop_6_17[24] , 
        \ScanLink192[3] , \wRegOut_7_127[23] , \wRegInBot_5_30[9] , 
        \wRegOut_6_7[11] , \wRegInBot_6_54[16] , \wRegInTop_6_62[14] , 
        \wRegInTop_7_19[14] , \ScanLink189[18] , \wRegOut_7_104[12] , 
        \wRegInBot_6_21[26] , \wRegInTop_6_34[15] , \wRegOut_7_1[6] , 
        \wRegInTop_6_41[25] , \wRegEnTop_6_2[0] , \wRegInTop_6_21[21] , 
        \ScanLink191[0] , \wRegInBot_6_41[22] , \wRegInTop_6_54[11] , 
        \wRegOut_7_111[26] , \wRegInBot_3_1[18] , \wRegOut_4_0[15] , 
        \wRegInBot_6_17[23] , \wRegInBot_6_34[12] , \wRegInBot_6_62[13] , 
        \wRegInTop_7_79[10] , \wRegOut_3_3[10] , \wRegInTop_3_4[12] , 
        \wRegOut_6_23[9] , \ScanLink223[3] , \wRegInTop_6_31[1] , 
        \wRegOut_7_126[5] , \wRegInTop_7_10[7] , \ScanLink143[6] , 
        \wRegInTop_3_6[2] , \wRegInBot_3_7[4] , \wRegInTop_5_6[6] , 
        \wRegOut_5_13[2] , \wRegOut_7_21[26] , \wRegOut_7_54[16] , 
        \wRegInBot_5_7[0] , \wRegOut_7_77[27] , \wRegOut_7_17[23] , 
        \wRegOut_7_62[13] , \wRegInTop_5_8[14] , \wRegOut_6_19[13] , 
        \wRegOut_7_34[12] , \wRegInTop_5_11[19] , \ScanLink81[17] , 
        \wRegOut_7_41[22] , \ScanLink94[23] , \wRegOut_6_42[0] , 
        \wRegOut_7_63[6] , \ScanLink179[15] , \wRegOut_6_41[3] , 
        \wRegInTop_6_50[8] , \ScanLink119[11] , \wRegOut_7_60[5] , 
        \wRegInTop_7_67[28] , \ScanLink252[23] , \ScanLink241[9] , 
        \wRegInTop_7_12[18] , \wRegInBot_3_4[7] , \wRegInTop_4_7[17] , 
        \ScanLink39[23] , \ScanLink59[27] , \wRegInTop_7_31[30] , 
        \wRegInTop_7_44[19] , \ScanLink182[14] , \ScanLink227[13] , 
        \wRegInTop_7_67[31] , \wRegInTop_7_31[29] , \ScanLink204[22] , 
        \wRegInBot_5_4[3] , \wRegInTop_5_5[5] , \ScanLink197[20] , 
        \ScanLink211[16] , \ScanLink232[27] , \ScanLink247[17] , 
        \wRegOut_5_10[1] , \wRegOut_5_14[22] , \wRegEnTop_7_21[0] , 
        \wRegOut_5_22[27] , \wRegInBot_6_5[19] , \wRegInTop_6_0[13] , 
        \wRegOut_7_99[12] , \wRegInTop_3_5[1] , \wRegOut_4_3[9] , 
        \wRegInTop_7_119[12] , \wRegInBot_4_14[2] , \wRegOut_5_4[30] , 
        \wRegInBot_5_27[31] , \ScanLink119[22] , \wRegInBot_5_27[28] , 
        \ScanLink78[9] , \wRegOut_6_26[4] , \ScanLink94[10] , \ScanLink189[2] , 
        \wRegInTop_7_109[8] , \wRegOut_7_123[8] , \wRegOut_5_4[29] , 
        \ScanLink65[6] , \ScanLink81[24] , \wRegOut_6_19[20] , 
        \ScanLink179[26] , \wRegOut_7_62[20] , \wRegOut_7_17[10] , 
        \wRegOut_7_41[11] , \wRegInTop_7_114[7] , \wRegInTop_5_8[27] , 
        \wRegOut_7_34[21] , \wRegOut_5_22[14] , \wRegInTop_6_2[7] , 
        \wRegInBot_6_3[1] , \wRegInTop_6_29[3] , \wRegOut_7_21[15] , 
        \wRegOut_7_54[25] , \wRegOut_7_77[14] , \wRegOut_1_0[16] , 
        \wRegOut_3_3[23] , \wRegInTop_4_7[24] , \ScanLink39[10] , 
        \wRegOut_5_14[11] , \wRegInTop_6_0[20] , \ScanLink66[5] , 
        \wRegOut_6_38[8] , \wRegOut_7_7[8] , \ScanLink238[2] , 
        \wRegInTop_7_117[4] , \wRegOut_7_99[21] , \wRegInTop_7_119[21] , 
        \wRegInBot_6_0[2] , \wRegInTop_6_1[4] , \ScanLink158[7] , 
        \ScanLink211[25] , \wRegOut_6_25[7] , \ScanLink197[13] , 
        \ScanLink232[14] , \ScanLink247[24] , \wRegOut_5_10[20] , 
        \wRegOut_5_26[25] , \ScanLink59[14] , \wRegInTop_7_16[9] , 
        \ScanLink182[27] , \ScanLink227[20] , \ScanLink252[10] , 
        \ScanLink145[8] , \ScanLink204[11] , \wRegInTop_6_4[11] , 
        \wRegOut_7_88[24] , \wRegInTop_7_108[24] , \ScanLink42[3] , 
        \wRegInBot_5_12[1] , \wRegOut_7_119[2] , \wRegInTop_4_3[15] , 
        \wRegInTop_6_13[9] , \ScanLink48[11] , \ScanLink215[14] , 
        \ScanLink243[15] , \wRegOut_1_0[25] , \wRegInBot_2_1[15] , 
        \wRegOut_3_7[12] , \wRegOut_7_20[7] , \ScanLink193[22] , 
        \ScanLink236[25] , \ScanLink28[15] , \wRegInBot_6_43[3] , 
        \ScanLink186[16] , \ScanLink223[11] , \wRegOut_5_0[18] , 
        \wRegInBot_5_23[19] , \ScanLink90[21] , \ScanLink90[5] , 
        \ScanLink168[23] , \ScanLink200[20] , \wRegOut_6_9[1] , 
        \ScanLink93[6] , \ScanLink85[15] , \wRegOut_7_23[4] , \ScanLink202[8] , 
        \wRegOut_3_7[21] , \ScanLink41[0] , \wRegInBot_6_40[0] , 
        \ScanLink108[27] , \wRegOut_7_13[21] , \wRegOut_7_30[10] , 
        \wRegOut_7_66[11] , \wRegOut_7_45[20] , \wRegInBot_5_11[2] , 
        \wRegOut_7_25[24] , \wRegOut_7_50[14] , \wRegOut_7_73[25] , 
        \wRegInTop_4_3[26] , \ScanLink28[26] , \wRegInTop_6_18[19] , 
        \wRegInTop_7_16[29] , \wRegInTop_7_40[31] , \ScanLink186[25] , 
        \wRegInTop_7_63[19] , \ScanLink223[22] , \wRegInTop_7_16[30] , 
        \wRegInTop_7_35[18] , \ScanLink200[13] , \wRegInTop_7_99[2] , 
        \ScanLink48[22] , \wRegOut_5_29[8] , \wRegInTop_7_40[28] , 
        \ScanLink215[27] , \wRegInBot_4_9[9] , \wRegOut_7_44[3] , 
        \ScanLink236[16] , \ScanLink193[11] , \wRegOut_5_10[13] , 
        \wRegInBot_6_1[31] , \wRegInBot_6_27[7] , \ScanLink243[26] , 
        \wRegInBot_6_1[28] , \wRegOut_7_88[17] , \wRegInTop_7_108[17] , 
        \wRegOut_1_1[0] , \ScanLink3[21] , \wRegInBot_2_1[26] , 
        \ScanLink25[4] , \ScanLink26[7] , \wRegOut_4_15[1] , \ScanLink118[5] , 
        \wRegOut_5_26[16] , \wRegEnTop_6_24[0] , \wRegInTop_6_4[22] , 
        \wRegOut_7_96[5] , \wRegOut_7_13[12] , \wRegOut_7_25[17] , 
        \wRegInTop_7_48[7] , \wRegOut_7_50[27] , \wRegOut_7_66[22] , 
        \wRegOut_7_73[16] , \wRegOut_7_95[6] , \wRegOut_7_45[13] , 
        \ScanLink106[9] , \wRegOut_7_30[23] , \ScanLink108[14] , 
        \wRegInTop_7_55[8] , \wRegInTop_7_98[18] , \ScanLink5[1] , 
        \wRegInTop_5_15[31] , \wRegInTop_5_15[28] , \ScanLink85[26] , 
        \wRegInBot_6_24[4] , \wRegOut_7_47[0] , \wRegOut_7_88[9] , 
        \ScanLink168[10] , \ScanLink90[12] , \wRegOut_6_3[20] , 
        \wRegInTop_6_13[15] , \wRegInTop_7_68[15] , \wRegOut_7_123[12] , 
        \wRegEnBot_6_16[0] , \wRegInBot_6_25[17] , \wRegInTop_6_45[14] , 
        \wRegInBot_6_13[12] , \wRegInTop_6_25[10] , \wRegInTop_6_30[24] , 
        \wRegInBot_6_50[27] , \wRegOut_7_100[23] , \wRegInBot_6_30[23] , 
        \wRegInTop_6_50[20] , \wRegInBot_6_45[13] , \wRegOut_7_115[17] , 
        \ScanLink6[2] , \ScanLink7[21] , \wRegInTop_3_0[23] , 
        \wRegInBot_3_5[30] , \wRegInBot_3_5[29] , \wRegInBot_6_58[2] , 
        \wRegOut_4_4[24] , \wRegInTop_6_15[7] , \wRegInTop_7_34[1] , 
        \ScanLink167[0] , \ScanLink59[2] , \wRegInBot_5_2[23] , 
        \wRegInTop_6_16[4] , \wRegOut_7_26[9] , \wRegOut_7_102[3] , 
        \wRegInTop_7_37[2] , \ScanLink207[5] , \wRegInTop_7_9[3] , 
        \ScanLink164[3] , \wRegInTop_4_10[14] , \wRegInBot_4_10[13] , 
        \wRegInTop_5_7[30] , \ScanLink204[6] , \wRegInTop_5_7[29] , 
        \ScanLink95[8] , \wRegEnTop_7_79[0] , \wRegOut_7_101[0] , 
        \wRegInTop_5_28[21] , \ScanLink120[29] , \ScanLink103[18] , 
        \ScanLink120[30] , \ScanLink155[19] , \ScanLink176[31] , 
        \wRegInTop_7_93[14] , \wRegOut_7_38[5] , \ScanLink176[28] , 
        \ScanLink219[9] , \wRegOut_6_19[3] , \wRegInTop_7_86[20] , 
        \ScanLink7[12] , \wRegInTop_3_0[10] , \wRegInBot_5_28[26] , 
        \ScanLink88[7] , \ScanLink103[4] , \wRegInTop_7_50[5] , 
        \wRegOut_4_4[17] , \ScanLink20[9] , \ScanLink23[19] , 
        \wRegInTop_4_8[19] , \wRegInBot_6_21[9] , \wRegOut_7_83[28] , 
        \wRegInTop_7_103[28] , \wRegInTop_6_25[23] , \wRegOut_7_83[31] , 
        \wRegInTop_7_103[31] , \wRegInTop_7_120[19] , \wRegInBot_6_45[20] , 
        \wRegInTop_7_82[3] , \wRegInTop_5_20[1] , \wRegInBot_6_30[10] , 
        \wRegInTop_6_50[13] , \wRegOut_7_115[24] , \ScanLink56[30] , 
        \ScanLink75[18] , \wRegInTop_6_13[26] , \wRegInBot_6_13[21] , 
        \ScanLink248[19] , \wRegInTop_7_68[26] , \wRegOut_7_123[21] , 
        \wRegOut_7_100[10] , \wRegOut_6_3[13] , \wRegInTop_6_30[17] , 
        \wRegInBot_6_50[14] , \wRegInTop_4_10[27] , \wRegInTop_5_23[2] , 
        \ScanLink56[29] , \wRegInBot_6_25[24] , \wRegInTop_6_45[27] , 
        \wRegInBot_4_10[20] , \wRegInTop_5_28[12] , \wRegInBot_5_28[15] , 
        \wRegInTop_7_81[0] , \wRegInTop_7_86[13] , \wRegOut_7_93[8] , 
        \wRegOut_6_20[18] , \ScanLink100[7] , \wRegInTop_7_93[27] , 
        \wRegOut_6_55[28] , \wRegInTop_7_53[6] , \wRegOut_7_78[30] , 
        \wRegInBot_3_1[30] , \wRegInBot_3_1[29] , \wRegOut_4_5[5] , 
        \wRegInBot_4_9[20] , \wRegInBot_5_2[10] , \wRegOut_6_55[31] , 
        \wRegOut_6_60[8] , \wRegInTop_6_17[15] , \wRegEnBot_6_56[0] , 
        \wRegOut_7_78[29] , \wRegOut_7_127[12] , \wRegInTop_6_62[25] , 
        \wRegInTop_7_19[25] , \wRegInTop_5_3[9] , \wRegOut_6_7[20] , 
        \ScanLink189[29] , \wRegOut_7_104[23] , \wRegInBot_6_18[2] , 
        \wRegInTop_6_21[10] , \wRegInBot_6_21[17] , \wRegInTop_6_34[24] , 
        \wRegInBot_6_54[27] , \wRegInTop_6_41[14] , \wRegInTop_6_48[8] , 
        \ScanLink189[30] , \wRegInBot_6_34[23] , \wRegInBot_6_41[13] , 
        \wRegInTop_6_54[20] , \wRegOut_7_111[17] , \wRegInBot_6_62[22] , 
        \wRegInTop_7_79[21] , \wRegInBot_6_17[12] , \wRegOut_4_0[24] , 
        \wRegInTop_3_4[23] , \ScanLink19[2] , \wRegInTop_6_55[7] , 
        \ScanLink127[0] , \wRegInTop_7_74[1] , \wRegInTop_6_56[4] , 
        \wRegOut_7_8[23] , \wRegOut_7_66[9] , \ScanLink247[5] , 
        \ScanLink124[3] , \wRegInTop_7_77[2] , \wRegInBot_3_1[8] , 
        \wRegOut_4_6[6] , \wRegInBot_4_14[13] , \wRegInTop_5_3[30] , 
        \wRegInBot_5_6[23] , \wRegInTop_5_3[29] , \ScanLink244[6] , 
        \ScanLink124[29] , \ScanLink151[19] , \wRegEnTop_7_39[0] , 
        \ScanLink172[31] , \ScanLink172[28] , \wRegInTop_3_4[10] , 
        \wRegInTop_4_14[14] , \ScanLink107[18] , \wRegInTop_7_97[14] , 
        \ScanLink124[30] , \wRegEnTop_5_5[0] , \wRegOut_6_59[3] , 
        \wRegOut_7_78[5] , \wRegInTop_7_82[20] , \wRegOut_5_29[29] , 
        \wRegOut_4_0[17] , \wRegOut_5_29[30] , \wRegInTop_6_31[3] , 
        \wRegInTop_7_10[5] , \ScanLink143[4] , \wRegInBot_6_61[9] , 
        \wRegEnTop_7_106[0] , \ScanLink223[1] , \wRegInTop_7_107[28] , 
        \wRegOut_7_87[31] , \wRegOut_7_87[28] , \wRegInTop_7_107[31] , 
        \wRegOut_7_126[7] , \wRegInTop_7_124[19] , \wRegInBot_4_9[13] , 
        \ScanLink52[30] , \wRegInTop_6_7[8] , \wRegInTop_6_21[23] , 
        \wRegInBot_6_34[10] , \wRegInTop_6_54[13] , \ScanLink239[30] , 
        \ScanLink191[2] , \wRegOut_7_111[24] , \wRegInBot_6_17[21] , 
        \wRegInBot_6_41[20] , \ScanLink239[29] , \wRegInBot_6_62[11] , 
        \wRegInTop_7_79[12] , \wRegInTop_7_19[16] , \ScanLink27[19] , 
        \ScanLink52[29] , \ScanLink71[18] , \wRegInTop_6_17[26] , 
        \wRegInTop_6_62[16] , \wRegOut_7_127[21] , \wRegOut_6_7[13] , 
        \wRegInBot_6_21[24] , \wRegInTop_6_41[27] , \wRegInTop_7_111[8] , 
        \wRegInBot_6_54[14] , \wRegInTop_4_14[27] , \ScanLink60[9] , 
        \wRegInTop_6_34[17] , \wRegOut_7_104[10] , \wRegOut_7_1[4] , 
        \wRegInTop_7_82[13] , \wRegOut_0_0[19] , \ScanLink192[1] , 
        \wRegInBot_0_0[4] , \ScanLink3[12] , \wRegInBot_4_14[20] , 
        \wRegOut_7_2[7] , \wRegInTop_7_97[27] , \wRegInBot_5_6[10] , 
        \wRegOut_6_24[18] , \wRegInTop_6_32[0] , \ScanLink140[7] , 
        \wRegInTop_7_13[6] , \wRegOut_7_125[4] , \wRegOut_6_51[28] , 
        \wRegOut_7_8[10] , \wRegOut_6_51[31] , \wRegOut_3_3[21] , 
        \wRegOut_3_3[12] , \wRegInBot_3_4[5] , \wRegInTop_3_5[3] , 
        \wRegOut_5_22[25] , \wRegOut_6_20[8] , \ScanLink220[2] , 
        \wRegOut_7_99[10] , \wRegInTop_7_119[10] , \wRegInTop_4_7[15] , 
        \wRegInBot_5_4[1] , \wRegInTop_6_0[11] , \wRegInTop_5_5[7] , 
        \wRegOut_5_14[20] , \wRegOut_5_10[3] , \ScanLink211[14] , 
        \ScanLink39[21] , \wRegInTop_6_53[9] , \ScanLink197[22] , 
        \ScanLink232[25] , \ScanLink247[15] , \wRegInTop_3_6[0] , 
        \wRegOut_5_4[18] , \wRegInBot_5_27[19] , \ScanLink59[25] , 
        \wRegOut_6_41[1] , \ScanLink182[16] , \ScanLink227[11] , 
        \wRegOut_7_60[7] , \ScanLink252[21] , \ScanLink94[21] , 
        \ScanLink119[13] , \ScanLink204[20] , \ScanLink81[15] , 
        \wRegOut_6_42[2] , \wRegOut_7_63[4] , \ScanLink242[8] , 
        \wRegOut_6_19[11] , \ScanLink179[17] , \wRegOut_7_62[11] , 
        \wRegInBot_3_7[6] , \wRegOut_7_17[21] , \wRegOut_4_0[8] , 
        \wRegInTop_5_6[4] , \wRegInBot_5_7[2] , \wRegInTop_5_8[16] , 
        \wRegOut_7_34[10] , \wRegOut_7_41[20] , \wRegOut_5_13[0] , 
        \wRegOut_7_54[14] , \wRegOut_7_21[24] , \wRegOut_7_77[25] , 
        \wRegInTop_7_12[29] , \wRegInTop_7_44[31] , \wRegInTop_7_67[19] , 
        \ScanLink252[12] , \wRegInTop_4_7[26] , \ScanLink59[16] , 
        \wRegInTop_7_12[30] , \wRegInTop_7_44[28] , \ScanLink182[25] , 
        \ScanLink227[22] , \wRegInTop_7_31[18] , \ScanLink204[13] , 
        \ScanLink39[12] , \wRegOut_5_14[13] , \wRegInBot_6_5[31] , 
        \wRegOut_6_25[5] , \ScanLink197[11] , \ScanLink211[27] , 
        \wRegEnTop_7_97[0] , \wRegOut_7_120[9] , \ScanLink247[26] , 
        \ScanLink232[16] , \wRegOut_5_22[16] , \wRegInBot_6_0[0] , 
        \wRegInTop_6_1[6] , \wRegInBot_6_5[28] , \ScanLink158[5] , 
        \wRegInTop_7_117[6] , \ScanLink66[7] , \wRegOut_1_0[27] , 
        \wRegOut_1_0[14] , \wRegInBot_2_1[17] , \wRegInBot_4_14[0] , 
        \wRegInTop_6_0[22] , \wRegOut_7_99[23] , \wRegInTop_7_119[23] , 
        \wRegInTop_6_2[5] , \wRegInBot_6_3[3] , \ScanLink238[0] , 
        \wRegOut_7_21[17] , \wRegOut_6_19[22] , \wRegInTop_6_29[1] , 
        \wRegOut_7_54[27] , \wRegOut_7_17[12] , \wRegOut_7_77[16] , 
        \wRegOut_7_62[22] , \wRegOut_7_34[23] , \wRegInTop_5_8[25] , 
        \wRegInTop_7_114[5] , \ScanLink41[2] , \wRegInTop_5_11[31] , 
        \wRegInTop_5_11[28] , \ScanLink65[4] , \wRegOut_7_4[9] , 
        \ScanLink81[26] , \wRegInTop_7_15[8] , \ScanLink146[9] , 
        \wRegOut_7_41[13] , \ScanLink189[0] , \ScanLink179[24] , 
        \wRegInBot_5_28[9] , \wRegOut_6_26[6] , \ScanLink94[12] , 
        \ScanLink119[20] , \wRegInBot_5_11[0] , \wRegOut_7_25[26] , 
        \wRegOut_7_50[16] , \wRegOut_6_9[3] , \wRegOut_7_13[23] , 
        \wRegOut_7_66[13] , \wRegOut_7_73[27] , \wRegOut_7_30[12] , 
        \wRegOut_7_45[22] , \wRegInTop_7_98[30] , \ScanLink93[4] , 
        \wRegInBot_6_40[2] , \wRegInTop_7_98[29] , \ScanLink108[25] , 
        \wRegOut_3_7[10] , \wRegInTop_5_15[19] , \ScanLink85[17] , 
        \ScanLink90[23] , \wRegOut_7_23[6] , \ScanLink168[21] , 
        \wRegInTop_6_10[8] , \wRegInBot_6_43[1] , \wRegInTop_7_35[30] , 
        \wRegInTop_4_3[17] , \ScanLink28[17] , \wRegInTop_6_18[28] , 
        \wRegInTop_7_16[18] , \ScanLink186[14] , \ScanLink223[13] , 
        \wRegInTop_7_63[28] , \wRegOut_7_20[5] , \wRegInTop_7_35[29] , 
        \ScanLink201[9] , \wRegInTop_7_40[19] , \wRegInTop_7_63[31] , 
        \ScanLink200[22] , \ScanLink48[13] , \wRegInTop_6_18[31] , 
        \ScanLink90[7] , \ScanLink215[16] , \wRegOut_5_10[22] , 
        \ScanLink193[20] , \ScanLink236[27] , \ScanLink243[17] , 
        \wRegOut_7_88[26] , \wRegInTop_7_108[26] , \wRegInBot_2_1[24] , 
        \wRegOut_5_0[30] , \ScanLink38[9] , \ScanLink42[1] , 
        \wRegInBot_5_12[3] , \wRegInBot_6_1[19] , \wRegOut_7_119[0] , 
        \wRegInBot_5_23[31] , \wRegOut_5_26[27] , \wRegEnTop_7_61[0] , 
        \wRegInTop_6_4[13] , \wRegInBot_6_24[6] , \ScanLink168[12] , 
        \ScanLink90[10] , \wRegInBot_5_23[28] , \wRegOut_7_47[2] , 
        \ScanLink85[24] , \ScanLink25[6] , \wRegOut_5_0[29] , 
        \wRegInBot_6_39[9] , \ScanLink108[16] , \wRegOut_7_13[10] , 
        \wRegOut_7_30[21] , \wRegOut_7_66[20] , \wRegOut_7_95[4] , 
        \ScanLink26[5] , \wRegOut_4_15[3] , \wRegOut_5_26[14] , 
        \wRegOut_7_25[15] , \wRegOut_7_45[11] , \wRegInTop_7_48[5] , 
        \wRegOut_7_50[25] , \wRegOut_7_73[14] , \wRegOut_5_10[11] , 
        \wRegInTop_6_4[20] , \wRegOut_7_88[15] , \wRegOut_7_96[7] , 
        \wRegInTop_7_108[15] , \wRegEnBot_2_1[0] , \ScanLink5[3] , 
        \ScanLink6[0] , \wRegOut_3_7[23] , \wRegInTop_4_3[24] , 
        \ScanLink118[7] , \ScanLink48[20] , \ScanLink215[25] , 
        \wRegInBot_6_27[5] , \ScanLink243[24] , \wRegOut_7_44[1] , 
        \ScanLink193[13] , \ScanLink236[14] , \ScanLink28[24] , 
        \ScanLink186[27] , \ScanLink223[20] , \ScanLink105[8] , 
        \wRegInTop_7_56[9] , \ScanLink200[11] , \wRegInTop_7_99[0] , 
        \ScanLink7[23] , \wRegInTop_4_10[16] , \wRegOut_6_19[1] , 
        \wRegInBot_4_10[11] , \wRegInTop_5_28[23] , \wRegInBot_5_28[24] , 
        \wRegOut_7_38[7] , \wRegInTop_7_86[22] , \ScanLink88[5] , 
        \wRegInTop_6_16[6] , \wRegOut_6_20[29] , \wRegOut_6_55[19] , 
        \wRegOut_7_25[8] , \wRegInTop_7_93[16] , \ScanLink204[4] , 
        \wRegOut_7_101[2] , \wRegInTop_7_9[1] , \ScanLink164[1] , 
        \wRegInTop_7_37[0] , \wRegInTop_3_0[21] , \wRegInBot_5_2[21] , 
        \wRegOut_6_20[30] , \ScanLink59[0] , \wRegOut_7_78[18] , 
        \wRegOut_7_102[1] , \ScanLink96[9] , \wRegOut_4_4[26] , 
        \ScanLink207[7] , \wRegInTop_4_8[28] , \wRegInTop_6_15[5] , 
        \ScanLink167[2] , \wRegOut_7_83[19] , \wRegInTop_7_103[19] , 
        \wRegInTop_7_120[31] , \wRegInTop_7_120[28] , \wRegInTop_6_25[12] , 
        \wRegInTop_7_34[3] , \wRegInBot_6_45[11] , \ScanLink248[31] , 
        \wRegOut_7_115[15] , \wRegInBot_6_30[21] , \wRegInTop_6_50[22] , 
        \wRegInBot_6_58[0] , \ScanLink248[28] , \ScanLink7[10] , 
        \ScanLink23[31] , \wRegInTop_4_8[31] , \wRegInBot_6_13[10] , 
        \ScanLink23[28] , \ScanLink75[29] , \wRegInTop_6_13[17] , 
        \wRegInTop_7_68[17] , \wRegOut_7_123[10] , \wRegOut_7_100[21] , 
        \wRegInBot_5_2[12] , \ScanLink56[18] , \wRegOut_6_3[22] , 
        \wRegInBot_6_50[25] , \ScanLink75[30] , \wRegInTop_6_30[26] , 
        \wRegInBot_6_25[15] , \wRegInBot_6_22[8] , \wRegInTop_6_45[16] , 
        \wRegInTop_3_0[12] , \wRegInBot_3_5[18] , \wRegOut_4_4[15] , 
        \ScanLink23[8] , \wRegInTop_5_7[18] , \ScanLink100[5] , 
        \wRegInTop_7_53[4] , \wRegInTop_5_28[10] , \ScanLink103[30] , 
        \ScanLink120[18] , \wRegInTop_4_10[25] , \wRegInBot_4_10[22] , 
        \wRegOut_5_31[8] , \ScanLink103[29] , \ScanLink155[28] , 
        \wRegInTop_7_93[25] , \ScanLink155[31] , \ScanLink176[19] , 
        \wRegInTop_5_20[3] , \wRegInTop_5_23[0] , \wRegInTop_7_86[11] , 
        \wRegInBot_5_28[17] , \wRegOut_6_3[11] , \wRegInTop_6_13[24] , 
        \wRegInTop_7_68[24] , \wRegInTop_7_81[2] , \wRegOut_7_123[23] , 
        \wRegInBot_6_25[26] , \wRegOut_7_90[9] , \wRegInTop_6_45[25] , 
        \wRegInBot_6_50[16] , \wRegInBot_6_13[23] , \wRegInTop_6_25[21] , 
        \wRegInTop_6_30[15] , \wRegOut_7_100[12] , \wRegInBot_6_30[12] , 
        \wRegInTop_6_50[11] , \wRegInBot_6_45[22] , \wRegInTop_7_82[1] , 
        \wRegOut_7_115[26] , \wRegOut_6_63[9] , \wRegOut_3_3[0] , 
        \wRegOut_3_6[30] , \wRegOut_6_9[24] , \wRegInBot_6_19[16] , 
        \ScanLink103[6] , \wRegInTop_7_50[7] , \ScanLink192[19] , 
        \wRegInTop_7_77[25] , \wRegInTop_7_21[24] , \wRegInTop_7_54[14] , 
        \wRegInTop_7_34[10] , \wRegInTop_7_41[20] , \wRegInTop_7_46[3] , 
        \wRegOut_3_6[29] , \wRegInBot_4_7[24] , \wRegInTop_6_19[11] , 
        \ScanLink115[2] , \wRegInTop_7_62[11] , \wRegInTop_4_5[8] , 
        \wRegInTop_7_17[21] , \wRegOut_7_49[4] , \wRegOut_5_3[4] , 
        \wRegInBot_6_0[20] , \wRegInTop_7_94[5] , \wRegOut_3_0[3] , 
        \wRegInBot_6_29[3] , \wRegInTop_3_1[18] , \wRegInBot_3_4[12] , 
        \wRegInBot_4_7[17] , \ScanLink28[3] , \wRegInTop_4_14[2] , 
        \wRegOut_5_0[7] , \wRegInBot_5_8[27] , \wRegOut_7_6[27] , 
        \wRegInTop_7_97[6] , \wRegOut_5_1[23] , \wRegInTop_5_14[20] , 
        \wRegInBot_5_22[22] , \ScanLink169[18] , \wRegOut_7_57[8] , 
        \wRegOut_7_98[1] , \wRegOut_5_11[31] , \wRegInBot_5_14[27] , 
        \wRegInTop_7_99[10] , \wRegInTop_5_22[25] , \wRegInBot_6_0[13] , 
        \wRegOut_6_7[5] , \ScanLink116[1] , \wRegInTop_7_45[0] , 
        \wRegOut_5_11[28] , \wRegInTop_6_5[19] , \wRegOut_6_9[17] , 
        \wRegInTop_7_1[9] , \wRegInTop_7_34[23] , \wRegInTop_7_41[13] , 
        \ScanLink201[28] , \wRegOut_7_114[5] , \wRegInTop_7_17[12] , 
        \wRegOut_5_1[10] , \wRegInBot_5_14[14] , \ScanLink49[19] , 
        \wRegOut_6_11[9] , \wRegInTop_6_19[22] , \wRegInTop_7_62[22] , 
        \ScanLink201[31] , \ScanLink222[19] , \ScanLink211[3] , 
        \wRegInBot_6_19[25] , \wRegInTop_7_21[17] , \wRegInTop_7_77[16] , 
        \wRegInTop_7_22[7] , \ScanLink171[6] , \wRegInTop_7_54[27] , 
        \wRegInTop_7_99[23] , \wRegInBot_6_50[8] , \ScanLink212[0] , 
        \wRegInBot_5_8[14] , \wRegInTop_5_14[13] , \wRegInTop_5_22[16] , 
        \wRegOut_7_117[6] , \wRegInBot_5_22[11] , \ScanLink91[30] , 
        \wRegInTop_7_21[4] , \ScanLink172[5] , \ScanLink91[29] , 
        \ScanLink51[8] , \wRegOut_6_4[6] , \wRegInTop_7_120[9] , 
        \wRegOut_7_6[14] , \wRegInBot_6_31[1] , \wRegEnTop_7_7[0] , 
        \wRegOut_7_12[30] , \wRegOut_7_31[18] , \wRegOut_7_44[28] , 
        \wRegOut_7_12[29] , \wRegOut_7_44[31] , \wRegOut_7_67[19] , 
        \wRegInTop_7_121[11] , \wRegOut_4_14[14] , \wRegOut_7_52[5] , 
        \wRegOut_7_82[20] , \wRegInTop_7_102[20] , \wRegOut_7_97[14] , 
        \wRegInTop_7_117[14] , \ScanLink2[18] , \wRegInTop_2_0[1] , 
        \wRegInBot_2_1[7] , \wRegInBot_2_2[4] , \wRegInBot_4_2[0] , 
        \wRegInTop_4_3[6] , \ScanLink22[11] , \ScanLink57[21] , 
        \wRegOut_7_101[18] , \ScanLink30[1] , \wRegOut_5_22[1] , 
        \wRegEnTop_7_13[0] , \wRegOut_7_122[30] , \ScanLink74[10] , 
        \wRegOut_7_80[3] , \ScanLink229[15] , \wRegOut_7_122[29] , 
        \ScanLink199[26] , \wRegInTop_2_3[2] , \ScanLink14[14] , 
        \ScanLink61[24] , \wRegInBot_6_12[29] , \wRegInTop_5_30[9] , 
        \ScanLink249[11] , \wRegInBot_6_44[31] , \wRegInTop_4_0[5] , 
        \wRegInTop_4_9[11] , \ScanLink42[15] , \wRegInBot_6_12[30] , 
        \wRegInBot_6_31[18] , \wRegInBot_6_44[28] , \ScanLink37[25] , 
        \ScanLink102[23] , \wRegInBot_4_1[3] , \wRegInBot_4_11[28] , 
        \wRegOut_7_83[0] , \wRegInBot_4_11[31] , \ScanLink33[2] , 
        \ScanLink121[12] , \ScanLink177[13] , \wRegOut_5_6[9] , 
        \wRegOut_5_21[2] , \ScanLink154[22] , \ScanLink117[17] , 
        \ScanLink134[26] , \ScanLink141[16] , \wRegInTop_7_91[8] , 
        \ScanLink162[27] , \wRegOut_2_2[26] , \wRegOut_2_2[15] , 
        \wRegInTop_7_1[16] , \ScanLink6[29] , \ScanLink8[6] , \ScanLink14[27] , 
        \wRegInBot_5_3[18] , \wRegInTop_5_6[12] , \wRegOut_6_21[10] , 
        \wRegInBot_6_32[2] , \wRegOut_7_51[6] , \wRegOut_7_79[21] , 
        \wRegOut_6_34[24] , \wRegOut_6_54[20] , \wRegOut_6_41[14] , 
        \wRegInTop_6_62[8] , \wRegOut_6_17[15] , \wRegOut_6_62[25] , 
        \wRegOut_7_19[25] , \ScanLink249[22] , \ScanLink22[22] , 
        \wRegInTop_4_9[22] , \ScanLink61[17] , \wRegInTop_6_51[31] , 
        \ScanLink199[15] , \wRegInTop_6_24[18] , \wRegInTop_7_125[4] , 
        \ScanLink37[16] , \ScanLink42[26] , \ScanLink54[5] , 
        \wRegInTop_6_51[28] , \wRegOut_6_2[28] , \wRegInTop_7_7[7] , 
        \ScanLink57[12] , \wRegOut_6_2[31] , \wRegInTop_6_18[0] , 
        \wRegInTop_7_39[6] , \ScanLink74[23] , \wRegInBot_6_55[5] , 
        \ScanLink229[26] , \wRegOut_7_97[27] , \wRegInBot_3_4[21] , 
        \wRegOut_4_14[27] , \wRegInBot_5_19[8] , \wRegOut_6_17[7] , 
        \wRegInTop_7_117[27] , \wRegOut_7_36[1] , \ScanLink86[3] , 
        \wRegInTop_7_24[9] , \ScanLink177[8] , \wRegInTop_7_121[22] , 
        \wRegInTop_7_102[13] , \wRegInTop_5_6[21] , \wRegOut_7_82[13] , 
        \wRegOut_7_111[8] , \wRegOut_6_14[4] , \ScanLink85[0] , 
        \wRegOut_6_41[27] , \wRegOut_6_34[17] , \wRegInBot_6_56[6] , 
        \wRegOut_6_62[16] , \wRegOut_7_19[16] , \wRegOut_6_17[26] , 
        \wRegOut_7_35[2] , \ScanLink6[30] , \wRegOut_6_54[13] , 
        \wRegOut_7_79[12] , \wRegInTop_5_2[10] , \ScanLink57[6] , 
        \wRegOut_6_2[8] , \wRegOut_6_21[23] , \ScanLink141[25] , 
        \ScanLink134[15] , \wRegInTop_7_126[7] , \wRegInTop_7_87[31] , 
        \wRegInTop_5_29[30] , \ScanLink117[24] , \wRegInTop_7_1[25] , 
        \ScanLink162[14] , \ScanLink209[1] , \wRegInTop_7_87[28] , 
        \wRegInTop_5_29[29] , \ScanLink102[10] , \ScanLink177[20] , 
        \wRegInBot_6_8[8] , \ScanLink121[21] , \wRegInTop_7_4[4] , 
        \ScanLink154[11] , \ScanLink169[4] , \wRegOut_6_30[26] , 
        \wRegOut_6_45[16] , \wRegOut_6_13[17] , \wRegOut_7_68[17] , 
        \wRegInTop_2_1[26] , \wRegInBot_3_0[23] , \wRegInBot_3_0[10] , 
        \ScanLink10[16] , \wRegInBot_5_23[2] , \wRegOut_6_25[12] , 
        \wRegOut_6_30[2] , \wRegOut_7_11[4] , \ScanLink230[8] , 
        \ScanLink106[21] , \ScanLink113[15] , \wRegOut_6_50[22] , 
        \ScanLink130[24] , \ScanLink145[14] , \wRegInTop_7_5[14] , 
        \ScanLink166[25] , \wRegInTop_7_83[19] , \ScanLink173[11] , 
        \wRegInTop_7_102[1] , \ScanLink65[26] , \ScanLink73[0] , 
        \ScanLink125[10] , \ScanLink150[20] , \ScanLink238[23] , 
        \wRegInTop_6_20[30] , \wRegInTop_7_78[18] , \wRegInBot_4_8[19] , 
        \ScanLink26[13] , \ScanLink33[27] , \ScanLink46[17] , 
        \wRegInTop_6_55[19] , \wRegInTop_6_20[29] , \ScanLink181[8] , 
        \wRegInBot_5_20[1] , \ScanLink53[23] , \wRegInTop_7_101[2] , 
        \wRegOut_6_6[19] , \ScanLink70[12] , \ScanLink70[3] , 
        \wRegOut_5_28[23] , \ScanLink188[10] , \wRegOut_7_93[16] , 
        \wRegInTop_7_113[16] , \wRegInTop_6_21[9] , \wRegInTop_7_125[13] , 
        \ScanLink17[4] , \wRegOut_4_10[16] , \wRegOut_6_33[1] , 
        \wRegOut_7_12[7] , \wRegInTop_7_106[22] , \wRegInBot_4_15[19] , 
        \wRegOut_7_86[22] , \ScanLink106[12] , \ScanLink173[22] , 
        \ScanLink125[23] , \ScanLink129[6] , \ScanLink150[13] , 
        \ScanLink130[17] , \ScanLink145[27] , \wRegOut_4_10[25] , 
        \wRegInTop_5_2[23] , \wRegInBot_5_7[30] , \wRegInBot_5_7[29] , 
        \wRegOut_6_49[9] , \ScanLink113[26] , \wRegInTop_7_5[27] , 
        \ScanLink166[16] , \ScanLink249[3] , \wRegOut_7_9[30] , 
        \wRegOut_6_50[11] , \wRegOut_7_9[29] , \wRegInTop_7_67[8] , 
        \wRegOut_6_25[21] , \ScanLink134[9] , \wRegOut_6_13[24] , 
        \wRegInBot_6_16[4] , \wRegOut_6_30[15] , \wRegOut_6_45[25] , 
        \wRegOut_6_54[6] , \wRegOut_7_68[24] , \wRegOut_7_75[0] , 
        \wRegInTop_7_106[11] , \wRegInTop_7_125[20] , \ScanLink10[25] , 
        \wRegInTop_3_5[30] , \wRegOut_4_8[0] , \wRegOut_7_86[11] , 
        \wRegInBot_6_15[7] , \wRegOut_7_93[25] , \wRegInTop_7_113[25] , 
        \wRegInTop_3_5[29] , \wRegOut_5_28[10] , \wRegOut_6_57[5] , 
        \wRegOut_7_76[3] , \ScanLink26[20] , \ScanLink53[10] , 
        \wRegOut_7_105[29] , \ScanLink70[21] , \wRegInTop_6_58[2] , 
        \wRegInTop_7_79[4] , \wRegOut_7_105[30] , \wRegOut_7_126[18] , 
        \wRegInBot_6_63[28] , \ScanLink188[23] , \ScanLink14[7] , 
        \ScanLink33[14] , \ScanLink65[15] , \ScanLink238[10] , 
        \wRegInBot_6_16[18] , \wRegInBot_6_35[30] , \wRegEnTop_6_16[0] , 
        \wRegInBot_6_40[19] , \wRegInBot_6_63[31] , \wRegOut_5_5[21] , 
        \ScanLink46[24] , \wRegInBot_6_35[29] , \wRegInBot_5_10[25] , 
        \wRegInTop_5_26[27] , \wRegInBot_5_26[20] , \ScanLink68[1] , 
        \wRegInTop_6_24[4] , \ScanLink156[3] , \wRegInTop_7_119[0] , 
        \wRegInTop_2_1[15] , \ScanLink9[27] , \wRegInTop_5_10[22] , 
        \ScanLink95[18] , \wRegInTop_7_88[26] , \ScanLink236[6] , 
        \ScanLink9[14] , \wRegInBot_4_3[26] , \wRegOut_5_15[19] , 
        \wRegInBot_6_4[22] , \wRegOut_6_18[31] , \wRegOut_7_2[25] , 
        \wRegOut_7_35[29] , \ScanLink184[5] , \wRegOut_7_40[19] , 
        \wRegOut_7_63[31] , \wRegOut_6_18[28] , \wRegOut_7_16[18] , 
        \wRegOut_7_35[30] , \wRegOut_7_63[28] , \wRegEnBot_6_24[0] , 
        \ScanLink187[6] , \wRegInTop_6_1[31] , \wRegInTop_6_1[28] , 
        \wRegOut_7_98[29] , \wRegOut_6_28[0] , \wRegInTop_7_118[29] , 
        \wRegOut_7_98[30] , \wRegInTop_6_27[7] , \wRegInTop_7_30[12] , 
        \wRegInTop_7_45[22] , \wRegInTop_7_118[30] , \ScanLink155[0] , 
        \ScanLink205[19] , \ScanLink226[31] , \wRegInTop_7_66[13] , 
        \ScanLink253[18] , \ScanLink38[18] , \wRegInTop_7_13[23] , 
        \wRegOut_7_14[9] , \wRegInTop_7_73[27] , \ScanLink226[28] , 
        \ScanLink235[5] , \wRegInTop_7_50[16] , \wRegInTop_5_11[2] , 
        \wRegInTop_7_25[26] , \wRegInBot_5_26[13] , \wRegOut_7_2[16] , 
        \ScanLink6[20] , \wRegInTop_3_1[22] , \wRegOut_3_2[18] , 
        \wRegOut_5_5[12] , \wRegInTop_5_10[11] , \wRegInTop_6_40[0] , 
        \ScanLink118[19] , \ScanLink132[7] , \wRegInTop_7_61[6] , 
        \wRegInTop_7_88[15] , \wRegInBot_5_10[16] , \wRegOut_6_52[8] , 
        \ScanLink252[2] , \wRegInTop_5_26[14] , \wRegInTop_6_43[3] , 
        \ScanLink131[4] , \wRegInTop_7_25[15] , \ScanLink196[31] , 
        \ScanLink196[28] , \wRegInTop_7_73[14] , \wRegInTop_7_13[10] , 
        \wRegInTop_7_30[21] , \wRegInTop_7_50[25] , \wRegInTop_7_62[5] , 
        \wRegInTop_7_45[11] , \wRegInBot_3_4[31] , \ScanLink12[9] , 
        \wRegInBot_4_3[15] , \wRegInTop_5_8[2] , \wRegInBot_5_9[4] , 
        \wRegInBot_6_13[9] , \wRegInTop_7_66[20] , \ScanLink251[1] , 
        \wRegInTop_5_12[1] , \wRegInBot_6_4[11] , \wRegOut_6_1[2] , 
        \wRegOut_6_2[21] , \wRegInBot_6_51[26] , \wRegOut_7_101[22] , 
        \wRegInTop_6_12[14] , \wRegInTop_6_18[9] , \wRegInBot_6_24[16] , 
        \wRegInTop_6_31[25] , \wRegInTop_6_44[15] , \wRegInTop_7_69[14] , 
        \wRegOut_7_122[13] , \wRegInBot_6_12[13] , \wRegInBot_6_48[3] , 
        \wRegInTop_6_24[11] , \wRegInBot_6_31[22] , \wRegInBot_6_44[12] , 
        \wRegInTop_6_51[21] , \wRegOut_7_114[16] , \wRegInBot_3_4[28] , 
        \wRegInTop_7_24[0] , \ScanLink177[1] , \wRegOut_4_5[25] , 
        \ScanLink49[3] , \wRegInBot_5_19[1] , \wRegOut_7_36[8] , 
        \ScanLink217[4] , \wRegOut_7_112[2] , \wRegInTop_3_1[11] , 
        \wRegInTop_4_11[15] , \wRegInBot_4_11[12] , \wRegInBot_5_3[22] , 
        \wRegInTop_5_6[31] , \wRegInTop_5_6[28] , \wRegInTop_7_27[3] , 
        \ScanLink174[2] , \ScanLink85[9] , \wRegOut_7_111[1] , 
        \ScanLink214[7] , \wRegInTop_5_29[20] , \ScanLink102[19] , 
        \ScanLink177[29] , \wRegInTop_7_92[15] , \ScanLink121[31] , 
        \wRegInBot_5_29[27] , \wRegOut_6_2[1] , \ScanLink121[28] , 
        \ScanLink154[18] , \ScanLink177[30] , \ScanLink98[6] , 
        \wRegOut_7_28[4] , \ScanLink209[8] , \wRegInTop_7_87[21] , 
        \wRegOut_4_5[16] , \wRegInBot_6_31[8] , \ScanLink113[5] , 
        \wRegInTop_6_61[2] , \wRegInTop_7_40[4] , \wRegOut_7_82[30] , 
        \wRegInTop_7_102[30] , \wRegInTop_7_121[18] , \wRegInTop_7_102[29] , 
        \wRegInTop_4_9[18] , \wRegInTop_4_11[6] , \wRegOut_5_5[3] , 
        \wRegOut_7_82[29] , \wRegInBot_6_12[20] , \wRegInTop_5_30[0] , 
        \ScanLink249[18] , \wRegInTop_6_24[22] , \wRegInBot_6_31[11] , 
        \wRegInTop_6_51[12] , \wRegInTop_7_92[2] , \wRegOut_7_114[25] , 
        \ScanLink57[28] , \wRegInBot_6_44[21] , \wRegInBot_6_24[25] , 
        \wRegInBot_1_0[2] , \wRegInTop_2_0[8] , \wRegOut_3_5[7] , 
        \wRegInBot_4_2[9] , \ScanLink22[18] , \wRegOut_5_22[8] , 
        \wRegOut_6_2[12] , \wRegInTop_6_44[26] , \wRegInBot_6_51[15] , 
        \wRegOut_7_101[11] , \ScanLink30[8] , \ScanLink57[31] , 
        \wRegInTop_6_31[16] , \ScanLink74[19] , \wRegInTop_6_12[27] , 
        \wRegInTop_7_69[27] , \wRegOut_7_122[20] , \wRegInTop_4_11[26] , 
        \wRegInBot_5_29[14] , \wRegInTop_7_91[1] , \wRegOut_5_6[0] , 
        \wRegInTop_7_87[12] , \ScanLink6[13] , \wRegOut_3_6[4] , 
        \wRegInTop_4_12[5] , \wRegInTop_7_92[26] , \wRegEnBot_4_4[0] , 
        \wRegInBot_4_11[21] , \wRegOut_7_83[9] , \wRegInBot_5_3[11] , 
        \wRegInTop_5_29[13] , \ScanLink110[6] , \wRegInTop_6_62[1] , 
        \wRegInTop_7_43[7] , \wRegOut_6_54[30] , \wRegOut_7_79[28] , 
        \wRegOut_5_27[24] , \wRegInTop_6_5[10] , \wRegOut_6_21[19] , 
        \wRegOut_6_54[29] , \wRegOut_7_79[31] , \wRegInTop_7_1[0] , 
        \wRegOut_1_1[17] , \wRegInTop_1_1[4] , \ScanLink52[2] , 
        \wRegOut_7_109[3] , \wRegInTop_7_123[3] , \wRegInBot_2_0[14] , 
        \wRegOut_3_6[13] , \wRegInTop_4_2[14] , \wRegOut_5_11[21] , 
        \ScanLink49[10] , \ScanLink192[23] , \wRegOut_7_89[25] , 
        \wRegInTop_7_109[25] , \ScanLink237[24] , \ScanLink214[15] , 
        \ScanLink242[14] , \ScanLink29[14] , \ScanLink201[21] , 
        \ScanLink80[4] , \wRegInBot_6_53[2] , \wRegOut_5_1[19] , 
        \wRegInBot_5_22[18] , \wRegOut_6_11[0] , \ScanLink187[17] , 
        \ScanLink222[10] , \wRegOut_7_30[6] , \wRegOut_6_12[3] , 
        \ScanLink91[20] , \ScanLink169[22] , \ScanLink109[26] , 
        \wRegInBot_6_50[1] , \wRegOut_3_6[20] , \ScanLink29[27] , 
        \ScanLink51[1] , \ScanLink83[7] , \ScanLink84[14] , \wRegOut_7_33[5] , 
        \ScanLink212[9] , \wRegInTop_7_2[3] , \wRegOut_7_44[21] , 
        \wRegOut_7_12[20] , \wRegOut_7_31[11] , \wRegOut_7_67[10] , 
        \wRegOut_7_24[25] , \wRegOut_7_51[15] , \wRegOut_7_72[24] , 
        \wRegInTop_7_120[0] , \wRegEnTop_7_72[0] , \wRegInTop_7_41[29] , 
        \wRegInTop_6_19[18] , \wRegInTop_7_17[31] , \wRegInTop_7_34[19] , 
        \wRegInTop_7_41[30] , \ScanLink201[12] , \wRegInTop_7_89[3] , 
        \wRegInTop_7_62[18] , \wRegInTop_7_17[28] , \ScanLink187[24] , 
        \ScanLink222[23] , \ScanLink242[27] , \ScanLink2[22] , 
        \wRegOut_1_1[24] , \wRegInTop_4_2[27] , \wRegInBot_6_37[6] , 
        \wRegOut_7_54[2] , \ScanLink237[17] , \ScanLink192[10] , 
        \ScanLink49[23] , \ScanLink214[26] , \wRegInBot_6_0[29] , 
        \wRegInBot_2_0[27] , \wRegOut_3_3[9] , \wRegInTop_4_5[1] , 
        \wRegOut_5_11[12] , \wRegInBot_6_0[30] , \ScanLink108[4] , 
        \wRegOut_7_89[16] , \wRegInTop_7_109[16] , \wRegInTop_6_5[23] , 
        \wRegOut_7_86[4] , \wRegInBot_4_4[7] , \wRegInTop_4_6[2] , 
        \ScanLink35[5] , \ScanLink36[6] , \wRegOut_5_24[6] , 
        \wRegOut_5_27[17] , \wRegOut_7_24[16] , \wRegOut_7_72[17] , 
        \wRegOut_7_31[22] , \wRegOut_7_51[26] , \wRegInTop_7_58[6] , 
        \wRegOut_5_27[5] , \wRegOut_7_44[12] , \wRegOut_7_12[13] , 
        \wRegInBot_4_7[4] , \wRegOut_7_67[23] , \wRegOut_7_85[7] , 
        \ScanLink84[27] , \wRegOut_3_2[22] , \wRegOut_3_2[11] , 
        \ScanLink11[3] , \wRegInTop_5_14[30] , \wRegInTop_5_28[2] , 
        \ScanLink109[15] , \wRegInTop_7_99[19] , \ScanLink116[8] , 
        \wRegInTop_7_45[9] , \wRegInTop_5_14[29] , \ScanLink91[13] , 
        \wRegInBot_6_34[5] , \ScanLink169[11] , \wRegOut_7_20[27] , 
        \wRegOut_7_55[17] , \wRegOut_7_57[1] , \wRegOut_7_98[8] , 
        \wRegOut_7_76[26] , \wRegInTop_5_9[15] , \wRegOut_7_35[13] , 
        \wRegOut_7_40[23] , \wRegInTop_5_10[18] , \wRegInBot_6_10[3] , 
        \wRegOut_6_18[12] , \wRegOut_7_63[12] , \wRegOut_7_16[22] , 
        \ScanLink80[16] , \wRegOut_6_52[1] , \wRegOut_7_73[7] , 
        \wRegInTop_6_40[9] , \ScanLink178[14] , \ScanLink118[10] , 
        \ScanLink58[26] , \ScanLink95[22] , \wRegInTop_7_30[28] , 
        \wRegInBot_6_13[0] , \wRegInTop_7_30[31] , \wRegInTop_7_45[18] , 
        \wRegInTop_7_66[30] , \ScanLink205[23] , \wRegInTop_7_13[19] , 
        \ScanLink12[0] , \wRegInTop_4_6[16] , \wRegOut_6_51[2] , 
        \ScanLink183[15] , \wRegInTop_7_66[29] , \ScanLink226[12] , 
        \ScanLink196[21] , \wRegOut_7_70[4] , \ScanLink251[8] , 
        \ScanLink233[26] , \ScanLink253[22] , \ScanLink210[17] , 
        \ScanLink246[16] , \ScanLink38[22] , \wRegInBot_6_4[18] , 
        \wRegInTop_4_6[25] , \wRegOut_5_5[31] , \wRegOut_5_5[28] , 
        \wRegInTop_5_12[8] , \wRegOut_5_15[23] , \wRegInTop_6_1[12] , 
        \wRegOut_7_98[13] , \wRegInTop_7_118[13] , \wRegOut_5_23[26] , 
        \wRegInBot_5_26[30] , \wRegInBot_5_26[29] , \wRegInTop_7_119[9] , 
        \ScanLink68[8] , \ScanLink95[11] , \wRegOut_7_9[5] , 
        \wRegEnTop_7_84[0] , \ScanLink80[25] , \wRegOut_6_36[5] , 
        \ScanLink118[23] , \wRegOut_7_17[3] , \ScanLink178[27] , 
        \wRegInTop_5_9[26] , \wRegInBot_5_25[5] , \wRegOut_7_35[20] , 
        \ScanLink199[3] , \wRegInTop_7_104[6] , \wRegOut_5_15[10] , 
        \wRegOut_5_23[15] , \wRegInBot_5_26[6] , \wRegInTop_6_1[21] , 
        \ScanLink75[7] , \wRegOut_6_18[21] , \wRegOut_7_16[11] , 
        \wRegOut_7_40[10] , \wRegOut_7_63[21] , \wRegInTop_6_39[2] , 
        \wRegInTop_7_18[4] , \wRegOut_7_20[14] , \wRegOut_7_76[15] , 
        \wRegOut_7_55[24] , \wRegOut_7_98[20] , \wRegInTop_7_118[20] , 
        \wRegOut_6_28[9] , \ScanLink228[3] , \wRegInTop_7_107[5] , 
        \ScanLink76[4] , \ScanLink148[6] , \wEnable_0[0] , \wRegOut_6_35[6] , 
        \wRegOut_7_14[0] , \ScanLink246[25] , \ScanLink196[12] , 
        \ScanLink233[15] , \ScanLink38[11] , \ScanLink58[15] , 
        \wRegEnTop_6_9[0] , \ScanLink210[24] , \ScanLink155[9] , 
        \ScanLink205[10] , \ScanLink253[11] , \wRegInTop_4_15[17] , 
        \ScanLink183[26] , \ScanLink226[21] , \wRegInBot_4_15[10] , 
        \wRegEnBot_6_45[0] , \wRegOut_6_49[0] , \wRegOut_7_68[6] , 
        \wRegInTop_7_83[23] , \wRegInTop_5_17[5] , \wRegOut_5_18[2] , 
        \wRegInTop_7_96[17] , \wRegOut_7_75[9] , \ScanLink254[5] , 
        \ScanLink2[11] , \wRegInTop_3_5[20] , \wRegInBot_5_7[20] , 
        \wRegOut_6_25[31] , \wRegOut_5_28[19] , \wRegOut_6_25[28] , 
        \wRegInTop_6_46[7] , \wRegOut_6_50[18] , \wRegOut_7_9[20] , 
        \ScanLink134[0] , \wRegInTop_7_67[1] , \wRegOut_4_1[27] , 
        \wRegInTop_6_45[4] , \ScanLink137[3] , \wRegInTop_7_125[29] , 
        \wRegInTop_7_64[2] , \wRegInTop_7_125[30] , \wRegOut_4_8[9] , 
        \wRegOut_7_86[18] , \wRegInTop_7_106[18] , \wRegInBot_4_8[23] , 
        \ScanLink26[30] , \ScanLink26[29] , \wRegInBot_6_16[11] , 
        \wRegInBot_6_63[21] , \wRegInTop_7_78[22] , \ScanLink238[19] , 
        \wRegInTop_6_20[13] , \wRegInBot_6_35[20] , \wRegInBot_6_40[10] , 
        \wRegInTop_6_55[23] , \wRegOut_7_110[14] , \ScanLink53[19] , 
        \wRegOut_6_6[23] , \wRegOut_7_105[20] , \ScanLink70[31] , 
        \wRegInBot_6_20[14] , \wRegInTop_6_35[27] , \wRegInBot_6_55[24] , 
        \wRegInTop_6_40[17] , \wRegInTop_6_16[16] , \wRegOut_7_126[11] , 
        \wRegInTop_7_18[26] , \wRegInBot_5_7[13] , \wRegInTop_5_14[6] , 
        \ScanLink70[28] , \wRegInTop_6_63[26] , \wRegOut_2_0[5] , 
        \wRegInTop_2_0[25] , \wRegInBot_3_0[19] , \wRegOut_4_1[14] , 
        \wRegInBot_4_8[10] , \wRegInTop_4_15[24] , \wRegInBot_4_15[23] , 
        \wRegInTop_5_2[19] , \wRegInBot_6_8[1] , \wRegOut_7_9[13] , 
        \ScanLink230[1] , \wRegInTop_6_9[7] , \wRegInTop_6_22[3] , 
        \ScanLink150[4] , \ScanLink106[28] , \wRegInTop_7_96[24] , 
        \wRegEnTop_7_115[0] , \ScanLink73[9] , \ScanLink106[31] , 
        \ScanLink125[19] , \ScanLink150[30] , \ScanLink173[18] , 
        \wRegInTop_7_102[8] , \ScanLink150[29] , \ScanLink182[2] , 
        \wRegInBot_5_20[8] , \wRegInBot_6_20[27] , \wRegInTop_7_83[10] , 
        \wRegOut_6_6[10] , \wRegInTop_6_40[24] , \wRegInTop_6_35[14] , 
        \wRegInBot_6_55[17] , \wRegOut_7_105[13] , \wRegInTop_6_16[25] , 
        \wRegInTop_6_63[15] , \wRegInTop_7_18[15] , \ScanLink188[19] , 
        \wRegOut_7_126[22] , \wRegInBot_6_16[22] , \wRegInTop_6_20[20] , 
        \wRegInBot_6_35[13] , \wRegInTop_6_55[10] , \wRegInBot_6_63[12] , 
        \wRegInTop_7_78[11] , \wRegOut_6_33[8] , \wRegInBot_6_40[23] , 
        \ScanLink181[1] , \wRegOut_7_110[27] , \ScanLink233[2] , 
        \ScanLink8[24] , \wRegOut_3_3[31] , \wRegOut_3_3[28] , 
        \wRegInTop_3_5[13] , \wRegInBot_4_2[25] , \wRegInTop_6_21[0] , 
        \wRegInTop_7_12[20] , \wRegInTop_7_24[25] , \ScanLink153[7] , 
        \wRegInTop_7_51[15] , \wRegOut_7_120[0] , \wRegEnTop_7_58[0] , 
        \wRegInTop_7_67[10] , \ScanLink197[18] , \wRegInTop_7_72[24] , 
        \ScanLink225[6] , \wRegInTop_7_16[2] , \wRegInTop_7_44[21] , 
        \wRegInTop_7_31[11] , \wRegInBot_4_14[9] , \wRegInBot_6_0[9] , 
        \wRegInTop_6_37[4] , \wRegOut_6_38[3] , \wRegOut_7_7[3] , 
        \ScanLink145[3] , \wRegOut_7_19[5] , \ScanLink238[9] , 
        \wRegInBot_6_5[21] , \ScanLink197[5] , \wRegEnBot_6_6[0] , 
        \wRegOut_7_4[0] , \wRegInTop_6_29[8] , \wRegOut_7_3[26] , 
        \ScanLink194[6] , \wRegInTop_5_11[21] , \wRegEnBot_6_37[0] , 
        \wRegInBot_5_27[23] , \wRegInBot_5_28[0] , \ScanLink119[29] , 
        \wRegInTop_7_89[25] , \ScanLink226[5] , \wRegInTop_7_109[3] , 
        \wRegOut_7_123[3] , \ScanLink78[2] , \ScanLink119[30] , 
        \wRegInTop_2_0[16] , \wRegOut_2_3[6] , \wRegOut_5_4[22] , 
        \wRegInTop_5_27[24] , \wRegInTop_6_34[7] , \wRegInTop_7_15[1] , 
        \ScanLink146[0] , \ScanLink189[9] , \wRegInBot_5_11[26] , 
        \wRegEnTop_3_0[0] , \wRegInBot_5_4[8] , \wRegOut_5_14[30] , 
        \wRegOut_5_14[29] , \wRegInBot_6_5[12] , \wRegInBot_4_2[16] , 
        \wRegOut_4_3[2] , \wRegInTop_6_0[18] , \wRegOut_7_99[19] , 
        \wRegInTop_7_119[19] , \wRegOut_5_4[11] , \ScanLink39[31] , 
        \ScanLink39[28] , \wRegOut_6_41[8] , \wRegInTop_7_12[13] , 
        \wRegInTop_7_67[23] , \ScanLink204[30] , \ScanLink227[18] , 
        \ScanLink241[2] , \ScanLink252[28] , \wRegInTop_6_53[0] , 
        \ScanLink121[7] , \wRegInTop_7_24[16] , \wRegInTop_7_31[22] , 
        \wRegInTop_7_44[12] , \ScanLink204[29] , \ScanLink252[31] , 
        \wRegInTop_7_51[26] , \wRegInTop_7_72[17] , \wRegInTop_7_72[6] , 
        \wRegInBot_5_11[15] , \wRegInTop_5_27[17] , \ScanLink242[1] , 
        \wRegInTop_5_11[12] , \ScanLink94[28] , \wRegInTop_7_89[16] , 
        \wRegInBot_5_27[10] , \wRegOut_5_13[9] , \ScanLink94[31] , 
        \wRegInTop_6_50[3] , \ScanLink122[4] , \wRegInTop_7_71[5] , 
        \wRegOut_7_3[15] , \ScanLink8[17] , \wRegInBot_3_1[13] , 
        \wRegInTop_3_6[9] , \wRegOut_7_41[30] , \wRegOut_7_62[18] , 
        \wRegOut_4_0[1] , \wRegOut_6_19[18] , \wRegInBot_6_61[0] , 
        \wRegOut_7_17[31] , \wRegOut_7_17[28] , \wRegOut_7_34[19] , 
        \wRegOut_7_41[29] , \wRegOut_4_11[15] , \wRegOut_6_23[2] , 
        \ScanLink223[8] , \wRegInTop_7_107[21] , \wRegOut_5_29[20] , 
        \wRegOut_7_87[21] , \wRegInTop_7_124[10] , \wRegOut_0_0[10] , 
        \wRegOut_1_1[9] , \wRegInTop_3_4[19] , \wRegInBot_4_11[4] , 
        \ScanLink52[20] , \ScanLink71[11] , \wRegOut_7_92[15] , 
        \wRegInTop_7_112[15] , \ScanLink189[13] , \wRegOut_7_127[28] , 
        \wRegInTop_7_111[1] , \ScanLink27[10] , \wRegInBot_5_30[2] , 
        \ScanLink60[0] , \wRegOut_7_104[19] , \wRegOut_7_127[31] , 
        \wRegInBot_6_6[7] , \ScanLink11[15] , \ScanLink32[24] , 
        \ScanLink47[14] , \wRegInBot_6_17[31] , \wRegInTop_6_7[1] , 
        \wRegInBot_6_34[19] , \wRegInBot_6_41[29] , \ScanLink64[25] , 
        \wRegInBot_6_17[28] , \ScanLink239[20] , \wRegInBot_6_41[30] , 
        \wRegInBot_4_12[7] , \wRegInBot_6_62[18] , \wRegInBot_3_2[2] , 
        \wRegInTop_3_3[4] , \ScanLink11[26] , \wRegEnTop_4_11[0] , 
        \wRegInBot_4_14[30] , \ScanLink63[3] , \ScanLink124[13] , 
        \wRegInTop_7_112[2] , \wRegInBot_4_14[29] , \ScanLink107[22] , 
        \ScanLink151[23] , \wRegInBot_5_6[19] , \wRegInTop_6_4[2] , 
        \wRegInBot_6_5[4] , \ScanLink112[16] , \ScanLink172[12] , 
        \ScanLink131[27] , \wRegInTop_7_4[17] , \ScanLink167[26] , 
        \wRegOut_6_24[11] , \ScanLink144[17] , \ScanLink192[8] , 
        \wRegOut_6_51[21] , \wRegOut_7_8[19] , \wRegInBot_6_62[3] , 
        \ScanLink32[17] , \wRegInTop_5_3[13] , \wRegOut_6_12[14] , 
        \wRegOut_6_20[1] , \wRegOut_7_69[14] , \wRegOut_6_31[25] , 
        \wRegInTop_6_21[19] , \wRegInTop_6_32[9] , \wRegOut_6_44[15] , 
        \wRegInBot_5_2[6] , \ScanLink47[27] , \wRegOut_5_16[4] , 
        \wRegInTop_6_54[29] , \wRegInTop_7_79[31] , \wRegInTop_7_79[28] , 
        \wRegInTop_5_3[0] , \ScanLink64[16] , \wRegInTop_6_54[30] , 
        \ScanLink239[13] , \wRegOut_6_7[30] , \wRegInBot_4_9[29] , 
        \ScanLink71[22] , \ScanLink189[20] , \wRegInBot_4_9[30] , 
        \ScanLink27[23] , \wRegOut_6_7[29] , \ScanLink52[13] , 
        \wRegOut_5_29[13] , \wRegInTop_6_48[1] , \wRegInTop_7_69[7] , 
        \wRegOut_0_0[23] , \ScanLink3[31] , \wRegInBot_3_1[20] , 
        \wRegOut_4_11[26] , \wRegOut_6_47[6] , \wRegOut_7_92[26] , 
        \wRegInTop_7_112[26] , \wRegOut_7_66[0] , \wRegInTop_7_107[12] , 
        \wRegInTop_5_3[20] , \wRegInTop_5_19[3] , \wRegOut_7_87[12] , 
        \wRegOut_6_12[27] , \wRegOut_6_44[5] , \ScanLink127[9] , 
        \wRegInTop_7_124[23] , \wRegInTop_7_74[8] , \wRegOut_7_65[3] , 
        \wRegOut_7_69[27] , \wRegOut_6_44[26] , \wRegOut_6_31[16] , 
        \wRegOut_6_51[12] , \ScanLink3[28] , \wRegOut_6_24[22] , 
        \wRegInTop_5_0[3] , \wRegInBot_5_1[5] , \wRegInTop_7_4[24] , 
        \ScanLink167[15] , \ScanLink112[25] , \wRegOut_5_15[7] , 
        \ScanLink144[24] , \wRegInTop_7_82[29] , \ScanLink131[14] , 
        \ScanLink151[10] , \wRegInTop_7_82[30] , \wRegInBot_0_0[0] , 
        \ScanLink0[7] , \ScanLink6[9] , \wRegOut_2_3[16] , \wRegInTop_3_0[7] , 
        \ScanLink124[20] , \ScanLink139[5] , \ScanLink172[21] , 
        \wRegInBot_3_1[1] , \wRegInTop_5_7[11] , \wRegOut_6_16[16] , 
        \ScanLink107[11] , \wRegOut_6_35[27] , \wRegOut_6_63[26] , 
        \wRegOut_7_18[26] , \wRegOut_6_20[13] , \wRegOut_6_40[17] , 
        \wRegInBot_6_22[1] , \wRegOut_6_55[23] , \ScanLink7[19] , 
        \wRegOut_7_78[22] , \wRegInBot_3_5[11] , \ScanLink15[17] , 
        \ScanLink23[1] , \wRegInTop_5_23[9] , \ScanLink116[14] , 
        \wRegOut_6_60[3] , \wRegOut_7_41[5] , \ScanLink163[24] , 
        \wRegInTop_7_86[18] , \ScanLink120[11] , \wRegInTop_7_0[15] , 
        \ScanLink135[25] , \ScanLink140[15] , \wRegInTop_4_8[12] , 
        \wRegOut_4_10[7] , \wRegInTop_5_28[19] , \ScanLink155[21] , 
        \ScanLink43[16] , \wRegOut_5_31[1] , \ScanLink103[20] , 
        \wRegInTop_6_50[18] , \ScanLink176[10] , \wRegOut_7_93[3] , 
        \wRegInTop_6_25[28] , \ScanLink36[26] , \wRegInTop_7_82[8] , 
        \ScanLink60[27] , \ScanLink198[25] , \wRegInTop_6_25[31] , 
        \ScanLink248[12] , \ScanLink20[2] , \ScanLink23[12] , 
        \wRegOut_4_13[4] , \ScanLink56[22] , \ScanLink75[13] , 
        \wRegOut_7_90[0] , \ScanLink228[16] , \wRegOut_6_3[18] , 
        \wRegOut_5_8[6] , \wRegInBot_6_21[2] , \wRegOut_7_96[17] , 
        \wRegInTop_7_116[17] , \wRegOut_7_42[6] , \wRegInBot_4_10[18] , 
        \wRegOut_4_15[17] , \ScanLink120[22] , \wRegOut_6_63[0] , 
        \wRegInTop_7_103[23] , \ScanLink155[12] , \wRegOut_7_83[23] , 
        \wRegInTop_7_120[12] , \ScanLink179[7] , \ScanLink103[13] , 
        \ScanLink176[23] , \wRegInTop_7_0[26] , \ScanLink163[17] , 
        \wRegOut_2_3[25] , \wRegInBot_5_2[31] , \ScanLink47[5] , 
        \wRegInBot_5_17[7] , \wRegOut_6_19[8] , \ScanLink116[27] , 
        \ScanLink219[2] , \ScanLink140[26] , \ScanLink135[16] , 
        \wRegOut_6_55[10] , \wRegInTop_7_9[8] , \wRegInBot_5_2[28] , 
        \wRegOut_6_20[20] , \wRegInTop_7_37[9] , \ScanLink164[8] , 
        \wRegInTop_3_0[31] , \wRegInTop_3_0[28] , \wRegInBot_3_5[22] , 
        \wRegOut_4_15[24] , \wRegInTop_5_7[22] , \wRegEnTop_5_14[0] , 
        \wRegInBot_6_46[5] , \wRegOut_6_63[15] , \wRegOut_7_18[15] , 
        \wRegOut_7_78[11] , \wRegOut_7_25[1] , \wRegOut_6_16[25] , 
        \wRegOut_6_40[24] , \ScanLink95[3] , \wRegOut_6_35[14] , 
        \wRegInTop_7_103[10] , \ScanLink59[9] , \wRegOut_7_83[10] , 
        \wRegOut_7_102[8] , \wRegInTop_7_120[21] , \ScanLink96[0] , 
        \wRegInBot_6_45[6] , \wRegOut_7_96[24] , \wRegInTop_7_116[24] , 
        \ScanLink15[24] , \ScanLink23[21] , \ScanLink75[20] , 
        \wRegOut_7_26[2] , \wRegOut_7_100[31] , \wRegOut_7_123[19] , 
        \wRegOut_7_100[28] , \ScanLink228[25] , \wRegInTop_4_8[21] , 
        \wRegInBot_5_14[4] , \ScanLink56[11] , \wRegInTop_7_29[5] , 
        \ScanLink36[15] , \ScanLink43[25] , \ScanLink44[6] , 
        \wRegInBot_6_45[18] , \wRegInBot_6_30[28] , \wRegInBot_6_58[9] , 
        \ScanLink248[21] , \wRegInBot_4_6[27] , \wRegOut_5_0[20] , 
        \wRegInTop_5_23[26] , \ScanLink60[14] , \wRegInBot_6_30[31] , 
        \ScanLink198[16] , \wRegInBot_6_13[19] , \wRegEnBot_5_26[0] , 
        \ScanLink106[2] , \wRegInTop_7_55[3] , \ScanLink38[0] , 
        \wRegInTop_5_15[23] , \wRegInBot_5_15[24] , \wRegInTop_7_98[13] , 
        \ScanLink90[19] , \wRegOut_7_88[2] , \wRegInBot_5_9[24] , 
        \wRegInBot_5_23[21] , \wRegOut_7_7[24] , \wRegInTop_7_87[5] , 
        \wRegOut_5_10[18] , \wRegInTop_5_25[7] , \wRegInTop_5_26[4] , 
        \wRegInBot_6_39[0] , \wRegOut_7_13[19] , \wRegOut_7_30[31] , 
        \wRegOut_7_30[28] , \wRegOut_7_66[29] , \wRegOut_7_45[18] , 
        \wRegOut_7_66[30] , \wRegInBot_6_1[23] , \wRegInTop_6_4[30] , 
        \wRegInTop_7_84[6] , \wRegInTop_6_4[29] , \wRegInTop_6_18[12] , 
        \wRegOut_7_59[7] , \wRegInTop_7_63[12] , \wRegInTop_7_16[22] , 
        \wRegInTop_4_8[4] , \ScanLink48[29] , \wRegOut_5_29[3] , 
        \wRegOut_6_8[27] , \ScanLink223[29] , \ScanLink105[1] , 
        \wRegInTop_7_35[13] , \wRegInTop_7_40[23] , \wRegInTop_7_56[0] , 
        \ScanLink223[30] , \wRegInTop_7_55[17] , \ScanLink200[18] , 
        \wRegInTop_7_99[9] , \wRegInTop_7_20[27] , \wRegInBot_4_9[2] , 
        \wRegOut_7_44[8] , \wRegInTop_7_76[26] , \wRegInBot_5_9[17] , 
        \wRegInBot_5_11[9] , \ScanLink48[30] , \wRegInBot_6_18[15] , 
        \wRegOut_7_7[17] , \wRegOut_1_0[23] , \wRegOut_1_0[10] , 
        \wRegOut_1_1[30] , \ScanLink3[4] , \wRegOut_3_7[19] , 
        \wRegOut_5_0[13] , \wRegInTop_5_15[10] , \ScanLink168[28] , 
        \wRegInBot_5_15[17] , \wRegInTop_5_23[15] , \wRegInBot_5_23[12] , 
        \wRegInTop_6_10[1] , \ScanLink168[31] , \wRegInTop_7_31[7] , 
        \ScanLink162[6] , \wRegOut_7_107[5] , \wRegInTop_7_98[20] , 
        \ScanLink202[3] , \wRegInTop_6_13[2] , \wRegInTop_7_20[14] , 
        \ScanLink193[30] , \ScanLink161[5] , \wRegInBot_6_18[26] , 
        \wRegInTop_7_32[4] , \wRegInTop_7_55[24] , \ScanLink193[29] , 
        \wRegInTop_7_76[15] , \wRegInBot_4_6[14] , \wRegOut_6_8[14] , 
        \wRegInTop_6_18[21] , \wRegInBot_6_43[8] , \wRegInTop_7_16[11] , 
        \wRegInTop_7_63[21] , \ScanLink201[0] , \wRegInTop_7_35[20] , 
        \wRegInTop_7_40[10] , \wRegOut_7_104[6] , \wRegInTop_2_0[5] , 
        \wRegInTop_2_1[22] , \ScanLink9[23] , \wRegInBot_4_3[22] , 
        \wRegInTop_4_6[31] , \wRegInTop_4_6[28] , \ScanLink42[8] , 
        \wRegInBot_6_1[10] , \wRegOut_7_119[9] , \ScanLink246[31] , 
        \wRegInTop_7_25[22] , \wRegInTop_7_50[12] , \ScanLink210[29] , 
        \ScanLink246[28] , \wRegInTop_7_13[27] , \wRegInTop_7_66[17] , 
        \wRegInTop_7_73[23] , \ScanLink210[30] , \ScanLink233[18] , 
        \ScanLink235[1] , \wRegOut_5_23[18] , \ScanLink58[18] , 
        \wRegInTop_7_30[16] , \wRegInTop_7_45[26] , \wRegEnTop_7_110[0] , 
        \wRegInTop_6_27[3] , \ScanLink155[4] , \wRegInTop_7_107[8] , 
        \wRegInBot_5_25[8] , \wRegInBot_6_4[26] , \ScanLink76[9] , 
        \wRegOut_6_28[4] , \ScanLink187[2] , \wRegOut_7_2[21] , 
        \wRegInTop_7_18[9] , \wRegOut_7_20[19] , \wRegOut_7_55[29] , 
        \ScanLink184[1] , \wRegInTop_5_10[26] , \wRegOut_7_55[30] , 
        \wRegOut_7_76[18] , \wRegInBot_5_26[24] , \ScanLink68[5] , 
        \wRegOut_6_36[8] , \wRegOut_7_9[8] , \wRegInTop_7_88[22] , 
        \ScanLink236[2] , \wRegInTop_7_119[4] , \wRegInTop_2_1[11] , 
        \wRegInBot_4_3[11] , \wRegOut_5_5[25] , \wRegInTop_5_26[23] , 
        \ScanLink80[31] , \wRegInTop_6_24[0] , \ScanLink156[7] , 
        \wRegInBot_5_10[21] , \ScanLink80[28] , \wRegInTop_5_12[5] , 
        \wRegInBot_6_4[15] , \wRegEnBot_6_40[0] , \wRegOut_5_5[16] , 
        \wRegInTop_5_8[6] , \wRegInBot_5_9[0] , \wRegInTop_7_13[14] , 
        \ScanLink183[18] , \wRegInTop_7_66[24] , \wRegOut_7_70[9] , 
        \ScanLink251[5] , \wRegInBot_5_10[12] , \wRegInTop_5_26[10] , 
        \wRegInTop_6_43[7] , \ScanLink131[0] , \wRegInTop_7_25[11] , 
        \wRegInTop_7_30[25] , \wRegInTop_7_45[15] , \wRegInTop_7_50[21] , 
        \wRegInTop_7_62[1] , \wRegInTop_7_73[10] , \ScanLink252[6] , 
        \wRegInTop_5_10[15] , \ScanLink178[19] , \wRegInTop_7_88[11] , 
        \wRegInBot_5_26[17] , \wRegInBot_2_1[3] , \wRegOut_2_2[11] , 
        \wRegInBot_3_0[27] , \wRegInBot_3_0[14] , \ScanLink9[10] , 
        \wRegInTop_6_40[4] , \wRegOut_7_2[12] , \ScanLink132[3] , 
        \wRegInTop_7_61[2] , \wRegOut_4_1[19] , \wRegInTop_5_9[18] , 
        \wRegInTop_5_11[6] , \wRegOut_7_12[3] , \ScanLink10[21] , 
        \ScanLink10[12] , \wRegOut_4_10[12] , \ScanLink26[17] , 
        \wRegInBot_5_20[5] , \ScanLink53[27] , \wRegOut_5_28[27] , 
        \wRegOut_6_33[5] , \wRegEnTop_7_81[0] , \wRegOut_7_86[26] , 
        \wRegInTop_7_106[26] , \wRegInTop_7_125[17] , \ScanLink70[16] , 
        \wRegInTop_7_18[18] , \wRegOut_7_93[12] , \wRegInTop_7_113[12] , 
        \wRegInTop_6_16[28] , \wRegInTop_6_40[30] , \wRegInTop_6_63[18] , 
        \ScanLink188[14] , \wRegInTop_7_101[6] , \wRegInTop_6_40[29] , 
        \ScanLink33[23] , \ScanLink46[13] , \ScanLink70[7] , 
        \wRegInTop_6_35[19] , \wRegInTop_6_16[31] , \ScanLink65[22] , 
        \ScanLink238[27] , \ScanLink14[3] , \wRegInTop_4_15[30] , 
        \wRegInTop_4_15[29] , \wRegInBot_5_23[6] , \wRegInTop_7_96[30] , 
        \wRegInTop_7_102[5] , \ScanLink73[4] , \ScanLink125[14] , 
        \ScanLink106[25] , \ScanLink150[24] , \wRegInTop_7_96[29] , 
        \ScanLink173[15] , \ScanLink113[11] , \ScanLink130[20] , 
        \wRegInTop_7_5[10] , \ScanLink166[21] , \ScanLink33[10] , 
        \wRegInTop_5_2[14] , \wRegOut_6_13[13] , \wRegOut_6_25[16] , 
        \ScanLink145[10] , \wEnable_5[0] , \wRegOut_6_30[6] , 
        \wRegOut_6_50[26] , \wRegOut_7_11[0] , \wRegOut_7_68[13] , 
        \wRegOut_6_30[22] , \ScanLink150[9] , \wRegOut_6_45[12] , 
        \wRegOut_7_110[19] , \ScanLink46[20] , \wRegOut_4_10[21] , 
        \ScanLink26[24] , \ScanLink65[11] , \ScanLink238[14] , 
        \ScanLink70[25] , \wRegInBot_6_55[30] , \wRegInBot_6_55[29] , 
        \ScanLink188[27] , \ScanLink53[14] , \wRegOut_5_28[14] , 
        \wRegInBot_6_20[19] , \wRegInTop_6_58[6] , \wRegInTop_7_79[0] , 
        \wRegInBot_6_15[3] , \wRegOut_6_57[1] , \wRegOut_7_93[21] , 
        \wRegInTop_7_113[21] , \wRegOut_7_76[7] , \wRegInTop_7_106[15] , 
        \ScanLink17[0] , \wRegOut_4_8[4] , \wRegOut_7_86[15] , 
        \wRegInTop_5_2[27] , \wRegOut_6_13[20] , \wRegInBot_6_16[0] , 
        \wRegInTop_6_45[9] , \wRegInTop_7_125[24] , \wRegOut_6_54[2] , 
        \wRegOut_7_68[20] , \wRegOut_7_75[4] , \ScanLink254[8] , 
        \wRegOut_6_45[21] , \wRegOut_6_25[25] , \wRegOut_6_30[11] , 
        \wRegOut_6_50[15] , \ScanLink113[22] , \wRegInTop_7_5[23] , 
        \ScanLink166[12] , \ScanLink249[7] , \ScanLink130[13] , 
        \ScanLink145[23] , \wRegInTop_5_6[16] , \wRegInTop_5_17[8] , 
        \ScanLink125[27] , \ScanLink150[17] , \ScanLink129[2] , 
        \ScanLink173[26] , \wRegOut_6_17[11] , \ScanLink106[16] , 
        \wRegOut_6_34[20] , \wRegOut_6_62[21] , \wRegOut_7_19[21] , 
        \wRegOut_6_21[14] , \wRegOut_6_41[10] , \wRegInBot_6_32[6] , 
        \wRegOut_6_54[24] , \ScanLink117[13] , \wRegOut_7_51[2] , 
        \wRegOut_7_79[25] , \ScanLink162[23] , \wRegOut_2_2[22] , 
        \wRegInBot_2_2[0] , \wRegOut_3_6[9] , \wRegInTop_4_0[1] , 
        \wRegInTop_4_12[8] , \wRegInTop_7_1[12] , \ScanLink33[6] , 
        \wRegInBot_5_29[19] , \ScanLink134[22] , \ScanLink121[16] , 
        \ScanLink141[12] , \wRegOut_5_21[6] , \ScanLink154[26] , 
        \ScanLink102[27] , \wRegOut_7_83[4] , \wRegInBot_4_1[7] , 
        \wRegInTop_4_9[15] , \ScanLink42[11] , \ScanLink177[17] , 
        \ScanLink37[21] , \wRegOut_7_114[28] , \ScanLink199[22] , 
        \wRegInTop_2_3[6] , \ScanLink14[10] , \ScanLink61[20] , 
        \ScanLink249[15] , \wRegInBot_3_4[16] , \wRegInBot_4_2[4] , 
        \wRegInTop_4_3[2] , \ScanLink74[14] , \wRegOut_7_114[31] , 
        \wRegInBot_6_24[31] , \wRegOut_7_80[7] , \ScanLink229[11] , 
        \ScanLink22[15] , \ScanLink57[25] , \wRegInBot_6_24[28] , 
        \ScanLink30[5] , \wRegOut_5_22[5] , \wRegInBot_6_51[18] , 
        \wRegInBot_6_31[5] , \ScanLink113[8] , \wRegInTop_7_40[9] , 
        \wRegOut_7_97[10] , \wRegInTop_7_117[10] , \wRegOut_7_52[1] , 
        \wRegInTop_4_11[18] , \wRegOut_4_14[10] , \wRegInTop_7_102[24] , 
        \ScanLink102[14] , \ScanLink121[25] , \wRegInTop_7_4[0] , 
        \wRegOut_7_82[24] , \wRegInTop_7_121[15] , \ScanLink154[15] , 
        \ScanLink169[0] , \ScanLink177[24] , \wRegInTop_7_92[18] , 
        \ScanLink117[20] , \wRegInTop_7_1[21] , \ScanLink162[10] , 
        \wRegOut_7_28[9] , \ScanLink209[5] , \ScanLink57[2] , 
        \ScanLink134[11] , \ScanLink141[21] , \wRegInTop_7_126[3] , 
        \wRegEnBot_6_18[0] , \wRegOut_6_21[27] , \wRegOut_6_54[17] , 
        \wRegOut_3_0[7] , \ScanLink8[2] , \wRegInBot_3_4[25] , 
        \wRegOut_4_14[23] , \wRegInTop_5_6[25] , \wRegOut_6_14[0] , 
        \wRegInBot_6_56[2] , \wRegOut_7_19[12] , \wRegOut_7_79[16] , 
        \wRegOut_6_62[12] , \wRegOut_6_17[22] , \wRegOut_7_35[6] , 
        \wRegOut_6_41[23] , \ScanLink85[4] , \wRegOut_6_34[13] , 
        \wRegInTop_7_102[17] , \wRegOut_4_5[31] , \wRegOut_4_5[28] , 
        \wRegOut_7_82[17] , \ScanLink86[7] , \wRegInTop_7_121[26] , 
        \wRegInBot_6_55[1] , \wRegOut_7_97[23] , \ScanLink14[23] , 
        \ScanLink22[26] , \ScanLink74[27] , \wRegInTop_6_12[19] , 
        \wRegOut_6_17[3] , \wRegInTop_7_117[23] , \wRegOut_7_36[5] , 
        \ScanLink217[9] , \wRegInTop_7_69[19] , \wRegInTop_6_31[31] , 
        \wRegInTop_7_7[3] , \ScanLink229[22] , \wRegInTop_4_9[26] , 
        \ScanLink57[16] , \wRegInTop_6_31[28] , \wRegInTop_6_18[4] , 
        \wRegInTop_6_44[18] , \wRegInTop_7_39[2] , \wRegInTop_7_125[0] , 
        \ScanLink37[12] , \ScanLink42[22] , \ScanLink54[1] , 
        \wRegEnTop_7_77[0] , \ScanLink249[26] , \wRegInBot_4_7[9] , 
        \ScanLink28[7] , \wRegOut_5_1[27] , \wRegInTop_5_22[21] , 
        \ScanLink61[13] , \ScanLink199[11] , \ScanLink116[5] , 
        \wRegInTop_7_45[4] , \wRegInTop_5_14[24] , \wRegInBot_5_14[23] , 
        \wRegInTop_7_99[14] , \wRegInBot_6_34[8] , \ScanLink109[18] , 
        \wRegOut_7_98[5] , \wRegInTop_4_14[6] , \wRegOut_5_0[3] , 
        \wRegInBot_5_22[26] , \wRegOut_7_6[23] , \wRegInTop_7_97[2] , 
        \wRegInBot_5_8[23] , \wRegInBot_6_29[7] , \wRegOut_5_3[0] , 
        \ScanLink35[8] , \wRegOut_5_27[8] , \wRegOut_1_1[29] , 
        \wRegInBot_6_0[24] , \wRegInTop_1_1[9] , \wRegInBot_2_0[19] , 
        \wRegOut_3_3[4] , \wRegEnBot_4_1[0] , \ScanLink108[9] , 
        \wRegOut_7_49[0] , \wRegInTop_7_94[1] , \wRegInBot_4_7[20] , 
        \wRegInTop_6_19[15] , \wRegInTop_7_62[15] , \wRegOut_7_86[9] , 
        \wRegInTop_7_17[25] , \wRegOut_5_1[14] , \wRegInBot_5_8[10] , 
        \wRegOut_6_4[2] , \wRegOut_6_9[20] , \ScanLink187[29] , 
        \wRegInBot_6_19[12] , \ScanLink115[6] , \wRegInTop_7_34[14] , 
        \wRegInTop_7_41[24] , \wRegInTop_7_46[7] , \ScanLink187[30] , 
        \wRegInTop_7_21[20] , \wRegInTop_7_54[10] , \wRegInTop_7_77[21] , 
        \wRegOut_7_51[18] , \wRegOut_7_6[10] , \wRegOut_7_72[30] , 
        \wRegOut_7_24[28] , \wRegInTop_5_14[17] , \wRegOut_7_24[31] , 
        \wRegOut_7_72[29] , \wRegInBot_5_14[10] , \wRegInTop_5_22[12] , 
        \wRegInBot_5_22[15] , \wRegInTop_7_21[0] , \ScanLink172[1] , 
        \wRegOut_7_117[2] , \wRegInTop_7_99[27] , \ScanLink84[19] , 
        \ScanLink212[4] , \wRegOut_7_33[8] , \wRegInTop_4_2[19] , 
        \wRegInTop_7_21[13] , \ScanLink214[18] , \ScanLink237[30] , 
        \wRegInTop_7_22[3] , \ScanLink171[2] , \wRegInTop_7_54[23] , 
        \wRegInBot_4_7[13] , \wRegInBot_6_19[21] , \ScanLink237[29] , 
        \wRegInTop_7_77[12] , \ScanLink242[19] , \ScanLink29[19] , 
        \wRegInTop_6_19[26] , \wRegInTop_7_17[16] , \wRegInTop_7_62[26] , 
        \ScanLink211[7] , \wRegInTop_7_34[27] , \wRegInTop_7_41[17] , 
        \wRegOut_7_114[1] , \wRegOut_5_27[30] , \wRegOut_5_27[29] , 
        \wRegOut_6_9[13] , \ScanLink80[9] , \wRegInBot_6_0[17] , 
        \wRegOut_7_89[28] , \wRegInTop_7_109[28] , \wRegOut_6_7[1] , 
        \wRegOut_7_89[31] , \wRegInTop_7_109[31] , \ScanLink5[7] , 
        \wRegOut_6_3[26] , \wRegOut_7_100[25] , \wRegInTop_6_13[13] , 
        \wRegInBot_6_25[11] , \wRegInTop_6_30[22] , \wRegInBot_6_50[21] , 
        \wRegInTop_6_45[12] , \wRegInTop_7_29[8] , \wRegInTop_7_68[13] , 
        \ScanLink228[31] , \wRegOut_7_123[14] , \wRegInBot_6_58[4] , 
        \ScanLink228[28] , \ScanLink6[4] , \wRegOut_2_3[31] , 
        \wRegOut_2_3[28] , \ScanLink7[27] , \wRegInTop_3_0[25] , 
        \ScanLink15[30] , \ScanLink15[29] , \ScanLink43[31] , 
        \wRegInBot_5_14[9] , \ScanLink60[19] , \wRegInBot_6_13[14] , 
        \wRegInTop_6_25[16] , \wRegOut_4_4[22] , \wRegOut_4_15[30] , 
        \ScanLink36[18] , \wRegInBot_6_45[15] , \wRegOut_7_115[11] , 
        \ScanLink43[28] , \wRegInTop_6_50[26] , \wRegInBot_6_30[25] , 
        \wRegInTop_6_15[1] , \ScanLink167[6] , \wRegInTop_7_34[7] , 
        \wRegOut_4_15[29] , \ScanLink59[4] , \ScanLink207[3] , 
        \wRegOut_7_96[29] , \wRegInTop_7_116[29] , \wRegOut_7_96[30] , 
        \wRegOut_7_102[5] , \wRegInTop_7_116[30] , \wRegInBot_5_2[25] , 
        \wRegInTop_6_16[2] , \wRegInTop_7_9[5] , \wRegInTop_7_37[4] , 
        \wRegInBot_4_10[15] , \wRegOut_6_16[31] , \wRegOut_6_40[29] , 
        \ScanLink164[5] , \wRegEnTop_6_58[0] , \wRegOut_7_101[6] , 
        \wRegOut_6_16[28] , \wRegOut_6_35[19] , \wRegOut_6_40[30] , 
        \wRegOut_7_18[18] , \wRegInBot_6_46[8] , \wRegOut_6_63[18] , 
        \ScanLink204[0] , \ScanLink47[8] , \wRegInTop_5_28[27] , 
        \wRegInTop_7_93[12] , \wRegInBot_5_28[20] , \ScanLink88[1] , 
        \ScanLink7[14] , \wRegInTop_3_0[16] , \wRegInTop_4_10[12] , 
        \wRegEnBot_5_23[0] , \wRegOut_6_19[5] , \wRegOut_7_38[3] , 
        \wRegInTop_7_86[26] , \wRegOut_4_4[11] , \ScanLink103[2] , 
        \wRegInTop_7_50[3] , \wRegInTop_4_10[21] , \wRegOut_4_13[9] , 
        \wRegInTop_5_20[7] , \wRegInBot_6_13[27] , \ScanLink198[28] , 
        \wRegOut_6_3[15] , \wRegInTop_6_25[25] , \wRegInBot_6_30[16] , 
        \wRegInTop_6_50[15] , \ScanLink198[31] , \wRegInBot_6_25[22] , 
        \wRegInBot_6_45[26] , \wRegInTop_7_82[5] , \wRegOut_7_115[22] , 
        \wRegInTop_6_45[21] , \wRegInBot_6_50[12] , \wRegInBot_5_28[13] , 
        \wRegInTop_6_13[20] , \wRegInTop_6_30[11] , \wRegOut_7_100[16] , 
        \wRegInTop_7_68[20] , \wRegOut_7_123[27] , \ScanLink116[19] , 
        \ScanLink135[28] , \ScanLink140[18] , \wRegInTop_7_81[6] , 
        \ScanLink163[30] , \wRegInBot_4_10[26] , \wRegInTop_5_23[4] , 
        \wRegInTop_7_0[18] , \ScanLink135[31] , \ScanLink163[29] , 
        \wRegInTop_7_86[15] , \wRegInTop_7_93[21] , \wRegInBot_5_2[16] , 
        \wRegInTop_5_28[14] , \ScanLink100[1] , \wRegInTop_7_53[0] , 
        \wRegInBot_5_12[7] , \wRegOut_5_26[23] , \wRegInTop_6_4[17] , 
        \wRegOut_7_41[8] , \ScanLink3[9] , \ScanLink42[5] , \wRegOut_7_119[4] , 
        \wRegInBot_2_1[13] , \wRegOut_3_7[14] , \wRegInTop_4_3[13] , 
        \wRegOut_5_10[26] , \ScanLink48[17] , \wRegInTop_7_20[19] , 
        \wRegInTop_7_55[30] , \ScanLink193[24] , \wRegOut_7_88[22] , 
        \wRegInTop_7_108[22] , \ScanLink236[23] , \ScanLink243[13] , 
        \wRegInTop_7_76[18] , \ScanLink215[12] , \ScanLink161[8] , 
        \ScanLink28[13] , \wRegOut_6_8[19] , \wRegInTop_7_32[9] , 
        \wRegInTop_7_55[29] , \ScanLink200[26] , \ScanLink90[3] , 
        \wRegInBot_6_43[5] , \wRegInBot_4_6[19] , \wRegEnTop_5_11[0] , 
        \ScanLink186[10] , \ScanLink223[17] , \ScanLink90[27] , 
        \wRegOut_7_20[1] , \ScanLink168[25] , \wRegInBot_6_40[6] , 
        \ScanLink108[21] , \wRegOut_3_7[27] , \ScanLink28[20] , 
        \ScanLink41[6] , \wRegInBot_5_11[4] , \wRegInTop_5_23[18] , 
        \wRegOut_6_9[7] , \ScanLink85[13] , \wRegOut_7_23[2] , 
        \wRegOut_7_107[8] , \ScanLink93[0] , \wRegOut_7_13[27] , 
        \wRegOut_7_30[16] , \wRegOut_7_45[26] , \wRegOut_7_66[17] , 
        \wRegOut_7_73[23] , \wRegOut_7_25[22] , \wRegOut_7_50[12] , 
        \ScanLink200[15] , \wRegInTop_7_99[4] , \wRegInTop_4_3[20] , 
        \wRegInTop_4_8[9] , \ScanLink186[23] , \ScanLink223[24] , 
        \wRegInBot_6_18[18] , \wRegInBot_6_27[1] , \ScanLink243[20] , 
        \wRegOut_7_44[5] , \ScanLink193[17] , \ScanLink236[10] , 
        \ScanLink48[24] , \ScanLink215[21] , \wRegOut_2_0[8] , 
        \wRegInBot_2_1[20] , \ScanLink25[2] , \ScanLink26[1] , 
        \wRegOut_4_15[7] , \wRegOut_5_10[15] , \wRegInTop_5_26[9] , 
        \ScanLink118[3] , \wRegOut_7_88[11] , \wRegInTop_7_108[11] , 
        \wRegInTop_6_4[24] , \wRegOut_7_96[3] , \wRegOut_5_26[10] , 
        \wRegInBot_5_9[30] , \wRegInBot_5_9[29] , \wRegOut_7_7[30] , 
        \wRegOut_7_7[29] , \wRegOut_7_73[10] , \wRegOut_7_25[11] , 
        \wRegInTop_7_87[8] , \wRegOut_7_30[25] , \wRegInTop_7_48[1] , 
        \wRegOut_7_50[21] , \ScanLink85[20] , \wRegOut_7_13[14] , 
        \wRegOut_7_45[15] , \wRegOut_7_66[24] , \wRegOut_7_95[0] , 
        \wRegInBot_5_7[6] , \wRegInBot_5_15[30] , \wRegInBot_5_15[29] , 
        \ScanLink108[12] , \wRegInBot_6_24[2] , \ScanLink168[16] , 
        \ScanLink90[14] , \wRegOut_7_47[6] , \wRegOut_7_77[21] , 
        \wRegInTop_2_0[31] , \wRegInTop_2_0[28] , \wRegOut_3_3[16] , 
        \wRegInTop_3_6[4] , \wRegInTop_5_6[0] , \wRegInTop_5_8[12] , 
        \wRegOut_5_13[4] , \wRegOut_7_54[10] , \wRegOut_7_3[18] , 
        \wRegOut_7_21[20] , \wRegOut_7_34[14] , \wRegOut_7_41[24] , 
        \wRegOut_7_62[15] , \wRegInBot_3_7[2] , \wRegOut_6_19[15] , 
        \wRegOut_7_17[25] , \wRegInBot_5_11[18] , \ScanLink59[21] , 
        \ScanLink81[11] , \wRegOut_6_42[6] , \ScanLink94[25] , 
        \ScanLink119[17] , \ScanLink122[9] , \ScanLink179[13] , 
        \wRegOut_7_63[0] , \wRegInTop_7_71[8] , \ScanLink204[24] , 
        \wRegInBot_3_4[1] , \wRegInTop_3_5[7] , \wRegInTop_4_7[11] , 
        \wRegOut_6_41[5] , \ScanLink182[12] , \ScanLink227[15] , 
        \wRegOut_7_60[3] , \ScanLink197[26] , \ScanLink252[25] , 
        \ScanLink211[10] , \ScanLink232[21] , \ScanLink247[11] , 
        \wRegInBot_5_4[5] , \ScanLink39[25] , \wRegOut_5_10[7] , 
        \wRegInTop_5_5[3] , \wRegOut_5_14[24] , \wRegInTop_6_0[15] , 
        \wRegOut_7_99[14] , \wRegOut_5_22[21] , \wRegInTop_7_119[14] , 
        \wRegInTop_7_89[31] , \ScanLink94[16] , \ScanLink119[24] , 
        \wRegInTop_7_89[28] , \ScanLink8[30] , \ScanLink8[29] , 
        \wRegInBot_4_14[4] , \wRegInTop_5_27[30] , \ScanLink81[22] , 
        \wRegOut_6_26[2] , \ScanLink226[8] , \wRegInTop_5_27[29] , 
        \ScanLink179[20] , \wRegOut_7_34[27] , \ScanLink189[4] , 
        \wRegInTop_7_114[1] , \wRegInTop_5_8[21] , \ScanLink65[0] , 
        \wRegOut_6_19[26] , \wRegOut_7_17[16] , \wRegOut_7_41[17] , 
        \wRegOut_7_62[26] , \wRegOut_7_77[12] , \wRegOut_5_22[12] , 
        \wRegInTop_6_0[26] , \wRegInTop_6_2[1] , \wRegInBot_6_3[7] , 
        \wRegOut_7_21[13] , \wRegInTop_6_29[5] , \wRegOut_7_54[23] , 
        \wRegOut_7_99[27] , \wRegOut_7_19[8] , \ScanLink238[4] , 
        \wRegInTop_7_119[27] , \wRegInTop_7_117[2] , \ScanLink3[25] , 
        \wRegOut_3_3[25] , \wRegInBot_4_2[31] , \wRegInTop_4_7[22] , 
        \wRegEnTop_4_14[0] , \wRegOut_5_14[17] , \wRegInBot_6_0[4] , 
        \ScanLink66[3] , \wRegInTop_6_1[2] , \ScanLink197[8] , 
        \ScanLink158[1] , \wRegOut_6_25[1] , \ScanLink197[15] , 
        \wRegInTop_7_72[29] , \ScanLink247[22] , \ScanLink232[12] , 
        \wRegInTop_7_24[31] , \wRegInTop_7_51[18] , \wRegInTop_7_72[30] , 
        \ScanLink39[16] , \wRegInTop_6_37[9] , \wRegInTop_7_24[28] , 
        \ScanLink211[23] , \wRegInBot_4_2[28] , \ScanLink59[12] , 
        \ScanLink204[17] , \ScanLink252[16] , \wRegEnTop_3_5[0] , 
        \wRegInTop_4_14[10] , \wRegInBot_5_1[8] , \ScanLink112[31] , 
        \ScanLink131[19] , \wRegInTop_7_4[30] , \ScanLink144[29] , 
        \ScanLink182[21] , \ScanLink227[26] , \ScanLink144[30] , 
        \ScanLink167[18] , \wRegOut_6_59[7] , \wRegInTop_7_4[29] , 
        \wRegInBot_4_14[17] , \ScanLink112[28] , \wRegOut_7_78[1] , 
        \wRegInTop_7_82[24] , \wRegOut_4_6[2] , \wRegOut_6_44[8] , 
        \ScanLink139[8] , \wRegInTop_7_97[10] , \ScanLink244[2] , 
        \ScanLink3[16] , \wRegInTop_3_3[9] , \wRegInTop_3_4[27] , 
        \ScanLink19[6] , \wRegInBot_5_6[27] , \wRegInTop_6_56[0] , 
        \wRegOut_7_8[27] , \ScanLink124[7] , \wRegInTop_7_77[6] , 
        \ScanLink247[1] , \wRegOut_4_0[20] , \wRegInTop_6_55[3] , 
        \ScanLink127[4] , \wRegInTop_7_74[5] , \wRegOut_5_16[9] , 
        \wRegInBot_6_17[16] , \wRegInBot_6_18[6] , \wRegInBot_6_62[26] , 
        \wRegInTop_7_79[25] , \wRegInTop_6_21[14] , \wRegInBot_6_41[17] , 
        \wRegInTop_6_54[24] , \wRegOut_7_111[13] , \wRegOut_6_7[24] , 
        \wRegInBot_6_34[27] , \wRegInBot_6_54[23] , \wRegOut_7_104[27] , 
        \wRegInBot_6_21[13] , \wRegInTop_6_34[20] , \wRegInTop_6_41[10] , 
        \wRegOut_4_5[1] , \wRegInBot_4_9[24] , \wRegInTop_6_17[11] , 
        \wRegOut_7_127[16] , \wRegInTop_7_19[21] , \wRegInBot_5_6[14] , 
        \wRegInTop_6_62[21] , \wRegInTop_4_14[23] , \wRegInBot_4_14[24] , 
        \wRegOut_6_12[19] , \wRegOut_6_31[31] , \wRegOut_6_31[28] , 
        \wRegOut_7_8[14] , \ScanLink220[6] , \wRegOut_7_125[0] , 
        \wRegInTop_6_32[4] , \wRegOut_6_44[18] , \ScanLink140[3] , 
        \wRegInTop_7_13[2] , \wRegOut_7_69[19] , \wRegInTop_7_97[23] , 
        \wRegInBot_6_5[9] , \wRegOut_7_2[3] , \ScanLink192[5] , 
        \wRegInTop_7_82[17] , \wRegOut_1_1[4] , \ScanLink11[18] , 
        \wRegInBot_4_9[17] , \wRegInBot_4_11[9] , \wRegInBot_6_21[20] , 
        \wRegInTop_6_41[23] , \wRegOut_6_7[17] , \wRegInBot_6_54[10] , 
        \wRegInTop_6_34[13] , \wRegOut_7_1[0] , \wRegOut_7_104[14] , 
        \ScanLink32[30] , \ScanLink64[28] , \wRegInTop_6_17[22] , 
        \wRegInTop_6_62[12] , \wRegInTop_7_19[12] , \wRegOut_7_127[25] , 
        \wRegEnBot_6_32[0] , \wRegInBot_6_17[25] , \wRegInBot_6_62[15] , 
        \wRegInTop_7_79[16] , \wRegInTop_6_54[17] , \wRegOut_4_0[13] , 
        \wRegOut_4_11[18] , \ScanLink32[29] , \ScanLink47[19] , 
        \ScanLink64[31] , \wRegEnBot_6_3[0] , \wRegInBot_6_34[14] , 
        \wRegInTop_6_21[27] , \ScanLink191[6] , \wRegInBot_6_41[24] , 
        \wRegOut_7_111[20] , \wRegOut_7_126[3] , \ScanLink223[5] , 
        \wRegInTop_3_4[14] , \wRegOut_7_92[18] , \wRegInTop_7_112[18] , 
        \ScanLink0[3] , \wRegOut_1_0[19] , \wRegInBot_2_1[30] , 
        \wRegInBot_2_1[29] , \wRegInTop_4_3[30] , \wRegInTop_4_8[0] , 
        \wRegInTop_6_31[7] , \wRegInTop_7_10[1] , \ScanLink143[0] , 
        \ScanLink243[29] , \wRegInTop_4_3[29] , \wRegInBot_4_9[6] , 
        \wRegInBot_6_27[8] , \wRegInTop_7_76[22] , \ScanLink215[31] , 
        \ScanLink236[19] , \wRegInBot_6_18[11] , \wRegInTop_7_55[13] , 
        \ScanLink243[30] , \wRegInBot_4_6[23] , \ScanLink28[30] , 
        \ScanLink28[29] , \wRegOut_5_29[7] , \ScanLink215[28] , 
        \wRegOut_6_8[23] , \wRegEnTop_6_39[0] , \wRegInTop_7_20[23] , 
        \wRegInTop_7_40[27] , \ScanLink105[5] , \wRegInTop_7_35[17] , 
        \wRegInTop_7_56[4] , \wRegInTop_7_63[16] , \wRegInTop_6_18[16] , 
        \ScanLink26[8] , \wRegOut_5_26[19] , \wRegInTop_7_16[26] , 
        \wRegOut_7_59[3] , \ScanLink38[4] , \wRegInBot_5_9[20] , 
        \wRegInTop_5_26[0] , \wRegInBot_6_1[27] , \wRegInTop_7_84[2] , 
        \wRegOut_7_88[18] , \wRegInTop_7_108[18] , \wRegInBot_6_39[4] , 
        \wRegOut_7_95[9] , \wRegInTop_5_25[3] , \wRegOut_7_50[31] , 
        \wRegOut_7_73[19] , \wRegOut_7_7[20] , \wRegOut_7_25[18] , 
        \wRegInTop_7_48[8] , \wRegOut_7_50[28] , \wRegInTop_7_87[1] , 
        \wRegInTop_5_15[27] , \wRegInBot_5_23[25] , \wRegOut_7_88[6] , 
        \wRegOut_5_0[24] , \wRegInBot_5_15[20] , \ScanLink85[29] , 
        \wRegInTop_7_98[17] , \wRegInTop_5_23[22] , \ScanLink85[30] , 
        \ScanLink106[6] , \wRegInTop_7_55[7] , \ScanLink3[0] , 
        \wRegInBot_6_1[14] , \wRegInBot_4_6[10] , \wRegOut_6_8[10] , 
        \wRegInTop_7_35[24] , \wRegInTop_7_40[14] , \wRegOut_7_104[2] , 
        \wRegInTop_7_16[15] , \wRegOut_5_0[17] , \wRegInBot_5_15[13] , 
        \wRegInTop_6_13[6] , \wRegInTop_6_18[25] , \wRegOut_7_20[8] , 
        \ScanLink186[19] , \wRegInTop_7_63[25] , \ScanLink201[4] , 
        \wRegInBot_6_18[22] , \wRegInTop_7_20[10] , \wRegInTop_7_76[11] , 
        \ScanLink161[1] , \wRegInTop_7_32[0] , \wRegInTop_7_55[20] , 
        \wRegInTop_7_98[24] , \ScanLink108[28] , \ScanLink202[7] , 
        \wRegInBot_5_9[13] , \wRegInTop_5_15[14] , \wRegInTop_5_23[11] , 
        \ScanLink93[9] , \ScanLink108[31] , \wRegOut_7_107[1] , 
        \wRegInBot_5_23[16] , \wRegInTop_6_10[5] , \wRegInTop_7_31[3] , 
        \ScanLink162[2] , \wRegOut_2_3[21] , \wRegOut_2_3[12] , 
        \wRegInBot_3_5[15] , \wRegOut_4_4[18] , \wRegInBot_6_21[6] , 
        \wRegOut_7_7[13] , \wRegInTop_7_120[16] , \ScanLink15[13] , 
        \ScanLink20[6] , \ScanLink23[16] , \wRegOut_4_15[13] , 
        \wRegOut_6_63[4] , \wRegOut_7_42[2] , \wRegInTop_7_103[27] , 
        \wRegOut_5_8[2] , \wRegOut_7_83[27] , \ScanLink56[26] , 
        \wRegOut_7_96[13] , \wRegInTop_7_116[13] , \wRegInTop_6_45[28] , 
        \wRegOut_4_13[0] , \wRegInTop_7_68[30] , \ScanLink60[23] , 
        \ScanLink75[17] , \wRegInTop_6_13[30] , \wRegInTop_6_30[18] , 
        \wRegInTop_6_13[29] , \wRegInTop_6_45[31] , \ScanLink228[12] , 
        \wRegInTop_7_68[29] , \wRegOut_7_90[4] , \ScanLink198[21] , 
        \ScanLink248[16] , \ScanLink23[5] , \wRegInTop_4_8[16] , 
        \ScanLink43[12] , \ScanLink36[22] , \ScanLink103[24] , 
        \wRegInTop_7_93[28] , \ScanLink120[15] , \ScanLink176[14] , 
        \wRegOut_7_93[7] , \wRegInTop_7_93[31] , \wRegOut_4_10[3] , 
        \ScanLink155[25] , \wRegInTop_4_10[31] , \wRegOut_5_31[5] , 
        \wRegInTop_4_10[28] , \ScanLink135[21] , \ScanLink140[11] , 
        \ScanLink116[10] , \wRegInTop_7_0[11] , \ScanLink163[20] , 
        \wRegInBot_3_5[26] , \ScanLink15[20] , \wRegInTop_5_7[15] , 
        \wRegOut_6_20[17] , \wRegInBot_6_22[5] , \wRegOut_6_60[7] , 
        \wRegOut_7_41[1] , \wRegOut_7_78[26] , \wRegOut_6_35[23] , 
        \wRegOut_6_55[27] , \ScanLink100[8] , \wRegOut_6_40[13] , 
        \wRegOut_6_16[12] , \wRegInTop_7_53[9] , \wRegOut_6_63[22] , 
        \wRegOut_7_18[22] , \ScanLink248[25] , \ScanLink23[25] , 
        \wRegInTop_4_8[25] , \wRegInBot_5_14[0] , \ScanLink60[10] , 
        \ScanLink198[12] , \ScanLink36[11] , \wRegOut_7_115[18] , 
        \ScanLink43[21] , \ScanLink44[2] , \wRegInBot_6_50[28] , 
        \wRegOut_4_15[20] , \ScanLink56[15] , \ScanLink75[24] , 
        \wRegInBot_6_25[18] , \wRegInBot_6_50[31] , \wRegInTop_7_29[1] , 
        \wRegInTop_6_15[8] , \ScanLink96[4] , \wRegInBot_6_45[2] , 
        \ScanLink228[21] , \wRegOut_7_26[6] , \wRegOut_7_96[20] , 
        \wRegInTop_7_116[20] , \wRegInTop_7_120[25] , \wRegInTop_7_103[14] , 
        \wRegInTop_5_7[26] , \wRegOut_7_83[14] , \wRegOut_6_16[21] , 
        \ScanLink95[7] , \wRegOut_6_40[20] , \wRegOut_6_35[10] , 
        \wRegInBot_6_46[1] , \wRegOut_7_18[11] , \wRegOut_6_63[11] , 
        \wRegOut_7_25[5] , \ScanLink204[9] , \wRegInTop_5_3[17] , 
        \ScanLink47[1] , \wRegInBot_5_17[3] , \wRegOut_6_20[24] , 
        \wRegOut_6_55[14] , \wRegOut_7_78[15] , \ScanLink140[22] , 
        \wRegInBot_5_28[29] , \ScanLink88[8] , \ScanLink135[12] , 
        \wRegInBot_5_28[30] , \ScanLink116[23] , \wRegInTop_7_0[22] , 
        \ScanLink163[13] , \wRegEnTop_7_64[0] , \ScanLink219[6] , 
        \wRegOut_6_31[21] , \ScanLink103[17] , \ScanLink176[27] , 
        \ScanLink120[26] , \ScanLink155[16] , \ScanLink179[3] , 
        \wRegOut_6_44[11] , \wRegInTop_6_4[6] , \wRegInBot_6_5[0] , 
        \wRegOut_6_12[10] , \wRegOut_7_69[10] , \wRegOut_6_20[5] , 
        \wRegInBot_6_62[7] , \wRegOut_6_24[15] , \wRegOut_6_51[25] , 
        \wRegOut_7_125[9] , \ScanLink131[23] , \wRegEnTop_7_92[0] , 
        \ScanLink112[12] , \ScanLink144[13] , \wRegOut_0_0[14] , 
        \ScanLink107[26] , \wRegInTop_7_4[13] , \ScanLink167[22] , 
        \ScanLink172[16] , \ScanLink11[11] , \wRegInBot_4_12[3] , 
        \wRegInTop_7_112[6] , \ScanLink63[7] , \ScanLink124[17] , 
        \ScanLink64[21] , \wRegEnTop_6_61[0] , \ScanLink151[27] , 
        \ScanLink239[24] , \wRegInBot_4_11[0] , \ScanLink32[20] , 
        \ScanLink47[10] , \wRegInBot_6_6[3] , \wRegOut_7_111[30] , 
        \wRegInTop_6_7[5] , \ScanLink52[24] , \wRegInBot_6_21[29] , 
        \wRegOut_7_111[29] , \ScanLink27[14] , \wRegInBot_5_30[6] , 
        \wRegInTop_7_111[5] , \ScanLink60[4] , \wRegInBot_6_54[19] , 
        \wRegOut_5_29[24] , \ScanLink71[15] , \wRegInBot_6_21[30] , 
        \wRegOut_7_1[9] , \ScanLink189[17] , \wRegOut_7_92[11] , 
        \wRegInTop_7_112[11] , \wRegOut_0_0[27] , \wRegInTop_3_0[3] , 
        \wRegInBot_3_1[17] , \wRegInBot_6_61[4] , \wRegInTop_7_10[8] , 
        \ScanLink143[9] , \wRegInTop_7_124[14] , \wRegOut_4_11[11] , 
        \wRegOut_6_23[6] , \ScanLink172[25] , \wRegOut_7_87[25] , 
        \wRegInTop_7_107[25] , \wRegInBot_3_1[5] , \wRegInTop_7_97[19] , 
        \ScanLink107[15] , \ScanLink151[14] , \wRegInBot_3_1[24] , 
        \wRegOut_4_0[30] , \wRegInTop_4_14[19] , \wRegInBot_5_1[1] , 
        \wRegOut_5_15[3] , \ScanLink124[24] , \ScanLink139[1] , 
        \ScanLink144[20] , \ScanLink131[10] , \wRegInTop_7_4[20] , 
        \ScanLink167[11] , \ScanLink112[21] , \wRegOut_7_78[8] , 
        \wRegInTop_5_0[7] , \wRegInTop_5_3[24] , \wRegOut_6_24[26] , 
        \wRegOut_6_51[16] , \wRegInTop_6_56[9] , \wRegOut_6_12[23] , 
        \wRegOut_6_31[12] , \wRegOut_6_44[22] , \wRegOut_6_44[1] , 
        \wRegOut_7_65[7] , \wRegOut_7_69[23] , \wRegInTop_7_124[27] , 
        \wRegOut_4_11[22] , \wRegInTop_7_107[16] , \wRegOut_4_0[29] , 
        \wRegInTop_5_19[7] , \wRegOut_7_87[16] , \wRegOut_5_29[17] , 
        \wRegOut_6_47[2] , \wRegOut_7_92[22] , \wRegInTop_7_112[22] , 
        \wRegOut_7_66[4] , \ScanLink247[8] , \wRegInBot_0_0[9] , 
        \wRegInTop_2_0[21] , \wRegInBot_3_2[6] , \wRegInTop_3_3[0] , 
        \ScanLink27[27] , \ScanLink52[17] , \wRegInTop_6_34[29] , 
        \wRegInTop_6_41[19] , \wRegInTop_6_48[5] , \wRegInTop_7_19[31] , 
        \wRegInTop_6_62[31] , \wRegInTop_7_69[3] , \ScanLink71[26] , 
        \wRegInTop_6_17[18] , \wRegInTop_6_34[30] , \wRegInTop_7_19[28] , 
        \ScanLink189[24] , \ScanLink11[22] , \wRegOut_4_5[8] , 
        \wRegInTop_6_62[28] , \wRegInBot_5_2[2] , \ScanLink32[13] , 
        \wRegInTop_5_3[4] , \ScanLink64[12] , \ScanLink239[17] , 
        \wRegOut_5_4[26] , \ScanLink47[23] , \wRegOut_5_16[0] , 
        \wRegInBot_5_11[22] , \ScanLink179[29] , \wRegEnTop_7_103[0] , 
        \wRegInTop_5_27[20] , \wRegInBot_5_27[27] , \wRegInBot_5_28[4] , 
        \wRegInTop_6_34[3] , \wRegInTop_7_15[5] , \ScanLink146[4] , 
        \ScanLink179[30] , \wRegInTop_7_109[7] , \wRegOut_7_123[7] , 
        \ScanLink78[6] , \ScanLink8[20] , \wRegInTop_5_11[25] , 
        \wRegInTop_7_89[21] , \ScanLink226[1] , \wRegInTop_5_8[31] , 
        \wRegInTop_5_8[28] , \wRegInTop_6_2[8] , \wRegOut_7_3[22] , 
        \ScanLink194[2] , \wRegInTop_7_114[8] , \ScanLink65[9] , 
        \wRegOut_7_4[4] , \wRegEnTop_5_28[0] , \wRegInBot_6_5[25] , 
        \wRegOut_6_38[7] , \wRegOut_7_19[1] , \ScanLink158[8] , 
        \ScanLink197[1] , \wRegOut_7_7[7] , \wRegInBot_1_0[6] , 
        \ScanLink2[26] , \wRegOut_2_0[1] , \wRegOut_4_0[5] , 
        \wRegInBot_4_2[21] , \wRegInTop_6_37[0] , \wRegInTop_7_16[6] , 
        \wRegInTop_7_31[15] , \wRegInTop_7_44[25] , \ScanLink145[7] , 
        \ScanLink182[31] , \wRegInTop_7_67[14] , \wRegOut_6_25[8] , 
        \wRegInTop_7_12[24] , \ScanLink182[28] , \wRegInTop_7_72[20] , 
        \wRegEnBot_6_53[0] , \wRegInTop_7_24[21] , \wRegInTop_7_51[11] , 
        \ScanLink225[2] , \wRegOut_7_120[4] , \wRegInTop_2_0[12] , 
        \ScanLink8[13] , \wRegInTop_5_6[9] , \wRegOut_7_77[28] , 
        \wRegInBot_5_27[14] , \wRegOut_7_3[11] , \wRegOut_7_21[30] , 
        \wRegOut_7_54[19] , \wRegOut_7_77[31] , \wRegOut_7_21[29] , 
        \wRegOut_2_3[2] , \wRegInBot_3_4[8] , \wRegInBot_4_2[12] , 
        \wRegInTop_4_7[18] , \wRegOut_5_4[15] , \wRegInTop_5_11[16] , 
        \wRegInTop_6_50[7] , \ScanLink122[0] , \wRegInTop_7_71[1] , 
        \wRegInTop_7_89[12] , \wRegInBot_5_11[11] , \ScanLink81[18] , 
        \wRegOut_7_63[9] , \ScanLink242[5] , \wRegInTop_5_27[13] , 
        \wRegInTop_6_53[4] , \ScanLink121[3] , \wRegInTop_7_24[12] , 
        \wRegInTop_7_72[13] , \ScanLink232[28] , \ScanLink247[18] , 
        \ScanLink211[19] , \ScanLink232[31] , \ScanLink59[28] , 
        \wRegInTop_7_31[26] , \wRegInTop_7_51[22] , \wRegInTop_7_72[2] , 
        \wRegInTop_7_12[17] , \wRegInTop_7_44[16] , \wRegOut_4_3[6] , 
        \wRegOut_5_22[31] , \ScanLink59[31] , \wRegInTop_7_67[27] , 
        \ScanLink241[6] , \wRegOut_5_22[28] , \wRegInBot_6_5[16] , 
        \ScanLink10[31] , \wRegInBot_4_8[27] , \wRegEnTop_5_0[0] , 
        \wRegInTop_6_16[12] , \wRegOut_7_126[15] , \wRegInTop_5_14[2] , 
        \wRegInTop_6_63[22] , \wRegInTop_7_18[22] , \wRegOut_6_6[27] , 
        \wRegInBot_6_55[20] , \wRegOut_7_105[24] , \wRegInTop_6_20[17] , 
        \wRegInBot_6_20[10] , \wRegInTop_6_35[23] , \wRegInTop_6_40[13] , 
        \wRegInTop_7_79[9] , \wRegInBot_6_40[14] , \ScanLink10[28] , 
        \ScanLink33[19] , \ScanLink46[29] , \wRegInTop_6_55[27] , 
        \wRegOut_7_110[10] , \wRegInBot_6_35[24] , \wRegInTop_7_78[26] , 
        \wRegInTop_3_5[24] , \wRegOut_4_1[23] , \ScanLink46[30] , 
        \wRegInBot_6_16[15] , \wRegInBot_6_63[25] , \ScanLink65[18] , 
        \wRegOut_4_10[31] , \wRegOut_4_10[28] , \wRegInTop_6_45[0] , 
        \ScanLink137[7] , \wRegInTop_7_64[6] , \wRegOut_7_93[31] , 
        \wRegInTop_7_113[31] , \wRegInTop_6_46[3] , \wRegOut_6_57[8] , 
        \wRegOut_7_93[28] , \wRegInTop_7_113[28] , \wRegOut_7_9[24] , 
        \ScanLink134[4] , \wRegInTop_7_67[5] , \ScanLink2[15] , 
        \wRegInTop_3_5[17] , \ScanLink17[9] , \wRegInTop_4_15[13] , 
        \wRegInBot_4_15[14] , \wRegInBot_5_7[24] , \wRegOut_5_18[6] , 
        \wRegOut_6_13[29] , \wRegInBot_6_16[9] , \wRegOut_6_45[31] , 
        \wRegOut_7_68[29] , \ScanLink254[1] , \wRegOut_6_45[28] , 
        \wRegOut_7_68[30] , \wRegOut_6_13[30] , \wRegOut_6_30[18] , 
        \wRegInTop_5_17[1] , \wRegOut_6_49[4] , \wRegInTop_7_96[13] , 
        \wRegOut_7_68[2] , \wRegInTop_7_83[27] , \wRegOut_4_1[10] , 
        \wRegInTop_6_21[4] , \ScanLink153[3] , \wRegInBot_4_8[14] , 
        \wRegInBot_6_16[26] , \wRegInTop_6_20[24] , \wRegInBot_6_35[17] , 
        \wRegInTop_6_55[14] , \ScanLink233[6] , \wRegInBot_6_40[27] , 
        \ScanLink181[5] , \wRegOut_7_110[23] , \wRegInBot_6_63[16] , 
        \wRegInTop_7_18[11] , \wRegInTop_7_78[15] , \wRegInTop_4_15[20] , 
        \wRegOut_6_6[14] , \wRegInTop_6_16[21] , \wRegInTop_6_63[11] , 
        \wRegOut_7_126[26] , \wRegInBot_6_20[23] , \wRegInTop_6_40[20] , 
        \wRegInBot_6_55[13] , \wRegInTop_6_35[10] , \wRegOut_7_105[17] , 
        \ScanLink113[18] , \ScanLink130[30] , \wRegInBot_4_15[27] , 
        \wRegEnBot_6_21[0] , \wRegInTop_7_83[14] , \ScanLink130[29] , 
        \wRegInTop_7_5[19] , \ScanLink166[28] , \ScanLink145[19] , 
        \ScanLink166[31] , \ScanLink182[6] , \wRegInTop_7_96[20] , 
        \wRegInBot_5_7[17] , \wRegInBot_6_8[5] , \wRegInTop_6_9[3] , 
        \wRegInTop_6_22[7] , \ScanLink150[0] , \wRegOut_7_9[17] , 
        \wRegOut_1_1[13] , \wRegInBot_2_0[10] , \wRegInTop_2_1[18] , 
        \wRegOut_3_2[15] , \ScanLink12[4] , \wRegOut_5_15[27] , 
        \wRegOut_5_23[22] , \wRegOut_7_11[9] , \ScanLink230[5] , 
        \wRegInTop_6_1[16] , \wRegOut_7_98[17] , \wRegInTop_7_118[17] , 
        \wRegInTop_4_6[12] , \ScanLink131[9] , \wRegInTop_7_25[18] , 
        \ScanLink210[13] , \wRegInTop_7_50[28] , \wRegInTop_7_62[8] , 
        \ScanLink38[26] , \wRegInBot_5_9[9] , \wRegInBot_6_13[4] , 
        \wRegInTop_7_50[31] , \ScanLink196[25] , \ScanLink233[22] , 
        \ScanLink246[12] , \wRegInTop_7_73[19] , \wRegInBot_4_3[18] , 
        \ScanLink58[22] , \wRegOut_6_51[6] , \ScanLink183[11] , 
        \ScanLink226[16] , \wRegOut_7_70[0] , \ScanLink253[26] , 
        \ScanLink95[26] , \ScanLink118[14] , \ScanLink205[27] , 
        \wRegInTop_7_88[18] , \ScanLink9[19] , \ScanLink11[7] , 
        \wRegInTop_5_9[11] , \wRegInTop_5_26[19] , \wRegInBot_6_10[7] , 
        \ScanLink80[12] , \wRegOut_6_52[5] , \wRegOut_6_18[16] , 
        \ScanLink178[10] , \wRegOut_7_73[3] , \wRegOut_7_63[16] , 
        \wRegOut_7_16[26] , \wRegOut_7_35[17] , \wRegOut_7_40[27] , 
        \wRegEnTop_6_13[0] , \wRegOut_7_55[13] , \wRegOut_7_20[23] , 
        \wRegOut_7_76[22] , \wRegOut_3_2[26] , \ScanLink253[15] , 
        \wRegInTop_4_6[21] , \ScanLink58[11] , \ScanLink183[22] , 
        \ScanLink226[25] , \ScanLink205[14] , \ScanLink38[15] , 
        \wRegInBot_5_8[19] , \wRegInTop_5_9[22] , \wRegOut_5_15[14] , 
        \wRegOut_6_35[2] , \wRegOut_7_14[4] , \ScanLink210[20] , 
        \ScanLink233[11] , \ScanLink235[8] , \ScanLink246[21] , 
        \ScanLink196[16] , \wRegOut_5_23[11] , \wRegInBot_5_26[2] , 
        \ScanLink148[2] , \wRegInTop_7_107[1] , \wRegInBot_5_25[1] , 
        \wRegInTop_6_1[25] , \ScanLink76[0] , \wRegOut_7_98[24] , 
        \wRegOut_6_18[25] , \wRegInTop_6_39[6] , \wRegOut_7_2[28] , 
        \ScanLink228[7] , \wRegInTop_7_118[24] , \wRegInTop_7_18[0] , 
        \wRegOut_7_20[10] , \wRegOut_7_55[20] , \ScanLink184[8] , 
        \wRegOut_7_2[31] , \wRegOut_7_16[15] , \wRegOut_7_76[11] , 
        \wRegOut_7_63[25] , \wRegOut_7_35[24] , \wRegInTop_7_104[2] , 
        \wRegInBot_5_10[31] , \ScanLink75[3] , \wRegOut_7_40[14] , 
        \wRegInBot_5_10[28] , \ScanLink80[21] , \wRegInTop_6_24[9] , 
        \ScanLink199[7] , \ScanLink178[23] , \ScanLink51[5] , \ScanLink95[15] , 
        \wRegOut_6_36[1] , \ScanLink118[27] , \wRegOut_7_17[7] , 
        \wRegOut_7_6[19] , \wRegOut_7_9[1] , \wRegOut_7_51[11] , 
        \wRegInTop_7_120[4] , \wRegOut_7_24[21] , \wRegInBot_5_14[19] , 
        \ScanLink83[3] , \wRegInTop_7_2[7] , \wRegOut_7_12[24] , 
        \wRegOut_7_67[14] , \wRegOut_7_72[20] , \wRegOut_7_44[25] , 
        \wRegOut_7_31[15] , \ScanLink109[22] , \wRegInBot_6_50[5] , 
        \wRegOut_3_6[17] , \wRegOut_6_12[7] , \ScanLink84[10] , 
        \wRegOut_7_33[1] , \ScanLink91[24] , \ScanLink169[26] , 
        \wRegInBot_6_53[6] , \wRegInTop_7_21[9] , \ScanLink172[8] , 
        \wRegInTop_4_2[10] , \ScanLink29[10] , \wRegOut_6_11[4] , 
        \ScanLink187[13] , \ScanLink222[14] , \wRegOut_7_30[2] , 
        \ScanLink201[25] , \wRegOut_7_114[8] , \ScanLink49[14] , 
        \ScanLink80[0] , \wRegInBot_6_19[31] , \ScanLink214[11] , 
        \wRegOut_5_11[25] , \wRegInBot_6_19[28] , \ScanLink192[27] , 
        \ScanLink237[20] , \ScanLink242[10] , \wRegOut_7_89[21] , 
        \wRegInTop_7_109[21] , \wRegOut_6_7[8] , \wRegOut_1_1[20] , 
        \wRegInTop_1_1[0] , \ScanLink52[6] , \wRegOut_7_109[7] , 
        \wRegInTop_7_123[7] , \wRegInBot_2_0[23] , \wRegInTop_5_22[28] , 
        \wRegOut_5_27[20] , \wRegInTop_7_1[4] , \wRegInTop_6_5[14] , 
        \ScanLink91[17] , \wRegInBot_6_34[1] , \ScanLink169[15] , 
        \wRegOut_7_57[5] , \ScanLink84[23] , \wRegInBot_4_4[3] , 
        \wRegInTop_4_5[5] , \wRegInTop_4_6[6] , \wRegInTop_5_22[31] , 
        \wRegInTop_5_28[6] , \ScanLink109[11] , \wRegOut_7_12[17] , 
        \wRegInBot_4_7[0] , \wRegOut_7_67[27] , \wRegOut_7_85[3] , 
        \ScanLink35[1] , \wRegEnTop_7_16[0] , \wRegOut_7_31[26] , 
        \ScanLink36[2] , \wRegOut_5_24[2] , \wRegOut_5_27[13] , 
        \wRegOut_5_27[1] , \wRegOut_7_44[16] , \wRegOut_7_24[12] , 
        \wRegOut_7_51[22] , \wRegInTop_7_58[2] , \wRegOut_7_72[13] , 
        \wRegInTop_6_5[27] , \wRegOut_7_49[9] , \wRegOut_7_86[0] , 
        \wRegOut_5_3[9] , \wRegInTop_7_109[12] , \wRegOut_5_11[16] , 
        \wRegOut_7_89[12] , \wRegOut_2_2[18] , \ScanLink6[24] , 
        \wRegOut_3_6[24] , \wRegInTop_4_2[23] , \ScanLink108[0] , 
        \wRegInTop_7_77[31] , \wRegInTop_7_94[8] , \wRegInBot_4_7[29] , 
        \ScanLink49[27] , \wRegInTop_7_21[29] , \wRegInTop_7_54[19] , 
        \ScanLink214[22] , \wRegOut_6_9[30] , \wRegInBot_6_37[2] , 
        \wRegInTop_7_77[28] , \ScanLink242[23] , \wRegInTop_7_21[30] , 
        \wRegOut_7_54[6] , \ScanLink192[14] , \ScanLink237[13] , 
        \wRegInBot_4_7[30] , \ScanLink29[23] , \ScanLink187[20] , 
        \ScanLink222[27] , \wRegOut_6_9[29] , \wRegInTop_4_11[11] , 
        \wRegInTop_7_1[28] , \ScanLink141[31] , \ScanLink162[19] , 
        \ScanLink201[16] , \wRegInTop_7_89[7] , \wRegInBot_4_11[16] , 
        \wRegInTop_5_29[24] , \wRegInBot_5_29[23] , \wRegOut_6_2[5] , 
        \ScanLink117[29] , \wRegInTop_7_1[31] , \ScanLink141[28] , 
        \wRegOut_7_28[0] , \wRegInTop_7_87[25] , \ScanLink98[2] , 
        \ScanLink134[18] , \ScanLink117[30] , \wRegInTop_7_4[9] , 
        \ScanLink169[9] , \wRegOut_6_14[9] , \ScanLink214[3] , 
        \wRegInTop_7_92[11] , \wRegInTop_7_27[7] , \wRegOut_7_111[5] , 
        \ScanLink174[6] , \wRegInTop_3_1[26] , \wRegInBot_5_3[26] , 
        \ScanLink49[7] , \wRegInBot_5_19[5] , \wRegOut_7_112[6] , 
        \wRegOut_4_5[21] , \wRegInBot_6_55[8] , \ScanLink217[0] , 
        \ScanLink54[8] , \wRegOut_6_1[6] , \wRegInTop_6_24[15] , 
        \wRegInTop_7_24[4] , \ScanLink177[5] , \wRegInTop_7_125[9] , 
        \wRegInBot_6_44[16] , \wRegOut_7_114[12] , \wRegOut_6_2[25] , 
        \wRegInTop_6_12[10] , \wRegInBot_6_12[17] , \wRegInBot_6_31[26] , 
        \wRegInTop_6_51[25] , \wRegInBot_6_48[7] , \ScanLink199[18] , 
        \wRegInTop_7_69[10] , \wRegOut_7_122[17] , \wRegOut_7_101[26] , 
        \wRegInBot_6_24[12] , \wRegInTop_6_31[21] , \wRegInBot_6_51[22] , 
        \wRegEnTop_7_2[0] , \wRegInTop_6_44[11] , \ScanLink6[17] , 
        \wRegInBot_5_3[15] , \wRegOut_3_5[3] , \wRegOut_3_6[0] , 
        \wRegInTop_4_0[8] , \wRegInTop_5_29[17] , \wRegEnBot_5_30[0] , 
        \wRegOut_6_17[18] , \wRegOut_6_34[30] , \wRegOut_6_34[29] , 
        \wRegOut_6_62[28] , \wRegOut_7_19[28] , \wRegOut_6_41[19] , 
        \ScanLink110[2] , \wRegOut_7_19[31] , \wRegOut_6_62[31] , 
        \wRegInTop_6_62[5] , \wRegInTop_7_43[3] , \wRegInTop_7_92[22] , 
        \wRegInBot_4_11[25] , \wRegInTop_4_11[22] , \wRegInTop_4_12[1] , 
        \wRegOut_5_6[4] , \wRegInTop_7_87[16] , \wRegInBot_5_29[10] , 
        \wRegInTop_7_69[23] , \wRegInTop_7_91[5] , \ScanLink229[18] , 
        \wRegOut_7_122[24] , \wRegInTop_6_12[23] , \wRegInBot_6_24[21] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[11] , \wRegOut_1_1[31] , 
        \wRegOut_1_1[28] , \wRegInTop_2_1[23] , \wRegInBot_2_2[9] , 
        \ScanLink37[28] , \ScanLink42[18] , \ScanLink61[30] , 
        \wRegOut_6_2[16] , \wRegInTop_6_44[22] , \wRegInTop_6_31[12] , 
        \wRegInBot_6_51[11] , \wRegOut_7_101[15] , \wRegInBot_6_31[15] , 
        \wRegInTop_6_51[16] , \wRegInTop_6_24[26] , \wRegOut_7_114[21] , 
        \wRegInBot_6_44[25] , \wRegInTop_7_92[6] , \wRegInBot_3_0[26] , 
        \wRegInBot_3_0[15] , \wRegInTop_3_1[15] , \ScanLink14[19] , 
        \wRegInTop_4_11[2] , \wRegOut_5_5[7] , \ScanLink61[29] , 
        \wRegInBot_6_12[24] , \ScanLink37[31] , \wRegInTop_5_30[4] , 
        \wRegOut_4_5[12] , \wRegOut_4_14[19] , \wRegOut_7_52[8] , 
        \wRegInTop_4_15[31] , \ScanLink113[1] , \wRegInTop_6_61[6] , 
        \wRegInTop_7_40[0] , \wRegOut_7_97[19] , \wRegInTop_7_117[19] , 
        \wRegInTop_4_15[28] , \ScanLink130[21] , \ScanLink145[11] , 
        \wRegInTop_5_2[15] , \wRegInBot_5_23[7] , \ScanLink106[24] , 
        \ScanLink113[10] , \wRegInTop_7_5[11] , \ScanLink166[20] , 
        \ScanLink125[15] , \ScanLink173[14] , \wRegInTop_7_96[28] , 
        \wRegInTop_7_102[4] , \ScanLink73[5] , \ScanLink150[25] , 
        \wRegInTop_7_96[31] , \wRegOut_6_30[23] , \wRegOut_6_45[13] , 
        \wRegEnTop_5_20[0] , \wRegOut_6_13[12] , \ScanLink150[8] , 
        \wRegOut_6_30[7] , \wRegOut_7_11[1] , \wRegOut_7_68[12] , 
        \wRegOut_5_28[26] , \wRegOut_6_25[17] , \wRegOut_6_50[27] , 
        \wRegOut_7_93[13] , \wRegInTop_7_113[13] , \wRegOut_7_86[27] , 
        \wRegInTop_7_125[16] , \ScanLink10[20] , \ScanLink10[13] , 
        \wRegOut_4_1[18] , \wRegOut_4_10[13] , \wRegOut_6_33[4] , 
        \wRegOut_7_12[2] , \wRegInTop_7_106[27] , \ScanLink65[23] , 
        \ScanLink238[26] , \ScanLink17[1] , \ScanLink26[16] , \ScanLink33[22] , 
        \ScanLink46[12] , \wRegInBot_5_20[4] , \wRegInTop_6_40[28] , 
        \wRegInTop_7_101[7] , \ScanLink53[26] , \ScanLink70[6] , 
        \wRegInTop_6_16[30] , \wRegInTop_6_35[18] , \wRegInTop_5_2[26] , 
        \ScanLink70[17] , \wRegInTop_6_40[31] , \wRegInTop_6_63[19] , 
        \ScanLink188[15] , \wRegInTop_6_16[29] , \wRegInTop_7_18[19] , 
        \wRegOut_6_25[24] , \wRegOut_6_50[14] , \wRegEnTop_5_8[0] , 
        \wRegInBot_6_16[1] , \wRegOut_6_30[10] , \wRegOut_6_45[20] , 
        \wRegInTop_5_17[9] , \wRegOut_6_13[21] , \ScanLink106[17] , 
        \wRegOut_6_54[3] , \ScanLink173[27] , \wRegOut_7_68[21] , 
        \wRegOut_7_75[5] , \ScanLink254[9] , \ScanLink125[26] , 
        \ScanLink129[3] , \ScanLink150[16] , \ScanLink145[22] , 
        \ScanLink26[25] , \ScanLink113[23] , \ScanLink130[12] , 
        \wRegEnTop_7_34[0] , \wRegInTop_7_5[22] , \ScanLink166[13] , 
        \wRegInBot_6_55[28] , \ScanLink249[6] , \ScanLink53[15] , 
        \wRegInTop_6_58[7] , \wRegInTop_7_79[1] , \ScanLink70[24] , 
        \wRegInBot_6_20[18] , \wRegInBot_6_55[31] , \ScanLink188[26] , 
        \ScanLink14[2] , \ScanLink33[11] , \ScanLink65[10] , \wCtrlOut_3[0] , 
        \wRegOut_7_110[18] , \ScanLink238[15] , \ScanLink46[21] , 
        \wRegOut_4_10[20] , \wRegInTop_6_45[8] , \wRegInTop_7_125[25] , 
        \wRegOut_7_86[14] , \wRegInTop_7_106[14] , \ScanLink9[22] , 
        \wRegOut_4_8[5] , \wRegOut_5_28[15] , \wRegInBot_6_15[2] , 
        \wRegInTop_7_113[20] , \wRegOut_6_57[0] , \wRegOut_7_93[20] , 
        \wRegOut_7_76[6] , \wRegOut_5_5[24] , \wRegInBot_5_25[9] , 
        \wRegOut_7_2[20] , \wRegOut_7_20[18] , \wRegOut_7_55[31] , 
        \wRegOut_7_76[19] , \wRegInTop_7_18[8] , \wRegOut_7_55[28] , 
        \ScanLink184[0] , \wRegInBot_5_10[20] , \ScanLink80[29] , 
        \wRegInTop_5_26[22] , \ScanLink80[30] , \wRegInTop_6_24[1] , 
        \ScanLink156[6] , \wRegInTop_7_119[5] , \wRegInTop_2_1[10] , 
        \wRegInBot_4_3[23] , \wRegInTop_5_10[27] , \wRegInBot_5_26[25] , 
        \ScanLink68[4] , \wRegOut_7_9[9] , \ScanLink58[19] , \wRegOut_6_36[9] , 
        \ScanLink155[5] , \wRegInTop_7_45[27] , \wRegInTop_7_88[23] , 
        \ScanLink236[3] , \wRegInTop_6_27[2] , \wRegInTop_7_30[17] , 
        \wRegInTop_7_66[16] , \wRegInTop_4_6[30] , \wRegInTop_7_13[26] , 
        \wRegInTop_4_6[29] , \wRegInTop_7_50[13] , \wRegInTop_7_73[22] , 
        \ScanLink210[31] , \ScanLink246[29] , \ScanLink233[19] , 
        \ScanLink235[0] , \wRegOut_5_23[19] , \wRegInBot_6_4[27] , 
        \wRegInTop_7_25[23] , \ScanLink246[30] , \ScanLink210[28] , 
        \ScanLink76[8] , \wRegOut_6_28[5] , \ScanLink187[3] , 
        \wRegInTop_7_107[9] , \ScanLink9[11] , \wRegOut_5_5[17] , 
        \wRegInTop_5_10[14] , \wRegEnBot_5_12[0] , \wRegInBot_5_26[16] , 
        \wRegInTop_6_40[5] , \ScanLink132[2] , \wRegInTop_7_61[3] , 
        \wRegInTop_7_88[10] , \wRegInBot_5_10[13] , \ScanLink178[18] , 
        \ScanLink252[7] , \wRegInTop_5_9[19] , \wRegInTop_5_26[11] , 
        \wRegInTop_5_11[7] , \wRegOut_3_3[5] , \wRegInBot_4_3[10] , 
        \wRegInTop_5_12[4] , \wRegOut_7_2[13] , \wRegInBot_6_4[14] , 
        \wRegInTop_6_43[6] , \wRegInTop_7_25[10] , \wRegInTop_7_73[11] , 
        \ScanLink131[1] , \wRegInTop_7_50[20] , \wRegInTop_7_62[0] , 
        \wRegInTop_7_13[15] , \wRegInTop_7_30[24] , \wRegInTop_7_45[14] , 
        \ScanLink183[19] , \wRegInTop_5_8[7] , \wRegInBot_5_9[1] , 
        \wRegOut_7_70[8] , \ScanLink251[4] , \wRegInTop_7_66[25] , 
        \ScanLink108[8] , \wRegOut_7_49[1] , \wRegOut_7_86[8] , 
        \wRegInTop_7_94[0] , \wRegOut_5_3[1] , \wRegInBot_6_0[25] , 
        \wRegInTop_1_1[8] , \wRegEnTop_2_3[0] , \wRegOut_3_0[6] , 
        \wRegInBot_4_7[21] , \wRegOut_6_9[21] , \wRegInBot_6_19[13] , 
        \wRegInTop_7_77[20] , \wRegInTop_7_21[21] , \wRegInTop_7_54[11] , 
        \wRegInTop_6_19[14] , \ScanLink115[7] , \wRegInTop_7_41[25] , 
        \ScanLink187[31] , \wRegInTop_7_34[15] , \wRegInTop_7_46[6] , 
        \ScanLink187[28] , \wRegInTop_7_62[14] , \ScanLink28[6] , 
        \wRegInTop_7_17[24] , \wRegOut_5_1[26] , \wRegInTop_5_14[25] , 
        \wRegInBot_5_22[27] , \wRegInBot_6_34[9] , \wRegOut_7_98[4] , 
        \ScanLink35[9] , \wRegInBot_5_14[22] , \ScanLink109[19] , 
        \wRegInTop_5_22[20] , \wRegInTop_7_99[15] , \wRegOut_5_27[9] , 
        \ScanLink116[4] , \wRegInTop_7_45[5] , \wRegInBot_6_29[6] , 
        \wRegInBot_4_7[8] , \wRegInTop_4_14[7] , \wRegOut_5_0[2] , 
        \wRegInTop_4_2[18] , \wRegInBot_4_7[12] , \ScanLink29[18] , 
        \wRegInBot_5_8[22] , \ScanLink80[8] , \wRegOut_7_6[22] , 
        \wRegInTop_7_34[26] , \wRegInTop_7_97[3] , \wRegOut_7_114[0] , 
        \wRegOut_6_9[12] , \wRegInTop_7_41[16] , \wRegInTop_7_17[17] , 
        \wRegInTop_6_19[27] , \ScanLink211[6] , \wRegInBot_6_19[20] , 
        \wRegInTop_7_62[27] , \wRegInTop_7_21[12] , \wRegInTop_7_77[13] , 
        \ScanLink237[28] , \ScanLink242[18] , \ScanLink214[19] , 
        \ScanLink237[31] , \wRegInBot_6_0[16] , \wRegOut_6_7[0] , 
        \wRegInTop_7_22[2] , \ScanLink171[3] , \wRegInTop_7_54[22] , 
        \ScanLink3[8] , \wRegInTop_2_0[4] , \wRegInBot_2_0[18] , 
        \wRegInBot_5_8[11] , \wRegOut_5_27[31] , \wRegOut_7_89[30] , 
        \wRegOut_7_89[29] , \wRegInTop_7_109[30] , \wRegInTop_7_109[29] , 
        \wRegOut_5_27[28] , \wRegOut_7_72[28] , \wRegInBot_5_14[11] , 
        \wRegOut_6_4[3] , \wRegOut_7_24[30] , \wRegOut_7_51[19] , 
        \wRegOut_7_72[31] , \wRegOut_7_6[11] , \wRegOut_7_24[29] , 
        \ScanLink84[18] , \wRegOut_7_33[9] , \wRegInTop_7_99[26] , 
        \ScanLink212[5] , \wRegInBot_2_1[2] , \wRegOut_2_2[10] , 
        \wRegInBot_2_2[1] , \wRegInBot_4_2[5] , \wRegInTop_4_3[3] , 
        \ScanLink22[14] , \ScanLink30[4] , \wRegOut_5_1[15] , 
        \wRegInTop_5_14[16] , \wRegInTop_5_22[13] , \wRegOut_7_117[3] , 
        \wRegInBot_5_22[14] , \wRegInTop_7_21[1] , \ScanLink172[0] , 
        \ScanLink57[24] , \wRegInBot_6_24[29] , \wRegOut_5_22[4] , 
        \ScanLink74[15] , \wRegInBot_6_24[30] , \wRegInBot_6_51[19] , 
        \ScanLink229[10] , \wRegOut_7_80[6] , \ScanLink61[21] , 
        \ScanLink199[23] , \wRegInTop_2_3[7] , \ScanLink14[11] , 
        \wRegOut_7_114[30] , \wRegInBot_3_4[17] , \wRegInTop_4_9[14] , 
        \ScanLink37[20] , \ScanLink42[10] , \ScanLink249[14] , 
        \wRegOut_7_114[29] , \wRegInBot_6_31[4] , \wRegInTop_7_121[14] , 
        \wRegOut_7_82[25] , \wRegOut_4_14[11] , \wRegOut_7_52[0] , 
        \ScanLink113[9] , \wRegOut_7_97[11] , \wRegInTop_7_102[25] , 
        \wRegInTop_7_117[11] , \wRegInTop_7_40[8] , \wRegOut_7_79[24] , 
        \wRegOut_3_6[8] , \wRegInTop_4_0[0] , \wRegInTop_5_6[17] , 
        \wRegOut_6_21[15] , \wRegInBot_6_32[7] , \wRegOut_7_51[3] , 
        \wRegOut_6_34[21] , \wRegOut_6_54[25] , \wRegOut_6_41[11] , 
        \wRegOut_6_17[10] , \ScanLink102[26] , \wRegOut_6_62[20] , 
        \wRegOut_7_19[20] , \wRegInBot_4_1[6] , \ScanLink177[16] , 
        \wRegOut_7_83[5] , \ScanLink33[7] , \wRegOut_5_21[7] , 
        \ScanLink121[17] , \ScanLink154[27] , \wRegInBot_5_29[18] , 
        \wRegEnTop_6_31[0] , \ScanLink134[23] , \ScanLink141[13] , 
        \wRegInTop_4_12[9] , \ScanLink117[12] , \wRegInTop_7_1[13] , 
        \ScanLink162[22] , \wRegInBot_2_1[12] , \wRegOut_2_2[23] , 
        \ScanLink8[3] , \wRegInBot_6_55[0] , \wRegInTop_7_117[22] , 
        \wRegInBot_3_4[24] , \wRegOut_4_5[30] , \wRegOut_6_17[2] , 
        \wRegOut_7_97[22] , \ScanLink86[6] , \wRegOut_7_36[4] , 
        \ScanLink217[8] , \wRegInTop_7_121[27] , \wRegOut_4_5[29] , 
        \wRegOut_4_14[22] , \wRegOut_7_82[16] , \wRegInTop_7_102[16] , 
        \ScanLink14[22] , \ScanLink22[27] , \wRegInTop_4_9[27] , 
        \ScanLink37[13] , \ScanLink61[12] , \ScanLink249[27] , 
        \ScanLink199[10] , \ScanLink42[23] , \wRegInTop_7_125[1] , 
        \ScanLink54[0] , \wRegInTop_6_31[29] , \wRegInTop_7_7[2] , 
        \wRegInTop_4_11[19] , \ScanLink57[17] , \wRegInTop_6_18[5] , 
        \wRegInTop_6_44[19] , \wRegInTop_7_39[3] , \ScanLink57[3] , 
        \ScanLink74[26] , \wRegInTop_6_12[18] , \wRegInTop_6_31[30] , 
        \wRegInTop_7_69[18] , \ScanLink229[23] , \ScanLink141[20] , 
        \wRegInTop_7_126[2] , \ScanLink117[21] , \wRegInTop_7_1[20] , 
        \ScanLink134[10] , \ScanLink162[11] , \ScanLink209[4] , 
        \wRegOut_7_28[8] , \wRegInTop_5_6[24] , \ScanLink102[15] , 
        \ScanLink177[25] , \ScanLink121[24] , \wRegInTop_7_4[1] , 
        \wRegInTop_7_92[19] , \ScanLink154[14] , \ScanLink169[1] , 
        \wRegOut_6_14[1] , \wRegOut_6_17[23] , \ScanLink85[5] , 
        \wRegOut_6_34[12] , \wRegOut_6_41[22] , \wRegInBot_6_56[3] , 
        \wRegOut_6_62[13] , \wRegOut_7_19[13] , \wRegOut_7_35[7] , 
        \wRegOut_7_79[17] , \wRegInTop_5_23[19] , \wRegOut_6_9[6] , 
        \wRegOut_6_21[26] , \wRegOut_6_54[16] , \wRegOut_7_107[9] , 
        \ScanLink93[1] , \wRegInBot_6_40[7] , \ScanLink108[20] , 
        \ScanLink41[7] , \wRegInBot_5_11[5] , \ScanLink85[12] , 
        \ScanLink90[26] , \wRegOut_7_23[3] , \ScanLink168[24] , 
        \wRegEnTop_6_43[0] , \wRegOut_7_50[13] , \wRegOut_7_25[23] , 
        \wRegOut_5_10[27] , \wRegOut_7_13[26] , \wRegOut_7_66[16] , 
        \wRegOut_7_73[22] , \wRegOut_7_30[17] , \wRegOut_7_45[27] , 
        \wRegOut_7_88[23] , \wRegInTop_7_108[23] , \wRegInBot_2_1[21] , 
        \wRegOut_3_7[15] , \wRegInBot_4_6[18] , \ScanLink42[4] , 
        \wRegInBot_5_12[6] , \wRegOut_7_119[5] , \wRegOut_5_26[22] , 
        \wRegInTop_6_4[16] , \wRegInBot_6_43[4] , \ScanLink186[11] , 
        \ScanLink223[16] , \wRegInTop_4_3[12] , \ScanLink28[12] , 
        \wRegOut_6_8[18] , \ScanLink90[2] , \wRegOut_7_20[0] , 
        \ScanLink200[27] , \ScanLink48[16] , \wRegInTop_7_20[18] , 
        \wRegInTop_7_32[8] , \wRegInTop_7_55[28] , \ScanLink215[13] , 
        \ScanLink25[3] , \wRegOut_7_13[15] , \ScanLink161[9] , 
        \wRegInTop_7_55[31] , \ScanLink193[25] , \ScanLink236[22] , 
        \wRegInTop_7_76[19] , \ScanLink243[12] , \wRegOut_7_30[24] , 
        \wRegOut_7_66[25] , \wRegOut_7_95[1] , \wRegInBot_5_9[31] , 
        \wRegOut_7_7[28] , \wRegOut_7_25[10] , \wRegOut_7_45[14] , 
        \wRegInTop_7_48[0] , \wRegOut_7_50[20] , \wRegInBot_5_9[28] , 
        \wRegOut_7_7[31] , \wRegInTop_7_87[9] , \wRegOut_7_73[11] , 
        \wRegInBot_5_15[31] , \wRegInBot_6_24[3] , \ScanLink90[15] , 
        \ScanLink168[17] , \wRegOut_7_47[7] , \ScanLink85[21] , 
        \wRegOut_3_7[26] , \wRegInTop_4_3[21] , \wRegInBot_5_15[28] , 
        \ScanLink108[13] , \wRegInTop_4_8[8] , \ScanLink48[25] , 
        \wRegInBot_6_27[0] , \ScanLink215[20] , \wRegInBot_6_18[19] , 
        \ScanLink243[21] , \wRegOut_7_44[4] , \ScanLink186[22] , 
        \ScanLink193[16] , \ScanLink236[11] , \ScanLink223[25] , 
        \ScanLink26[0] , \ScanLink28[21] , \ScanLink200[14] , 
        \wRegInTop_7_99[5] , \wRegOut_4_15[6] , \wRegOut_5_26[11] , 
        \wRegOut_5_10[14] , \wRegInTop_6_4[25] , \wRegOut_7_88[10] , 
        \wRegOut_7_96[2] , \wRegInTop_7_108[10] , \wRegInTop_5_26[8] , 
        \ScanLink118[2] , \wRegOut_1_1[5] , \ScanLink3[24] , \ScanLink5[6] , 
        \ScanLink6[5] , \wRegOut_2_3[30] , \wRegOut_6_16[30] , 
        \wRegOut_6_16[29] , \wRegOut_6_40[31] , \wRegInBot_6_46[9] , 
        \wRegOut_6_63[19] , \wRegOut_7_18[19] , \wRegOut_6_40[28] , 
        \ScanLink204[1] , \wRegOut_7_101[7] , \wRegInTop_6_16[3] , 
        \wRegOut_6_35[18] , \wRegInTop_7_9[4] , \ScanLink164[4] , 
        \wRegOut_2_3[29] , \ScanLink7[26] , \wRegInTop_7_37[5] , 
        \wRegEnTop_7_121[0] , \wRegInBot_5_2[24] , \ScanLink15[31] , 
        \wRegInTop_4_10[13] , \wRegOut_6_19[4] , \wRegInTop_7_86[27] , 
        \wRegInBot_4_10[14] , \ScanLink47[9] , \wRegOut_7_38[2] , 
        \wRegInTop_5_28[26] , \wRegInBot_5_28[21] , \ScanLink88[0] , 
        \wRegInBot_6_45[14] , \wRegInTop_7_93[13] , \ScanLink15[28] , 
        \ScanLink36[19] , \ScanLink43[29] , \wRegInBot_5_14[8] , 
        \wRegOut_7_115[10] , \wRegInTop_6_25[17] , \wRegInBot_6_30[24] , 
        \wRegInTop_6_50[27] , \wRegInBot_6_58[5] , \ScanLink7[15] , 
        \wRegInTop_3_0[24] , \ScanLink43[30] , \wRegInBot_6_13[15] , 
        \ScanLink60[18] , \wRegOut_6_3[27] , \wRegInTop_6_13[12] , 
        \wRegInTop_6_30[23] , \wRegInTop_7_68[12] , \ScanLink228[29] , 
        \wRegOut_7_123[15] , \wRegInBot_6_50[20] , \wRegOut_7_100[24] , 
        \wRegInBot_6_25[10] , \wRegInTop_6_45[13] , \wRegInTop_7_29[9] , 
        \ScanLink228[30] , \wRegOut_7_96[31] , \wRegInTop_7_116[31] , 
        \wRegOut_7_102[4] , \wRegOut_4_4[23] , \ScanLink59[5] , 
        \ScanLink207[2] , \wRegOut_7_96[28] , \wRegInTop_7_116[28] , 
        \wRegInTop_4_10[20] , \wRegInBot_4_10[27] , \wRegOut_4_15[31] , 
        \wRegOut_4_15[28] , \wRegInTop_5_28[15] , \wRegInTop_6_15[0] , 
        \wRegInTop_7_34[6] , \ScanLink167[7] , \wRegInTop_7_93[20] , 
        \ScanLink116[18] , \wRegInTop_7_86[14] , \ScanLink135[30] , 
        \wRegInBot_5_2[17] , \wRegInTop_5_23[5] , \wRegInTop_7_0[19] , 
        \wRegInBot_5_28[12] , \ScanLink135[29] , \ScanLink163[28] , 
        \ScanLink140[19] , \ScanLink163[31] , \wRegInTop_7_81[7] , 
        \wRegOut_7_41[9] , \wRegInTop_3_0[17] , \wRegOut_4_4[10] , 
        \ScanLink100[0] , \wRegInTop_7_53[1] , \wRegInTop_3_3[8] , 
        \wRegInTop_3_4[26] , \wRegOut_4_0[21] , \wRegOut_4_13[8] , 
        \wRegOut_6_3[14] , \wRegInTop_6_13[21] , \ScanLink103[3] , 
        \wRegInTop_7_50[2] , \wRegInBot_6_25[23] , \wRegInTop_6_45[20] , 
        \wRegInTop_7_68[21] , \wRegOut_7_123[26] , \wRegInTop_6_30[10] , 
        \wRegInBot_6_50[13] , \wRegOut_7_100[17] , \wRegInTop_5_20[6] , 
        \wRegInBot_6_13[26] , \wRegInTop_6_25[24] , \wRegInBot_6_30[17] , 
        \wRegInBot_6_45[27] , \wRegInTop_6_50[14] , \ScanLink198[30] , 
        \wRegInTop_7_82[4] , \wRegOut_7_115[23] , \ScanLink198[29] , 
        \wRegInTop_6_55[2] , \ScanLink127[5] , \wRegInTop_7_74[4] , 
        \ScanLink19[7] , \wRegInTop_6_17[10] , \ScanLink247[0] , 
        \wRegOut_4_5[0] , \wRegInTop_6_62[20] , \wRegOut_7_127[17] , 
        \wRegOut_4_6[3] , \wRegInBot_4_9[25] , \wRegInBot_4_14[16] , 
        \wRegEnBot_5_7[0] , \wRegOut_5_16[8] , \wRegOut_6_7[25] , 
        \wRegInTop_6_34[21] , \wRegInTop_7_19[20] , \wRegOut_7_104[26] , 
        \wRegInTop_6_21[15] , \wRegInBot_6_21[12] , \wRegInTop_6_41[11] , 
        \wRegInBot_6_54[22] , \wRegInBot_6_41[16] , \wRegOut_7_111[12] , 
        \wRegInBot_6_34[26] , \wRegInTop_6_54[25] , \wRegInBot_6_62[27] , 
        \wRegInTop_7_79[24] , \wRegInBot_6_17[17] , \wRegInBot_6_18[7] , 
        \ScanLink139[9] , \wRegInTop_4_14[11] , \wRegInBot_5_1[9] , 
        \wRegInTop_7_97[11] , \wRegInTop_7_4[28] , \ScanLink144[31] , 
        \ScanLink167[19] , \wRegInTop_7_82[25] , \ScanLink112[30] , 
        \ScanLink112[29] , \wRegOut_6_59[6] , \ScanLink131[18] , 
        \wRegInTop_7_4[31] , \wRegOut_7_78[0] , \ScanLink144[28] , 
        \wRegInTop_6_56[1] , \ScanLink124[6] , \wRegOut_7_8[26] , 
        \wRegInTop_7_77[7] , \wRegInBot_5_6[26] , \ScanLink47[18] , 
        \ScanLink64[30] , \wRegInBot_6_34[15] , \wRegOut_6_44[9] , 
        \ScanLink244[3] , \ScanLink11[19] , \ScanLink32[31] , \ScanLink32[28] , 
        \wRegInTop_6_54[16] , \wRegOut_7_111[21] , \ScanLink64[29] , 
        \wRegInTop_6_21[26] , \wRegInBot_6_41[25] , \ScanLink191[7] , 
        \wRegInBot_6_17[24] , \wRegInBot_6_62[14] , \wRegInTop_3_4[15] , 
        \wRegInBot_4_9[16] , \wRegInTop_6_62[13] , \wRegInTop_7_79[17] , 
        \wRegInTop_7_19[13] , \wRegInBot_4_11[8] , \wRegInTop_6_17[23] , 
        \wRegInTop_6_41[22] , \wRegOut_7_127[24] , \wRegOut_6_7[16] , 
        \wRegInBot_6_21[21] , \wRegInTop_6_34[12] , \wRegOut_7_1[1] , 
        \wRegInBot_6_54[11] , \wRegOut_7_104[15] , \wRegInTop_6_31[6] , 
        \wRegInTop_7_10[0] , \ScanLink143[1] , \ScanLink3[17] , 
        \wRegOut_4_0[12] , \wRegOut_4_11[19] , \wRegOut_7_92[19] , 
        \wRegInTop_7_112[19] , \ScanLink223[4] , \wRegInBot_5_6[15] , 
        \wRegOut_6_12[18] , \wRegOut_6_31[30] , \wRegOut_7_126[2] , 
        \wRegOut_6_31[29] , \wRegOut_7_69[18] , \wRegInTop_6_32[5] , 
        \wRegOut_6_44[19] , \wRegInTop_7_13[3] , \wRegOut_7_8[15] , 
        \ScanLink140[2] , \wRegOut_7_125[1] , \ScanLink220[7] , 
        \wRegInTop_4_14[22] , \wRegInTop_7_82[16] , \wRegInBot_0_0[8] , 
        \wRegInBot_0_0[1] , \wRegOut_2_0[9] , \wRegOut_3_3[17] , 
        \wRegInTop_4_7[10] , \wRegInBot_4_14[25] , \wRegInBot_6_5[8] , 
        \wRegOut_7_2[2] , \ScanLink192[4] , \wRegInTop_7_97[22] , 
        \ScanLink39[24] , \ScanLink211[11] , \ScanLink182[13] , 
        \ScanLink197[27] , \ScanLink232[20] , \ScanLink247[10] , 
        \ScanLink227[14] , \wRegInBot_3_4[0] , \wRegInTop_3_5[6] , 
        \wRegOut_5_22[20] , \ScanLink59[20] , \wRegOut_6_41[4] , 
        \wRegOut_7_60[2] , \ScanLink252[24] , \ScanLink204[25] , 
        \wRegInTop_7_119[15] , \wRegInTop_3_6[5] , \wRegInBot_5_4[4] , 
        \wRegOut_5_14[25] , \wRegInTop_6_0[14] , \wRegOut_7_99[15] , 
        \wRegInTop_5_5[2] , \wRegOut_5_10[6] , \wRegOut_6_19[14] , 
        \wRegInBot_3_7[3] , \wRegOut_7_17[24] , \wRegOut_7_62[14] , 
        \wRegInTop_5_8[13] , \wRegOut_7_41[25] , \wRegOut_5_13[5] , 
        \wRegOut_7_21[21] , \wRegOut_7_34[15] , \wRegOut_7_54[11] , 
        \wRegOut_7_3[19] , \wRegOut_7_77[20] , \wRegInTop_5_6[1] , 
        \wRegInBot_5_7[7] , \wRegInBot_5_11[19] , \ScanLink94[24] , 
        \ScanLink119[16] , \ScanLink122[8] , \wRegInTop_7_71[9] , 
        \wRegOut_5_14[16] , \ScanLink81[10] , \wRegOut_6_42[7] , 
        \ScanLink179[12] , \wRegOut_7_63[1] , \wRegInBot_6_0[5] , 
        \wRegInTop_6_1[3] , \ScanLink66[2] , \ScanLink158[0] , 
        \ScanLink197[9] , \wRegInTop_7_117[3] , \ScanLink0[2] , 
        \wRegInTop_2_0[30] , \wRegOut_3_3[24] , \wRegOut_5_22[13] , 
        \wRegInTop_6_0[27] , \wRegInTop_7_119[26] , \wRegEnBot_6_29[0] , 
        \wRegOut_7_19[9] , \wRegOut_7_99[26] , \ScanLink238[5] , 
        \ScanLink252[17] , \ScanLink182[20] , \ScanLink227[27] , 
        \wRegInBot_4_2[30] , \wRegInBot_4_2[29] , \ScanLink204[16] , 
        \wRegInTop_4_7[23] , \ScanLink39[17] , \ScanLink59[13] , 
        \wRegInTop_6_37[8] , \wRegInTop_7_72[31] , \wRegInTop_5_27[31] , 
        \wRegInTop_5_27[28] , \wRegOut_6_25[0] , \wRegInTop_7_24[30] , 
        \wRegInTop_7_24[29] , \wRegInTop_7_51[19] , \wRegInTop_7_72[28] , 
        \ScanLink211[22] , \ScanLink247[23] , \ScanLink197[14] , 
        \ScanLink232[13] , \ScanLink81[23] , \ScanLink179[21] , 
        \ScanLink189[5] , \ScanLink94[17] , \ScanLink226[9] , 
        \wRegInTop_2_0[29] , \wRegOut_6_26[3] , \wRegInTop_7_89[29] , 
        \ScanLink119[25] , \wRegInBot_2_1[31] , \wRegOut_2_3[20] , 
        \wRegOut_2_3[13] , \ScanLink8[31] , \wRegInBot_6_3[6] , 
        \wRegInTop_7_89[30] , \wRegOut_7_21[12] , \ScanLink8[28] , 
        \wRegInTop_6_2[0] , \wRegInTop_6_29[4] , \wRegOut_7_54[22] , 
        \ScanLink23[4] , \wRegOut_4_10[2] , \wRegInTop_4_10[30] , 
        \wRegInTop_4_10[29] , \wRegInBot_4_14[5] , \wRegInTop_5_8[20] , 
        \wRegOut_6_19[27] , \wRegOut_7_17[17] , \wRegOut_7_77[13] , 
        \wRegOut_7_62[27] , \ScanLink65[1] , \wRegOut_7_34[26] , 
        \wRegInTop_7_114[0] , \wRegEnTop_7_46[0] , \wRegOut_7_41[16] , 
        \ScanLink116[11] , \wRegInTop_7_0[10] , \ScanLink135[20] , 
        \ScanLink163[21] , \ScanLink120[14] , \ScanLink140[10] , 
        \wRegInTop_7_93[30] , \wRegOut_5_31[4] , \ScanLink155[24] , 
        \wRegInTop_5_7[14] , \wRegOut_6_16[13] , \ScanLink103[25] , 
        \ScanLink176[15] , \wRegInTop_7_93[29] , \wRegOut_7_93[6] , 
        \wRegOut_6_35[22] , \wRegOut_6_63[23] , \wRegOut_7_18[23] , 
        \wRegOut_6_20[16] , \ScanLink100[9] , \wRegOut_6_40[12] , 
        \wRegInTop_7_53[8] , \wRegInBot_6_22[4] , \wRegOut_6_55[26] , 
        \wRegOut_7_78[27] , \wRegInBot_3_5[14] , \wRegEnBot_4_9[0] , 
        \wRegOut_6_60[6] , \wRegOut_7_41[0] , \wRegOut_5_8[3] , 
        \wRegInBot_6_21[7] , \wRegOut_7_96[12] , \wRegInTop_7_116[12] , 
        \wRegOut_7_42[3] , \wRegOut_7_83[26] , \ScanLink15[12] , 
        \wRegOut_4_4[19] , \wRegInTop_4_8[17] , \wRegOut_4_15[12] , 
        \ScanLink36[23] , \ScanLink43[13] , \wRegOut_6_63[5] , 
        \wRegInTop_7_103[26] , \wRegInTop_7_120[17] , \ScanLink60[22] , 
        \ScanLink198[20] , \ScanLink20[7] , \ScanLink56[27] , \ScanLink75[16] , 
        \wRegInTop_6_45[30] , \ScanLink248[17] , \ScanLink228[13] , 
        \wRegInTop_6_13[28] , \wRegOut_7_90[5] , \wRegInTop_6_45[29] , 
        \wRegInTop_7_68[28] , \wRegInTop_6_30[19] , \ScanLink23[17] , 
        \wRegOut_4_13[1] , \wRegInTop_6_13[31] , \wRegEnTop_6_22[0] , 
        \wRegOut_6_20[25] , \wRegOut_6_55[15] , \wRegInTop_7_68[31] , 
        \wRegOut_7_78[14] , \wRegInBot_3_5[27] , \ScanLink15[21] , 
        \ScanLink23[24] , \wRegInTop_5_7[27] , \wRegOut_6_16[20] , 
        \wRegInBot_6_46[0] , \wRegOut_6_63[10] , \wRegOut_7_18[10] , 
        \wRegOut_6_40[21] , \wRegOut_7_25[4] , \ScanLink204[8] , 
        \ScanLink47[0] , \wRegInBot_5_17[2] , \wRegInBot_5_28[31] , 
        \ScanLink95[6] , \wRegOut_6_35[11] , \ScanLink103[16] , 
        \ScanLink120[27] , \ScanLink155[17] , \ScanLink176[26] , 
        \ScanLink179[2] , \ScanLink116[22] , \wRegInTop_7_0[23] , 
        \ScanLink163[12] , \ScanLink219[7] , \ScanLink140[23] , 
        \wRegInBot_5_28[28] , \ScanLink88[9] , \ScanLink75[25] , 
        \wRegInBot_6_50[30] , \ScanLink135[13] , \ScanLink228[20] , 
        \wRegInBot_6_50[29] , \wRegInTop_4_8[24] , \ScanLink36[10] , 
        \ScanLink56[14] , \wRegInTop_7_29[0] , \wRegInBot_6_25[19] , 
        \wRegOut_7_115[19] , \ScanLink43[20] , \wRegInBot_5_14[1] , 
        \ScanLink44[3] , \wRegOut_4_15[21] , \ScanLink60[11] , 
        \ScanLink248[24] , \ScanLink198[13] , \wRegOut_7_83[15] , 
        \wRegInTop_7_103[15] , \wRegInBot_5_9[21] , \wRegInTop_5_25[2] , 
        \wRegInTop_6_15[9] , \wRegInTop_7_120[24] , \ScanLink96[5] , 
        \wRegInBot_6_45[3] , \wRegInTop_7_116[21] , \wRegOut_7_7[21] , 
        \wRegOut_7_25[19] , \wRegOut_7_26[7] , \wRegOut_7_96[21] , 
        \wRegInTop_7_48[9] , \wRegOut_7_50[29] , \wRegOut_7_73[18] , 
        \wRegInTop_7_87[0] , \wRegOut_7_50[30] , \wRegInBot_6_39[5] , 
        \wRegOut_7_95[8] , \wRegInBot_2_1[28] , \wRegOut_5_0[25] , 
        \wRegInTop_5_23[23] , \ScanLink85[31] , \ScanLink106[7] , 
        \wRegInTop_7_55[6] , \wRegInTop_4_3[31] , \wRegInTop_4_3[28] , 
        \wRegInBot_4_6[22] , \ScanLink28[31] , \ScanLink38[5] , 
        \wRegInTop_5_15[26] , \wRegInBot_5_15[21] , \ScanLink85[28] , 
        \wRegInTop_7_98[16] , \wRegOut_7_88[7] , \wRegInBot_5_23[24] , 
        \wRegInTop_6_18[17] , \wRegInTop_7_63[17] , \wRegInTop_7_16[27] , 
        \ScanLink28[28] , \wRegOut_6_8[22] , \ScanLink105[4] , 
        \wRegInTop_7_40[26] , \wRegInTop_7_35[16] , \wRegInTop_7_56[5] , 
        \wRegOut_5_29[6] , \wRegInTop_7_20[22] , \wRegInTop_7_55[12] , 
        \ScanLink243[31] , \ScanLink215[29] , \wRegInBot_6_27[9] , 
        \wRegInTop_4_8[1] , \wRegInTop_7_76[23] , \ScanLink243[28] , 
        \wRegInBot_4_9[7] , \wRegInBot_6_18[10] , \ScanLink26[9] , 
        \wRegInTop_5_26[1] , \ScanLink215[30] , \wRegOut_7_88[19] , 
        \ScanLink236[18] , \wRegInTop_7_108[19] , \wRegInBot_6_1[26] , 
        \wRegInTop_7_84[3] , \wRegOut_5_0[16] , \wRegInTop_5_15[15] , 
        \wRegOut_5_26[18] , \wRegOut_7_59[2] , \wRegInBot_5_15[12] , 
        \wRegInTop_5_23[10] , \wRegInBot_5_23[17] , \wRegInTop_6_10[4] , 
        \ScanLink162[3] , \ScanLink93[8] , \ScanLink108[30] , 
        \wRegInTop_7_31[2] , \wRegOut_7_107[0] , \ScanLink108[29] , 
        \ScanLink202[6] , \wRegInTop_7_98[25] , \wRegOut_7_7[12] , 
        \wRegOut_1_0[18] , \ScanLink3[1] , \wRegInBot_5_9[12] , 
        \wRegEnBot_6_10[0] , \wRegInBot_6_1[15] , \wRegInBot_4_6[11] , 
        \wRegInTop_6_13[7] , \wRegInTop_7_20[11] , \wRegInBot_6_18[23] , 
        \wRegInTop_7_32[1] , \ScanLink161[0] , \wRegInTop_7_55[21] , 
        \ScanLink186[18] , \wRegInTop_7_76[10] , \wRegOut_6_8[11] , 
        \wRegInTop_6_18[24] , \wRegInTop_7_16[14] , \wRegOut_7_20[9] , 
        \ScanLink201[5] , \wRegInTop_7_35[25] , \wRegInTop_7_63[24] , 
        \wRegOut_7_104[3] , \wRegInTop_7_40[15] , \wRegOut_2_0[0] , 
        \wRegInTop_2_0[20] , \wRegInBot_4_2[20] , \wRegEnTop_6_4[0] , 
        \wRegOut_6_38[6] , \wRegOut_7_7[6] , \wRegOut_7_19[0] , 
        \ScanLink158[9] , \wRegInBot_6_5[24] , \wRegOut_6_25[9] , 
        \wRegInTop_7_24[20] , \wRegInTop_7_51[10] , \ScanLink197[0] , 
        \wRegOut_7_120[5] , \wRegInTop_7_72[21] , \wRegInTop_7_12[25] , 
        \ScanLink182[29] , \wRegInTop_7_67[15] , \ScanLink225[3] , 
        \wRegInTop_5_11[24] , \wRegInTop_6_37[1] , \wRegInTop_7_16[7] , 
        \ScanLink145[6] , \wRegInTop_7_44[24] , \ScanLink182[30] , 
        \wRegInTop_7_31[14] , \wRegInBot_5_28[5] , \wRegInTop_7_89[20] , 
        \ScanLink226[0] , \wRegInTop_7_109[6] , \wRegOut_7_123[6] , 
        \wRegOut_2_3[3] , \ScanLink8[21] , \wRegOut_5_4[27] , 
        \wRegInTop_5_27[21] , \wRegInBot_5_27[26] , \ScanLink78[7] , 
        \ScanLink179[31] , \wRegInTop_6_34[2] , \wRegInTop_7_15[4] , 
        \ScanLink146[5] , \ScanLink179[28] , \wRegInTop_5_8[30] , 
        \wRegInBot_5_11[23] , \wRegInTop_5_8[29] , \ScanLink65[8] , 
        \wRegOut_7_4[5] , \wRegEnTop_7_89[0] , \wRegInTop_7_114[9] , 
        \wRegInTop_6_2[9] , \wRegOut_7_3[23] , \ScanLink194[3] , 
        \wRegInBot_4_2[13] , \wRegInTop_4_7[19] , \ScanLink59[30] , 
        \wRegInTop_7_12[16] , \ScanLink59[29] , \wRegInTop_7_67[26] , 
        \ScanLink241[7] , \wRegInTop_6_53[5] , \wRegInTop_7_24[13] , 
        \wRegInTop_7_31[27] , \wRegInTop_7_44[17] , \ScanLink211[18] , 
        \ScanLink232[30] , \wRegInTop_7_51[23] , \wRegInTop_7_72[3] , 
        \ScanLink121[2] , \wRegInTop_7_72[12] , \ScanLink232[29] , 
        \ScanLink247[19] , \wRegInBot_3_4[9] , \wRegOut_5_22[30] , 
        \wRegOut_5_22[29] , \wRegInBot_6_5[17] , \wRegOut_4_3[7] , 
        \wRegOut_7_3[10] , \wRegOut_7_21[28] , \wRegOut_7_54[18] , 
        \wRegOut_7_77[30] , \wRegInTop_2_0[13] , \ScanLink8[12] , 
        \wRegOut_7_21[31] , \wRegOut_7_77[29] , \wRegEnBot_3_2[0] , 
        \wRegInTop_5_6[8] , \wRegOut_4_0[4] , \wRegOut_5_4[14] , 
        \wRegInBot_5_11[10] , \wRegInTop_5_27[12] , \ScanLink81[19] , 
        \ScanLink242[4] , \wRegOut_7_63[8] , \wRegInTop_5_11[17] , 
        \wRegInTop_7_89[13] , \wRegInBot_3_1[16] , \ScanLink11[10] , 
        \wRegInBot_4_11[1] , \wRegInBot_5_27[15] , \ScanLink71[14] , 
        \wRegInTop_6_50[6] , \ScanLink122[1] , \ScanLink189[16] , 
        \wRegInTop_7_71[0] , \wRegInBot_6_21[31] , \wRegInTop_7_111[4] , 
        \ScanLink27[15] , \ScanLink52[25] , \wRegInBot_5_30[7] , 
        \wRegInBot_6_21[28] , \ScanLink60[5] , \wRegOut_7_1[8] , 
        \ScanLink32[21] , \ScanLink47[11] , \wRegInBot_6_54[18] , 
        \wRegInBot_6_6[2] , \wRegInTop_6_7[4] , \wRegOut_7_111[28] , 
        \ScanLink64[20] , \ScanLink239[25] , \wRegInBot_6_61[5] , 
        \wRegOut_7_111[31] , \wRegOut_7_87[24] , \wRegOut_4_11[10] , 
        \wRegOut_6_23[7] , \wRegInTop_7_107[24] , \wRegInTop_7_124[15] , 
        \wRegOut_0_0[15] , \wRegInBot_4_12[2] , \wRegInTop_5_3[16] , 
        \wRegOut_5_29[25] , \wRegOut_6_12[11] , \wRegOut_6_20[4] , 
        \wRegOut_6_24[14] , \wRegInTop_7_10[9] , \ScanLink143[8] , 
        \wRegOut_7_92[10] , \wRegInTop_7_112[10] , \wRegOut_6_51[24] , 
        \wRegOut_7_125[8] , \wRegInBot_6_62[6] , \wRegOut_6_31[20] , 
        \wRegOut_7_69[11] , \wRegOut_6_44[10] , \ScanLink124[16] , 
        \wRegInTop_7_112[7] , \ScanLink63[6] , \ScanLink151[26] , 
        \ScanLink107[27] , \ScanLink112[13] , \ScanLink172[17] , 
        \wRegInTop_7_4[12] , \ScanLink167[23] , \wRegEnTop_7_118[0] , 
        \wRegInTop_6_4[7] , \wRegInBot_6_5[1] , \ScanLink131[22] , 
        \ScanLink144[12] , \wRegOut_0_0[26] , \wRegInBot_3_1[25] , 
        \wRegOut_4_0[28] , \wRegOut_4_11[23] , \wRegOut_5_29[16] , 
        \wRegOut_6_47[3] , \wRegOut_7_92[23] , \wRegInTop_7_112[23] , 
        \wRegOut_7_66[5] , \ScanLink247[9] , \wRegOut_7_87[17] , 
        \wRegInTop_7_107[17] , \wRegInBot_3_2[7] , \wRegInTop_3_3[1] , 
        \ScanLink11[23] , \wRegOut_4_0[31] , \wRegInTop_5_19[6] , 
        \ScanLink32[12] , \wRegInTop_7_124[26] , \ScanLink47[22] , 
        \wRegOut_5_16[1] , \wRegEnTop_7_27[0] , \wRegInBot_5_2[3] , 
        \wRegInTop_5_3[5] , \ScanLink64[13] , \wRegInTop_6_17[19] , 
        \ScanLink239[16] , \wRegInTop_6_34[31] , \wRegOut_4_5[9] , 
        \ScanLink189[25] , \wRegInTop_6_62[29] , \ScanLink27[26] , 
        \ScanLink71[27] , \wRegInTop_6_34[28] , \wRegInTop_7_19[29] , 
        \wRegInTop_4_14[18] , \wRegInTop_5_0[6] , \wRegInBot_5_1[0] , 
        \ScanLink52[16] , \wRegInTop_6_41[18] , \wRegInTop_6_48[4] , 
        \wRegInTop_6_62[30] , \wRegInTop_7_69[2] , \wRegInTop_7_4[21] , 
        \wRegInTop_7_19[30] , \ScanLink112[20] , \ScanLink167[10] , 
        \wRegOut_7_78[9] , \wRegOut_5_15[2] , \ScanLink144[21] , 
        \ScanLink124[25] , \ScanLink131[11] , \ScanLink139[0] , 
        \ScanLink151[15] , \wRegEnBot_1_0[0] , \ScanLink2[27] , 
        \wRegInTop_2_1[19] , \wRegInTop_3_0[2] , \ScanLink172[24] , 
        \wRegInBot_3_1[4] , \ScanLink107[14] , \wRegInTop_7_97[18] , 
        \wRegInTop_5_3[25] , \wRegOut_6_12[22] , \wRegOut_6_44[23] , 
        \wRegOut_6_44[0] , \wRegOut_7_65[6] , \wRegOut_7_69[22] , 
        \wRegInTop_5_26[18] , \wRegInBot_6_10[6] , \wRegOut_6_24[27] , 
        \wRegOut_6_31[13] , \wRegOut_6_51[17] , \wRegInTop_6_56[8] , 
        \wRegEnBot_6_48[0] , \ScanLink80[13] , \wRegOut_6_52[4] , 
        \ScanLink178[11] , \wRegOut_7_73[2] , \ScanLink9[18] , 
        \ScanLink95[27] , \ScanLink118[15] , \wRegInTop_7_88[19] , 
        \wRegOut_7_76[23] , \wRegOut_3_2[27] , \wRegOut_3_2[14] , 
        \ScanLink11[6] , \wRegOut_7_20[22] , \wRegOut_7_55[12] , 
        \ScanLink12[5] , \wRegInTop_5_9[10] , \wRegOut_7_40[26] , 
        \wRegOut_6_18[17] , \wRegOut_7_35[16] , \wRegOut_7_16[27] , 
        \wRegOut_7_63[17] , \wRegInBot_4_3[19] , \wRegInBot_5_9[8] , 
        \wRegOut_5_15[26] , \wRegOut_5_23[23] , \wRegInTop_6_1[17] , 
        \wRegInTop_7_118[16] , \wRegOut_7_98[16] , \ScanLink58[23] , 
        \ScanLink205[26] , \ScanLink183[10] , \ScanLink226[17] , 
        \wRegInBot_6_13[5] , \wRegInTop_4_6[20] , \wRegInTop_4_6[13] , 
        \ScanLink38[27] , \wRegOut_6_51[7] , \wRegInTop_7_25[19] , 
        \wRegInTop_7_50[30] , \ScanLink196[24] , \wRegOut_7_70[1] , 
        \ScanLink253[27] , \ScanLink233[23] , \wRegInTop_7_73[18] , 
        \ScanLink246[13] , \ScanLink210[12] , \ScanLink38[14] , 
        \wRegInTop_5_9[23] , \ScanLink131[8] , \wRegInTop_7_50[29] , 
        \wRegInTop_7_62[9] , \wRegInBot_5_10[30] , \wRegInBot_5_10[29] , 
        \wRegInBot_5_25[0] , \wRegOut_7_35[25] , \wRegInTop_7_104[3] , 
        \ScanLink75[2] , \ScanLink80[20] , \wRegOut_6_18[24] , 
        \wRegOut_7_16[14] , \wRegOut_7_40[15] , \ScanLink95[14] , 
        \wRegInTop_6_39[7] , \wRegOut_7_2[30] , \wRegOut_7_63[24] , 
        \wRegOut_7_2[29] , \wRegOut_7_20[11] , \wRegOut_7_76[10] , 
        \wRegInTop_7_18[1] , \ScanLink184[9] , \wRegOut_7_55[21] , 
        \wRegOut_7_9[0] , \wRegOut_6_36[0] , \wRegOut_7_17[6] , 
        \ScanLink118[26] , \ScanLink178[22] , \wRegInTop_6_24[8] , 
        \wRegOut_6_35[3] , \wRegOut_7_14[5] , \ScanLink196[17] , 
        \ScanLink199[6] , \ScanLink246[20] , \ScanLink233[10] , 
        \ScanLink235[9] , \ScanLink58[10] , \ScanLink205[15] , 
        \ScanLink210[21] , \ScanLink183[23] , \ScanLink226[24] , 
        \ScanLink253[14] , \wRegOut_5_15[15] , \wRegOut_5_23[10] , 
        \wRegInBot_5_26[3] , \wRegInTop_6_1[24] , \wRegInTop_7_118[25] , 
        \wRegOut_7_98[25] , \ScanLink228[6] , \wRegInTop_7_107[0] , 
        \ScanLink76[1] , \wRegEnTop_7_55[0] , \ScanLink148[3] , 
        \wRegOut_5_18[7] , \wRegOut_6_13[31] , \wRegOut_6_45[29] , 
        \wRegOut_6_30[19] , \wRegOut_6_13[28] , \wRegInBot_6_16[8] , 
        \wRegOut_6_45[30] , \wRegOut_7_68[31] , \wRegOut_7_68[28] , 
        \ScanLink254[0] , \ScanLink2[14] , \ScanLink10[30] , \ScanLink10[29] , 
        \ScanLink17[8] , \wRegInBot_5_7[25] , \wRegInTop_6_46[2] , 
        \ScanLink134[5] , \wRegOut_7_9[25] , \wRegInTop_7_67[4] , 
        \wRegInTop_4_15[12] , \wRegInTop_7_83[26] , \wRegInBot_4_15[15] , 
        \wRegOut_6_49[5] , \wRegOut_7_68[3] , \wRegInTop_5_17[0] , 
        \wRegInTop_7_96[12] , \ScanLink46[31] , \wRegInBot_6_63[24] , 
        \wRegInTop_7_78[27] , \ScanLink65[19] , \wRegInBot_6_16[14] , 
        \wRegInTop_3_5[25] , \wRegInBot_4_8[26] , \ScanLink33[18] , 
        \wRegInBot_6_40[15] , \wRegOut_7_110[11] , \wRegInTop_5_14[3] , 
        \ScanLink46[28] , \wRegInTop_6_20[16] , \wRegOut_6_6[26] , 
        \wRegInTop_6_35[22] , \wRegInBot_6_35[25] , \wRegInTop_6_55[26] , 
        \wRegOut_7_105[25] , \wRegInTop_6_16[13] , \wRegInBot_6_20[11] , 
        \wRegInTop_6_40[12] , \wRegInBot_6_55[21] , \wRegInTop_7_79[8] , 
        \wRegOut_7_126[14] , \wRegInTop_6_63[23] , \wRegInTop_7_18[23] , 
        \wRegOut_6_57[9] , \wRegOut_7_93[29] , \wRegInTop_7_113[29] , 
        \wRegOut_7_93[30] , \wRegInTop_7_113[30] , \wRegOut_4_1[22] , 
        \wRegOut_4_10[30] , \wRegInTop_6_45[1] , \ScanLink137[6] , 
        \wRegInTop_7_64[7] , \wRegOut_4_10[29] , \wRegInTop_4_15[21] , 
        \wRegInBot_4_15[26] , \wRegInTop_7_96[21] , \ScanLink113[19] , 
        \ScanLink130[28] , \ScanLink145[18] , \ScanLink182[7] , 
        \ScanLink166[30] , \wRegInTop_7_83[15] , \wRegInBot_5_7[16] , 
        \ScanLink130[31] , \wRegInTop_7_5[18] , \ScanLink166[29] , 
        \wRegOut_7_11[8] , \ScanLink230[4] , \wRegInTop_3_1[27] , 
        \wRegInTop_3_5[16] , \wRegOut_4_1[11] , \wRegInBot_6_8[4] , 
        \wRegOut_7_9[16] , \wRegInTop_6_9[2] , \wRegInTop_6_22[6] , 
        \ScanLink150[1] , \ScanLink233[7] , \wRegOut_4_5[20] , 
        \wRegInBot_4_8[15] , \wRegOut_6_6[15] , \wRegInBot_6_20[22] , 
        \wRegInTop_6_21[5] , \ScanLink153[2] , \wRegInTop_6_40[21] , 
        \wRegInTop_6_35[11] , \wRegInBot_6_55[12] , \wRegInTop_6_63[10] , 
        \wRegOut_7_105[16] , \wRegInTop_6_16[20] , \wRegInTop_7_18[10] , 
        \wRegInBot_6_16[27] , \wRegOut_7_126[27] , \wRegInTop_6_20[25] , 
        \wRegInBot_6_35[16] , \wRegInBot_6_63[17] , \wRegInTop_7_78[14] , 
        \wRegInBot_6_40[26] , \wRegInTop_6_55[15] , \wRegOut_7_110[22] , 
        \wRegInTop_7_24[5] , \ScanLink181[4] , \ScanLink177[4] , 
        \wRegInBot_5_19[4] , \wRegInBot_6_55[9] , \ScanLink217[1] , 
        \wRegOut_7_112[7] , \wRegInBot_4_11[17] , \ScanLink49[6] , 
        \ScanLink54[9] , \wRegOut_6_1[7] , \wRegOut_6_2[24] , 
        \wRegInTop_6_31[20] , \wRegInBot_6_51[23] , \wRegOut_7_101[27] , 
        \wRegInTop_6_12[11] , \wRegInBot_6_24[13] , \wRegInTop_6_44[10] , 
        \wRegInBot_6_12[16] , \wRegInBot_6_48[6] , \wRegInTop_7_69[11] , 
        \wRegOut_7_122[16] , \wRegInBot_6_44[17] , \ScanLink199[19] , 
        \wRegOut_7_114[13] , \wRegInTop_7_125[8] , \wRegInTop_6_24[14] , 
        \wRegInBot_6_31[27] , \wRegInTop_6_51[24] , \wRegInTop_5_29[25] , 
        \wRegInTop_7_4[8] , \wRegInTop_7_92[10] , \wRegOut_6_2[4] , 
        \ScanLink169[8] , \wRegInTop_7_1[30] , \wRegInBot_2_2[8] , 
        \ScanLink6[25] , \wRegInTop_4_11[10] , \wRegEnTop_5_19[0] , 
        \wRegInBot_5_29[22] , \ScanLink134[19] , \ScanLink141[29] , 
        \ScanLink98[3] , \ScanLink117[31] , \wRegInTop_7_1[29] , 
        \ScanLink141[30] , \ScanLink162[18] , \wRegInTop_7_87[24] , 
        \ScanLink117[28] , \wRegOut_7_28[1] , \wRegInBot_5_3[27] , 
        \wRegOut_5_5[6] , \ScanLink61[28] , \wRegOut_6_14[8] , 
        \wRegInTop_7_27[6] , \ScanLink174[7] , \ScanLink214[2] , 
        \wRegOut_7_111[4] , \wRegInBot_6_12[25] , \ScanLink14[18] , 
        \ScanLink37[30] , \wRegEnBot_6_62[0] , \wRegInTop_4_11[3] , 
        \ScanLink37[29] , \ScanLink42[19] , \ScanLink61[31] , 
        \wRegInTop_5_30[5] , \wRegInBot_6_31[14] , \wRegInTop_6_51[17] , 
        \wRegInTop_7_92[7] , \wRegInTop_6_24[27] , \wRegInBot_6_44[24] , 
        \wRegOut_7_114[20] , \wRegInTop_6_44[23] , \wRegOut_0_0[18] , 
        \wRegInBot_0_0[5] , \wRegInBot_1_0[7] , \wRegOut_2_2[19] , 
        \wRegInTop_3_1[14] , \wRegOut_3_5[2] , \wRegEnTop_4_6[0] , 
        \wRegOut_6_2[17] , \wRegInBot_6_24[20] , \wRegInTop_6_31[13] , 
        \wRegInBot_6_51[10] , \wRegOut_7_101[14] , \ScanLink229[19] , 
        \wRegInTop_6_12[22] , \wRegInTop_7_69[22] , \wRegOut_7_97[18] , 
        \wRegInTop_7_117[18] , \wRegOut_7_122[25] , \wRegOut_4_5[13] , 
        \wRegOut_4_14[18] , \ScanLink113[0] , \wRegInTop_6_61[7] , 
        \wRegInTop_7_40[1] , \wRegInBot_5_3[14] , \wRegOut_6_17[19] , 
        \wRegOut_6_34[31] , \wRegOut_6_34[28] , \wRegOut_7_52[9] , 
        \wRegOut_6_41[18] , \wRegOut_6_62[30] , \wRegInTop_7_43[2] , 
        \wRegInTop_6_62[4] , \ScanLink110[3] , \wRegOut_7_19[30] , 
        \wRegOut_6_62[29] , \wRegOut_7_19[29] , \ScanLink6[16] , 
        \wRegOut_3_6[16] , \wRegOut_3_6[1] , \wRegInTop_4_0[9] , 
        \wRegInTop_4_11[23] , \wRegOut_5_6[5] , \wRegInBot_5_29[11] , 
        \wRegInTop_7_91[4] , \wRegInTop_7_87[17] , \wRegInTop_4_12[0] , 
        \wRegInTop_7_92[23] , \wRegInTop_4_2[11] , \wRegInBot_4_11[24] , 
        \ScanLink49[15] , \wRegInTop_5_29[16] , \wRegInBot_6_19[29] , 
        \ScanLink192[26] , \ScanLink237[21] , \ScanLink242[11] , 
        \wRegInBot_6_19[30] , \ScanLink214[10] , \ScanLink29[11] , 
        \ScanLink80[1] , \ScanLink201[24] , \wRegOut_7_114[9] , 
        \wRegInBot_6_53[7] , \ScanLink187[12] , \ScanLink222[15] , 
        \wRegOut_5_27[21] , \wRegInTop_6_5[15] , \wRegOut_6_11[5] , 
        \wRegOut_7_30[3] , \wRegInTop_7_1[5] , \wRegOut_1_1[21] , 
        \wRegOut_1_1[12] , \wRegOut_6_7[9] , \wRegInTop_1_1[1] , 
        \wRegOut_7_109[6] , \wRegInTop_7_123[6] , \wRegInBot_2_0[11] , 
        \wRegInBot_5_8[18] , \wRegOut_5_11[24] , \ScanLink52[7] , 
        \wRegEnTop_6_50[0] , \wRegInTop_7_2[6] , \wRegOut_7_89[20] , 
        \wRegInTop_7_109[20] , \wRegOut_7_12[25] , \wRegOut_7_31[14] , 
        \wRegOut_7_44[24] , \wRegOut_7_67[15] , \wRegOut_7_72[21] , 
        \wRegInBot_5_14[18] , \ScanLink51[4] , \wRegOut_7_24[20] , 
        \wRegOut_7_51[10] , \wRegInTop_7_120[5] , \ScanLink91[25] , 
        \wRegOut_7_6[18] , \wRegInTop_7_21[8] , \ScanLink172[9] , 
        \wRegInBot_6_50[4] , \ScanLink169[27] , \wRegOut_6_12[6] , 
        \ScanLink109[23] , \ScanLink83[2] , \ScanLink84[11] , 
        \wRegOut_7_33[0] , \ScanLink108[1] , \wRegInTop_7_94[9] , 
        \wRegInBot_2_0[22] , \wRegOut_3_6[25] , \wRegInBot_4_4[2] , 
        \wRegInTop_4_5[4] , \wRegOut_5_3[8] , \wRegOut_7_89[13] , 
        \wRegOut_5_11[17] , \wRegInTop_7_109[13] , \wRegInTop_6_5[26] , 
        \wRegOut_7_86[1] , \wRegInBot_4_7[31] , \ScanLink29[22] , 
        \ScanLink36[3] , \wRegOut_7_49[8] , \wRegOut_5_24[3] , 
        \wRegOut_5_27[12] , \wRegOut_6_9[28] , \ScanLink201[17] , 
        \wRegInTop_7_89[6] , \wRegOut_6_9[31] , \ScanLink187[21] , 
        \ScanLink222[26] , \wRegInTop_4_2[22] , \wRegInBot_4_7[28] , 
        \wRegInBot_6_37[3] , \wRegInTop_7_77[29] , \wRegInTop_7_21[31] , 
        \ScanLink242[22] , \wRegOut_7_54[7] , \ScanLink192[15] , 
        \wRegInTop_7_54[18] , \wRegInTop_7_77[30] , \ScanLink237[12] , 
        \ScanLink49[26] , \wRegInTop_5_22[30] , \ScanLink84[22] , 
        \wRegInTop_7_21[28] , \ScanLink214[23] , \wRegOut_3_3[20] , 
        \wRegOut_3_3[13] , \wRegInBot_3_4[4] , \wRegInTop_3_5[2] , 
        \wRegInTop_3_6[1] , \wRegInTop_4_6[7] , \ScanLink35[0] , 
        \wRegInTop_5_22[29] , \wRegInTop_5_28[7] , \ScanLink109[10] , 
        \wRegOut_5_27[0] , \ScanLink91[16] , \wRegInBot_6_34[0] , 
        \ScanLink169[14] , \wRegOut_7_24[13] , \wRegOut_7_57[4] , 
        \wRegOut_7_72[12] , \wRegOut_7_31[27] , \wRegOut_7_51[23] , 
        \wRegInTop_7_58[3] , \wRegOut_7_44[17] , \wRegInBot_4_7[1] , 
        \wRegOut_7_12[16] , \wRegOut_7_67[26] , \wRegOut_7_85[2] , 
        \wRegOut_5_4[19] , \wRegOut_6_42[3] , \ScanLink179[16] , 
        \wRegInTop_5_6[5] , \wRegInBot_5_7[3] , \wRegInBot_5_27[18] , 
        \ScanLink81[14] , \wRegOut_7_63[5] , \ScanLink242[9] , 
        \ScanLink94[20] , \ScanLink119[12] , \wRegOut_7_77[24] , 
        \wRegInTop_5_8[17] , \wRegOut_5_13[1] , \wRegOut_7_21[25] , 
        \wRegOut_7_54[15] , \wRegEnTop_7_22[0] , \wRegOut_7_41[21] , 
        \wRegOut_7_34[11] , \wRegInBot_3_7[7] , \wRegOut_4_0[9] , 
        \wRegOut_6_19[10] , \wRegOut_7_17[20] , \wRegOut_7_62[10] , 
        \wRegInBot_5_4[0] , \wRegOut_5_10[2] , \wRegOut_5_14[21] , 
        \wRegInTop_5_5[6] , \wRegInTop_6_0[10] , \wRegOut_5_22[24] , 
        \wRegOut_7_99[11] , \wRegInTop_7_119[11] , \ScanLink59[24] , 
        \ScanLink204[21] , \ScanLink182[17] , \ScanLink227[10] , 
        \wRegInTop_4_7[27] , \wRegInTop_4_7[14] , \ScanLink39[20] , 
        \wRegOut_6_41[0] , \wRegOut_7_60[6] , \ScanLink252[20] , 
        \ScanLink197[23] , \ScanLink232[24] , \ScanLink211[15] , 
        \ScanLink247[14] , \wRegInBot_4_14[1] , \wRegInTop_5_8[24] , 
        \wRegInTop_6_53[8] , \wRegInTop_7_114[4] , \ScanLink39[13] , 
        \wRegInTop_5_11[30] , \ScanLink65[5] , \wRegOut_7_34[22] , 
        \wRegInTop_6_2[4] , \wRegInBot_6_3[2] , \wRegOut_6_19[23] , 
        \wRegOut_7_4[8] , \wRegOut_7_17[13] , \wRegOut_7_41[12] , 
        \wRegOut_7_62[23] , \wRegOut_7_77[17] , \wRegInTop_6_29[0] , 
        \wRegOut_7_21[16] , \wRegOut_7_54[26] , \wRegInTop_5_11[29] , 
        \wRegInBot_5_28[8] , \ScanLink94[13] , \ScanLink81[27] , 
        \wRegOut_6_26[7] , \ScanLink119[21] , \ScanLink179[25] , 
        \wRegOut_6_25[4] , \wRegInTop_7_15[9] , \ScanLink189[1] , 
        \ScanLink146[8] , \ScanLink197[10] , \ScanLink232[17] , 
        \ScanLink247[27] , \wRegOut_7_120[8] , \ScanLink59[17] , 
        \wRegInTop_7_12[31] , \wRegInTop_7_44[29] , \ScanLink211[26] , 
        \ScanLink204[12] , \wRegInTop_7_31[19] , \wRegInTop_7_44[30] , 
        \ScanLink252[13] , \ScanLink182[24] , \wRegInTop_7_67[18] , 
        \ScanLink227[23] , \wRegInTop_6_0[23] , \wRegInTop_7_12[28] , 
        \wRegOut_7_99[22] , \wRegInTop_7_119[22] , \ScanLink238[1] , 
        \wRegInTop_7_117[7] , \ScanLink3[20] , \wRegInTop_5_3[31] , 
        \wRegInTop_5_3[28] , \wRegOut_5_14[12] , \wRegOut_5_22[17] , 
        \ScanLink66[6] , \wRegInBot_6_0[1] , \wRegInTop_6_1[7] , 
        \wRegInBot_6_5[29] , \ScanLink158[4] , \wRegInBot_6_5[30] , 
        \ScanLink244[7] , \wRegInBot_3_1[31] , \wRegInBot_3_1[9] , 
        \wRegInTop_4_14[15] , \wRegInBot_5_6[22] , \wRegInTop_6_56[5] , 
        \ScanLink124[2] , \wRegOut_7_8[22] , \wRegOut_6_59[2] , 
        \wRegInTop_7_77[3] , \wRegInTop_7_82[21] , \wRegInBot_4_14[12] , 
        \ScanLink172[29] , \wRegOut_7_78[4] , \ScanLink107[19] , 
        \ScanLink124[31] , \wRegInTop_3_4[22] , \wRegEnBot_3_7[0] , 
        \wRegOut_4_5[4] , \wRegOut_4_6[7] , \wRegInTop_5_3[8] , 
        \wRegInBot_6_17[13] , \wRegInBot_6_18[3] , \ScanLink124[28] , 
        \ScanLink151[18] , \wRegInTop_7_97[15] , \ScanLink172[30] , 
        \wRegInBot_6_62[23] , \wRegInTop_7_79[20] , \wRegOut_6_7[21] , 
        \wRegInTop_6_21[11] , \wRegInBot_6_41[12] , \wRegOut_7_111[16] , 
        \wRegInTop_6_34[25] , \wRegInBot_6_34[22] , \wRegInTop_6_54[21] , 
        \wRegInBot_6_54[26] , \wRegOut_7_104[22] , \wRegInTop_6_17[14] , 
        \wRegInBot_6_21[16] , \wRegInTop_6_41[15] , \wRegInTop_6_48[9] , 
        \ScanLink189[31] , \wRegOut_7_127[13] , \wRegInBot_4_9[21] , 
        \wRegInTop_6_62[24] , \wRegInTop_7_19[24] , \ScanLink189[28] , 
        \wRegOut_7_66[8] , \ScanLink247[4] , \ScanLink19[3] , 
        \wRegInBot_3_1[28] , \wRegOut_4_0[25] , \wRegInTop_6_55[6] , 
        \ScanLink127[1] , \wRegInTop_7_74[0] , \wRegInBot_4_14[21] , 
        \wRegInTop_7_97[26] , \wRegInTop_4_14[26] , \wRegEnTop_6_1[0] , 
        \wRegOut_7_2[6] , \ScanLink192[0] , \wRegInTop_7_82[12] , 
        \wRegOut_1_0[26] , \wRegOut_1_0[15] , \wRegOut_1_1[1] , 
        \ScanLink3[13] , \wRegInBot_5_6[11] , \wRegOut_6_20[9] , 
        \wRegOut_6_51[30] , \ScanLink220[3] , \wRegInTop_3_4[11] , 
        \wRegOut_4_0[16] , \wRegOut_6_24[19] , \wRegOut_7_125[5] , 
        \wRegInTop_6_32[1] , \wRegOut_6_51[29] , \wRegOut_7_8[11] , 
        \wRegInTop_7_13[7] , \wRegInBot_6_61[8] , \ScanLink140[6] , 
        \wRegOut_7_87[30] , \wRegOut_7_126[6] , \wRegInTop_7_107[30] , 
        \wRegInTop_7_124[18] , \wRegOut_7_87[29] , \wRegInTop_7_107[29] , 
        \wRegOut_5_29[31] , \ScanLink223[0] , \wRegInBot_4_9[12] , 
        \ScanLink27[18] , \ScanLink52[28] , \wRegOut_5_29[28] , 
        \wRegInTop_6_31[2] , \wRegInTop_7_10[4] , \ScanLink143[5] , 
        \wRegInTop_6_41[26] , \wRegInTop_7_111[9] , \ScanLink60[8] , 
        \wRegInBot_6_21[25] , \wRegOut_6_7[12] , \wRegInTop_6_34[16] , 
        \wRegOut_7_1[5] , \wRegInBot_6_54[15] , \wRegOut_7_104[11] , 
        \ScanLink52[31] , \wRegInTop_6_62[17] , \ScanLink71[19] , 
        \wRegInTop_6_17[27] , \wRegInTop_7_19[17] , \wRegInBot_6_17[20] , 
        \wRegOut_7_127[20] , \wRegInBot_6_34[11] , \wRegInBot_6_62[10] , 
        \ScanLink239[28] , \wRegInTop_7_79[13] , \wRegInTop_6_54[12] , 
        \ScanLink239[31] , \ScanLink5[2] , \wRegInTop_3_0[20] , 
        \wRegOut_4_4[27] , \wRegInTop_6_7[9] , \wRegInBot_6_41[21] , 
        \wRegOut_7_111[25] , \wRegInTop_6_15[4] , \wRegInTop_6_21[22] , 
        \ScanLink191[3] , \wRegInTop_7_120[29] , \wRegInTop_7_34[2] , 
        \ScanLink167[3] , \wRegOut_7_83[18] , \wRegInTop_7_120[30] , 
        \ScanLink96[8] , \ScanLink207[6] , \wRegInTop_7_103[18] , 
        \wRegOut_7_102[0] , \ScanLink23[30] , \ScanLink23[29] , 
        \ScanLink59[1] , \wRegInTop_6_30[27] , \ScanLink56[19] , 
        \wRegOut_6_3[23] , \wRegOut_7_100[20] , \ScanLink75[31] , 
        \wRegInBot_6_25[14] , \wRegInTop_6_45[17] , \wRegInBot_6_50[24] , 
        \wRegInTop_6_13[16] , \wRegInTop_4_8[30] , \ScanLink75[28] , 
        \wRegInTop_7_68[16] , \wRegOut_7_123[11] , \wRegInBot_6_58[1] , 
        \ScanLink6[1] , \wRegInTop_4_8[29] , \wRegInBot_6_13[11] , 
        \ScanLink248[29] , \wRegInBot_6_45[10] , \wRegInBot_4_10[10] , 
        \wRegEnBot_6_15[0] , \wRegInTop_6_25[13] , \wRegOut_7_115[14] , 
        \ScanLink248[30] , \wRegInBot_6_30[20] , \wRegInTop_6_50[23] , 
        \wRegInTop_5_28[22] , \wRegInTop_7_93[17] , \wRegInBot_5_28[25] , 
        \ScanLink88[4] , \ScanLink7[22] , \wRegInTop_4_10[17] , 
        \wRegInTop_7_86[23] , \wRegOut_6_19[0] , \wRegOut_7_38[6] , 
        \ScanLink7[11] , \wRegInTop_3_0[13] , \wRegInBot_5_2[20] , 
        \wRegOut_6_20[31] , \wRegOut_7_78[19] , \wRegInTop_5_20[2] , 
        \wRegInBot_6_13[22] , \wRegInTop_6_16[7] , \wRegOut_6_55[18] , 
        \wRegInTop_7_9[0] , \ScanLink164[0] , \wRegOut_6_20[28] , 
        \wRegOut_7_25[9] , \wRegInTop_7_37[1] , \ScanLink204[5] , 
        \wRegOut_7_101[3] , \wRegOut_6_3[10] , \wRegInTop_6_25[20] , 
        \wRegInBot_6_30[13] , \wRegInBot_6_45[23] , \wRegInTop_6_50[10] , 
        \wRegInTop_7_82[0] , \wRegOut_7_115[27] , \wRegInBot_6_25[27] , 
        \wRegInTop_6_45[24] , \wRegInTop_6_30[14] , \wRegInTop_6_13[25] , 
        \wRegInBot_6_50[17] , \wRegOut_7_100[13] , \wRegInTop_7_68[25] , 
        \wRegOut_7_90[8] , \wRegOut_7_123[22] , \wRegInBot_3_5[19] , 
        \ScanLink103[7] , \wRegOut_6_63[8] , \wRegInTop_7_50[6] , 
        \wRegOut_4_4[14] , \wRegInBot_5_2[13] , \wRegInTop_5_7[19] , 
        \wRegInTop_7_53[5] , \ScanLink100[4] , \wRegInBot_6_22[9] , 
        \wRegOut_3_7[11] , \wRegInTop_4_3[16] , \ScanLink23[9] , 
        \wRegInTop_4_10[24] , \wRegInBot_5_28[16] , \wRegInTop_7_81[3] , 
        \wRegInTop_7_86[10] , \wRegInBot_4_10[23] , \wRegInTop_5_23[1] , 
        \ScanLink103[28] , \ScanLink155[30] , \ScanLink176[18] , 
        \wRegInTop_7_93[24] , \wRegInTop_5_28[11] , \wRegOut_5_31[9] , 
        \ScanLink103[31] , \ScanLink120[19] , \ScanLink155[29] , 
        \ScanLink48[12] , \ScanLink193[21] , \ScanLink236[26] , 
        \ScanLink243[16] , \ScanLink215[17] , \ScanLink28[16] , 
        \wRegInTop_6_18[30] , \wRegInTop_7_35[28] , \ScanLink200[23] , 
        \ScanLink90[6] , \wRegInTop_7_63[30] , \wRegInBot_6_43[0] , 
        \wRegInTop_7_35[31] , \wRegInTop_7_40[18] , \ScanLink186[15] , 
        \ScanLink223[12] , \wRegInTop_7_16[19] , \wRegInBot_5_12[2] , 
        \wRegOut_5_26[26] , \wRegInTop_6_4[12] , \wRegInTop_6_18[29] , 
        \wRegOut_7_20[4] , \ScanLink201[8] , \wRegInTop_7_63[29] , 
        \wRegInBot_6_1[18] , \wRegInBot_2_1[16] , \ScanLink41[3] , 
        \wRegOut_5_10[23] , \ScanLink42[0] , \wRegOut_7_119[1] , 
        \wRegInBot_5_11[1] , \wRegOut_7_13[22] , \wRegOut_7_30[13] , 
        \wRegOut_7_45[23] , \wRegOut_7_88[27] , \wRegInTop_7_108[27] , 
        \wRegOut_7_66[12] , \wRegOut_7_73[26] , \wRegOut_7_25[27] , 
        \wRegOut_7_50[17] , \wRegInTop_5_15[18] , \wRegInTop_6_10[9] , 
        \ScanLink90[22] , \wRegInBot_6_40[3] , \ScanLink168[20] , 
        \ScanLink108[24] , \wRegInTop_7_98[28] , \wRegOut_6_9[2] , 
        \ScanLink85[16] , \wRegOut_7_23[7] , \ScanLink93[5] , 
        \wRegInTop_7_98[31] , \ScanLink118[6] , \wRegInTop_2_0[0] , 
        \wRegInBot_2_1[25] , \wRegOut_3_7[22] , \ScanLink26[4] , 
        \wRegOut_5_10[10] , \wRegOut_7_88[14] , \wRegInTop_7_108[14] , 
        \wRegInTop_6_4[21] , \wRegOut_7_96[6] , \ScanLink28[25] , 
        \wRegOut_4_15[2] , \wRegOut_5_26[15] , \ScanLink105[9] , 
        \wRegInTop_7_99[1] , \wRegInTop_7_56[8] , \ScanLink200[10] , 
        \ScanLink186[26] , \ScanLink223[21] , \wRegInTop_4_3[25] , 
        \wRegInBot_6_27[4] , \wRegOut_7_44[0] , \ScanLink236[15] , 
        \ScanLink243[25] , \ScanLink193[12] , \wRegOut_5_0[28] , 
        \ScanLink48[21] , \ScanLink85[25] , \ScanLink215[24] , 
        \wRegInBot_2_1[6] , \ScanLink25[7] , \wRegOut_5_0[31] , 
        \ScanLink108[17] , \ScanLink38[8] , \wRegInBot_5_23[29] , 
        \wRegInBot_5_23[30] , \wRegInBot_6_24[7] , \ScanLink90[11] , 
        \ScanLink168[13] , \wRegOut_7_47[3] , \wRegOut_7_25[14] , 
        \wRegOut_7_73[15] , \wRegOut_7_30[20] , \wRegInTop_7_48[4] , 
        \wRegOut_7_50[24] , \wRegEnTop_6_27[0] , \wRegInBot_6_39[8] , 
        \wRegOut_7_45[10] , \wRegOut_7_13[11] , \wRegOut_7_66[21] , 
        \wRegOut_7_95[5] , \wRegOut_5_6[8] , \ScanLink117[16] , 
        \wRegInTop_7_1[17] , \ScanLink162[26] , \wRegOut_2_2[14] , 
        \wRegInTop_4_0[4] , \wRegInBot_4_11[30] , \ScanLink33[3] , 
        \wRegOut_5_21[3] , \ScanLink121[13] , \ScanLink134[27] , 
        \ScanLink141[17] , \wRegInTop_7_91[9] , \ScanLink154[23] , 
        \ScanLink102[22] , \wRegInBot_4_1[2] , \ScanLink177[12] , 
        \wRegOut_7_83[1] , \wRegInBot_4_11[29] , \wRegInBot_5_3[19] , 
        \wRegInTop_5_6[13] , \wRegOut_6_17[14] , \wRegOut_6_34[25] , 
        \wRegOut_6_62[24] , \wRegOut_7_19[24] , \wRegOut_6_21[11] , 
        \wRegOut_6_41[15] , \wRegInTop_6_62[9] , \wRegInBot_6_32[3] , 
        \wRegOut_6_54[21] , \wRegOut_7_79[20] , \wRegInBot_2_2[5] , 
        \wRegInTop_3_1[19] , \wRegOut_7_51[7] , \wRegInBot_3_4[13] , 
        \wRegInBot_6_31[0] , \wRegOut_7_97[15] , \wRegInTop_7_117[15] , 
        \wRegOut_7_52[4] , \wRegOut_7_82[21] , \wRegInTop_4_9[10] , 
        \wRegOut_4_14[15] , \wRegInTop_7_102[21] , \ScanLink37[24] , 
        \ScanLink42[14] , \wRegInBot_6_12[31] , \wRegInTop_7_121[10] , 
        \wRegInBot_6_31[19] , \wRegInBot_6_44[29] , \ScanLink61[25] , 
        \wRegInBot_6_12[28] , \ScanLink199[27] , \wRegInTop_2_3[3] , 
        \ScanLink14[15] , \wRegInBot_6_44[30] , \wRegInBot_4_2[1] , 
        \wRegInTop_4_3[7] , \wRegInTop_5_30[8] , \ScanLink74[11] , 
        \ScanLink229[14] , \ScanLink249[10] , \wRegOut_7_80[2] , 
        \wRegOut_7_122[28] , \wRegInBot_1_0[3] , \ScanLink2[19] , 
        \wRegInTop_2_1[27] , \wRegOut_2_2[27] , \ScanLink6[31] , 
        \ScanLink22[10] , \ScanLink30[0] , \ScanLink57[20] , \wRegOut_5_22[0] , 
        \wRegOut_7_101[19] , \wRegOut_7_122[31] , \wRegOut_6_54[12] , 
        \ScanLink6[28] , \wRegOut_6_21[22] , \wRegOut_7_79[13] , 
        \wRegOut_3_0[2] , \ScanLink8[7] , \wRegInBot_3_4[20] , 
        \ScanLink14[26] , \ScanLink22[23] , \wRegInTop_5_6[20] , 
        \wRegOut_6_14[5] , \wRegOut_6_17[27] , \wRegInBot_6_56[7] , 
        \wRegOut_6_62[17] , \wRegOut_7_19[17] , \wRegOut_6_41[26] , 
        \wRegOut_7_35[3] , \wRegOut_7_111[9] , \ScanLink57[7] , 
        \wRegInTop_5_29[31] , \wRegInTop_5_29[28] , \ScanLink85[1] , 
        \wRegOut_6_34[16] , \wRegInTop_7_4[5] , \ScanLink154[10] , 
        \ScanLink121[20] , \ScanLink169[5] , \ScanLink177[21] , 
        \wRegOut_6_2[9] , \ScanLink102[11] , \ScanLink117[25] , 
        \wRegInTop_7_1[24] , \ScanLink162[15] , \wRegInTop_7_87[29] , 
        \ScanLink209[0] , \wRegEnTop_6_55[0] , \ScanLink141[24] , 
        \wRegInTop_7_126[6] , \wRegOut_6_2[30] , \ScanLink134[14] , 
        \wRegInTop_7_87[30] , \wRegOut_6_2[29] , \ScanLink74[22] , 
        \ScanLink229[27] , \wRegInTop_7_7[6] , \wRegInTop_4_9[23] , 
        \ScanLink37[17] , \ScanLink57[13] , \wRegInTop_6_18[1] , 
        \wRegInTop_7_39[7] , \ScanLink42[27] , \wRegInTop_6_24[19] , 
        \wRegInTop_7_125[5] , \ScanLink54[4] , \wRegInTop_6_51[29] , 
        \wRegOut_4_14[26] , \ScanLink61[16] , \ScanLink249[23] , 
        \wRegInTop_6_51[30] , \ScanLink199[14] , \wRegOut_7_82[12] , 
        \wRegInTop_7_102[12] , \wRegInBot_5_19[9] , \wRegInTop_7_24[8] , 
        \wRegInTop_7_121[23] , \ScanLink177[9] , \ScanLink86[2] , 
        \wRegInBot_6_55[4] , \wRegInTop_7_117[26] , \wRegEnTop_4_3[0] , 
        \wRegInTop_4_14[3] , \wRegOut_5_0[6] , \wRegOut_6_17[6] , 
        \wRegOut_7_97[26] , \wRegOut_7_6[26] , \wRegOut_7_36[0] , 
        \wRegInTop_7_97[7] , \wRegInBot_5_8[26] , \wRegInBot_6_29[2] , 
        \wRegOut_3_3[1] , \wRegOut_3_6[31] , \wRegOut_3_6[28] , 
        \ScanLink28[2] , \wRegOut_5_1[22] , \wRegInTop_5_22[24] , 
        \ScanLink116[0] , \wRegInTop_7_45[1] , \wRegInTop_5_14[21] , 
        \wRegInBot_5_14[26] , \wRegInTop_7_99[11] , \ScanLink169[19] , 
        \wRegOut_7_57[9] , \wRegOut_7_98[0] , \wRegInBot_5_22[23] , 
        \wRegInTop_6_19[10] , \wRegInTop_7_17[20] , \wRegInTop_7_62[10] , 
        \wRegInBot_4_7[25] , \wRegOut_6_9[25] , \ScanLink115[3] , 
        \wRegInTop_7_41[21] , \wRegInTop_7_34[11] , \wRegInTop_7_46[2] , 
        \wRegInTop_4_5[9] , \wRegOut_5_3[5] , \wRegInBot_6_19[17] , 
        \wRegInTop_7_21[25] , \wRegInTop_7_54[15] , \wRegInTop_7_77[24] , 
        \ScanLink192[18] , \wRegInBot_6_0[21] , \wRegInTop_7_94[4] , 
        \wRegInBot_4_3[27] , \wRegInBot_4_7[16] , \wRegOut_5_1[11] , 
        \wRegInTop_5_14[12] , \ScanLink91[28] , \wRegOut_7_49[5] , 
        \wRegInBot_5_14[15] , \wRegInTop_5_22[17] , \wRegInBot_5_22[10] , 
        \ScanLink91[31] , \ScanLink172[4] , \wRegInTop_7_21[5] , 
        \wRegOut_7_117[7] , \wRegInBot_6_50[9] , \ScanLink212[1] , 
        \wRegInTop_7_99[22] , \wRegInBot_5_8[15] , \ScanLink51[9] , 
        \wRegOut_6_4[7] , \wRegOut_7_12[31] , \wRegOut_7_12[28] , 
        \wRegOut_7_44[30] , \wRegOut_7_67[18] , \wRegOut_7_31[19] , 
        \wRegOut_7_44[29] , \wRegInTop_7_120[8] , \wRegOut_7_6[15] , 
        \wRegOut_5_11[30] , \wRegOut_5_11[29] , \wRegInTop_6_5[18] , 
        \wRegInTop_7_1[8] , \ScanLink49[18] , \wRegInBot_6_0[12] , 
        \wRegOut_6_7[4] , \wRegInBot_6_19[24] , \wRegInTop_7_21[16] , 
        \wRegInTop_7_22[6] , \wRegInTop_7_54[26] , \ScanLink171[7] , 
        \ScanLink201[30] , \wRegInTop_7_77[17] , \ScanLink222[18] , 
        \ScanLink38[19] , \wRegOut_5_15[18] , \wRegInTop_6_1[30] , 
        \wRegOut_6_9[16] , \wRegOut_6_11[8] , \wRegInTop_7_17[13] , 
        \ScanLink211[2] , \wRegInTop_6_19[23] , \wRegInTop_7_34[22] , 
        \wRegInTop_7_62[23] , \ScanLink201[29] , \wRegOut_7_114[4] , 
        \wRegInTop_7_41[12] , \wRegInTop_7_118[31] , \wRegInTop_6_1[29] , 
        \wRegOut_7_98[31] , \wRegInTop_7_118[28] , \wRegOut_6_28[1] , 
        \wRegOut_7_98[28] , \wRegInBot_6_4[23] , \ScanLink187[7] , 
        \wRegInTop_7_13[22] , \wRegOut_7_14[8] , \wRegInTop_7_25[27] , 
        \wRegInTop_7_50[17] , \wRegInTop_7_73[26] , \wRegInTop_7_66[12] , 
        \ScanLink235[4] , \ScanLink253[19] , \ScanLink226[29] , 
        \wRegInTop_5_10[23] , \wRegInTop_6_27[6] , \ScanLink155[1] , 
        \wRegInTop_7_45[23] , \ScanLink226[30] , \wRegInTop_7_30[13] , 
        \ScanLink205[18] , \ScanLink95[19] , \wRegInTop_7_88[27] , 
        \ScanLink236[7] , \wRegInTop_7_119[1] , \wRegInTop_2_1[14] , 
        \ScanLink9[26] , \wRegOut_5_5[20] , \wRegInTop_5_26[26] , 
        \wRegInBot_5_26[21] , \ScanLink68[0] , \wRegInTop_6_24[5] , 
        \ScanLink156[2] , \wRegInBot_5_10[24] , \wRegOut_6_18[30] , 
        \wRegOut_6_18[29] , \wRegOut_7_16[19] , \wRegOut_7_35[31] , 
        \wRegOut_7_35[28] , \wRegOut_7_63[29] , \wRegOut_7_2[24] , 
        \wRegOut_7_40[18] , \wRegOut_7_63[30] , \ScanLink184[4] , 
        \ScanLink9[15] , \wRegOut_3_2[19] , \wRegInBot_4_3[14] , 
        \ScanLink12[8] , \wRegInTop_5_8[3] , \wRegInBot_5_9[5] , 
        \wRegInTop_7_13[11] , \wRegInBot_6_13[8] , \ScanLink251[0] , 
        \wRegInBot_6_4[10] , \wRegInTop_6_43[2] , \wRegInTop_7_25[14] , 
        \wRegInTop_7_30[20] , \wRegInTop_7_66[21] , \wRegInTop_7_45[10] , 
        \ScanLink196[30] , \ScanLink131[5] , \wRegInTop_7_50[24] , 
        \wRegInTop_7_62[4] , \ScanLink196[29] , \wRegInTop_7_73[15] , 
        \wRegInTop_5_12[0] , \wRegOut_7_2[17] , \wRegOut_5_5[13] , 
        \wRegInBot_5_10[17] , \wRegInTop_5_11[3] , \wRegInTop_5_26[15] , 
        \ScanLink252[3] , \wRegInTop_5_10[10] , \wRegOut_6_52[9] , 
        \ScanLink118[18] , \wRegInTop_7_88[14] , \wRegInBot_3_0[11] , 
        \ScanLink10[17] , \wRegInBot_4_8[18] , \wRegInBot_5_26[12] , 
        \wRegInTop_6_40[1] , \ScanLink132[6] , \ScanLink188[11] , 
        \wRegInTop_7_61[7] , \ScanLink26[12] , \wRegInBot_5_20[0] , 
        \ScanLink70[13] , \wRegInTop_7_101[3] , \ScanLink53[22] , 
        \ScanLink70[2] , \ScanLink33[26] , \ScanLink46[16] , \wRegOut_6_6[18] , 
        \wRegInTop_6_55[18] , \ScanLink65[27] , \wRegInTop_6_20[28] , 
        \ScanLink181[9] , \ScanLink238[22] , \wRegInTop_6_20[31] , 
        \wRegInTop_7_78[19] , \wRegOut_7_12[6] , \wRegOut_7_86[23] , 
        \wRegOut_4_10[17] , \wRegOut_5_28[22] , \wRegOut_6_33[0] , 
        \wRegInTop_7_106[23] , \wRegInTop_7_125[12] , \wRegInTop_6_21[8] , 
        \wRegOut_6_25[13] , \wRegOut_7_93[17] , \wRegInTop_7_113[17] , 
        \wRegOut_6_30[3] , \wRegOut_6_50[23] , \wRegOut_7_11[5] , 
        \ScanLink230[9] , \wRegOut_1_1[16] , \wRegInBot_2_0[15] , 
        \wRegInBot_3_0[22] , \wRegInTop_3_5[31] , \wRegInTop_3_5[28] , 
        \wRegInTop_5_2[11] , \wRegInBot_6_8[9] , \wRegOut_6_13[16] , 
        \wRegOut_6_30[27] , \wRegOut_7_68[16] , \wRegInBot_5_23[3] , 
        \wRegOut_6_45[17] , \ScanLink125[11] , \wRegInTop_7_102[0] , 
        \ScanLink73[1] , \ScanLink150[21] , \ScanLink106[20] , 
        \wRegEnTop_7_50[0] , \ScanLink113[14] , \ScanLink173[10] , 
        \wRegInTop_7_83[18] , \ScanLink130[25] , \wRegInTop_7_5[15] , 
        \ScanLink166[24] , \ScanLink145[15] , \wRegOut_5_28[11] , 
        \wRegInBot_6_15[6] , \wRegInTop_7_113[24] , \wRegOut_6_57[4] , 
        \wRegOut_7_93[24] , \wRegOut_4_10[24] , \wRegOut_7_76[2] , 
        \wRegOut_7_86[10] , \wRegInTop_7_106[10] , \ScanLink10[24] , 
        \ScanLink14[6] , \wRegOut_4_8[1] , \ScanLink33[15] , 
        \wRegInBot_6_63[30] , \wRegInTop_7_125[21] , \ScanLink46[25] , 
        \wRegInBot_6_35[28] , \wRegInBot_6_40[18] , \wRegInBot_6_63[29] , 
        \ScanLink17[5] , \ScanLink26[21] , \ScanLink65[14] , 
        \wRegInBot_6_35[31] , \ScanLink70[20] , \wRegInBot_6_16[19] , 
        \ScanLink188[22] , \wRegOut_7_105[31] , \ScanLink238[11] , 
        \wRegOut_7_126[19] , \wRegOut_7_105[28] , \ScanLink53[11] , 
        \wRegInTop_6_58[3] , \wRegInTop_7_79[5] , \wRegOut_6_49[8] , 
        \ScanLink113[27] , \wRegInTop_7_5[26] , \ScanLink166[17] , 
        \ScanLink249[2] , \ScanLink145[26] , \wRegInBot_4_15[18] , 
        \ScanLink125[22] , \ScanLink130[16] , \ScanLink150[12] , 
        \ScanLink129[7] , \ScanLink173[23] , \wRegInTop_5_2[22] , 
        \wRegOut_6_13[25] , \wRegInBot_6_16[5] , \ScanLink106[13] , 
        \wRegOut_6_45[24] , \wRegOut_6_54[7] , \wRegOut_7_68[25] , 
        \wRegOut_7_75[1] , \wRegInBot_5_7[31] , \wRegOut_6_30[14] , 
        \wRegOut_6_50[10] , \ScanLink134[8] , \wRegOut_7_9[28] , 
        \wRegInBot_5_7[28] , \wRegOut_6_25[20] , \wRegInTop_7_67[9] , 
        \wRegOut_7_9[31] , \ScanLink83[6] , \ScanLink109[27] , 
        \wRegInBot_6_50[0] , \wRegOut_5_1[18] , \wRegOut_5_11[20] , 
        \ScanLink51[0] , \wRegInBot_5_22[19] , \wRegOut_6_12[2] , 
        \ScanLink84[15] , \wRegOut_7_33[4] , \ScanLink212[8] , 
        \ScanLink91[21] , \ScanLink169[23] , \wRegOut_7_24[24] , 
        \wRegOut_7_51[14] , \wRegInTop_7_120[1] , \wRegInTop_7_2[2] , 
        \wRegOut_7_12[21] , \wRegOut_7_67[11] , \wRegOut_7_72[25] , 
        \wRegOut_7_31[10] , \wRegOut_7_44[20] , \wRegOut_7_89[24] , 
        \wRegInTop_7_109[24] , \wRegOut_1_1[25] , \wRegInTop_1_1[5] , 
        \wRegOut_7_109[2] , \wRegInTop_7_123[2] , \wRegInBot_2_0[26] , 
        \wRegOut_3_6[12] , \ScanLink52[3] , \wRegOut_5_27[25] , 
        \wRegInTop_7_1[1] , \wRegInTop_6_5[11] , \wRegInBot_6_53[3] , 
        \ScanLink187[16] , \ScanLink222[11] , \wRegInTop_4_2[15] , 
        \ScanLink29[15] , \wRegOut_6_11[1] , \ScanLink80[5] , 
        \wRegOut_7_30[7] , \ScanLink201[20] , \ScanLink49[11] , 
        \ScanLink214[14] , \wRegInTop_4_6[3] , \ScanLink192[22] , 
        \ScanLink237[25] , \ScanLink242[15] , \wRegInBot_4_7[5] , 
        \wRegOut_7_12[12] , \wRegOut_7_67[22] , \wRegOut_7_85[6] , 
        \ScanLink35[4] , \wRegOut_5_27[4] , \wRegOut_7_31[23] , 
        \wRegInTop_5_14[31] , \wRegInTop_5_14[28] , \wRegOut_7_24[17] , 
        \wRegOut_7_44[13] , \wRegOut_7_51[27] , \wRegInTop_7_58[7] , 
        \wRegOut_7_72[16] , \ScanLink91[12] , \wRegInBot_6_34[4] , 
        \ScanLink169[10] , \wRegOut_7_57[0] , \wRegOut_7_98[9] , 
        \ScanLink84[26] , \ScanLink116[9] , \wRegInTop_7_45[8] , 
        \wRegOut_3_3[8] , \wRegOut_3_6[21] , \wRegInTop_4_2[26] , 
        \wRegInTop_5_28[3] , \ScanLink109[14] , \wRegInTop_7_99[18] , 
        \ScanLink49[22] , \wRegInTop_6_19[19] , \wRegInBot_6_37[7] , 
        \ScanLink214[27] , \wRegOut_7_54[3] , \ScanLink192[11] , 
        \ScanLink242[26] , \ScanLink237[16] , \wRegInTop_7_17[29] , 
        \wRegInTop_7_41[31] , \ScanLink187[25] , \wRegInTop_7_62[19] , 
        \ScanLink222[22] , \wRegInBot_4_4[6] , \wRegInTop_4_5[0] , 
        \ScanLink29[26] , \ScanLink36[7] , \wRegInTop_7_17[30] , 
        \wRegInTop_7_41[28] , \ScanLink201[13] , \wRegInTop_7_89[2] , 
        \wRegInTop_7_34[18] , \wRegOut_5_24[7] , \wRegOut_5_27[16] , 
        \wRegEnTop_6_34[0] , \wRegInTop_6_5[22] , \wRegOut_7_86[5] , 
        \wRegOut_5_11[13] , \wRegOut_7_89[17] , \wRegInTop_7_109[17] , 
        \wRegInBot_6_0[31] , \ScanLink108[5] , \wRegInTop_2_0[9] , 
        \ScanLink6[21] , \wRegInTop_5_6[30] , \wRegInBot_6_0[28] , 
        \wRegInTop_5_6[29] , \ScanLink214[6] , \ScanLink85[8] , 
        \wRegEnTop_7_69[0] , \wRegOut_7_111[0] , \wRegInTop_7_27[2] , 
        \ScanLink174[3] , \wRegInTop_3_1[23] , \wRegInTop_4_11[14] , 
        \wRegInBot_5_3[23] , \wRegInTop_7_87[20] , \wRegInBot_4_11[13] , 
        \wRegInTop_5_29[21] , \wRegInBot_5_29[26] , \wRegOut_6_2[0] , 
        \wRegOut_7_28[5] , \ScanLink209[9] , \ScanLink98[7] , 
        \ScanLink154[19] , \ScanLink177[31] , \ScanLink121[29] , 
        \ScanLink177[28] , \wRegInBot_5_19[0] , \wRegOut_6_1[3] , 
        \wRegInTop_6_24[10] , \ScanLink102[18] , \wRegInBot_6_44[13] , 
        \ScanLink121[30] , \wRegInTop_7_92[14] , \wRegOut_7_114[17] , 
        \wRegOut_6_2[20] , \wRegInTop_6_12[15] , \wRegInBot_6_12[12] , 
        \wRegInBot_6_31[23] , \wRegInBot_6_48[2] , \wRegInTop_6_51[20] , 
        \wRegInTop_6_31[24] , \wRegInTop_7_69[15] , \wRegOut_7_122[12] , 
        \wRegOut_7_101[23] , \wRegInTop_6_18[8] , \wRegInTop_6_44[14] , 
        \wRegInBot_6_51[27] , \wRegInBot_6_24[17] , \wRegOut_7_112[3] , 
        \wRegInBot_3_4[30] , \wRegInBot_3_4[29] , \wRegOut_4_5[24] , 
        \ScanLink49[2] , \wRegOut_7_36[9] , \ScanLink217[5] , \wRegOut_3_6[5] , 
        \wRegInBot_4_11[20] , \wRegInTop_5_29[12] , \wRegInTop_7_24[1] , 
        \ScanLink177[0] , \wRegInTop_7_92[27] , \wRegInTop_4_11[27] , 
        \wRegOut_5_6[1] , \wRegOut_7_83[8] , \wRegInTop_7_87[13] , 
        \wRegInTop_4_12[4] , \ScanLink6[12] , \wRegInBot_5_3[10] , 
        \wRegInBot_5_29[15] , \wRegOut_6_21[18] , \wRegOut_7_79[30] , 
        \wRegInTop_7_91[0] , \wRegOut_6_54[28] , \wRegOut_7_79[29] , 
        \wRegOut_6_54[31] , \wRegInTop_3_1[10] , \wRegOut_4_5[17] , 
        \wRegInBot_6_31[9] , \ScanLink110[7] , \wRegInTop_6_62[0] , 
        \wRegInTop_7_43[6] , \wRegOut_7_82[28] , \wRegInTop_7_102[28] , 
        \wRegOut_7_82[31] , \wRegInTop_7_102[31] , \wRegInTop_7_121[19] , 
        \wRegOut_3_5[6] , \wRegEnBot_4_12[0] , \ScanLink57[30] , 
        \ScanLink113[4] , \wRegInTop_6_61[3] , \wRegInTop_7_40[5] , 
        \ScanLink74[18] , \wRegInBot_4_2[8] , \ScanLink57[29] , 
        \wRegInTop_6_12[26] , \wRegInTop_6_44[27] , \wRegInTop_7_69[26] , 
        \wRegOut_7_122[21] , \wRegOut_0_0[11] , \ScanLink2[23] , 
        \wRegInTop_3_5[21] , \wRegOut_4_1[26] , \ScanLink22[19] , 
        \ScanLink30[9] , \wRegInBot_6_24[24] , \wRegInTop_6_31[17] , 
        \wRegOut_5_22[9] , \wRegOut_6_2[13] , \wRegInBot_6_51[14] , 
        \wRegInTop_4_9[19] , \wRegInBot_6_31[10] , \wRegOut_7_101[10] , 
        \wRegInTop_6_51[13] , \wRegInTop_4_11[7] , \wRegOut_5_5[2] , 
        \wRegInBot_6_12[21] , \wRegInTop_6_24[23] , \wRegInBot_6_44[20] , 
        \wRegInTop_7_92[3] , \wRegOut_7_114[24] , \ScanLink249[19] , 
        \wRegInTop_5_30[1] , \wRegOut_7_86[19] , \wRegOut_4_8[8] , 
        \wRegInTop_7_106[19] , \wRegInTop_7_125[31] , \wRegEnBot_5_17[0] , 
        \wRegInTop_6_45[5] , \wRegInTop_7_125[28] , \ScanLink137[2] , 
        \wRegInTop_7_64[3] , \wRegInBot_4_8[22] , \ScanLink26[31] , 
        \wRegOut_5_28[18] , \wRegInTop_6_16[17] , \wRegInTop_5_14[7] , 
        \wRegOut_7_126[10] , \ScanLink70[29] , \wRegInTop_6_63[27] , 
        \ScanLink26[28] , \wRegInTop_6_35[26] , \wRegInTop_7_18[27] , 
        \wRegOut_7_105[21] , \wRegInTop_4_15[16] , \wRegInBot_4_15[11] , 
        \ScanLink53[18] , \wRegOut_6_6[22] , \wRegInBot_6_55[25] , 
        \ScanLink70[30] , \wRegInTop_6_40[16] , \wRegInBot_6_20[15] , 
        \wRegInBot_6_16[10] , \wRegInTop_6_20[12] , \wRegInBot_6_40[11] , 
        \wRegOut_7_110[15] , \wRegInBot_6_35[21] , \wRegInTop_6_55[22] , 
        \wRegInBot_6_63[20] , \wRegInTop_7_78[23] , \ScanLink238[18] , 
        \wRegInTop_5_17[4] , \wRegOut_6_49[1] , \wRegInTop_7_83[22] , 
        \wRegInTop_7_96[16] , \wRegOut_6_25[29] , \wRegOut_6_50[19] , 
        \wRegOut_7_9[21] , \wRegOut_7_68[7] , \ScanLink134[1] , 
        \wRegInTop_6_46[6] , \wRegInTop_7_67[0] , \ScanLink2[10] , 
        \wRegInBot_3_0[18] , \wRegInTop_3_5[12] , \wRegInBot_4_8[11] , 
        \wRegInBot_5_7[21] , \wRegOut_6_25[30] , \wRegOut_5_18[3] , 
        \wRegOut_7_75[8] , \ScanLink254[4] , \wRegInBot_6_16[23] , 
        \wRegInTop_6_20[21] , \wRegInBot_6_35[12] , \wRegInBot_6_40[22] , 
        \wRegInTop_6_55[11] , \wRegOut_7_110[26] , \ScanLink181[0] , 
        \wRegInTop_6_63[14] , \wRegInBot_6_63[13] , \ScanLink188[18] , 
        \wRegInTop_7_78[10] , \wRegInTop_7_18[14] , \wRegInBot_5_20[9] , 
        \wRegInTop_6_16[24] , \wRegInTop_6_40[25] , \wRegOut_7_126[23] , 
        \wRegOut_6_6[11] , \wRegInBot_6_20[26] , \wRegInTop_6_35[15] , 
        \wRegInBot_6_55[16] , \wRegOut_7_105[12] , \wRegInTop_6_21[1] , 
        \ScanLink153[6] , \wRegOut_6_33[9] , \wRegOut_4_1[15] , 
        \wRegInTop_5_2[18] , \wRegInBot_6_8[0] , \ScanLink233[3] , 
        \wRegInBot_5_7[12] , \wRegInTop_6_9[6] , \wRegInTop_6_22[2] , 
        \wRegOut_7_9[12] , \ScanLink150[5] , \ScanLink230[0] , 
        \wRegOut_3_2[23] , \wRegOut_3_2[10] , \wRegInTop_4_6[17] , 
        \wRegInTop_4_15[25] , \wRegInTop_7_83[11] , \wRegInBot_4_15[22] , 
        \ScanLink73[8] , \ScanLink106[30] , \ScanLink125[18] , 
        \ScanLink182[3] , \ScanLink150[28] , \wRegInTop_7_102[9] , 
        \ScanLink106[29] , \ScanLink150[31] , \ScanLink173[19] , 
        \wRegInTop_7_96[25] , \ScanLink38[23] , \ScanLink210[16] , 
        \wRegInBot_6_13[1] , \ScanLink183[14] , \ScanLink196[20] , 
        \ScanLink226[13] , \ScanLink233[27] , \ScanLink246[17] , 
        \wRegInTop_7_30[30] , \ScanLink11[2] , \ScanLink12[1] , 
        \wRegInTop_5_12[9] , \wRegOut_5_23[27] , \ScanLink58[27] , 
        \wRegOut_6_51[3] , \wRegInTop_7_13[18] , \wRegInTop_7_66[28] , 
        \wRegOut_7_70[5] , \ScanLink253[23] , \ScanLink251[9] , 
        \ScanLink205[22] , \wRegInTop_7_30[29] , \wRegInTop_7_45[19] , 
        \wRegInTop_7_66[31] , \wRegOut_5_15[22] , \wRegInTop_6_1[13] , 
        \wRegOut_7_98[12] , \wRegInTop_7_118[12] , \wRegInBot_6_4[19] , 
        \wRegInTop_5_9[14] , \wRegOut_6_18[13] , \wRegEnTop_7_31[0] , 
        \wRegOut_7_16[23] , \wRegOut_7_63[13] , \wRegOut_7_40[22] , 
        \wRegOut_7_20[26] , \wRegOut_7_35[12] , \wRegOut_7_55[16] , 
        \wRegInTop_5_10[19] , \ScanLink95[23] , \ScanLink118[11] , 
        \wRegOut_7_76[27] , \wCtrlOut_6[0] , \wRegOut_5_15[11] , 
        \wRegInBot_6_10[2] , \wRegInTop_6_40[8] , \ScanLink80[17] , 
        \wRegOut_6_52[0] , \ScanLink178[15] , \wRegOut_7_73[6] , 
        \wRegOut_5_23[14] , \wRegInBot_5_26[7] , \ScanLink148[7] , 
        \wRegInTop_7_107[4] , \ScanLink76[5] , \wRegInTop_6_1[20] , 
        \wRegOut_6_28[8] , \wRegOut_7_98[21] , \wRegInTop_7_118[21] , 
        \ScanLink183[27] , \ScanLink226[20] , \ScanLink228[2] , 
        \ScanLink253[10] , \wRegInTop_4_6[24] , \ScanLink38[10] , 
        \ScanLink58[14] , \ScanLink155[8] , \ScanLink205[11] , 
        \wRegInBot_4_14[28] , \wRegOut_5_5[30] , \wRegEnTop_5_25[0] , 
        \ScanLink210[25] , \ScanLink246[24] , \wRegOut_6_35[7] , 
        \wRegOut_7_14[1] , \ScanLink196[13] , \ScanLink233[14] , 
        \wRegOut_5_5[29] , \ScanLink80[24] , \ScanLink178[26] , 
        \ScanLink199[2] , \wRegInTop_5_9[27] , \wRegInBot_5_26[31] , 
        \ScanLink95[10] , \wRegOut_6_36[4] , \wRegOut_7_17[2] , 
        \wRegInBot_5_26[28] , \ScanLink118[22] , \wRegInTop_7_119[8] , 
        \ScanLink68[9] , \wRegOut_7_9[4] , \wRegOut_6_18[20] , 
        \wRegInTop_6_39[3] , \wRegInTop_7_18[5] , \wRegOut_7_20[15] , 
        \wRegOut_7_55[25] , \wRegOut_7_16[10] , \wRegOut_7_76[14] , 
        \wRegOut_7_63[20] , \wRegInBot_5_25[4] , \wRegOut_7_35[21] , 
        \wRegInTop_7_104[7] , \wRegInTop_6_4[3] , \wRegInBot_6_5[5] , 
        \ScanLink75[6] , \wRegOut_7_40[11] , \ScanLink131[26] , 
        \ScanLink192[9] , \ScanLink107[23] , \ScanLink112[17] , 
        \ScanLink144[16] , \wRegInTop_7_4[16] , \ScanLink167[27] , 
        \ScanLink172[13] , \ScanLink124[12] , \wRegInTop_7_112[3] , 
        \wRegInBot_4_12[6] , \wRegInBot_4_14[31] , \ScanLink63[2] , 
        \ScanLink151[22] , \wRegInTop_5_3[12] , \wRegOut_6_31[24] , 
        \wRegInTop_6_32[8] , \wRegOut_6_44[14] , \wRegInBot_5_6[18] , 
        \wRegOut_6_12[15] , \wRegOut_7_69[15] , \wRegOut_6_20[0] , 
        \wRegInBot_6_62[2] , \wRegOut_6_24[10] , \wRegOut_6_51[20] , 
        \wRegOut_7_8[18] , \wRegOut_7_92[14] , \wRegInTop_7_112[14] , 
        \wRegOut_0_0[22] , \wRegOut_1_1[8] , \wRegInBot_3_1[12] , 
        \wRegInTop_3_4[18] , \wRegOut_5_29[21] , \wRegInBot_6_61[1] , 
        \wRegInTop_7_124[11] , \wRegOut_7_87[20] , \ScanLink223[9] , 
        \ScanLink11[14] , \wRegOut_4_11[14] , \ScanLink64[24] , 
        \wRegInBot_6_17[29] , \wRegOut_6_23[3] , \wRegInTop_7_107[20] , 
        \ScanLink239[21] , \ScanLink47[15] , \wRegInBot_6_41[31] , 
        \wRegInBot_6_62[19] , \wRegInBot_6_17[30] , \wRegInBot_6_34[18] , 
        \ScanLink3[30] , \ScanLink3[29] , \wRegInBot_4_11[5] , 
        \ScanLink32[25] , \wRegInBot_6_6[6] , \wRegInTop_6_7[0] , 
        \wRegInBot_6_41[28] , \ScanLink27[11] , \ScanLink52[21] , 
        \wRegInBot_5_30[3] , \wRegInTop_7_111[0] , \ScanLink60[1] , 
        \wRegEnTop_7_43[0] , \wRegOut_7_104[18] , \ScanLink71[10] , 
        \ScanLink189[12] , \wRegOut_7_127[30] , \wRegOut_7_127[29] , 
        \wRegOut_6_51[13] , \wRegInTop_3_0[6] , \wRegInTop_5_3[21] , 
        \wRegOut_6_24[23] , \wRegOut_6_12[26] , \wRegOut_6_31[17] , 
        \wRegOut_6_44[27] , \wRegOut_6_44[4] , \ScanLink172[20] , 
        \wRegOut_7_65[2] , \wRegOut_7_69[26] , \wRegInBot_3_1[0] , 
        \ScanLink107[10] , \ScanLink124[21] , \ScanLink151[11] , 
        \ScanLink139[4] , \wRegInBot_3_1[21] , \wRegInBot_3_2[3] , 
        \wRegInTop_3_3[5] , \wRegInBot_4_9[31] , \ScanLink27[22] , 
        \wRegInTop_5_0[2] , \wRegInBot_5_1[4] , \wRegOut_5_15[6] , 
        \ScanLink144[25] , \wRegInTop_7_82[31] , \ScanLink131[15] , 
        \wRegInTop_7_4[25] , \ScanLink112[24] , \ScanLink167[14] , 
        \wRegInTop_7_82[28] , \wRegOut_6_7[28] , \ScanLink52[12] , 
        \wRegInTop_6_48[0] , \wRegInTop_7_69[6] , \wRegOut_6_7[31] , 
        \ScanLink189[21] , \ScanLink11[27] , \wRegInBot_4_9[28] , 
        \ScanLink71[23] , \wRegOut_4_11[27] , \ScanLink32[16] , 
        \wRegInBot_5_2[7] , \wRegInTop_7_79[29] , \wRegInTop_5_3[1] , 
        \ScanLink64[17] , \wRegInTop_6_54[31] , \ScanLink239[12] , 
        \ScanLink47[26] , \wRegOut_5_16[5] , \wRegInTop_6_21[18] , 
        \wRegInTop_7_79[30] , \wRegInTop_6_54[28] , \ScanLink127[8] , 
        \wRegInTop_7_74[9] , \wRegInTop_7_124[22] , \wRegOut_7_87[13] , 
        \wRegInTop_7_107[13] , \wRegInTop_5_19[2] , \wRegOut_6_47[7] , 
        \wRegOut_7_92[27] , \wRegInTop_7_112[27] , \wRegOut_7_66[1] , 
        \ScanLink0[6] , \ScanLink3[5] , \wRegOut_2_0[4] , \wRegInTop_2_0[24] , 
        \ScanLink8[25] , \wRegOut_5_29[12] , \wRegInBot_4_14[8] , 
        \wRegInTop_6_29[9] , \wRegOut_7_3[27] , \ScanLink194[7] , 
        \wRegOut_5_4[23] , \wRegOut_7_4[1] , \wRegInBot_5_11[27] , 
        \wRegInTop_5_27[25] , \wRegInBot_5_28[1] , \wRegInTop_6_34[6] , 
        \wRegInTop_7_15[0] , \ScanLink189[8] , \ScanLink146[1] , 
        \wRegInTop_7_109[2] , \wRegOut_7_123[2] , \wRegInTop_2_0[17] , 
        \wRegOut_3_3[30] , \wRegInTop_5_11[20] , \wRegInBot_5_27[22] , 
        \ScanLink78[3] , \ScanLink119[31] , \wRegInTop_6_37[5] , 
        \ScanLink119[28] , \wRegInTop_7_89[24] , \ScanLink226[4] , 
        \wRegInTop_7_16[3] , \ScanLink145[2] , \wRegInTop_7_44[20] , 
        \wRegInTop_7_31[10] , \wRegOut_3_3[29] , \wRegInTop_7_67[11] , 
        \wRegInBot_4_2[24] , \wRegInBot_6_0[8] , \wRegInTop_7_12[21] , 
        \wRegInTop_7_24[24] , \wRegInTop_7_51[14] , \ScanLink197[19] , 
        \wRegInTop_7_72[25] , \ScanLink225[7] , \wRegOut_7_120[1] , 
        \wRegInBot_6_5[20] , \wRegOut_6_38[2] , \wRegOut_7_19[4] , 
        \ScanLink197[4] , \ScanLink238[8] , \wRegOut_7_7[2] , 
        \wRegInTop_3_6[8] , \wRegOut_5_4[10] , \wRegInTop_5_11[13] , 
        \wRegInBot_5_27[11] , \ScanLink94[30] , \ScanLink122[5] , 
        \wRegInTop_6_50[2] , \wRegInTop_7_71[4] , \wRegInTop_7_89[17] , 
        \wRegInBot_5_11[14] , \ScanLink94[29] , \ScanLink242[0] , 
        \wRegInTop_5_27[16] , \wRegOut_6_19[19] , \wRegOut_7_17[30] , 
        \wRegOut_7_34[18] , \wRegOut_7_41[28] , \wRegOut_4_0[0] , 
        \wRegOut_7_41[31] , \wRegOut_7_62[19] , \wRegOut_7_17[29] , 
        \wRegOut_2_3[7] , \ScanLink8[16] , \wRegEnBot_5_2[0] , 
        \wRegOut_4_3[3] , \wRegOut_5_13[8] , \wRegOut_7_3[14] , 
        \wRegInBot_5_4[9] , \wRegOut_5_14[31] , \wRegInTop_6_0[19] , 
        \wRegInTop_7_119[18] , \wRegOut_7_99[18] , \wRegOut_5_14[28] , 
        \wRegInBot_6_5[13] , \wRegOut_3_7[18] , \wRegInBot_4_2[17] , 
        \ScanLink39[30] , \wRegInTop_7_72[16] , \ScanLink39[29] , 
        \wRegInTop_6_53[1] , \wRegInTop_7_24[17] , \wRegInTop_7_72[7] , 
        \ScanLink121[6] , \wRegInTop_7_51[27] , \wRegInTop_7_12[12] , 
        \wRegInTop_7_31[23] , \ScanLink204[28] , \wRegInTop_7_44[13] , 
        \ScanLink252[30] , \ScanLink204[31] , \ScanLink227[19] , 
        \wRegInBot_4_6[26] , \wRegInTop_4_8[5] , \wRegOut_5_10[19] , 
        \wRegInBot_6_1[22] , \wRegInTop_6_4[31] , \wRegInTop_6_4[28] , 
        \wRegOut_6_41[9] , \ScanLink241[3] , \ScanLink252[29] , 
        \wRegInTop_7_67[22] , \wRegOut_7_59[6] , \wRegInTop_7_84[7] , 
        \wRegInTop_5_26[5] , \wRegInTop_7_76[27] , \wRegInBot_4_9[3] , 
        \ScanLink48[31] , \wRegInBot_6_18[14] , \ScanLink48[28] , 
        \wRegOut_7_44[9] , \wRegInTop_7_55[16] , \wRegOut_5_29[2] , 
        \wRegInTop_7_20[26] , \wRegOut_6_8[26] , \wRegInTop_6_18[13] , 
        \ScanLink105[0] , \wRegInTop_7_40[22] , \ScanLink200[19] , 
        \ScanLink223[31] , \wRegInTop_7_99[8] , \wRegInTop_7_35[12] , 
        \wRegInTop_7_56[1] , \wRegInTop_7_63[13] , \ScanLink223[28] , 
        \wRegInBot_4_6[15] , \wRegOut_5_0[21] , \ScanLink38[1] , 
        \wRegInTop_7_16[23] , \wRegInTop_5_15[22] , \wRegInBot_5_23[20] , 
        \ScanLink90[18] , \wRegOut_7_88[3] , \wRegInBot_5_9[25] , 
        \wRegInBot_5_15[25] , \wRegInTop_5_23[27] , \wRegInTop_7_98[12] , 
        \wRegInTop_5_25[6] , \wRegInBot_6_39[1] , \ScanLink106[3] , 
        \wRegInTop_7_55[2] , \wRegOut_7_13[18] , \wRegOut_7_30[29] , 
        \wRegOut_7_45[19] , \wRegOut_7_66[31] , \wRegOut_7_30[30] , 
        \wRegOut_7_66[28] , \wRegOut_6_8[15] , \wRegOut_7_7[25] , 
        \wRegInTop_7_35[21] , \wRegInTop_7_87[4] , \wRegOut_7_104[7] , 
        \wRegInTop_7_40[11] , \wRegInTop_7_16[10] , \ScanLink42[9] , 
        \wRegInBot_6_1[11] , \wRegInTop_6_13[3] , \wRegInTop_6_18[20] , 
        \wRegInBot_6_43[9] , \ScanLink201[1] , \wRegInBot_6_18[27] , 
        \wRegInTop_7_63[20] , \wRegInTop_7_20[15] , \ScanLink193[28] , 
        \wRegInTop_7_76[14] , \wRegEnTop_7_124[0] , \ScanLink193[31] , 
        \wRegInTop_7_32[5] , \wRegInTop_7_55[25] , \ScanLink161[4] , 
        \wRegOut_7_119[8] , \ScanLink6[8] , \wRegOut_2_3[17] , 
        \wRegInBot_3_5[10] , \ScanLink15[16] , \ScanLink20[3] , 
        \wRegOut_5_0[12] , \wRegInBot_5_9[16] , \wRegInBot_5_11[8] , 
        \wRegInBot_5_15[16] , \wRegOut_7_7[16] , \ScanLink202[2] , 
        \wRegInTop_7_98[21] , \wRegInTop_5_15[11] , \wRegInTop_5_23[14] , 
        \wRegOut_7_107[4] , \wRegInBot_5_23[13] , \wRegInTop_6_10[0] , 
        \ScanLink162[7] , \wRegInTop_7_31[6] , \ScanLink168[30] , 
        \ScanLink56[23] , \ScanLink168[29] , \ScanLink23[13] , 
        \wRegOut_4_13[5] , \ScanLink60[26] , \wRegOut_6_3[19] , 
        \ScanLink75[12] , \ScanLink228[17] , \wRegOut_7_90[1] , 
        \ScanLink198[24] , \wRegInTop_4_8[13] , \ScanLink36[27] , 
        \ScanLink43[17] , \wRegInTop_6_25[30] , \ScanLink248[13] , 
        \wRegInTop_6_50[19] , \wRegInTop_7_82[9] , \wRegInBot_6_21[3] , 
        \wRegInTop_6_25[29] , \wRegInTop_7_120[13] , \wRegOut_7_83[22] , 
        \wRegOut_4_15[16] , \wRegOut_6_63[1] , \wRegOut_7_42[7] , 
        \wRegInTop_7_103[22] , \wRegOut_5_8[7] , \wRegOut_7_78[23] , 
        \wRegOut_7_96[16] , \wRegInTop_7_116[16] , \ScanLink7[18] , 
        \wRegInBot_6_22[0] , \wRegOut_6_60[2] , \wRegOut_7_41[4] , 
        \wRegInTop_3_0[30] , \ScanLink23[0] , \wRegOut_4_10[6] , 
        \wRegInTop_5_7[10] , \wRegOut_6_20[12] , \wRegOut_6_35[26] , 
        \wRegOut_6_55[22] , \wRegOut_6_40[16] , \wRegOut_6_16[17] , 
        \ScanLink103[21] , \wRegOut_6_63[27] , \wRegOut_7_18[27] , 
        \ScanLink120[10] , \ScanLink176[11] , \wRegOut_7_93[2] , 
        \wRegOut_5_31[0] , \ScanLink155[20] , \wRegInTop_5_23[8] , 
        \wRegInTop_5_28[18] , \ScanLink116[15] , \ScanLink135[24] , 
        \ScanLink140[14] , \wRegInTop_7_86[19] , \wRegInBot_6_45[7] , 
        \wRegInTop_7_0[14] , \ScanLink163[25] , \wRegInTop_7_116[25] , 
        \wRegOut_7_96[25] , \wRegInTop_3_0[29] , \wRegOut_7_26[3] , 
        \wRegOut_7_102[9] , \wRegInBot_3_5[23] , \wRegOut_4_15[25] , 
        \ScanLink59[8] , \ScanLink96[1] , \wRegOut_7_83[11] , 
        \wRegInTop_7_120[20] , \wRegInTop_7_103[11] , \ScanLink15[25] , 
        \ScanLink23[20] , \wRegInTop_4_8[20] , \ScanLink36[14] , 
        \ScanLink60[15] , \wRegInBot_6_58[8] , \ScanLink248[20] , 
        \wRegInBot_6_13[18] , \wRegInBot_6_30[30] , \ScanLink198[17] , 
        \ScanLink43[24] , \wRegInBot_5_14[5] , \wRegInBot_6_45[19] , 
        \wRegInBot_6_30[29] , \ScanLink44[7] , \wRegEnTop_6_46[0] , 
        \ScanLink47[4] , \wRegInBot_5_17[6] , \ScanLink56[10] , 
        \wRegInTop_7_29[4] , \wRegOut_7_100[29] , \ScanLink75[21] , 
        \wRegOut_7_100[30] , \wRegOut_7_123[18] , \ScanLink228[24] , 
        \ScanLink140[27] , \ScanLink135[17] , \wRegOut_2_3[24] , 
        \wRegInBot_4_10[19] , \wRegOut_6_19[9] , \ScanLink116[26] , 
        \wRegInTop_7_0[27] , \ScanLink163[16] , \ScanLink219[3] , 
        \ScanLink176[22] , \wRegInTop_5_7[23] , \ScanLink103[12] , 
        \ScanLink120[23] , \ScanLink155[13] , \ScanLink179[6] , 
        \wRegOut_6_16[24] , \ScanLink95[2] , \wRegOut_6_35[15] , 
        \wRegOut_6_40[25] , \wRegInBot_6_46[4] , \wRegOut_6_63[14] , 
        \wRegOut_7_18[14] , \wRegOut_7_25[0] , \wRegOut_7_78[10] , 
        \wRegInBot_3_1[10] , \ScanLink11[16] , \wRegInBot_4_9[19] , 
        \wRegInBot_4_11[7] , \ScanLink27[13] , \wRegInBot_5_2[30] , 
        \wRegInBot_5_2[29] , \wRegOut_6_55[11] , \wRegInTop_7_9[9] , 
        \ScanLink164[9] , \wRegInTop_7_37[8] , \ScanLink60[3] , 
        \wRegOut_6_20[21] , \wRegOut_6_7[19] , \wRegInBot_5_30[1] , 
        \wRegInTop_7_111[2] , \ScanLink52[23] , \ScanLink71[12] , 
        \ScanLink189[10] , \wRegInTop_7_79[18] , \wRegOut_4_11[16] , 
        \wRegEnTop_4_12[0] , \ScanLink32[27] , \ScanLink64[26] , 
        \wRegInTop_6_21[30] , \ScanLink239[23] , \ScanLink47[17] , 
        \wRegInTop_6_7[2] , \wRegInTop_6_21[29] , \ScanLink191[8] , 
        \wRegInBot_6_6[4] , \wRegInTop_6_54[19] , \wRegOut_7_87[22] , 
        \wRegInTop_7_124[13] , \wRegOut_6_23[1] , \wRegInTop_7_107[22] , 
        \wRegInTop_6_31[9] , \wRegInBot_6_61[3] , \wRegOut_7_92[16] , 
        \wRegInTop_7_112[16] , \wRegOut_0_0[13] , \ScanLink3[18] , 
        \wRegOut_5_29[23] , \wRegOut_6_20[2] , \ScanLink220[8] , 
        \wRegInBot_4_12[4] , \wRegInTop_5_3[10] , \wRegOut_6_24[12] , 
        \wRegOut_6_51[22] , \wRegInBot_6_62[0] , \ScanLink63[0] , 
        \wRegOut_6_12[17] , \wRegOut_6_31[26] , \wRegOut_6_44[16] , 
        \ScanLink107[21] , \ScanLink172[11] , \wRegOut_7_69[17] , 
        \ScanLink151[20] , \ScanLink124[10] , \wRegInTop_7_112[1] , 
        \wRegInTop_3_4[30] , \wRegInTop_6_4[1] , \ScanLink144[14] , 
        \wRegInBot_6_5[7] , \ScanLink112[15] , \ScanLink131[24] , 
        \wRegInTop_7_4[14] , \ScanLink167[25] , \wRegInTop_7_82[19] , 
        \wRegOut_7_66[3] , \wRegOut_6_47[5] , \wRegOut_7_92[25] , 
        \wRegInTop_7_112[25] , \wRegOut_0_0[20] , \wRegInTop_3_0[4] , 
        \wRegInBot_3_1[23] , \wRegInTop_3_4[29] , \ScanLink19[8] , 
        \wRegOut_5_29[10] , \wRegInTop_5_19[0] , \wRegInTop_7_124[20] , 
        \wRegOut_7_87[11] , \wRegInBot_3_1[2] , \wRegInBot_3_2[1] , 
        \ScanLink11[25] , \wRegOut_4_11[25] , \wRegInTop_7_107[11] , 
        \wRegInTop_5_3[3] , \wRegInBot_6_17[18] , \ScanLink64[15] , 
        \wRegInBot_6_34[30] , \ScanLink239[10] , \ScanLink27[20] , 
        \ScanLink32[14] , \wRegInBot_5_2[5] , \wRegInBot_6_62[28] , 
        \ScanLink47[24] , \wRegInBot_6_18[8] , \wRegOut_5_16[7] , 
        \wRegInBot_6_34[29] , \wRegInBot_6_41[19] , \ScanLink52[10] , 
        \wRegInTop_6_48[2] , \wRegInBot_6_62[31] , \wRegInTop_7_69[4] , 
        \wRegOut_7_104[29] , \wRegInTop_3_3[7] , \ScanLink71[21] , 
        \ScanLink189[23] , \wRegInTop_5_0[0] , \wRegOut_5_15[4] , 
        \ScanLink131[17] , \wRegOut_7_104[30] , \wRegOut_7_127[18] , 
        \wRegOut_6_59[9] , \ScanLink144[27] , \wRegInBot_5_1[6] , 
        \ScanLink112[26] , \ScanLink107[12] , \wRegInTop_7_4[27] , 
        \ScanLink167[16] , \wRegInBot_4_14[19] , \ScanLink172[22] , 
        \ScanLink124[23] , \ScanLink139[6] , \ScanLink0[4] , \wRegOut_2_0[6] , 
        \wRegInTop_2_0[26] , \wRegInBot_4_2[26] , \wRegInTop_5_3[23] , 
        \wRegOut_6_31[15] , \ScanLink151[13] , \wRegOut_6_44[25] , 
        \wRegInBot_5_6[30] , \wRegInBot_5_6[29] , \wRegOut_6_12[24] , 
        \wRegOut_6_44[6] , \wRegOut_7_65[0] , \wRegOut_7_69[24] , 
        \wRegOut_6_24[21] , \ScanLink124[9] , \wRegOut_7_8[30] , 
        \wRegInTop_7_77[8] , \ScanLink39[18] , \wRegOut_5_14[19] , 
        \wRegInTop_6_0[31] , \wRegInTop_6_0[28] , \wRegOut_6_38[0] , 
        \wRegOut_6_51[11] , \wRegOut_7_8[29] , \wRegOut_7_19[6] , 
        \wRegOut_7_7[0] , \wRegOut_7_99[29] , \wRegInTop_7_119[29] , 
        \wRegEnBot_6_5[0] , \wRegInBot_6_5[22] , \ScanLink197[6] , 
        \wRegOut_7_99[30] , \wRegInTop_7_119[30] , \wRegEnBot_6_34[0] , 
        \wRegInTop_7_24[26] , \wRegInTop_7_72[27] , \ScanLink225[5] , 
        \wRegInTop_7_51[16] , \wRegOut_7_120[3] , \wRegInTop_6_37[7] , 
        \ScanLink145[0] , \ScanLink204[19] , \ScanLink227[31] , 
        \wRegInTop_7_12[23] , \wRegInTop_7_16[1] , \wRegInTop_7_31[12] , 
        \wRegInTop_7_44[22] , \ScanLink227[28] , \wRegInTop_7_67[13] , 
        \ScanLink252[18] , \wRegOut_2_3[5] , \ScanLink8[27] , 
        \wRegOut_5_4[21] , \wRegInTop_5_11[22] , \wRegInBot_5_27[20] , 
        \wRegInBot_5_28[3] , \ScanLink78[1] , \ScanLink94[18] , 
        \wRegInTop_7_89[26] , \wRegInTop_7_109[0] , \wRegOut_7_123[0] , 
        \ScanLink226[6] , \wRegInBot_5_11[25] , \wRegInTop_5_27[27] , 
        \wRegInTop_6_34[4] , \wRegInTop_7_15[2] , \ScanLink146[3] , 
        \wRegOut_6_19[31] , \wRegOut_6_19[28] , \wRegOut_7_4[3] , 
        \wRegOut_7_34[29] , \wRegOut_7_41[19] , \wRegOut_7_62[31] , 
        \wRegOut_7_17[18] , \wRegOut_7_34[30] , \wRegOut_7_62[28] , 
        \wRegOut_3_3[18] , \wRegInBot_4_2[15] , \wRegInBot_6_3[9] , 
        \ScanLink194[5] , \wRegOut_7_3[25] , \wRegInTop_7_31[21] , 
        \wRegInTop_7_44[11] , \wRegInTop_7_67[20] , \ScanLink241[1] , 
        \wRegOut_5_10[9] , \wRegInTop_6_53[3] , \wRegInTop_7_12[10] , 
        \wRegInTop_7_51[25] , \ScanLink197[28] , \wRegInTop_7_72[14] , 
        \wRegInTop_7_72[5] , \ScanLink121[4] , \wRegInTop_7_24[15] , 
        \ScanLink197[31] , \wRegInBot_6_5[11] , \ScanLink8[14] , 
        \wRegInTop_3_5[9] , \wRegOut_4_3[1] , \wRegInBot_5_7[8] , 
        \wRegInTop_2_0[15] , \wRegEnTop_3_3[0] , \wRegOut_4_0[2] , 
        \wRegOut_7_3[16] , \wRegOut_5_4[12] , \wRegInBot_5_11[16] , 
        \wRegOut_6_42[8] , \ScanLink242[2] , \wRegInTop_5_27[14] , 
        \wRegInTop_6_50[0] , \ScanLink122[7] , \wRegInTop_7_71[6] , 
        \wRegOut_3_7[30] , \wRegOut_5_0[23] , \wRegInBot_5_9[27] , 
        \wRegInTop_5_11[11] , \wRegInBot_5_27[13] , \wRegInTop_5_25[4] , 
        \ScanLink119[19] , \wRegInTop_7_89[15] , \wRegInBot_5_15[27] , 
        \wRegInBot_6_39[3] , \wRegOut_7_7[27] , \wRegInTop_7_87[6] , 
        \wRegInTop_7_98[10] , \ScanLink38[3] , \wRegInTop_5_23[25] , 
        \ScanLink106[1] , \wRegInTop_7_55[0] , \wRegInBot_5_23[22] , 
        \wRegInTop_5_15[20] , \wRegOut_7_47[8] , \wRegOut_7_88[1] , 
        \ScanLink105[2] , \ScanLink168[18] , \wRegOut_3_7[29] , 
        \wRegEnBot_5_25[0] , \wRegInTop_7_35[10] , \wRegInTop_7_40[20] , 
        \wRegInTop_7_56[3] , \wRegOut_6_8[24] , \wRegInTop_7_16[21] , 
        \wRegInBot_4_6[24] , \wRegInTop_4_8[7] , \wRegInBot_4_9[1] , 
        \wRegInTop_6_18[11] , \wRegInTop_7_63[11] , \wRegInBot_6_18[16] , 
        \ScanLink193[19] , \wRegInTop_7_76[25] , \wRegOut_4_15[9] , 
        \wRegInTop_5_26[7] , \wRegOut_5_29[0] , \wRegInTop_7_20[24] , 
        \wRegInBot_6_1[20] , \wRegInTop_7_55[14] , \wRegInTop_7_84[5] , 
        \wRegOut_7_59[4] , \wRegOut_5_0[10] , \wRegInTop_5_15[13] , 
        \wRegInBot_5_23[11] , \wRegInTop_6_10[2] , \ScanLink90[30] , 
        \wRegInTop_7_31[4] , \ScanLink162[5] , \ScanLink90[29] , 
        \wRegInBot_5_15[14] , \wRegInBot_6_40[8] , \ScanLink202[0] , 
        \wRegInTop_5_23[16] , \wRegInTop_7_98[23] , \wRegOut_6_9[9] , 
        \wRegOut_7_107[6] , \wRegOut_7_13[30] , \wRegOut_7_13[29] , 
        \wRegOut_7_30[18] , \wRegOut_7_45[28] , \wRegOut_7_45[31] , 
        \wRegOut_7_66[19] , \wRegInBot_1_0[1] , \wRegInTop_1_1[7] , 
        \ScanLink3[7] , \wRegInBot_5_9[14] , \ScanLink41[8] , 
        \wRegOut_5_10[31] , \wRegInTop_6_4[19] , \wRegOut_7_7[14] , 
        \wRegOut_5_10[28] , \wRegInBot_5_12[9] , \wRegInBot_6_1[13] , 
        \ScanLink5[9] , \wRegOut_2_3[26] , \wRegOut_2_3[15] , 
        \wRegInBot_4_6[17] , \ScanLink48[19] , \wRegInTop_6_13[1] , 
        \wRegInBot_6_18[25] , \wRegInTop_7_76[16] , \wRegInTop_7_32[7] , 
        \wRegInTop_7_55[27] , \wRegInTop_7_20[17] , \ScanLink161[6] , 
        \wRegOut_6_8[17] , \wRegInTop_6_18[22] , \wRegInTop_7_35[23] , 
        \wRegInTop_7_40[13] , \ScanLink200[28] , \wRegOut_7_104[5] , 
        \wRegInTop_7_63[22] , \ScanLink201[3] , \ScanLink200[31] , 
        \ScanLink223[19] , \ScanLink23[2] , \wRegOut_4_10[4] , 
        \wRegInBot_4_10[28] , \ScanLink116[17] , \wRegInTop_7_0[16] , 
        \ScanLink135[26] , \ScanLink140[16] , \wRegInTop_7_16[12] , 
        \wRegInTop_7_81[8] , \ScanLink163[27] , \ScanLink176[13] , 
        \wRegOut_5_31[2] , \ScanLink103[23] , \wRegOut_7_93[0] , 
        \ScanLink155[22] , \wRegInBot_4_10[31] , \wRegInBot_5_2[18] , 
        \wRegInTop_5_7[12] , \ScanLink120[12] , \wRegOut_6_16[15] , 
        \wRegOut_6_35[24] , \wRegOut_6_40[14] , \wRegOut_6_63[25] , 
        \wRegOut_7_18[25] , \wRegInBot_6_22[2] , \wRegOut_6_60[0] , 
        \wRegOut_7_41[6] , \wRegOut_7_78[21] , \wRegInTop_3_0[18] , 
        \wRegEnTop_4_8[0] , \wRegOut_5_8[5] , \wRegOut_6_20[10] , 
        \wRegOut_6_55[20] , \wRegOut_7_96[14] , \wRegInTop_7_116[14] , 
        \wRegInBot_3_5[12] , \wRegOut_4_15[14] , \wRegOut_7_83[20] , 
        \wRegInTop_7_120[11] , \wRegOut_6_63[3] , \wRegInTop_7_103[20] , 
        \wRegOut_7_42[5] , \ScanLink15[14] , \wRegInBot_6_21[1] , 
        \ScanLink20[1] , \wRegInTop_4_8[11] , \wRegInTop_5_20[9] , 
        \wRegInBot_6_45[31] , \ScanLink248[11] , \ScanLink60[24] , 
        \wRegInBot_6_13[29] , \ScanLink198[26] , \ScanLink36[25] , 
        \ScanLink43[15] , \wRegInBot_6_30[18] , \wRegInBot_6_45[28] , 
        \wRegInBot_6_13[30] , \ScanLink23[11] , \wRegOut_4_13[7] , 
        \wRegOut_7_123[30] , \ScanLink56[21] , \wRegOut_7_100[18] , 
        \ScanLink75[10] , \wRegOut_7_90[3] , \ScanLink228[15] , 
        \wRegOut_7_123[29] , \wRegOut_7_78[12] , \ScanLink7[30] , 
        \ScanLink7[29] , \wRegOut_6_20[23] , \ScanLink15[27] , 
        \ScanLink23[22] , \wRegInTop_5_7[21] , \ScanLink95[0] , 
        \wRegOut_6_35[17] , \wRegOut_6_55[13] , \wRegOut_6_40[27] , 
        \ScanLink47[6] , \wRegInTop_5_28[30] , \wRegOut_6_16[26] , 
        \wRegOut_7_101[8] , \ScanLink103[10] , \wRegInBot_6_46[6] , 
        \wRegOut_6_63[16] , \wRegOut_7_25[2] , \wRegOut_7_18[16] , 
        \ScanLink176[20] , \wRegInTop_5_28[29] , \ScanLink120[21] , 
        \ScanLink155[11] , \ScanLink179[4] , \wRegInTop_7_86[31] , 
        \wRegInBot_5_17[4] , \ScanLink135[15] , \ScanLink56[12] , 
        \ScanLink116[24] , \ScanLink140[25] , \wRegInTop_7_86[28] , 
        \ScanLink219[1] , \wRegInTop_7_0[25] , \wRegInTop_7_29[6] , 
        \ScanLink163[14] , \ScanLink60[17] , \wRegOut_6_3[31] , 
        \wRegOut_6_3[28] , \ScanLink75[23] , \ScanLink228[26] , 
        \wRegInTop_6_50[31] , \ScanLink198[15] , \wRegInBot_3_5[21] , 
        \wRegInTop_4_8[22] , \ScanLink43[26] , \ScanLink248[22] , 
        \ScanLink44[5] , \wRegInTop_6_50[28] , \ScanLink36[16] , 
        \wRegInBot_5_14[7] , \wRegInTop_6_25[18] , \wRegInTop_7_34[9] , 
        \ScanLink167[8] , \wRegOut_7_83[13] , \wRegInTop_7_120[22] , 
        \wRegOut_3_6[10] , \wRegInTop_4_2[17] , \wRegOut_4_15[27] , 
        \wRegEnTop_5_17[0] , \wRegOut_7_26[1] , \wRegInTop_7_103[13] , 
        \ScanLink96[3] , \wRegInBot_6_45[5] , \wRegOut_7_96[27] , 
        \wRegInTop_7_116[27] , \ScanLink49[13] , \wRegOut_6_11[3] , 
        \wRegOut_7_30[5] , \ScanLink192[20] , \ScanLink214[16] , 
        \ScanLink237[27] , \ScanLink242[17] , \ScanLink211[9] , 
        \wRegInTop_6_19[28] , \wRegInTop_7_17[18] , \ScanLink187[14] , 
        \wRegInTop_7_62[28] , \ScanLink222[13] , \ScanLink29[17] , 
        \ScanLink80[7] , \wRegInBot_6_53[1] , \wRegInTop_7_34[30] , 
        \wRegInTop_6_19[31] , \wRegInTop_7_41[19] , \wRegOut_5_11[22] , 
        \wRegOut_5_27[27] , \wRegInTop_7_34[29] , \wRegInTop_7_62[31] , 
        \ScanLink201[22] , \wRegInTop_6_5[13] , \wRegInTop_7_1[3] , 
        \wRegOut_7_89[26] , \wRegInTop_7_109[26] , \ScanLink52[1] , 
        \wRegEnTop_7_71[0] , \wRegOut_7_109[0] , \wRegInTop_7_123[0] , 
        \wRegOut_1_1[27] , \wRegOut_1_1[14] , \wRegInBot_6_0[19] , 
        \wRegInBot_2_0[17] , \wRegInTop_5_14[19] , \ScanLink51[2] , 
        \wRegInTop_7_2[0] , \wRegOut_7_12[23] , \wRegOut_7_31[12] , 
        \wRegOut_7_67[13] , \wRegOut_7_44[22] , \ScanLink91[23] , 
        \wRegOut_7_24[26] , \wRegOut_7_51[16] , \wRegOut_7_72[27] , 
        \wRegInTop_7_120[3] , \wRegOut_6_12[0] , \ScanLink83[4] , 
        \ScanLink169[21] , \ScanLink84[17] , \wRegInTop_7_99[30] , 
        \wRegOut_7_33[6] , \wRegOut_5_11[11] , \ScanLink109[25] , 
        \wRegInBot_6_50[2] , \wRegInTop_7_99[29] , \ScanLink108[7] , 
        \wRegOut_7_89[15] , \wRegInTop_7_109[15] , \wRegEnTop_1_1[0] , 
        \wRegInBot_2_0[24] , \wRegOut_3_6[23] , \wRegInBot_4_4[4] , 
        \ScanLink36[5] , \wRegOut_5_24[5] , \wRegOut_5_27[14] , 
        \wRegInTop_4_5[2] , \wRegInTop_6_5[20] , \wRegOut_7_86[7] , 
        \ScanLink187[27] , \ScanLink222[20] , \wRegInTop_4_2[24] , 
        \ScanLink29[24] , \ScanLink115[8] , \ScanLink201[11] , 
        \wRegInTop_7_89[0] , \wRegInTop_7_46[9] , \ScanLink49[20] , 
        \ScanLink214[25] , \wRegOut_5_1[30] , \wRegInBot_6_37[5] , 
        \wRegOut_7_54[1] , \ScanLink237[14] , \ScanLink192[13] , 
        \ScanLink242[24] , \wRegOut_5_1[29] , \wRegInTop_5_28[1] , 
        \ScanLink109[16] , \wRegOut_3_0[9] , \wRegInBot_4_7[7] , 
        \ScanLink28[9] , \wRegInBot_5_22[31] , \ScanLink84[24] , 
        \wRegOut_7_57[2] , \ScanLink91[10] , \wRegInBot_6_34[6] , 
        \ScanLink169[12] , \wRegInTop_4_14[8] , \wRegInBot_5_22[28] , 
        \wRegOut_7_24[15] , \wRegOut_7_51[25] , \wRegInTop_7_58[5] , 
        \wRegOut_7_72[14] , \wRegInTop_3_1[21] , \wRegOut_4_5[26] , 
        \wRegInTop_4_6[1] , \wRegOut_7_67[20] , \wRegOut_7_85[4] , 
        \ScanLink35[6] , \wRegOut_5_27[6] , \wRegInBot_6_29[9] , 
        \wRegOut_7_12[10] , \wRegOut_7_44[11] , \wRegOut_7_31[21] , 
        \wRegOut_7_82[19] , \wRegInTop_7_102[19] , \wRegInTop_7_24[3] , 
        \wRegInTop_7_121[31] , \ScanLink177[2] , \wRegInTop_7_121[28] , 
        \ScanLink22[31] , \ScanLink49[0] , \ScanLink86[9] , 
        \wRegInBot_5_19[2] , \wRegOut_7_112[1] , \ScanLink74[29] , 
        \ScanLink217[7] , \wRegInTop_6_12[17] , \wRegInTop_7_69[17] , 
        \wRegOut_7_122[10] , \ScanLink22[28] , \ScanLink57[18] , 
        \wRegInTop_6_44[16] , \wRegOut_6_2[22] , \ScanLink74[30] , 
        \wRegInBot_6_24[15] , \wRegInTop_6_31[26] , \wRegInBot_6_51[25] , 
        \wRegInTop_4_9[31] , \wRegInTop_4_9[28] , \wRegInBot_6_31[21] , 
        \wRegOut_7_101[21] , \wRegInTop_6_51[22] , \wRegOut_7_114[15] , 
        \wRegOut_6_1[1] , \wRegInBot_6_44[11] , \wRegInBot_6_12[10] , 
        \wRegInTop_6_24[12] , \ScanLink249[31] , \wRegInTop_4_11[16] , 
        \wRegInBot_4_11[11] , \wRegInTop_5_29[23] , \wRegInBot_6_48[0] , 
        \ScanLink249[28] , \wRegInTop_7_92[16] , \wRegOut_7_28[7] , 
        \wRegInTop_7_87[22] , \ScanLink6[23] , \wRegInBot_5_3[21] , 
        \wRegInBot_5_29[24] , \ScanLink98[5] , \wRegOut_6_2[2] , 
        \wRegOut_6_21[29] , \wRegInTop_7_27[0] , \ScanLink174[1] , 
        \wRegOut_6_54[19] , \wRegOut_7_79[18] , \wRegOut_6_21[30] , 
        \wRegInTop_2_3[8] , \wRegInTop_6_24[21] , \wRegInBot_6_44[22] , 
        \wRegOut_7_35[8] , \ScanLink214[4] , \wRegOut_7_111[2] , 
        \wRegInTop_7_92[1] , \wRegOut_7_114[26] , \wRegInBot_6_31[12] , 
        \wRegInTop_6_51[11] , \wRegOut_3_5[4] , \wRegInTop_4_11[5] , 
        \wRegInTop_5_30[3] , \wRegOut_5_5[0] , \wRegInBot_6_12[23] , 
        \wRegInTop_6_12[24] , \wRegOut_7_80[9] , \wRegEnBot_4_7[0] , 
        \wRegOut_6_2[11] , \wRegInTop_6_31[15] , \wRegInTop_7_69[24] , 
        \wRegOut_7_122[23] , \wRegInBot_6_51[16] , \wRegOut_7_101[12] , 
        \wRegInBot_6_24[26] , \wRegInTop_6_44[25] , \wRegInBot_1_0[8] , 
        \ScanLink2[21] , \ScanLink6[10] , \wRegInTop_3_1[12] , 
        \ScanLink113[6] , \wRegInTop_6_61[1] , \wRegInTop_7_40[7] , 
        \wRegInBot_3_4[18] , \wRegOut_4_5[15] , \wRegInTop_5_6[18] , 
        \wRegInTop_6_62[2] , \ScanLink110[5] , \wRegInTop_7_43[4] , 
        \wRegOut_3_6[7] , \wRegInTop_4_11[25] , \wRegInTop_4_12[6] , 
        \wRegInBot_5_3[12] , \wRegInBot_6_32[8] , \wRegOut_5_6[3] , 
        \wRegInTop_7_87[11] , \ScanLink33[8] , \wRegOut_5_21[8] , 
        \wRegInBot_5_29[17] , \wRegInTop_7_91[2] , \ScanLink154[28] , 
        \wRegInTop_5_29[10] , \ScanLink102[30] , \ScanLink121[18] , 
        \ScanLink154[31] , \ScanLink177[19] , \wRegInBot_4_1[9] , 
        \wRegInBot_4_11[22] , \wRegInTop_5_2[30] , \ScanLink102[29] , 
        \wRegInTop_7_92[25] , \ScanLink254[6] , \wRegInTop_5_2[29] , 
        \wRegOut_5_18[1] , \wRegEnTop_7_29[0] , \wRegInBot_5_7[23] , 
        \wRegInTop_6_46[4] , \ScanLink134[3] , \wRegInTop_7_67[2] , 
        \wRegOut_7_9[23] , \ScanLink2[12] , \wRegInBot_3_0[30] , 
        \wRegInBot_3_0[29] , \wRegInTop_3_5[23] , \wRegInBot_4_8[20] , 
        \wRegInTop_4_15[14] , \wRegOut_7_68[5] , \wRegInTop_7_83[20] , 
        \ScanLink249[9] , \wRegInBot_4_15[13] , \wRegInTop_5_17[6] , 
        \ScanLink106[18] , \wRegOut_6_49[3] , \ScanLink125[30] , 
        \ScanLink125[29] , \ScanLink150[19] , \ScanLink173[31] , 
        \wRegInTop_7_96[14] , \ScanLink173[28] , \wRegInTop_5_14[5] , 
        \wRegInBot_6_16[12] , \wRegInTop_6_20[10] , \wRegInBot_6_35[23] , 
        \wRegInBot_6_40[13] , \wRegInTop_6_55[20] , \wRegOut_7_110[17] , 
        \wRegInTop_6_63[25] , \wRegInBot_6_63[22] , \ScanLink188[29] , 
        \wRegInTop_7_78[21] , \wRegInTop_7_18[25] , \wRegOut_6_6[20] , 
        \wRegInTop_6_16[15] , \wRegInBot_6_20[17] , \wRegInTop_6_40[14] , 
        \wRegEnBot_6_46[0] , \ScanLink188[30] , \wRegOut_7_126[12] , 
        \wRegInTop_6_58[8] , \wRegInTop_6_35[24] , \wRegInBot_6_55[27] , 
        \wRegOut_7_105[23] , \wRegOut_4_1[24] , \wRegOut_7_76[9] , 
        \wRegInTop_6_45[7] , \wRegInTop_7_64[1] , \ScanLink137[0] , 
        \wRegInTop_4_15[27] , \wRegInBot_4_15[20] , \wRegInBot_5_23[8] , 
        \wRegInTop_7_83[13] , \wRegInTop_7_96[27] , \wRegOut_6_25[18] , 
        \wRegOut_6_50[28] , \wRegOut_7_9[10] , \ScanLink182[1] , 
        \wRegOut_6_30[8] , \ScanLink230[2] , \wRegInTop_2_0[2] , 
        \wRegOut_2_2[16] , \wRegInBot_2_2[7] , \wRegInTop_2_3[1] , 
        \wRegOut_3_2[21] , \wRegOut_3_2[12] , \ScanLink11[0] , 
        \wRegInTop_3_5[10] , \wRegOut_4_1[17] , \wRegInBot_5_7[10] , 
        \wRegOut_6_50[31] , \wRegInBot_6_8[2] , \wRegInTop_6_9[4] , 
        \wRegInTop_6_22[0] , \ScanLink150[7] , \wRegOut_7_86[28] , 
        \ScanLink233[1] , \wRegInTop_6_21[3] , \ScanLink153[4] , 
        \wRegOut_7_86[31] , \wRegInTop_7_106[28] , \wRegInTop_7_106[31] , 
        \wRegInTop_7_125[19] , \wRegInBot_4_8[13] , \wRegOut_5_28[30] , 
        \wRegOut_5_28[29] , \wRegEnTop_7_116[0] , \wRegInTop_6_16[26] , 
        \wRegInTop_6_63[16] , \wRegOut_7_126[21] , \ScanLink26[19] , 
        \ScanLink53[30] , \ScanLink70[18] , \wRegInTop_7_18[16] , 
        \ScanLink70[9] , \wRegInTop_6_35[17] , \wRegOut_7_105[10] , 
        \wRegOut_5_5[18] , \ScanLink53[29] , \wRegOut_6_6[13] , 
        \wRegInBot_6_20[24] , \wRegInTop_6_40[27] , \wRegInBot_6_55[14] , 
        \wRegInTop_7_101[8] , \wRegInBot_6_16[21] , \wRegInTop_6_20[23] , 
        \wRegInBot_6_40[20] , \ScanLink181[2] , \wRegOut_7_110[24] , 
        \wRegInBot_6_35[10] , \wRegInTop_6_55[13] , \wRegInBot_6_63[11] , 
        \wRegInTop_7_78[12] , \ScanLink238[30] , \ScanLink80[15] , 
        \ScanLink178[17] , \ScanLink238[29] , \wRegOut_7_73[4] , 
        \wRegOut_6_52[2] , \ScanLink252[8] , \wRegInBot_5_26[19] , 
        \wRegInBot_6_10[0] , \ScanLink95[21] , \ScanLink118[13] , 
        \ScanLink12[3] , \wRegInTop_5_9[16] , \wRegInTop_5_11[8] , 
        \wRegOut_7_20[24] , \wRegOut_7_55[14] , \wRegOut_7_76[25] , 
        \wRegOut_6_18[11] , \wRegOut_7_16[21] , \wRegOut_7_63[11] , 
        \wRegOut_5_15[20] , \wRegOut_7_35[10] , \wRegOut_7_40[20] , 
        \wRegInTop_5_8[8] , \wRegOut_5_23[25] , \wRegInTop_6_1[11] , 
        \wRegInTop_7_118[10] , \wRegOut_7_70[7] , \wRegOut_7_98[10] , 
        \ScanLink253[21] , \wRegOut_6_51[1] , \ScanLink183[16] , 
        \ScanLink226[11] , \wRegInTop_4_6[26] , \wRegInTop_4_6[15] , 
        \ScanLink58[25] , \wRegInBot_6_13[3] , \ScanLink205[20] , 
        \wRegInTop_6_43[9] , \ScanLink38[21] , \wRegInTop_5_9[25] , 
        \ScanLink75[4] , \wRegOut_6_18[22] , \ScanLink196[22] , 
        \ScanLink210[14] , \ScanLink233[25] , \ScanLink246[15] , 
        \wRegOut_7_16[12] , \wRegOut_7_63[22] , \wRegOut_7_40[13] , 
        \wRegInTop_5_10[31] , \wRegInTop_5_10[28] , \wRegInBot_5_25[6] , 
        \wRegOut_6_36[6] , \wRegInTop_6_39[1] , \wRegOut_7_35[23] , 
        \wRegInTop_7_104[5] , \wRegInTop_7_18[7] , \wEnable_3[0] , 
        \wRegOut_7_20[17] , \wRegOut_7_55[27] , \wRegOut_7_76[16] , 
        \ScanLink118[20] , \wRegOut_7_17[0] , \ScanLink95[12] , 
        \wRegOut_7_9[6] , \ScanLink80[26] , \ScanLink156[9] , \ScanLink199[0] , 
        \ScanLink178[24] , \ScanLink210[27] , \wRegEnTop_7_87[0] , 
        \ScanLink38[12] , \wRegOut_6_35[5] , \wRegOut_7_14[3] , 
        \ScanLink183[25] , \ScanLink196[11] , \ScanLink233[16] , 
        \ScanLink246[26] , \ScanLink226[22] , \wRegInBot_4_2[3] , 
        \wRegOut_5_15[13] , \wRegOut_5_23[16] , \ScanLink58[16] , 
        \wRegInTop_7_13[29] , \wRegInTop_7_30[18] , \wRegInTop_7_45[31] , 
        \wRegInTop_7_66[19] , \ScanLink253[12] , \ScanLink205[13] , 
        \ScanLink76[7] , \wRegInTop_7_13[30] , \wRegInTop_7_45[28] , 
        \wRegInBot_5_26[5] , \wRegInTop_6_1[22] , \ScanLink228[0] , 
        \wRegInTop_7_107[6] , \wRegInTop_7_118[23] , \wRegOut_7_98[23] , 
        \wRegInBot_6_4[31] , \wRegInBot_6_4[28] , \ScanLink148[5] , 
        \wRegInTop_4_3[5] , \wRegOut_7_80[0] , \ScanLink229[16] , 
        \ScanLink22[12] , \ScanLink30[2] , \ScanLink74[13] , \wRegOut_5_22[2] , 
        \wRegOut_6_2[18] , \wRegInTop_4_9[12] , \ScanLink57[22] , 
        \wRegInTop_7_92[8] , \ScanLink37[26] , \ScanLink42[16] , 
        \wRegInTop_6_24[28] , \wRegInTop_6_51[18] , \ScanLink14[17] , 
        \ScanLink61[27] , \wRegInTop_6_24[31] , \ScanLink249[12] , 
        \ScanLink6[19] , \wRegInBot_3_4[11] , \wRegOut_4_14[17] , 
        \wRegOut_5_5[9] , \ScanLink199[25] , \wRegOut_7_82[23] , 
        \wRegInTop_7_102[23] , \wRegOut_6_21[13] , \wRegInBot_6_31[2] , 
        \wRegOut_7_52[6] , \wRegOut_6_54[23] , \wRegInTop_6_61[8] , 
        \wRegInTop_7_121[12] , \wRegOut_7_97[17] , \wRegInTop_7_117[17] , 
        \wRegOut_7_51[5] , \wRegOut_7_79[22] , \wRegInTop_4_0[6] , 
        \wRegInBot_4_1[0] , \ScanLink33[1] , \wRegInTop_5_6[11] , 
        \wRegOut_6_17[16] , \wRegInBot_6_32[1] , \wRegOut_6_62[26] , 
        \wRegOut_7_19[26] , \wRegOut_6_41[17] , \wRegOut_5_21[1] , 
        \wRegOut_6_34[27] , \wRegInTop_5_29[19] , \ScanLink154[21] , 
        \ScanLink121[11] , \wRegEnTop_7_10[0] , \ScanLink177[10] , 
        \wRegOut_7_83[3] , \ScanLink102[20] , \wRegInTop_7_1[15] , 
        \wRegInBot_2_1[4] , \ScanLink162[24] , \wRegOut_2_2[25] , 
        \ScanLink8[5] , \wRegInTop_3_1[31] , \wRegInTop_3_1[28] , 
        \ScanLink86[0] , \ScanLink117[14] , \wRegInTop_7_87[18] , 
        \ScanLink134[25] , \ScanLink141[15] , \ScanLink49[9] , 
        \wRegOut_6_17[4] , \wRegOut_7_36[2] , \wRegOut_7_112[8] , 
        \wRegOut_7_97[24] , \wRegInTop_7_117[24] , \wRegInBot_3_4[22] , 
        \wRegInBot_6_55[6] , \wRegOut_7_82[10] , \ScanLink14[24] , 
        \wRegInTop_4_9[21] , \wRegOut_4_14[24] , \ScanLink42[25] , 
        \wRegInTop_7_102[10] , \wRegInTop_7_121[21] , \ScanLink54[6] , 
        \wRegInBot_6_31[28] , \wRegInBot_6_44[18] , \ScanLink37[15] , 
        \ScanLink61[14] , \wRegOut_6_1[8] , \wRegInTop_7_125[7] , 
        \wRegInBot_6_12[19] , \wRegInBot_6_31[31] , \ScanLink199[16] , 
        \ScanLink22[21] , \ScanLink57[11] , \ScanLink74[20] , 
        \wRegInBot_6_48[9] , \ScanLink229[25] , \ScanLink249[21] , 
        \wRegInTop_6_18[3] , \wRegInTop_7_39[5] , \wRegOut_7_101[31] , 
        \wRegOut_7_122[19] , \wRegInBot_4_11[18] , \ScanLink57[5] , 
        \ScanLink117[27] , \wRegInTop_7_7[4] , \wRegOut_7_101[28] , 
        \ScanLink209[2] , \wRegInTop_7_1[26] , \ScanLink162[17] , 
        \ScanLink102[13] , \ScanLink121[22] , \ScanLink134[16] , 
        \ScanLink141[26] , \wRegInTop_7_126[4] , \wRegInTop_7_4[7] , 
        \ScanLink154[12] , \ScanLink169[7] , \ScanLink177[23] , 
        \wRegInBot_5_3[31] , \wRegInTop_5_6[22] , \wRegOut_6_14[7] , 
        \wRegOut_6_17[25] , \wRegOut_7_35[1] , \ScanLink85[3] , 
        \wRegOut_6_34[14] , \wRegInBot_6_56[5] , \wRegOut_6_62[15] , 
        \wRegOut_7_19[15] , \wRegOut_6_21[20] , \wRegOut_6_41[24] , 
        \ScanLink174[8] , \wRegOut_6_54[10] , \wRegInTop_7_27[9] , 
        \wRegOut_7_79[11] , \wRegEnBot_2_2[0] , \wRegOut_3_0[0] , 
        \wRegOut_3_3[3] , \wRegInBot_5_3[28] , \wRegInTop_6_5[30] , 
        \wRegInBot_4_7[27] , \wRegOut_5_3[7] , \wRegOut_5_11[18] , 
        \wRegInTop_6_5[29] , \wRegOut_7_49[7] , \ScanLink49[30] , 
        \ScanLink49[29] , \wRegInBot_6_0[23] , \wRegInTop_7_94[6] , 
        \wRegInTop_7_21[27] , \wRegInBot_6_19[15] , \wRegInTop_7_54[17] , 
        \wRegOut_7_54[8] , \wRegInTop_7_77[26] , \ScanLink222[29] , 
        \ScanLink28[0] , \wRegInTop_5_14[23] , \wRegOut_6_9[27] , 
        \wRegInTop_6_19[12] , \wRegInTop_7_17[22] , \ScanLink115[1] , 
        \wRegInTop_7_62[12] , \wRegInTop_7_89[9] , \wRegInTop_7_34[13] , 
        \ScanLink201[18] , \ScanLink222[30] , \wRegInTop_7_41[23] , 
        \wRegInTop_7_46[0] , \wRegOut_7_98[2] , \wRegInBot_5_22[21] , 
        \ScanLink91[19] , \wRegOut_5_1[20] , \wRegInBot_5_14[24] , 
        \wRegInTop_5_22[26] , \ScanLink116[2] , \wRegInTop_7_45[3] , 
        \wRegInTop_5_28[8] , \wRegInTop_7_99[13] , \wRegOut_7_67[29] , 
        \wRegInTop_4_6[8] , \wRegInTop_4_14[1] , \wRegInBot_6_29[0] , 
        \wRegOut_7_31[31] , \wRegOut_7_6[24] , \wRegOut_7_12[19] , 
        \wRegOut_7_31[28] , \wRegOut_7_44[18] , \wRegOut_7_67[30] , 
        \wRegInTop_7_97[5] , \wRegOut_5_0[4] , \wRegInBot_5_8[24] , 
        \wRegOut_3_6[19] , \wRegInBot_4_7[14] , \wRegInTop_6_19[21] , 
        \wRegInBot_6_53[8] , \wRegInTop_7_62[21] , \ScanLink211[0] , 
        \wRegInTop_7_17[11] , \ScanLink52[8] , \wRegOut_6_9[14] , 
        \wRegInBot_6_19[26] , \wRegInTop_7_21[14] , \wRegInTop_7_22[4] , 
        \wRegInTop_7_34[20] , \wRegInTop_7_41[10] , \wRegOut_7_114[6] , 
        \ScanLink171[5] , \wRegInTop_7_54[24] , \ScanLink192[30] , 
        \wRegInTop_7_77[15] , \ScanLink192[29] , \wRegInBot_6_0[10] , 
        \wRegOut_6_7[6] , \ScanLink2[31] , \wRegInTop_2_1[25] , 
        \ScanLink9[24] , \wRegOut_5_1[13] , \wRegInBot_5_8[17] , 
        \wRegOut_6_4[5] , \wRegEnTop_7_4[0] , \wRegOut_7_109[9] , 
        \wRegInTop_7_123[9] , \wRegOut_7_6[17] , \wRegInTop_5_22[15] , 
        \wRegInTop_7_2[9] , \wRegOut_6_12[9] , \wRegOut_7_117[5] , 
        \wRegInTop_5_14[10] , \wRegInBot_5_14[17] , \ScanLink212[3] , 
        \wRegInTop_7_99[20] , \wRegInBot_5_22[12] , \wRegInTop_7_21[7] , 
        \ScanLink169[28] , \ScanLink172[6] , \ScanLink169[31] , 
        \wRegEnBot_6_27[0] , \wRegInTop_6_39[8] , \ScanLink184[6] , 
        \wRegOut_7_2[26] , \wRegOut_5_5[22] , \wRegInBot_5_10[26] , 
        \wRegInTop_5_26[24] , \wRegInTop_6_24[7] , \ScanLink156[0] , 
        \ScanLink199[9] , \wRegInTop_5_10[21] , \ScanLink118[29] , 
        \wRegOut_7_17[9] , \wRegInTop_7_88[25] , \ScanLink236[5] , 
        \wRegInTop_2_1[16] , \wRegOut_3_2[31] , \wRegOut_3_2[28] , 
        \wRegInBot_5_26[23] , \ScanLink68[2] , \ScanLink118[30] , 
        \wRegInTop_7_119[3] , \wRegInBot_4_3[25] , \wRegInTop_7_13[20] , 
        \ScanLink155[3] , \wRegInTop_7_66[10] , \wRegInTop_5_10[12] , 
        \wRegInBot_6_4[21] , \wRegInTop_6_27[4] , \wRegInTop_7_25[25] , 
        \wRegInTop_7_30[11] , \wRegInTop_7_45[21] , \wRegEnTop_7_48[0] , 
        \wRegInTop_7_50[15] , \ScanLink187[5] , \ScanLink196[18] , 
        \ScanLink235[6] , \wRegInTop_7_73[24] , \wRegOut_6_28[3] , 
        \ScanLink95[28] , \ScanLink228[9] , \ScanLink95[31] , 
        \wRegInTop_7_88[16] , \wRegInTop_6_40[3] , \ScanLink132[4] , 
        \wRegInTop_7_61[5] , \wRegInBot_3_0[13] , \ScanLink9[17] , 
        \ScanLink11[9] , \wRegOut_5_5[11] , \wRegInTop_5_26[17] , 
        \wRegInBot_5_26[10] , \wRegInBot_5_10[15] , \wRegInBot_6_10[9] , 
        \ScanLink252[1] , \wRegInTop_5_11[1] , \wRegOut_7_16[28] , 
        \wRegOut_6_18[18] , \wRegOut_7_16[31] , \wRegOut_7_40[30] , 
        \wRegOut_7_63[18] , \wRegOut_7_35[19] , \wRegOut_7_40[29] , 
        \wRegOut_7_2[15] , \wRegInTop_3_5[19] , \wRegInBot_4_3[16] , 
        \ScanLink38[31] , \ScanLink38[28] , \wRegInTop_5_12[2] , 
        \wRegInTop_6_1[18] , \wRegOut_5_15[30] , \wRegOut_5_15[29] , 
        \wRegOut_7_98[19] , \wRegInTop_7_118[19] , \wRegInBot_6_4[12] , 
        \wRegInTop_7_50[26] , \wRegInTop_6_43[0] , \wRegInTop_7_62[6] , 
        \ScanLink131[7] , \wRegInTop_7_25[16] , \wRegInTop_5_8[1] , 
        \wRegInTop_7_73[17] , \wRegInBot_5_9[7] , \wRegOut_6_51[8] , 
        \wRegInTop_7_66[23] , \ScanLink251[2] , \ScanLink253[28] , 
        \ScanLink205[30] , \ScanLink226[18] , \wRegInTop_7_13[13] , 
        \wRegInBot_4_15[30] , \ScanLink113[16] , \wRegInTop_7_5[17] , 
        \wRegInTop_7_30[22] , \wRegInTop_7_45[12] , \ScanLink253[31] , 
        \ScanLink205[29] , \ScanLink166[26] , \ScanLink130[27] , 
        \ScanLink145[17] , \ScanLink182[8] , \ScanLink150[23] , 
        \wRegInBot_4_15[29] , \wRegInBot_5_23[1] , \ScanLink73[3] , 
        \ScanLink125[13] , \ScanLink173[12] , \wRegInTop_7_102[2] , 
        \wRegInTop_5_2[13] , \wRegOut_6_13[14] , \ScanLink106[22] , 
        \wRegInTop_6_22[9] , \wRegOut_6_45[15] , \wRegOut_7_68[14] , 
        \wRegInBot_5_7[19] , \wRegOut_6_25[11] , \wRegOut_6_30[25] , 
        \wRegOut_6_50[21] , \wRegOut_7_9[19] , \wRegOut_6_30[1] , 
        \wRegOut_7_11[7] , \wRegOut_4_10[15] , \wRegOut_5_28[20] , 
        \wRegOut_6_33[2] , \wRegOut_7_86[21] , \wRegOut_7_93[15] , 
        \wRegInTop_7_113[15] , \wRegInTop_7_106[21] , \ScanLink10[15] , 
        \ScanLink33[24] , \wRegOut_7_12[4] , \ScanLink233[8] , 
        \wRegInTop_7_125[10] , \ScanLink46[14] , \wRegInBot_6_16[31] , 
        \wRegInBot_6_35[19] , \wRegInBot_6_40[29] , \wRegInBot_6_40[30] , 
        \wRegInBot_6_63[18] , \ScanLink26[10] , \ScanLink65[25] , 
        \ScanLink70[11] , \wRegInBot_6_16[28] , \ScanLink188[13] , 
        \ScanLink238[20] , \wRegOut_7_126[28] , \ScanLink70[0] , 
        \wRegOut_7_105[19] , \wRegOut_7_126[31] , \wRegInBot_5_20[2] , 
        \ScanLink53[20] , \wRegInTop_7_101[1] , \wRegOut_6_25[22] , 
        \ScanLink2[28] , \wRegOut_6_50[12] , \wRegInBot_3_0[20] , 
        \ScanLink10[26] , \ScanLink14[4] , \ScanLink17[7] , 
        \wRegInTop_5_2[20] , \wRegEnBot_5_9[0] , \wRegOut_6_13[27] , 
        \wRegInBot_6_16[7] , \wRegOut_6_54[5] , \wRegOut_7_68[27] , 
        \wRegOut_7_75[3] , \wRegOut_5_18[8] , \wRegOut_6_30[16] , 
        \ScanLink106[11] , \wRegOut_6_45[26] , \ScanLink125[20] , 
        \ScanLink129[5] , \ScanLink150[10] , \ScanLink113[25] , 
        \ScanLink173[21] , \wRegInTop_7_83[29] , \wRegInTop_7_5[24] , 
        \ScanLink249[0] , \ScanLink166[15] , \wRegInBot_4_8[30] , 
        \wRegInBot_4_8[29] , \ScanLink70[22] , \wRegEnTop_6_15[0] , 
        \wRegInTop_7_83[30] , \ScanLink130[14] , \ScanLink145[24] , 
        \ScanLink188[20] , \wRegOut_6_6[30] , \wRegInTop_6_58[1] , 
        \wRegInTop_7_79[7] , \ScanLink26[23] , \ScanLink53[13] , 
        \ScanLink46[27] , \wRegOut_6_6[29] , \wRegInTop_6_55[29] , 
        \ScanLink33[17] , \wRegInTop_7_78[31] , \ScanLink65[16] , 
        \wRegInTop_6_20[19] , \wRegInTop_6_55[30] , \ScanLink238[13] , 
        \wRegInTop_7_78[28] , \wRegOut_4_8[3] , \wRegOut_7_86[12] , 
        \wRegOut_3_3[11] , \wRegInTop_4_7[16] , \wRegOut_4_10[26] , 
        \wRegInTop_7_106[12] , \wRegOut_5_28[13] , \ScanLink137[9] , 
        \wRegInTop_7_64[8] , \wRegInTop_7_125[23] , \wRegInBot_6_15[4] , 
        \wRegOut_6_57[6] , \wRegOut_7_76[0] , \wRegOut_7_93[26] , 
        \wRegInTop_7_113[26] , \ScanLink197[21] , \ScanLink247[16] , 
        \ScanLink232[26] , \ScanLink39[22] , \ScanLink59[26] , 
        \wRegInTop_7_31[28] , \wRegInTop_7_44[18] , \ScanLink211[17] , 
        \wRegInTop_7_67[30] , \ScanLink204[23] , \wRegOut_6_41[2] , 
        \wRegOut_7_60[4] , \ScanLink241[8] , \ScanLink252[22] , 
        \ScanLink182[15] , \wRegInTop_7_67[29] , \ScanLink227[12] , 
        \wRegInBot_3_4[6] , \wRegOut_4_3[8] , \wRegInTop_7_12[19] , 
        \wRegInTop_7_31[31] , \wRegInTop_7_119[13] , \wRegInTop_3_5[0] , 
        \wRegInTop_6_0[12] , \wRegOut_7_99[13] , \wRegInTop_3_6[3] , 
        \wRegInBot_3_7[5] , \wRegInBot_5_4[2] , \wRegInTop_5_5[4] , 
        \wRegOut_5_10[0] , \wRegOut_5_22[26] , \wRegInBot_6_5[18] , 
        \wRegOut_5_14[23] , \wRegInTop_5_8[15] , \wRegOut_7_34[13] , 
        \wRegOut_7_41[23] , \wRegOut_6_19[12] , \wRegOut_7_17[22] , 
        \wRegInTop_5_6[7] , \wRegOut_7_62[12] , \wRegInBot_5_7[1] , 
        \wRegOut_5_13[3] , \wRegOut_7_21[27] , \wRegOut_7_77[26] , 
        \wRegInTop_6_50[9] , \wRegOut_7_54[17] , \wRegOut_0_0[30] , 
        \wRegInBot_0_0[7] , \wRegInTop_5_11[18] , \wRegOut_5_14[10] , 
        \wRegInBot_6_0[3] , \wRegInTop_6_1[5] , \ScanLink81[16] , 
        \ScanLink94[22] , \ScanLink119[10] , \ScanLink179[14] , 
        \wRegOut_7_63[7] , \wRegOut_6_42[1] , \ScanLink158[6] , 
        \wRegInTop_6_0[21] , \wRegOut_6_38[9] , \ScanLink238[3] , 
        \wRegInTop_7_119[20] , \ScanLink66[4] , \wRegOut_7_7[9] , 
        \wRegOut_7_99[20] , \wRegInBot_3_2[8] , \wRegOut_3_3[22] , 
        \wRegOut_5_22[15] , \ScanLink59[15] , \ScanLink145[9] , 
        \wRegInTop_7_117[5] , \ScanLink204[10] , \wRegInTop_7_16[8] , 
        \ScanLink182[26] , \ScanLink227[21] , \wRegInTop_3_4[20] , 
        \wRegOut_4_0[27] , \wRegInTop_4_7[25] , \wRegOut_6_25[6] , 
        \ScanLink252[11] , \ScanLink197[12] , \ScanLink211[24] , 
        \ScanLink232[15] , \ScanLink247[25] , \wRegInBot_4_14[3] , 
        \wRegOut_5_4[31] , \wRegOut_5_4[28] , \ScanLink39[11] , 
        \ScanLink179[27] , \ScanLink81[25] , \ScanLink189[3] , 
        \wRegInTop_5_8[26] , \wRegInBot_5_27[30] , \wRegInBot_5_27[29] , 
        \ScanLink78[8] , \wRegEnTop_7_94[0] , \wRegOut_6_26[5] , 
        \wRegInTop_7_109[9] , \wRegOut_7_123[9] , \ScanLink119[23] , 
        \ScanLink65[7] , \wRegInTop_6_2[6] , \wRegInTop_6_29[2] , 
        \ScanLink94[11] , \wRegOut_7_77[15] , \wRegOut_7_54[24] , 
        \wRegInBot_6_3[0] , \wRegOut_7_21[14] , \wRegOut_7_41[10] , 
        \wRegOut_7_34[20] , \wRegInTop_5_19[9] , \wRegOut_6_19[21] , 
        \wRegInTop_7_114[6] , \wRegInTop_6_55[4] , \wRegOut_7_17[11] , 
        \wRegOut_7_62[21] , \wRegInTop_7_74[2] , \ScanLink127[3] , 
        \wRegInTop_7_124[29] , \wRegOut_7_87[18] , \wRegInTop_7_107[18] , 
        \wRegInTop_7_124[30] , \ScanLink247[6] , \ScanLink19[1] , 
        \ScanLink27[29] , \ScanLink52[19] , \wRegOut_5_29[19] , 
        \wRegInTop_6_41[17] , \wRegOut_6_7[23] , \ScanLink71[31] , 
        \wRegInBot_6_21[14] , \wRegInTop_6_34[27] , \wRegInBot_6_54[24] , 
        \wRegOut_7_104[20] , \wRegInTop_6_62[26] , \wRegOut_4_5[6] , 
        \wRegOut_4_6[5] , \wRegInBot_4_9[23] , \ScanLink27[30] , 
        \ScanLink71[28] , \wRegInTop_7_19[26] , \wRegInTop_6_17[16] , 
        \wRegOut_7_127[11] , \wRegEnTop_5_6[0] , \wRegInBot_6_17[11] , 
        \wRegInBot_6_18[1] , \wRegInBot_6_62[21] , \ScanLink239[19] , 
        \wRegInTop_7_79[22] , \wRegInTop_6_21[13] , \wRegInBot_6_34[20] , 
        \wRegInBot_6_41[10] , \wRegInTop_6_54[23] , \wRegOut_7_111[14] , 
        \wRegInTop_7_97[17] , \wRegOut_0_0[29] , \wRegInBot_4_14[10] , 
        \wRegEnBot_6_55[0] , \wRegOut_1_1[3] , \ScanLink3[22] , 
        \wRegInTop_4_14[17] , \wRegOut_7_78[6] , \wRegInTop_7_82[23] , 
        \wRegInTop_5_0[9] , \wRegOut_6_59[0] , \wRegInBot_5_6[20] , 
        \wRegOut_6_24[31] , \wRegInBot_6_17[22] , \wRegOut_6_24[28] , 
        \wRegInTop_6_56[7] , \ScanLink124[0] , \wRegInTop_7_77[1] , 
        \wRegOut_6_51[18] , \wRegInBot_6_62[12] , \wRegOut_7_8[20] , 
        \wRegOut_7_65[9] , \ScanLink244[5] , \wRegInTop_7_79[11] , 
        \wRegInTop_6_21[20] , \wRegInBot_6_41[23] , \ScanLink191[1] , 
        \wRegOut_7_111[27] , \wRegInBot_6_34[13] , \ScanLink3[11] , 
        \wRegInBot_3_1[19] , \wRegInTop_3_4[13] , \wRegInBot_4_9[10] , 
        \wRegInBot_5_30[8] , \wRegOut_6_7[10] , \wRegInTop_6_34[14] , 
        \wRegInTop_6_54[10] , \wRegOut_7_1[7] , \wRegOut_7_104[13] , 
        \wRegInBot_6_54[17] , \wRegInTop_6_17[25] , \wRegInBot_6_21[27] , 
        \wRegInTop_6_41[24] , \wRegInTop_6_62[15] , \wRegOut_7_127[22] , 
        \wRegInTop_7_19[15] , \ScanLink189[19] , \wRegInTop_6_31[0] , 
        \ScanLink143[7] , \wRegInTop_7_10[6] , \ScanLink223[2] , 
        \wRegOut_7_126[4] , \wRegOut_4_0[14] , \wRegInTop_5_3[19] , 
        \wRegOut_6_23[8] , \wRegInTop_6_32[3] , \ScanLink140[4] , 
        \wRegInTop_7_13[5] , \ScanLink220[1] , \wRegEnTop_7_105[0] , 
        \wRegInBot_5_6[13] , \wRegInBot_6_62[9] , \wRegInTop_6_4[8] , 
        \wRegOut_7_8[13] , \ScanLink192[2] , \wRegOut_7_125[7] , 
        \wRegEnBot_0_0[0] , \wRegInTop_4_14[24] , \wRegInTop_7_82[10] , 
        \wRegInBot_4_14[23] , \ScanLink151[30] , \ScanLink172[18] , 
        \ScanLink107[28] , \ScanLink151[29] , \wRegInTop_7_97[24] , 
        \wRegOut_1_0[24] , \wRegOut_1_0[17] , \wRegInBot_2_1[14] , 
        \ScanLink5[0] , \ScanLink6[3] , \ScanLink7[20] , \wRegInBot_5_2[22] , 
        \wRegInTop_5_7[31] , \wRegInTop_5_7[28] , \ScanLink63[9] , 
        \wRegOut_7_2[4] , \ScanLink95[9] , \ScanLink107[31] , 
        \ScanLink124[19] , \wRegInTop_7_112[8] , \wRegOut_7_101[1] , 
        \ScanLink204[7] , \wRegInTop_4_10[15] , \wRegInBot_5_28[27] , 
        \wRegInTop_6_16[5] , \ScanLink164[2] , \wRegInTop_7_37[3] , 
        \ScanLink88[6] , \wRegInTop_7_9[2] , \wRegOut_6_19[2] , 
        \wRegOut_7_38[4] , \wRegInTop_7_86[21] , \ScanLink219[8] , 
        \wRegInBot_4_10[12] , \ScanLink103[19] , \ScanLink120[31] , 
        \ScanLink176[29] , \wRegInTop_7_93[15] , \wRegInTop_5_28[20] , 
        \ScanLink120[28] , \ScanLink155[18] , \ScanLink176[30] , 
        \wRegInBot_6_13[13] , \ScanLink7[13] , \wRegInTop_3_0[22] , 
        \wRegOut_6_3[21] , \wRegInTop_6_25[11] , \wRegInBot_6_30[22] , 
        \wRegInBot_6_58[3] , \wRegInBot_6_45[12] , \wRegInTop_6_50[21] , 
        \wRegOut_7_115[16] , \wRegInBot_6_25[16] , \wRegInTop_6_45[15] , 
        \wRegInTop_6_30[25] , \wRegInBot_6_50[26] , \wRegInTop_6_13[14] , 
        \wRegOut_7_100[22] , \wRegOut_7_26[8] , \wRegInTop_7_68[14] , 
        \ScanLink207[4] , \wRegOut_7_123[13] , \wRegInBot_3_5[31] , 
        \ScanLink59[3] , \wRegInTop_6_15[6] , \wRegInTop_7_34[0] , 
        \wRegOut_7_102[2] , \ScanLink167[1] , \wRegInBot_3_5[28] , 
        \wRegOut_4_4[25] , \wRegInTop_4_10[26] , \wRegInBot_4_10[21] , 
        \wRegOut_7_93[9] , \wRegInTop_5_23[3] , \wRegInTop_5_28[13] , 
        \wRegInTop_7_93[26] , \wRegInBot_5_28[14] , \wRegInTop_7_81[1] , 
        \wRegInTop_7_86[12] , \wRegOut_6_60[9] , \wRegInTop_3_0[11] , 
        \wRegOut_4_4[16] , \wRegInBot_5_2[11] , \wRegOut_6_55[30] , 
        \wRegOut_7_78[28] , \wRegOut_6_20[19] , \wRegOut_6_55[29] , 
        \wRegOut_7_78[31] , \ScanLink100[6] , \wRegInTop_7_53[7] , 
        \wRegOut_7_83[30] , \wRegOut_7_83[29] , \wRegInTop_7_103[30] , 
        \wRegInTop_7_120[18] , \wRegInBot_6_21[8] , \wRegInTop_7_103[29] , 
        \ScanLink103[5] , \wRegInTop_7_50[4] , \ScanLink20[8] , 
        \ScanLink23[18] , \wRegInTop_6_30[16] , \wRegInTop_4_8[18] , 
        \wRegInTop_5_20[0] , \ScanLink56[31] , \ScanLink56[28] , 
        \wRegOut_6_3[12] , \wRegInBot_6_50[15] , \wRegOut_7_100[11] , 
        \wRegInBot_6_25[25] , \wRegInTop_6_45[26] , \ScanLink75[19] , 
        \wRegInTop_6_13[27] , \wRegInTop_7_68[27] , \wRegOut_7_123[20] , 
        \wRegInBot_6_13[20] , \ScanLink248[18] , \wRegInBot_6_45[21] , 
        \wRegOut_7_115[25] , \ScanLink85[14] , \wRegInTop_6_25[22] , 
        \wRegInTop_7_82[2] , \wRegInBot_6_30[11] , \wRegInTop_6_50[12] , 
        \ScanLink202[9] , \wRegOut_7_23[5] , \wRegOut_5_0[19] , 
        \ScanLink41[1] , \wRegInBot_5_23[18] , \wRegOut_6_9[0] , 
        \ScanLink93[7] , \wRegInBot_6_40[1] , \ScanLink108[26] , 
        \ScanLink90[20] , \ScanLink168[22] , \wRegEnTop_7_62[0] , 
        \wRegOut_7_73[24] , \ScanLink42[2] , \wRegInBot_5_11[3] , 
        \wRegOut_7_25[25] , \wRegOut_7_50[15] , \wRegOut_7_13[20] , 
        \wRegOut_7_30[11] , \wRegOut_7_45[21] , \wRegOut_7_66[10] , 
        \wRegOut_7_119[3] , \wRegInBot_2_1[27] , \wRegOut_3_7[13] , 
        \ScanLink28[14] , \wRegOut_5_10[21] , \wRegInBot_5_12[0] , 
        \wRegOut_7_88[25] , \wRegInTop_7_108[25] , \wRegOut_5_26[24] , 
        \wRegInTop_6_4[10] , \ScanLink90[4] , \wRegOut_7_20[6] , 
        \ScanLink200[21] , \ScanLink186[17] , \ScanLink223[10] , 
        \wRegInTop_4_3[14] , \wRegInTop_6_13[8] , \wRegInBot_6_43[2] , 
        \ScanLink193[23] , \ScanLink243[14] , \ScanLink236[24] , 
        \ScanLink25[5] , \ScanLink48[10] , \wRegOut_7_45[12] , 
        \ScanLink215[15] , \wRegInTop_5_15[30] , \wRegOut_7_13[13] , 
        \wRegOut_7_30[22] , \wRegOut_7_66[23] , \wRegOut_7_95[7] , 
        \wRegOut_7_25[16] , \wRegInTop_7_48[6] , \wRegOut_7_50[26] , 
        \wRegOut_7_73[17] , \wRegInTop_5_15[29] , \ScanLink90[13] , 
        \wRegOut_7_47[1] , \wRegOut_7_88[8] , \wRegInBot_6_24[5] , 
        \ScanLink108[15] , \ScanLink168[11] , \wRegInTop_7_98[19] , 
        \wRegOut_3_7[20] , \wRegInTop_4_3[27] , \wRegInBot_4_9[8] , 
        \ScanLink85[27] , \ScanLink106[8] , \wRegInTop_7_55[9] , 
        \ScanLink48[23] , \wRegInBot_6_27[6] , \wRegOut_7_44[2] , 
        \ScanLink193[10] , \ScanLink236[17] , \ScanLink243[27] , 
        \wRegOut_5_29[9] , \ScanLink215[26] , \ScanLink28[27] , 
        \wRegInTop_7_16[31] , \wRegInTop_7_35[19] , \ScanLink200[12] , 
        \wRegInTop_7_99[3] , \wRegInTop_7_40[29] , \wRegInTop_7_16[28] , 
        \ScanLink186[24] , \ScanLink223[23] , \ScanLink26[6] , 
        \wRegInTop_6_4[23] , \wRegInTop_6_18[18] , \wRegInTop_7_40[30] , 
        \wRegInTop_7_63[18] , \wRegOut_7_96[4] , \wRegOut_4_15[0] , 
        \wRegOut_5_26[17] , \ScanLink118[4] , \ScanLink2[25] , 
        \wRegInTop_2_1[31] , \wRegInTop_2_1[28] , \wRegOut_3_2[25] , 
        \wRegOut_3_2[16] , \wRegInTop_4_6[11] , \wRegOut_5_10[12] , 
        \wRegInBot_6_1[29] , \wRegInBot_6_1[30] , \ScanLink196[26] , 
        \wRegOut_7_88[16] , \ScanLink233[21] , \wRegInTop_7_108[16] , 
        \ScanLink246[11] , \ScanLink38[25] , \ScanLink58[21] , 
        \ScanLink205[24] , \ScanLink210[10] , \wRegOut_6_51[5] , 
        \wRegOut_7_70[3] , \ScanLink253[25] , \ScanLink183[12] , 
        \ScanLink226[15] , \ScanLink11[4] , \ScanLink12[7] , 
        \wRegOut_5_23[21] , \wRegInTop_6_1[15] , \wRegInBot_6_13[7] , 
        \wRegOut_7_98[14] , \wRegInTop_7_118[14] , \wRegInTop_5_9[12] , 
        \wRegOut_5_15[24] , \wRegEnTop_6_10[0] , \wRegOut_6_18[15] , 
        \wRegOut_7_16[25] , \wRegOut_7_35[14] , \wRegOut_7_40[24] , 
        \wRegOut_7_63[15] , \wRegOut_7_76[21] , \wRegInBot_4_3[31] , 
        \wRegInBot_5_10[18] , \ScanLink80[11] , \ScanLink95[25] , 
        \wRegOut_7_2[18] , \wRegOut_7_20[20] , \ScanLink132[9] , 
        \wRegOut_7_55[10] , \wRegInTop_7_61[8] , \ScanLink118[17] , 
        \ScanLink178[13] , \wRegOut_6_52[6] , \wRegOut_7_73[0] , 
        \wRegOut_5_15[17] , \wRegInBot_6_10[4] , \ScanLink148[1] , 
        \ScanLink187[8] , \wRegOut_5_23[12] , \wRegInTop_6_1[26] , 
        \ScanLink228[4] , \ScanLink76[3] , \wRegOut_7_98[27] , 
        \wRegInTop_7_118[27] , \wRegInBot_5_26[1] , \ScanLink58[12] , 
        \ScanLink205[17] , \wRegInTop_7_107[2] , \wRegInTop_6_27[9] , 
        \ScanLink183[21] , \ScanLink226[26] , \wRegInBot_4_3[28] , 
        \wRegInTop_4_6[22] , \wRegOut_6_35[1] , \wRegInTop_7_25[31] , 
        \ScanLink253[16] , \wRegOut_7_14[7] , \ScanLink233[12] , 
        \wRegInTop_7_25[28] , \ScanLink196[15] , \wRegInTop_7_73[29] , 
        \ScanLink246[22] , \wRegInTop_7_50[18] , \ScanLink210[23] , 
        \ScanLink38[16] , \wRegInTop_5_26[30] , \ScanLink178[20] , 
        \wRegInTop_7_73[30] , \wRegInTop_5_26[29] , \ScanLink80[22] , 
        \ScanLink199[4] , \wRegOut_6_36[2] , \wRegOut_7_9[2] , 
        \wRegInTop_7_88[31] , \ScanLink9[30] , \ScanLink9[29] , 
        \ScanLink95[16] , \ScanLink118[24] , \wRegOut_7_17[4] , 
        \wRegInTop_7_88[28] , \ScanLink236[8] , \wRegOut_7_76[12] , 
        \wRegInTop_6_39[5] , \wRegInTop_7_18[3] , \wRegOut_7_55[23] , 
        \wRegOut_7_20[13] , \wRegInTop_3_5[27] , \wRegOut_4_1[20] , 
        \wRegInTop_5_9[21] , \ScanLink75[0] , \wRegOut_7_40[17] , 
        \wRegInBot_5_25[2] , \wRegOut_6_18[26] , \wRegOut_7_35[27] , 
        \wRegInTop_7_104[1] , \wRegInTop_6_45[3] , \wRegOut_7_16[16] , 
        \wRegOut_7_63[26] , \wRegInTop_7_64[5] , \ScanLink137[4] , 
        \wRegInBot_6_15[9] , \ScanLink14[9] , \wRegInBot_4_8[24] , 
        \wRegInTop_5_14[1] , \wRegOut_6_6[24] , \wRegInBot_6_20[13] , 
        \wRegInTop_6_40[10] , \wRegInTop_6_35[20] , \wRegInBot_6_55[23] , 
        \wRegInTop_6_63[21] , \wRegOut_7_105[27] , \wRegInTop_6_16[11] , 
        \wRegInTop_7_18[21] , \wRegInBot_6_16[16] , \wRegOut_7_126[16] , 
        \wRegInBot_6_35[27] , \wRegInBot_6_63[26] , \wRegInTop_7_78[25] , 
        \wRegInTop_6_55[24] , \wRegInTop_4_15[10] , \wRegInBot_4_15[17] , 
        \wRegInTop_5_17[2] , \wRegInTop_6_20[14] , \wRegInBot_6_40[17] , 
        \wRegOut_7_110[13] , \wRegInTop_7_96[10] , \wRegOut_6_49[7] , 
        \ScanLink113[31] , \ScanLink129[8] , \ScanLink113[28] , 
        \ScanLink130[19] , \wRegInTop_7_5[30] , \ScanLink145[29] , 
        \wRegOut_7_68[1] , \wRegInTop_7_83[24] , \wRegInBot_5_7[27] , 
        \wRegInTop_7_5[29] , \ScanLink145[30] , \ScanLink166[18] , 
        \ScanLink2[16] , \ScanLink10[18] , \wRegOut_5_18[5] , 
        \wRegInTop_6_46[0] , \ScanLink134[7] , \wRegInTop_7_67[6] , 
        \wRegOut_7_9[27] , \wRegOut_6_54[8] , \wRegInTop_7_78[16] , 
        \ScanLink254[2] , \wRegInTop_3_5[14] , \wRegInBot_4_8[17] , 
        \ScanLink33[30] , \ScanLink33[29] , \ScanLink65[28] , 
        \wRegInBot_6_16[25] , \wRegInBot_6_63[15] , \wRegEnBot_6_22[0] , 
        \wRegInBot_6_40[24] , \wRegOut_7_110[20] , \ScanLink46[19] , 
        \wRegInTop_6_20[27] , \ScanLink181[6] , \ScanLink65[31] , 
        \wRegOut_6_6[17] , \wRegInTop_6_35[13] , \wRegInBot_6_35[14] , 
        \wRegInTop_6_55[17] , \wRegInBot_6_55[10] , \wRegOut_7_105[14] , 
        \wRegInTop_6_16[22] , \wRegInBot_6_20[20] , \wRegInTop_6_40[23] , 
        \wRegInTop_6_63[12] , \wRegOut_7_126[25] , \wRegInTop_7_18[12] , 
        \wRegInTop_6_21[7] , \ScanLink153[0] , \wRegOut_7_93[18] , 
        \wRegInTop_7_113[18] , \wRegOut_4_1[13] , \wRegOut_7_12[9] , 
        \wRegOut_4_10[18] , \ScanLink233[5] , \wRegInBot_6_8[6] , 
        \wRegInTop_6_9[0] , \wRegInTop_6_22[4] , \wRegOut_6_45[18] , 
        \ScanLink150[3] , \wRegOut_6_30[28] , \wRegOut_6_13[19] , 
        \wRegOut_6_30[31] , \wRegOut_7_68[19] , \ScanLink230[6] , 
        \wRegInBot_2_1[9] , \wRegOut_2_2[31] , \wRegOut_2_2[28] , 
        \wRegInTop_4_15[23] , \wRegInBot_5_7[14] , \wRegOut_7_9[14] , 
        \ScanLink182[5] , \wRegInTop_7_83[17] , \wRegInBot_4_15[24] , 
        \wRegOut_6_17[31] , \wRegOut_6_34[19] , \wRegInTop_7_96[23] , 
        \wRegEnTop_6_48[0] , \wRegOut_6_17[28] , \wRegOut_6_41[29] , 
        \wRegOut_7_111[6] , \wRegOut_6_41[30] , \wRegInBot_6_56[8] , 
        \wRegOut_6_62[18] , \ScanLink214[0] , \wRegOut_7_19[18] , 
        \ScanLink6[27] , \wRegInBot_5_3[25] , \wRegInTop_7_27[4] , 
        \ScanLink174[5] , \ScanLink8[8] , \ScanLink14[30] , \ScanLink14[29] , 
        \wRegInTop_4_11[12] , \ScanLink57[8] , \wRegInBot_5_29[20] , 
        \ScanLink98[1] , \wRegOut_6_2[6] , \wRegOut_7_28[3] , 
        \wRegInTop_7_87[26] , \wRegInTop_7_126[9] , \wRegInBot_4_11[15] , 
        \wRegInTop_7_92[12] , \ScanLink42[31] , \wRegInTop_5_29[27] , 
        \ScanLink61[19] , \wRegEnTop_7_1[0] , \wRegInBot_6_12[14] , 
        \ScanLink37[18] , \ScanLink42[28] , \wRegInBot_6_31[25] , 
        \wRegInBot_6_48[4] , \wRegInTop_6_51[26] , \wRegOut_7_114[11] , 
        \wRegOut_6_1[5] , \wRegInTop_6_24[16] , \wRegInBot_6_44[15] , 
        \wRegOut_6_2[26] , \wRegInBot_6_24[11] , \wRegInTop_6_44[12] , 
        \wRegInTop_7_39[8] , \ScanLink229[31] , \wRegInTop_6_31[22] , 
        \wRegInTop_7_7[9] , \wRegInTop_6_12[13] , \wRegInBot_6_51[21] , 
        \wRegOut_7_101[25] , \ScanLink229[28] , \wRegOut_6_17[9] , 
        \wRegInTop_7_69[13] , \wRegOut_7_122[14] , \ScanLink217[3] , 
        \wRegInTop_7_117[29] , \wRegInTop_3_1[25] , \wRegOut_7_97[29] , 
        \wRegOut_3_6[3] , \wRegOut_4_5[22] , \wRegOut_4_14[30] , 
        \ScanLink49[4] , \wRegInBot_5_19[6] , \wRegOut_7_97[30] , 
        \wRegOut_7_112[5] , \wRegInTop_7_117[30] , \wRegInTop_7_24[7] , 
        \ScanLink177[6] , \wRegOut_4_14[29] , \wRegInBot_4_11[26] , 
        \wRegInTop_4_12[2] , \wRegInTop_5_29[14] , \wRegInTop_7_92[21] , 
        \wRegInBot_5_29[13] , \ScanLink134[28] , \ScanLink141[18] , 
        \ScanLink162[30] , \wRegInTop_7_91[6] , \wRegInTop_7_1[18] , 
        \wRegOut_5_6[7] , \ScanLink162[29] , \wRegInTop_7_87[15] , 
        \ScanLink6[14] , \wRegInTop_4_11[21] , \ScanLink134[31] , 
        \ScanLink117[19] , \wRegOut_7_51[8] , \wRegInTop_3_1[16] , 
        \wRegOut_4_5[11] , \wRegInBot_5_3[16] , \ScanLink110[1] , 
        \wRegInTop_6_62[6] , \wRegInTop_7_43[0] , \ScanLink113[2] , 
        \wRegInTop_6_61[5] , \wRegInTop_7_40[3] , \wRegOut_6_2[15] , 
        \wRegInTop_6_31[11] , \wRegOut_7_101[16] , \wRegInBot_6_24[22] , 
        \wRegInTop_6_44[21] , \wRegInBot_6_51[12] , \wRegOut_0_0[17] , 
        \ScanLink0[0] , \wRegOut_1_0[30] , \wRegInBot_1_0[5] , 
        \wRegOut_1_1[10] , \wRegInTop_1_1[3] , \wRegInBot_2_0[13] , 
        \wRegOut_3_5[0] , \wRegInTop_4_3[8] , \wRegInTop_6_12[20] , 
        \wRegInTop_7_69[20] , \wRegOut_7_122[27] , \wRegInTop_4_11[1] , 
        \wRegInTop_5_30[7] , \wRegOut_5_5[4] , \wRegInBot_6_12[27] , 
        \ScanLink199[28] , \ScanLink84[13] , \wRegInTop_6_24[25] , 
        \wRegInBot_6_44[26] , \wRegInTop_7_92[5] , \wRegOut_7_114[22] , 
        \wRegInBot_6_31[16] , \wRegInTop_6_51[15] , \ScanLink199[31] , 
        \wRegOut_7_33[2] , \ScanLink51[6] , \wRegInTop_5_22[18] , 
        \wRegOut_6_12[4] , \ScanLink83[0] , \ScanLink109[21] , 
        \wRegInBot_6_50[6] , \ScanLink91[27] , \wRegOut_7_117[8] , 
        \ScanLink169[25] , \wRegOut_7_72[23] , \wRegOut_6_4[8] , 
        \wRegOut_7_24[22] , \wRegOut_7_51[12] , \wRegInTop_7_120[7] , 
        \wRegInTop_7_2[4] , \wRegOut_7_31[16] , \wRegOut_7_12[27] , 
        \wRegOut_7_44[26] , \wRegOut_7_67[17] , \ScanLink52[5] , 
        \wRegOut_7_109[4] , \wRegInTop_7_123[4] , \wRegOut_1_1[23] , 
        \wRegInBot_2_0[20] , \wRegOut_3_6[14] , \wRegInBot_4_7[19] , 
        \ScanLink29[13] , \wRegOut_5_11[26] , \wRegOut_7_89[22] , 
        \wRegInTop_7_109[22] , \wRegOut_5_27[23] , \wRegInTop_6_5[17] , 
        \ScanLink80[3] , \wRegInTop_7_1[7] , \wRegOut_6_9[19] , 
        \wRegOut_6_11[7] , \wRegOut_7_30[1] , \ScanLink201[26] , 
        \ScanLink187[10] , \ScanLink222[17] , \wRegInTop_4_2[13] , 
        \wRegInBot_6_53[5] , \wRegInTop_7_22[9] , \wRegInTop_7_54[30] , 
        \wRegInTop_7_77[18] , \ScanLink192[24] , \ScanLink237[23] , 
        \ScanLink242[13] , \wRegInTop_4_6[5] , \wRegInBot_4_7[3] , 
        \ScanLink35[2] , \ScanLink49[17] , \wRegInTop_7_21[19] , 
        \ScanLink171[8] , \wRegInTop_7_54[29] , \wRegOut_5_27[2] , 
        \ScanLink214[12] , \wRegOut_7_44[15] , \wRegOut_7_31[25] , 
        \wRegOut_7_67[24] , \wRegOut_7_85[0] , \wRegOut_5_0[9] , 
        \wRegInBot_5_8[29] , \wRegOut_7_12[14] , \wRegOut_7_72[10] , 
        \wRegInBot_5_8[30] , \wRegOut_7_6[30] , \wRegOut_7_51[21] , 
        \wRegInTop_7_58[1] , \wRegInTop_7_97[8] , \wRegInBot_5_14[29] , 
        \wRegInTop_5_28[5] , \ScanLink91[14] , \wRegOut_7_6[29] , 
        \wRegOut_7_24[11] , \wRegOut_7_57[6] , \wRegInBot_6_34[2] , 
        \ScanLink169[16] , \ScanLink109[12] , \wRegOut_3_6[27] , 
        \wRegInTop_4_2[20] , \wRegInBot_5_14[30] , \ScanLink84[20] , 
        \ScanLink49[24] , \wRegInBot_6_19[18] , \wRegInBot_6_37[1] , 
        \wRegOut_7_54[5] , \ScanLink192[17] , \ScanLink237[10] , 
        \ScanLink242[20] , \ScanLink214[21] , \ScanLink29[20] , 
        \ScanLink201[15] , \wRegInTop_7_89[4] , \ScanLink187[23] , 
        \ScanLink222[24] , \wRegInBot_4_4[0] , \wRegInTop_4_5[6] , 
        \wRegInTop_6_5[24] , \wRegOut_7_86[3] , \ScanLink36[1] , 
        \wRegOut_5_24[1] , \wRegEnTop_7_15[0] , \wRegOut_5_27[10] , 
        \ScanLink108[3] , \wRegOut_2_3[22] , \wRegOut_2_3[11] , 
        \wRegInBot_3_5[16] , \ScanLink15[10] , \ScanLink20[5] , 
        \wRegOut_5_11[15] , \ScanLink75[14] , \wRegOut_7_89[11] , 
        \wRegOut_7_90[7] , \wRegInTop_7_109[11] , \ScanLink228[11] , 
        \wRegInBot_6_25[31] , \ScanLink23[15] , \wRegInBot_6_50[18] , 
        \wRegInTop_4_8[15] , \wRegOut_4_13[3] , \ScanLink56[25] , 
        \wRegInBot_6_25[28] , \ScanLink36[21] , \ScanLink43[11] , 
        \wRegOut_7_115[28] , \wRegOut_7_115[31] , \wRegOut_4_15[10] , 
        \ScanLink60[20] , \ScanLink248[15] , \wRegOut_6_63[7] , 
        \ScanLink198[22] , \wRegOut_7_83[24] , \wRegInTop_7_103[24] , 
        \wRegOut_5_8[1] , \wRegInBot_6_21[5] , \wRegOut_7_42[1] , 
        \ScanLink103[8] , \wRegInTop_7_120[15] , \wRegInTop_7_50[9] , 
        \wRegOut_7_96[10] , \wRegInTop_7_116[10] , \wRegOut_6_20[14] , 
        \wRegOut_6_55[24] , \wRegOut_6_60[4] , \wRegOut_7_41[2] , 
        \wRegOut_7_78[25] , \wRegInBot_3_5[25] , \wRegOut_4_4[28] , 
        \ScanLink23[6] , \wRegOut_4_10[0] , \wRegInTop_5_7[16] , 
        \wRegOut_6_16[11] , \wRegInBot_6_22[6] , \wRegOut_6_63[21] , 
        \wRegOut_7_18[21] , \wRegOut_6_40[10] , \wRegOut_5_31[6] , 
        \wRegOut_6_35[20] , \ScanLink155[26] , \wRegInBot_5_28[19] , 
        \ScanLink103[27] , \ScanLink120[16] , \ScanLink176[17] , 
        \wRegOut_7_93[4] , \ScanLink116[13] , \wRegInTop_7_0[12] , 
        \ScanLink163[23] , \ScanLink140[12] , \ScanLink96[7] , 
        \ScanLink135[22] , \wRegInBot_6_45[1] , \wRegOut_7_26[5] , 
        \ScanLink207[9] , \wRegOut_7_96[23] , \wRegInTop_7_116[23] , 
        \wRegOut_7_83[17] , \ScanLink15[23] , \wRegOut_4_4[31] , 
        \wRegOut_4_15[23] , \wRegInTop_7_103[17] , \wRegInTop_4_8[26] , 
        \ScanLink43[22] , \wRegInTop_7_120[26] , \ScanLink44[1] , 
        \wRegEnTop_7_67[0] , \ScanLink36[12] , \wRegInBot_5_14[3] , 
        \ScanLink60[13] , \ScanLink198[11] , \ScanLink23[26] , 
        \ScanLink56[16] , \ScanLink75[27] , \ScanLink228[22] , 
        \ScanLink248[26] , \wRegInTop_6_13[19] , \wRegInTop_6_30[31] , 
        \wRegInTop_6_45[18] , \wRegInTop_7_29[2] , \wRegInTop_7_68[19] , 
        \wRegInTop_6_30[28] , \wRegInTop_4_10[18] , \wRegInTop_5_7[25] , 
        \ScanLink47[2] , \ScanLink116[20] , \wRegOut_7_38[9] , 
        \wRegInTop_7_0[21] , \ScanLink219[5] , \ScanLink163[10] , 
        \wRegInBot_5_17[0] , \ScanLink135[11] , \wRegOut_6_16[22] , 
        \ScanLink103[14] , \ScanLink120[25] , \ScanLink140[21] , 
        \ScanLink179[0] , \ScanLink155[15] , \ScanLink176[24] , 
        \wRegInTop_7_93[18] , \ScanLink95[4] , \wRegOut_6_35[13] , 
        \wRegInBot_6_46[2] , \wRegOut_7_25[6] , \wRegOut_6_63[12] , 
        \wRegOut_7_18[12] , \wRegInTop_6_16[8] , \wRegOut_6_40[23] , 
        \wRegOut_6_20[27] , \wRegOut_6_55[17] , \wRegOut_7_78[16] , 
        \wRegInTop_5_26[3] , \wRegOut_7_59[0] , \wRegOut_7_96[9] , 
        \wRegOut_1_0[29] , \ScanLink118[9] , \wRegInTop_7_84[1] , 
        \ScanLink3[3] , \wRegInTop_4_3[19] , \wRegInBot_4_6[20] , 
        \wRegInTop_4_8[3] , \wRegInBot_4_9[5] , \wRegOut_5_29[4] , 
        \wRegInBot_6_1[24] , \wRegInTop_7_20[20] , \wRegInTop_7_55[10] , 
        \wRegInBot_6_18[12] , \wRegInTop_7_76[21] , \ScanLink186[29] , 
        \wRegInBot_4_6[13] , \ScanLink25[8] , \wRegOut_5_0[27] , 
        \ScanLink38[7] , \wRegInTop_5_15[24] , \wRegOut_6_8[20] , 
        \wRegInTop_6_18[15] , \wRegInTop_7_16[25] , \ScanLink105[6] , 
        \wRegInTop_7_63[15] , \wRegInTop_7_35[14] , \wRegInTop_7_56[7] , 
        \ScanLink186[30] , \wRegInTop_7_40[24] , \wRegOut_7_88[5] , 
        \wRegInBot_5_23[26] , \wRegInBot_6_24[8] , \wRegInBot_5_15[23] , 
        \wRegInTop_5_23[21] , \ScanLink106[5] , \wRegInTop_7_55[4] , 
        \ScanLink108[18] , \wRegInTop_7_98[14] , \wRegInBot_6_39[7] , 
        \wRegInBot_5_9[23] , \wRegInTop_5_25[0] , \wRegOut_7_7[23] , 
        \wRegInTop_7_87[2] , \wRegInTop_6_18[26] , \wRegInTop_7_16[16] , 
        \wRegInTop_7_63[26] , \ScanLink201[7] , \ScanLink28[19] , 
        \wRegOut_6_8[13] , \ScanLink90[9] , \wRegInTop_7_40[17] , 
        \wRegInTop_7_35[27] , \wRegInTop_7_55[23] , \wRegOut_7_104[1] , 
        \wRegInTop_6_13[5] , \wRegInTop_7_32[3] , \wRegInBot_6_18[21] , 
        \wRegInTop_7_20[13] , \ScanLink161[2] , \wRegInTop_7_76[12] , 
        \ScanLink215[18] , \ScanLink236[30] , \ScanLink243[19] , 
        \wRegOut_7_88[28] , \ScanLink236[29] , \wRegInTop_7_108[28] , 
        \wRegOut_5_26[30] , \wRegOut_5_26[29] , \wRegInBot_6_1[17] , 
        \wRegOut_7_88[31] , \wRegInTop_7_108[31] , \wRegOut_7_7[10] , 
        \wRegOut_7_25[28] , \wRegOut_7_25[31] , \wRegOut_7_50[18] , 
        \wRegOut_7_73[30] , \wRegOut_2_0[2] , \wRegInTop_2_0[22] , 
        \wRegInBot_2_1[19] , \wRegInBot_5_9[10] , \wRegOut_7_73[29] , 
        \wRegInTop_5_23[12] , \wRegOut_7_107[2] , \ScanLink8[23] , 
        \wRegOut_5_0[14] , \wRegInTop_5_15[17] , \wRegInBot_5_15[10] , 
        \ScanLink85[19] , \wRegOut_7_23[8] , \ScanLink202[4] , 
        \wRegInTop_7_98[27] , \wRegInBot_5_23[15] , \wRegInTop_6_10[6] , 
        \wRegInTop_7_31[0] , \ScanLink162[1] , \wRegOut_7_3[21] , 
        \wRegOut_7_21[19] , \wRegOut_7_54[29] , \ScanLink194[1] , 
        \wRegOut_7_54[30] , \wRegOut_7_77[18] , \wRegOut_5_4[25] , 
        \wRegInBot_5_11[21] , \wRegInTop_5_27[23] , \ScanLink81[31] , 
        \wRegInTop_6_34[0] , \wRegOut_7_4[7] , \wRegInTop_7_15[6] , 
        \ScanLink146[7] , \ScanLink81[28] , \wRegInTop_5_11[26] , 
        \wRegOut_6_26[8] , \wRegInTop_7_89[22] , \ScanLink226[2] , 
        \wRegInTop_2_0[11] , \wRegInBot_4_2[22] , \wRegInBot_5_27[24] , 
        \wRegInBot_5_28[7] , \ScanLink78[5] , \wRegEnTop_7_100[0] , 
        \wRegInTop_7_109[4] , \wRegOut_7_123[4] , \wRegInTop_4_7[31] , 
        \wRegInTop_4_7[28] , \ScanLink59[18] , \wRegInTop_6_37[3] , 
        \wRegInTop_7_12[27] , \ScanLink145[4] , \wRegInTop_7_67[17] , 
        \wRegInTop_7_16[5] , \wRegInTop_7_31[16] , \wRegInTop_7_24[22] , 
        \wRegInTop_7_44[26] , \ScanLink211[29] , \wRegInTop_7_51[12] , 
        \wRegOut_7_120[7] , \wRegInTop_7_72[23] , \ScanLink211[30] , 
        \ScanLink225[1] , \ScanLink232[18] , \ScanLink247[31] , 
        \wRegInTop_5_11[15] , \wRegOut_5_22[18] , \wRegInTop_6_1[8] , 
        \ScanLink247[28] , \ScanLink66[9] , \wRegInBot_6_5[26] , 
        \ScanLink197[2] , \wRegOut_7_7[4] , \wRegOut_6_38[4] , 
        \wRegInTop_7_117[8] , \wRegOut_7_19[2] , \wRegInTop_6_50[4] , 
        \ScanLink122[3] , \wRegInTop_7_89[11] , \wRegInTop_7_71[2] , 
        \ScanLink8[10] , \wRegInBot_3_7[8] , \wRegOut_5_4[16] , 
        \wRegInTop_5_27[10] , \wRegInBot_5_27[17] , \ScanLink179[19] , 
        \wRegInBot_5_11[12] , \ScanLink242[6] , \wRegOut_4_0[6] , 
        \wRegEnTop_5_3[0] , \wRegInTop_5_8[18] , \wRegOut_7_3[12] , 
        \wRegOut_2_3[1] , \wRegOut_4_3[5] , \wRegInTop_5_5[9] , 
        \wRegEnBot_6_50[0] , \wRegInBot_4_2[11] , \wRegInBot_6_5[15] , 
        \wRegInTop_6_53[7] , \wRegInTop_7_51[21] , \wRegInTop_7_72[1] , 
        \ScanLink121[0] , \wRegInTop_7_12[14] , \wRegInTop_7_24[11] , 
        \ScanLink182[18] , \wRegOut_7_60[9] , \wRegInTop_7_72[10] , 
        \ScanLink241[5] , \wRegInTop_7_67[24] , \wRegInTop_4_14[30] , 
        \wRegInTop_4_14[29] , \ScanLink112[11] , \wRegInTop_7_4[10] , 
        \wRegInTop_7_31[25] , \wRegInTop_7_44[15] , \ScanLink167[21] , 
        \wRegInTop_6_4[5] , \ScanLink144[10] , \wRegInBot_6_5[3] , 
        \ScanLink63[4] , \ScanLink131[20] , \ScanLink151[24] , 
        \ScanLink124[14] , \wRegOut_7_2[9] , \wRegInTop_7_97[30] , 
        \wRegInTop_7_112[5] , \wRegInBot_4_12[0] , \wRegInTop_5_3[14] , 
        \wRegOut_6_12[13] , \ScanLink107[25] , \ScanLink172[15] , 
        \wRegInTop_7_97[29] , \wRegOut_6_44[12] , \wRegInTop_7_13[8] , 
        \wRegOut_7_69[13] , \wRegOut_6_20[6] , \wRegOut_6_24[16] , 
        \wRegOut_6_31[22] , \ScanLink140[9] , \wRegOut_6_51[26] , 
        \wRegInBot_6_62[4] , \wRegOut_0_0[24] , \wRegInBot_3_1[14] , 
        \wRegOut_4_11[12] , \wRegOut_5_29[27] , \wRegOut_7_87[26] , 
        \wRegOut_7_92[12] , \wRegInTop_7_112[12] , \wRegOut_6_23[5] , 
        \wRegInTop_7_107[26] , \ScanLink11[12] , \wRegOut_4_0[19] , 
        \ScanLink32[23] , \wRegInBot_6_61[7] , \wRegEnTop_7_91[0] , 
        \wRegInTop_7_124[17] , \wRegOut_7_126[9] , \ScanLink47[13] , 
        \wRegInTop_6_7[6] , \wRegInBot_6_6[0] , \wRegInBot_4_11[3] , 
        \ScanLink27[17] , \ScanLink60[7] , \ScanLink64[22] , \ScanLink71[16] , 
        \wRegInTop_6_17[28] , \ScanLink239[27] , \wRegInTop_6_41[30] , 
        \wRegInTop_6_62[18] , \ScanLink189[14] , \wRegInTop_7_19[18] , 
        \wRegInTop_6_17[31] , \wRegEnTop_6_62[0] , \wRegInTop_6_34[19] , 
        \wRegInBot_5_30[5] , \wRegInTop_6_41[29] , \wRegInTop_5_3[27] , 
        \ScanLink52[27] , \wRegInTop_7_111[6] , \wRegOut_6_12[20] , 
        \wRegOut_6_24[25] , \wRegOut_6_51[15] , \wRegOut_6_31[11] , 
        \wRegOut_6_44[2] , \wRegOut_7_65[4] , \ScanLink244[8] , 
        \wRegOut_7_69[20] , \wRegOut_6_44[21] , \ScanLink124[27] , 
        \ScanLink139[2] , \wRegInTop_3_0[0] , \wRegInBot_3_1[6] , 
        \wRegOut_4_6[8] , \wRegEnBot_5_19[0] , \ScanLink151[17] , 
        \ScanLink107[16] , \wRegInBot_3_1[27] , \wRegInBot_3_2[5] , 
        \wRegInTop_5_0[4] , \ScanLink172[26] , \wRegInBot_5_1[2] , 
        \ScanLink112[22] , \wRegOut_5_15[0] , \ScanLink131[13] , 
        \wRegInTop_7_4[23] , \ScanLink167[12] , \ScanLink144[23] , 
        \wRegInTop_3_3[3] , \ScanLink71[25] , \ScanLink189[27] , 
        \ScanLink11[21] , \ScanLink27[24] , \ScanLink52[14] , 
        \wRegInBot_6_21[19] , \wRegInTop_6_48[6] , \wRegInBot_6_54[30] , 
        \wRegInTop_7_69[0] , \ScanLink32[10] , \ScanLink47[20] , 
        \wRegInBot_6_54[29] , \wRegOut_5_16[3] , \wRegOut_7_111[19] , 
        \wRegInTop_5_3[7] , \ScanLink64[11] , \ScanLink239[14] , 
        \wRegInBot_5_2[1] , \wRegInTop_5_19[4] , \wRegOut_7_87[15] , 
        \wRegOut_4_11[21] , \wRegInTop_6_55[9] , \wRegInTop_7_107[15] , 
        \wRegInTop_7_124[24] , \ScanLink0[9] , \wRegOut_1_0[13] , 
        \wRegOut_3_7[17] , \wRegInTop_4_3[10] , \wRegOut_5_29[14] , 
        \wRegOut_6_47[1] , \wRegOut_7_66[7] , \wRegOut_7_92[21] , 
        \wRegInTop_7_112[21] , \ScanLink48[14] , \wRegInBot_6_18[31] , 
        \wRegInBot_6_18[28] , \ScanLink215[11] , \ScanLink243[10] , 
        \wRegOut_7_20[2] , \ScanLink193[27] , \ScanLink236[20] , 
        \ScanLink186[13] , \ScanLink223[14] , \ScanLink28[10] , 
        \ScanLink90[0] , \wRegInBot_6_43[6] , \wRegOut_5_10[25] , 
        \wRegOut_5_26[20] , \ScanLink200[25] , \wRegOut_7_104[8] , 
        \wRegInTop_6_4[14] , \wRegOut_7_88[21] , \wRegInTop_7_108[21] , 
        \ScanLink42[6] , \wRegInBot_5_12[4] , \wRegOut_7_119[7] , 
        \ScanLink41[5] , \wRegOut_7_13[24] , \wRegOut_7_30[15] , 
        \wRegOut_7_66[14] , \wRegOut_7_45[25] , \wRegInBot_5_11[7] , 
        \wRegOut_7_7[19] , \wRegOut_7_25[21] , \wRegOut_7_50[11] , 
        \wRegOut_1_0[20] , \wRegInBot_2_1[10] , \wRegInBot_5_9[19] , 
        \wRegOut_7_73[20] , \wRegEnTop_5_12[0] , \wRegOut_6_9[4] , 
        \ScanLink90[24] , \ScanLink93[3] , \wRegInTop_7_31[9] , 
        \ScanLink162[8] , \ScanLink168[26] , \ScanLink85[10] , 
        \wRegOut_7_23[1] , \wRegOut_5_10[16] , \wRegInBot_5_15[19] , 
        \wRegInBot_6_40[5] , \ScanLink108[22] , \ScanLink118[0] , 
        \wRegInTop_7_84[8] , \wRegOut_7_88[12] , \wRegInTop_7_108[12] , 
        \ScanLink3[26] , \wRegInBot_2_1[23] , \wRegOut_3_7[24] , 
        \ScanLink26[2] , \wRegOut_4_15[4] , \wRegOut_5_26[13] , 
        \wRegInTop_6_4[27] , \wRegOut_7_59[9] , \wRegOut_7_96[0] , 
        \ScanLink186[20] , \ScanLink223[27] , \wRegInTop_4_3[23] , 
        \wRegInBot_4_6[30] , \wRegInBot_4_6[29] , \wRegOut_6_8[30] , 
        \ScanLink200[16] , \wRegInTop_7_99[7] , \ScanLink28[23] , 
        \wRegOut_6_8[29] , \ScanLink48[27] , \wRegInTop_7_20[29] , 
        \ScanLink215[22] , \wRegInTop_5_23[28] , \wRegInBot_6_27[2] , 
        \wRegInTop_7_20[30] , \wRegInTop_7_55[19] , \wRegInTop_7_76[31] , 
        \wRegOut_7_44[6] , \ScanLink193[14] , \ScanLink236[13] , 
        \wRegInTop_7_76[28] , \ScanLink243[23] , \ScanLink108[11] , 
        \ScanLink5[4] , \wRegInTop_3_0[26] , \wRegOut_4_4[21] , 
        \ScanLink25[1] , \wRegInTop_5_23[31] , \wRegInTop_5_25[9] , 
        \ScanLink85[23] , \wRegInBot_6_24[1] , \ScanLink90[17] , 
        \wRegOut_7_47[5] , \wRegOut_7_25[12] , \ScanLink168[15] , 
        \wRegInTop_7_48[2] , \wRegOut_7_50[22] , \wRegOut_7_73[13] , 
        \wRegOut_7_13[17] , \wRegOut_7_66[27] , \wRegOut_7_95[3] , 
        \wRegOut_7_45[16] , \wRegOut_7_30[26] , \wRegInTop_6_15[2] , 
        \wRegInTop_7_34[4] , \ScanLink167[5] , \ScanLink44[8] , 
        \ScanLink59[7] , \wRegOut_6_3[25] , \wRegInTop_6_13[10] , 
        \wRegInBot_6_45[8] , \ScanLink207[0] , \wRegOut_7_102[6] , 
        \wRegInBot_6_25[12] , \wRegInTop_6_45[11] , \wRegInTop_7_68[10] , 
        \wRegOut_7_123[17] , \wRegInTop_6_30[21] , \wRegInBot_6_30[26] , 
        \wRegInBot_6_50[22] , \wRegOut_7_100[26] , \wRegInBot_6_13[17] , 
        \wRegInTop_6_25[15] , \wRegInBot_6_45[16] , \wRegInTop_6_50[25] , 
        \wRegOut_7_115[12] , \ScanLink198[18] , \ScanLink6[7] , 
        \wRegInTop_4_10[11] , \wRegInBot_4_10[16] , \wRegInTop_5_28[24] , 
        \wRegInBot_6_58[7] , \ScanLink179[9] , \wRegInTop_7_93[11] , 
        \ScanLink116[29] , \wRegInTop_7_86[25] , \wRegOut_7_38[0] , 
        \wRegOut_6_19[6] , \wRegInTop_7_0[28] , \wRegOut_2_3[18] , 
        \ScanLink7[24] , \wRegInBot_5_2[26] , \wRegInBot_5_17[9] , 
        \wRegInBot_5_28[23] , \ScanLink88[2] , \ScanLink140[31] , 
        \ScanLink163[19] , \ScanLink116[30] , \ScanLink135[18] , 
        \wRegInTop_7_0[31] , \wRegInTop_6_16[1] , \ScanLink140[28] , 
        \ScanLink164[6] , \wRegInTop_7_37[7] , \wRegInTop_7_9[6] , 
        \ScanLink7[17] , \wRegInTop_3_0[15] , \ScanLink15[19] , 
        \ScanLink36[28] , \wRegInBot_6_45[25] , \ScanLink204[3] , 
        \wRegOut_7_101[5] , \ScanLink43[18] , \wRegInTop_6_25[26] , 
        \wRegInTop_7_82[6] , \wRegOut_7_115[21] , \ScanLink60[30] , 
        \wRegInBot_6_30[15] , \wRegInTop_6_50[16] , \ScanLink36[31] , 
        \wRegInTop_5_20[4] , \ScanLink60[29] , \wRegInBot_6_13[24] , 
        \wRegOut_6_3[16] , \wRegInTop_6_13[23] , \wRegInTop_6_30[12] , 
        \wRegInTop_7_68[23] , \wRegOut_7_123[24] , \ScanLink228[18] , 
        \wRegOut_7_100[15] , \wRegInBot_6_25[21] , \wRegInTop_6_45[22] , 
        \wRegInBot_6_50[11] , \ScanLink103[1] , \wRegInTop_7_50[0] , 
        \wRegOut_4_4[12] , \wRegOut_5_8[8] , \wRegOut_7_96[19] , 
        \wRegInTop_7_116[19] , \wRegOut_4_15[19] , \wRegOut_7_42[8] , 
        \wRegEnBot_5_20[0] , \wRegOut_6_16[18] , \wRegOut_6_63[28] , 
        \wRegOut_7_18[28] , \wRegOut_6_35[30] , \ScanLink100[2] , 
        \wRegOut_6_40[19] , \wRegOut_6_63[31] , \wRegInTop_7_53[3] , 
        \wRegOut_7_18[31] , \wRegOut_6_35[29] , \wRegInBot_5_2[15] , 
        \wRegOut_4_10[9] , \wRegInTop_4_10[22] , \wRegInTop_5_23[7] , 
        \wRegInTop_7_86[16] , \wRegInBot_5_28[10] , \wRegInTop_7_81[5] , 
        \wRegInBot_4_10[25] , \wRegInTop_5_28[17] , \wRegInBot_5_6[24] , 
        \wRegOut_6_12[30] , \wRegOut_6_12[29] , \wRegInTop_7_93[22] , 
        \wRegOut_6_31[18] , \wRegOut_6_44[31] , \wRegOut_7_69[29] , 
        \ScanLink244[1] , \wRegOut_6_44[28] , \wRegOut_7_69[30] , 
        \wRegInTop_6_56[3] , \ScanLink124[4] , \wRegInTop_7_77[5] , 
        \wRegOut_7_8[24] , \wRegInTop_3_0[9] , \wRegOut_4_6[1] , 
        \wRegInTop_4_14[13] , \wRegOut_6_59[4] , \wRegOut_7_78[2] , 
        \wRegInTop_7_82[27] , \wRegOut_5_15[9] , \wRegInTop_7_97[13] , 
        \ScanLink11[31] , \wRegInBot_4_14[14] , \ScanLink32[19] , 
        \ScanLink47[29] , \wRegInBot_6_34[24] , \wRegInTop_6_54[27] , 
        \wRegOut_7_111[10] , \wRegInBot_6_41[14] , \ScanLink11[28] , 
        \ScanLink47[30] , \ScanLink64[18] , \wRegInTop_6_21[17] , 
        \wRegInBot_6_17[15] , \wRegInBot_6_62[25] , \wRegInTop_7_79[26] , 
        \wRegInTop_3_4[24] , \wRegEnTop_3_6[0] , \wRegOut_4_5[2] , 
        \wRegInBot_5_2[8] , \wRegInBot_6_18[5] , \wRegInBot_4_9[27] , 
        \wRegInTop_6_62[22] , \wRegInTop_7_19[22] , \wRegOut_6_7[27] , 
        \wRegInTop_6_17[12] , \wRegInBot_6_21[10] , \wRegInTop_6_41[13] , 
        \wRegOut_7_127[15] , \wRegInTop_7_69[9] , \wRegInTop_6_34[23] , 
        \wRegInBot_6_54[20] , \wRegOut_7_104[24] , \wRegOut_4_0[23] , 
        \ScanLink19[5] , \wRegOut_4_11[28] , \wRegOut_6_47[8] , 
        \wRegOut_7_92[31] , \wRegInTop_7_112[31] , \wRegOut_7_92[28] , 
        \wRegInTop_7_112[28] , \ScanLink247[2] , \wRegOut_4_11[31] , 
        \wRegInTop_6_55[0] , \wRegInTop_7_74[6] , \ScanLink127[7] , 
        \wRegInBot_4_12[9] , \wRegOut_7_2[0] , \wRegInBot_4_14[27] , 
        \wRegInTop_7_4[19] , \wRegInTop_7_97[20] , \ScanLink167[28] , 
        \wRegOut_0_0[5] , \wRegInBot_0_0[3] , \wRegOut_1_1[7] , 
        \ScanLink3[15] , \wRegInTop_4_14[20] , \wRegEnBot_6_31[0] , 
        \wRegInTop_7_82[14] , \wRegEnBot_6_0[0] , \ScanLink112[18] , 
        \ScanLink131[30] , \ScanLink131[29] , \ScanLink144[19] , 
        \ScanLink167[31] , \ScanLink192[6] , \wRegOut_7_8[17] , 
        \ScanLink220[5] , \wRegOut_7_125[3] , \wRegInTop_3_4[17] , 
        \wRegOut_4_0[10] , \wRegInBot_5_6[17] , \wRegInTop_6_32[7] , 
        \ScanLink140[0] , \wRegInTop_7_13[1] , \wRegInTop_6_31[4] , 
        \ScanLink143[3] , \ScanLink223[6] , \wRegOut_7_126[0] , 
        \wRegInTop_7_10[2] , \wRegInBot_4_9[14] , \wRegInTop_6_17[21] , 
        \wRegInTop_6_62[11] , \wRegOut_7_127[26] , \wRegInBot_6_6[9] , 
        \wRegOut_6_7[14] , \wRegInTop_6_34[10] , \wRegOut_7_1[3] , 
        \wRegInTop_7_19[11] , \wRegInBot_6_54[13] , \wRegOut_7_104[17] , 
        \wRegInTop_6_21[24] , \wRegInBot_6_21[23] , \wRegInTop_6_41[20] , 
        \wRegInBot_6_41[27] , \ScanLink191[5] , \wRegOut_7_111[23] , 
        \wRegInBot_6_34[17] , \wRegInTop_6_54[14] , \wRegInTop_2_0[18] , 
        \wRegInTop_5_27[19] , \wRegInBot_6_17[26] , \wRegInBot_6_62[16] , 
        \wRegInTop_7_79[15] , \ScanLink81[12] , \ScanLink179[10] , 
        \ScanLink94[26] , \wRegOut_6_42[5] , \wRegOut_7_63[3] , 
        \ScanLink119[14] , \wRegInTop_7_89[18] , \wRegOut_2_3[8] , 
        \ScanLink8[19] , \wRegOut_5_13[7] , \wRegOut_7_21[23] , 
        \wRegOut_7_54[13] , \wRegInTop_3_6[7] , \wRegInBot_3_7[1] , 
        \wRegInTop_5_6[3] , \wRegInBot_5_7[5] , \wRegOut_7_77[22] , 
        \wRegOut_7_17[26] , \wRegInTop_5_5[0] , \wRegInTop_5_8[11] , 
        \wRegOut_6_19[16] , \wRegOut_7_62[16] , \wRegOut_7_34[17] , 
        \wRegOut_7_41[27] , \wRegOut_5_14[27] , \wRegOut_3_3[26] , 
        \wRegOut_3_3[15] , \wRegInBot_3_4[2] , \wRegInBot_5_4[6] , 
        \wRegOut_5_10[4] , \wRegOut_5_22[22] , \wRegInTop_6_0[16] , 
        \wRegInTop_3_5[4] , \wRegOut_7_99[17] , \wRegInTop_7_119[17] , 
        \wRegInBot_4_2[18] , \wRegOut_6_41[6] , \wRegOut_7_60[0] , 
        \ScanLink252[26] , \ScanLink182[11] , \ScanLink227[16] , 
        \wRegInTop_4_7[21] , \wRegInTop_4_7[12] , \ScanLink59[22] , 
        \ScanLink204[27] , \wRegInTop_7_51[28] , \wRegInBot_4_14[7] , 
        \ScanLink39[26] , \wRegInTop_7_72[8] , \wRegInTop_5_8[22] , 
        \ScanLink65[3] , \wRegOut_6_19[25] , \ScanLink121[9] , 
        \wRegInTop_7_24[18] , \wRegInTop_7_51[31] , \wRegInTop_7_72[19] , 
        \ScanLink211[13] , \ScanLink197[25] , \ScanLink247[12] , 
        \ScanLink232[22] , \wRegOut_7_17[15] , \wRegOut_7_62[25] , 
        \wRegOut_7_41[14] , \wRegOut_7_34[24] , \wRegInTop_7_114[2] , 
        \wRegInBot_5_11[31] , \wRegInTop_6_2[2] , \wRegInTop_6_29[6] , 
        \wRegOut_7_54[20] , \ScanLink194[8] , \wRegInBot_6_3[4] , 
        \wRegOut_7_21[10] , \wRegOut_6_26[1] , \wRegOut_7_3[31] , 
        \wRegOut_7_3[28] , \wRegOut_7_77[11] , \ScanLink94[15] , 
        \ScanLink119[27] , \wRegInTop_6_34[9] , \ScanLink189[7] , 
        \wRegInBot_5_11[28] , \ScanLink81[21] , \ScanLink179[23] , 
        \ScanLink211[20] , \ScanLink39[15] , \wRegOut_6_25[2] , 
        \ScanLink182[22] , \ScanLink197[16] , \ScanLink225[8] , 
        \ScanLink227[25] , \ScanLink232[11] , \ScanLink247[21] , 
        \ScanLink59[11] , \ScanLink204[14] , \ScanLink252[15] , 
        \ScanLink0[19] , \wRegOut_1_1[19] , \wRegInBot_2_0[30] , 
        \wRegInBot_2_0[29] , \wRegInTop_2_1[21] , \wRegInBot_3_0[24] , 
        \wRegInBot_3_0[17] , \ScanLink10[11] , \ScanLink26[14] , 
        \wRegOut_5_14[14] , \wRegOut_5_22[11] , \ScanLink66[0] , 
        \wRegInTop_6_0[25] , \ScanLink238[7] , \wRegInTop_7_117[1] , 
        \wRegOut_7_99[24] , \wRegInTop_7_119[24] , \wRegInBot_6_0[7] , 
        \wRegInTop_6_1[1] , \ScanLink158[2] , \ScanLink70[4] , 
        \wRegInBot_6_55[19] , \wRegInBot_5_20[6] , \ScanLink53[24] , 
        \wRegInTop_7_101[5] , \ScanLink70[15] , \wRegInBot_6_20[30] , 
        \wRegInBot_6_20[29] , \ScanLink188[17] , \wRegOut_7_110[30] , 
        \wRegOut_4_10[11] , \ScanLink33[20] , \ScanLink65[21] , 
        \wRegOut_7_110[29] , \ScanLink238[24] , \ScanLink46[10] , 
        \wEnable_6[0] , \wRegOut_7_86[25] , \wRegInTop_7_125[14] , 
        \wRegOut_6_33[6] , \wRegOut_7_12[0] , \wRegInTop_7_106[25] , 
        \wRegOut_4_1[30] , \wRegInTop_5_2[17] , \wRegOut_5_28[24] , 
        \ScanLink153[9] , \wRegOut_7_93[11] , \wRegInTop_7_113[11] , 
        \wRegOut_6_25[15] , \wRegOut_6_30[5] , \wRegOut_6_50[25] , 
        \wRegOut_7_11[3] , \wRegEnTop_7_82[0] , \wRegInBot_5_23[5] , 
        \wRegInTop_6_9[9] , \wRegOut_6_45[11] , \ScanLink73[7] , 
        \wRegOut_6_13[10] , \wRegOut_6_30[21] , \ScanLink106[26] , 
        \ScanLink173[16] , \wRegOut_7_68[10] , \ScanLink150[27] , 
        \ScanLink125[17] , \wRegOut_5_28[17] , \wRegInBot_6_15[0] , 
        \ScanLink113[12] , \ScanLink130[23] , \ScanLink145[13] , 
        \wRegInTop_7_102[6] , \wRegInTop_7_5[13] , \ScanLink166[22] , 
        \wRegOut_6_57[2] , \wRegOut_7_76[4] , \wRegOut_7_93[22] , 
        \wRegInTop_7_113[22] , \wRegInTop_7_125[27] , \wRegOut_4_1[29] , 
        \wRegOut_4_8[7] , \wRegOut_7_86[16] , \ScanLink10[22] , 
        \wRegOut_4_10[22] , \ScanLink65[12] , \wRegInTop_7_106[16] , 
        \ScanLink238[17] , \ScanLink14[0] , \ScanLink46[23] , \ScanLink17[3] , 
        \ScanLink26[27] , \ScanLink33[13] , \ScanLink53[17] , 
        \wRegInTop_6_40[19] , \wRegInTop_6_63[31] , \wRegInTop_7_79[3] , 
        \wRegInTop_6_58[5] , \wRegInTop_7_18[31] , \wRegInTop_6_35[29] , 
        \wRegInTop_5_14[8] , \ScanLink70[26] , \wRegInTop_6_63[28] , 
        \wRegInTop_7_18[28] , \ScanLink188[24] , \wRegInTop_6_16[18] , 
        \wRegInTop_6_35[30] , \wRegInBot_4_3[21] , \wRegInTop_4_15[19] , 
        \ScanLink130[10] , \ScanLink145[20] , \wRegInTop_5_2[24] , 
        \wRegOut_6_30[12] , \ScanLink106[15] , \ScanLink113[21] , 
        \ScanLink249[4] , \wRegInTop_7_5[20] , \wRegOut_7_68[8] , 
        \ScanLink166[11] , \ScanLink125[24] , \ScanLink173[25] , 
        \wRegInTop_7_96[19] , \ScanLink129[1] , \ScanLink150[14] , 
        \wRegOut_6_45[22] , \wRegInBot_5_26[8] , \wRegOut_6_13[23] , 
        \wRegInBot_6_16[3] , \wRegOut_6_54[1] , \wRegOut_7_68[23] , 
        \wRegOut_7_75[7] , \wRegOut_6_25[26] , \wRegOut_6_28[7] , 
        \wRegInTop_6_46[9] , \wRegOut_6_50[16] , \wRegInBot_6_4[25] , 
        \ScanLink148[8] , \ScanLink187[1] , \wRegInTop_6_27[0] , 
        \wRegOut_6_35[8] , \ScanLink235[2] , \wRegInTop_7_25[21] , 
        \wRegInTop_7_73[20] , \ScanLink155[7] , \wRegInTop_7_50[11] , 
        \ScanLink183[31] , \wRegInTop_7_13[24] , \wRegInTop_7_30[15] , 
        \wRegInTop_7_45[25] , \ScanLink183[28] , \wRegInTop_7_66[14] , 
        \wRegInTop_2_1[12] , \ScanLink9[20] , \wRegOut_5_5[26] , 
        \wRegInTop_5_10[25] , \wRegInBot_5_26[27] , \ScanLink68[6] , 
        \wRegInTop_7_88[21] , \ScanLink236[1] , \wRegInTop_7_119[7] , 
        \wRegInBot_5_10[22] , \ScanLink178[29] , \wRegEnTop_7_113[0] , 
        \wRegInTop_5_9[31] , \wRegInTop_5_9[28] , \wRegInTop_5_26[20] , 
        \wRegInTop_6_24[3] , \ScanLink156[4] , \ScanLink178[30] , 
        \ScanLink75[9] , \wRegInTop_7_104[8] , \ScanLink9[13] , 
        \wRegInBot_4_3[12] , \wRegInTop_5_8[5] , \ScanLink58[28] , 
        \wRegOut_7_2[22] , \ScanLink184[2] , \wRegInTop_7_30[26] , 
        \wRegInTop_7_45[16] , \wRegInBot_5_9[3] , \wRegInTop_7_66[27] , 
        \ScanLink251[6] , \ScanLink58[31] , \wRegInTop_4_6[18] , 
        \wRegInTop_7_13[17] , \wRegInTop_7_62[2] , \wRegInTop_7_73[13] , 
        \ScanLink233[28] , \ScanLink246[18] , \wRegInTop_5_12[6] , 
        \wRegInBot_6_4[16] , \wRegInTop_6_43[4] , \wRegInTop_7_50[22] , 
        \ScanLink131[3] , \wRegInTop_7_25[12] , \ScanLink210[19] , 
        \ScanLink233[31] , \wRegOut_5_23[31] , \wRegOut_5_23[28] , 
        \wRegOut_7_20[30] , \wRegOut_5_5[15] , \wRegInTop_5_11[5] , 
        \wRegOut_7_2[11] , \wRegOut_7_20[29] , \wRegOut_7_76[28] , 
        \wRegOut_7_55[19] , \wRegOut_7_76[31] , \wRegEnBot_6_43[0] , 
        \wRegInBot_5_10[11] , \ScanLink80[18] , \wRegOut_7_73[9] , 
        \ScanLink252[5] , \wRegInTop_5_26[13] , \wRegInTop_6_40[7] , 
        \ScanLink132[0] , \wRegInTop_7_61[1] , \wRegOut_3_0[4] , 
        \wRegEnBot_4_2[0] , \wRegInTop_4_14[5] , \wRegInTop_5_10[16] , 
        \wRegInBot_5_26[14] , \wRegOut_7_51[31] , \wRegInTop_7_88[12] , 
        \wRegOut_5_0[0] , \wRegInBot_5_8[20] , \wRegOut_7_72[19] , 
        \wRegOut_7_6[20] , \wRegOut_7_24[18] , \wRegOut_7_51[28] , 
        \wRegInTop_7_58[8] , \wRegInTop_7_97[1] , \wRegOut_7_85[9] , 
        \wRegOut_5_1[24] , \wRegInBot_5_14[20] , \wRegInBot_6_29[4] , 
        \ScanLink84[29] , \wRegInTop_7_99[17] , \wRegInTop_5_22[22] , 
        \ScanLink84[30] , \ScanLink116[6] , \wRegInTop_7_45[7] , 
        \wRegOut_3_3[7] , \wRegInTop_4_2[30] , \wRegInBot_4_7[23] , 
        \ScanLink28[4] , \wRegInBot_5_22[25] , \ScanLink29[29] , 
        \wRegInTop_5_14[27] , \wRegOut_7_98[6] , \ScanLink115[5] , 
        \wRegInTop_7_34[17] , \wRegInTop_7_46[4] , \wRegInTop_7_41[27] , 
        \wRegOut_6_9[23] , \wRegInTop_7_17[26] , \ScanLink29[30] , 
        \wRegInTop_6_19[16] , \wRegInBot_6_19[11] , \wRegInTop_7_62[16] , 
        \wRegInTop_7_77[22] , \ScanLink214[31] , \ScanLink237[19] , 
        \wRegInTop_4_2[29] , \wRegEnTop_6_29[0] , \wRegInBot_6_37[8] , 
        \ScanLink242[29] , \wRegInTop_7_21[23] , \wRegInTop_7_54[13] , 
        \ScanLink214[28] , \wRegOut_5_3[3] , \wRegInBot_6_0[27] , 
        \wRegInTop_7_94[2] , \ScanLink242[30] , \wRegOut_7_89[18] , 
        \wRegInTop_7_109[18] , \wRegInBot_4_4[9] , \wRegOut_5_1[17] , 
        \ScanLink36[8] , \wRegOut_7_49[3] , \wRegInTop_5_14[14] , 
        \wRegInBot_5_22[16] , \wRegOut_5_24[8] , \wRegOut_5_27[19] , 
        \wRegInTop_7_21[3] , \ScanLink172[2] , \wRegInBot_5_8[13] , 
        \wRegInBot_5_14[13] , \ScanLink109[28] , \ScanLink212[7] , 
        \wRegInTop_5_22[11] , \wRegInTop_7_99[24] , \ScanLink83[9] , 
        \ScanLink109[31] , \wRegOut_7_117[1] , \wRegInBot_6_0[14] , 
        \wRegOut_6_4[1] , \wRegOut_7_6[13] , \wRegInTop_2_0[6] , 
        \wRegInBot_4_7[10] , \wRegOut_6_7[2] , \wRegOut_6_9[10] , 
        \wRegInBot_6_19[22] , \wRegInTop_7_77[11] , \wRegInTop_7_21[10] , 
        \wRegInTop_7_22[0] , \wRegInTop_7_54[20] , \ScanLink171[1] , 
        \wRegInTop_6_19[25] , \wRegInTop_7_34[24] , \wRegInTop_7_41[14] , 
        \wRegOut_7_114[2] , \wRegOut_7_30[8] , \ScanLink187[19] , 
        \wRegInTop_7_62[25] , \ScanLink211[4] , \wRegInTop_4_11[31] , 
        \ScanLink134[21] , \ScanLink141[11] , \wRegInTop_7_17[15] , 
        \wRegInTop_7_1[11] , \wRegInBot_2_1[0] , \ScanLink162[20] , 
        \wRegOut_2_2[21] , \wRegOut_2_2[12] , \wRegInTop_4_0[2] , 
        \wRegInBot_4_1[4] , \wRegInTop_4_11[28] , \ScanLink117[10] , 
        \ScanLink177[14] , \wRegOut_7_83[7] , \ScanLink33[5] , 
        \wRegOut_5_21[5] , \ScanLink102[24] , \wRegInTop_7_92[28] , 
        \ScanLink154[25] , \wRegInTop_5_6[15] , \ScanLink121[15] , 
        \wRegInTop_7_43[9] , \wRegInTop_7_92[31] , \wRegOut_6_17[12] , 
        \wRegOut_6_34[23] , \wRegOut_6_41[13] , \ScanLink110[8] , 
        \wRegOut_6_62[22] , \wRegOut_7_19[22] , \wRegInBot_6_32[5] , 
        \wRegOut_7_51[1] , \wRegOut_7_79[26] , \wRegInBot_2_2[3] , 
        \wRegInTop_2_3[5] , \wRegInBot_3_4[15] , \wRegOut_4_14[13] , 
        \wRegOut_6_21[17] , \wRegOut_6_54[27] , \wRegOut_7_82[27] , 
        \wRegOut_7_97[13] , \wRegInTop_7_117[13] , \wRegInTop_7_121[16] , 
        \wRegInTop_7_102[27] , \wRegOut_7_52[2] , \wRegOut_4_5[18] , 
        \wRegInBot_6_31[6] , \ScanLink14[13] , \wRegInTop_4_11[8] , 
        \ScanLink61[23] , \ScanLink249[16] , \wRegOut_3_5[9] , 
        \wRegInBot_4_2[7] , \ScanLink22[16] , \wRegInTop_4_9[16] , 
        \ScanLink199[21] , \ScanLink30[6] , \ScanLink37[22] , \ScanLink42[12] , 
        \wRegInTop_6_12[30] , \wRegOut_5_22[6] , \wRegInTop_6_31[18] , 
        \wRegInTop_7_69[30] , \ScanLink57[26] , \wRegInTop_6_44[28] , 
        \wRegInTop_6_12[29] , \wRegInTop_4_3[1] , \wRegInTop_6_44[31] , 
        \wRegInTop_7_69[29] , \wRegOut_7_80[4] , \ScanLink229[12] , 
        \ScanLink74[17] , \wRegOut_7_79[15] , \ScanLink8[1] , 
        \wRegInBot_3_4[26] , \ScanLink14[20] , \ScanLink22[25] , 
        \wRegInTop_5_6[26] , \wRegOut_6_21[24] , \ScanLink85[7] , 
        \wRegOut_6_34[10] , \wRegOut_6_54[14] , \wRegOut_6_41[20] , 
        \ScanLink57[15] , \ScanLink57[1] , \wRegOut_6_14[3] , 
        \wRegOut_6_17[21] , \wRegOut_7_35[5] , \ScanLink214[9] , 
        \ScanLink102[17] , \wRegInBot_6_56[1] , \wRegOut_6_62[11] , 
        \wRegOut_7_19[11] , \ScanLink121[26] , \ScanLink169[3] , 
        \ScanLink177[27] , \wRegInTop_7_4[3] , \ScanLink154[16] , 
        \wRegInBot_5_29[30] , \wRegInBot_5_29[29] , \wRegEnTop_7_74[0] , 
        \ScanLink98[8] , \ScanLink134[12] , \ScanLink141[22] , 
        \wRegInTop_7_126[0] , \wRegInTop_6_18[7] , \ScanLink117[23] , 
        \wRegInTop_7_1[22] , \ScanLink209[6] , \ScanLink162[13] , 
        \wRegInTop_7_39[1] , \wRegInBot_6_24[18] , \ScanLink61[10] , 
        \ScanLink74[24] , \wRegInBot_6_51[28] , \wRegInTop_7_7[0] , 
        \ScanLink229[21] , \wRegInBot_6_51[31] , \ScanLink199[12] , 
        \wRegInTop_4_9[25] , \ScanLink42[21] , \ScanLink249[25] , 
        \ScanLink54[2] , \ScanLink37[11] , \wRegOut_7_82[14] , 
        \wRegOut_7_114[18] , \wRegInTop_7_121[25] , \wRegInTop_7_125[3] , 
        \wRegOut_4_14[20] , \wRegInTop_7_102[14] , \wRegOut_6_17[0] , 
        \wRegOut_7_36[6] , \wRegOut_7_97[20] , \wRegInTop_7_117[20] , 
        \wRegOut_3_1[9] , \wRegInBot_3_2[22] , \wRegOut_4_12[24] , 
        \wRegInTop_5_29[1] , \ScanLink86[4] , \wRegInBot_6_55[2] , 
        \wRegInTop_7_127[21] , \wRegInTop_7_104[10] , \wRegInTop_3_7[31] , 
        \wRegOut_7_84[10] , \wRegInTop_3_7[28] , \ScanLink29[9] , 
        \wRegInTop_6_8[25] , \wRegInBot_6_35[6] , \wRegOut_7_56[2] , 
        \wRegOut_7_91[24] , \wRegInTop_7_111[24] , \wRegInBot_4_6[7] , 
        \ScanLink24[21] , \ScanLink51[11] , \wRegInTop_7_59[5] , 
        \wRegInTop_4_15[8] , \ScanLink72[20] , \wRegOut_7_107[28] , 
        \wRegOut_7_107[31] , \wRegOut_7_124[19] , \wRegInBot_3_2[11] , 
        \ScanLink12[24] , \wRegInTop_4_7[1] , \ScanLink67[14] , 
        \wRegInBot_6_37[31] , \wRegOut_7_84[4] , \wRegInBot_6_14[19] , 
        \wRegInBot_6_28[9] , \wRegInBot_6_61[29] , \ScanLink12[17] , 
        \wRegInTop_4_4[2] , \wRegInBot_4_5[4] , \ScanLink31[15] , 
        \ScanLink34[6] , \ScanLink219[20] , \ScanLink44[25] , 
        \wRegOut_5_26[6] , \wRegInBot_6_37[28] , \wRegInBot_6_61[30] , 
        \ScanLink37[5] , \wRegInBot_5_19[31] , \wRegInBot_5_19[28] , 
        \wRegInBot_6_42[18] , \ScanLink89[21] , \ScanLink104[13] , 
        \ScanLink109[7] , \ScanLink127[22] , \ScanLink171[23] , 
        \wRegOut_5_25[5] , \ScanLink152[12] , \ScanLink132[16] , 
        \ScanLink111[27] , \ScanLink147[26] , \wRegOut_7_87[7] , 
        \wRegInTop_5_0[22] , \wRegInBot_5_5[31] , \wRegInBot_5_5[28] , 
        \wRegInTop_7_7[26] , \ScanLink164[17] , \wRegOut_6_27[20] , 
        \wRegInTop_7_47[9] , \wRegOut_6_32[14] , \ScanLink114[8] , 
        \wRegOut_6_52[10] , \wRegInTop_7_88[0] , \wRegOut_7_29[10] , 
        \wRegOut_7_49[14] , \wRegOut_6_11[25] , \wRegOut_6_47[24] , 
        \wRegOut_7_55[1] , \wRegInTop_6_22[31] , \wRegInBot_6_36[5] , 
        \ScanLink24[12] , \ScanLink31[26] , \ScanLink67[27] , 
        \wRegInTop_7_59[31] , \wRegInTop_6_22[28] , \wRegInTop_7_59[28] , 
        \ScanLink44[16] , \wRegInTop_6_57[18] , \ScanLink219[13] , 
        \wRegInTop_7_3[0] , \ScanLink50[2] , \wRegOut_6_4[18] , 
        \ScanLink51[22] , \wRegInTop_6_8[16] , \ScanLink72[13] , 
        \wRegInTop_7_121[3] , \wRegOut_7_91[17] , \ScanLink82[4] , 
        \wRegInTop_7_111[17] , \wRegInTop_7_127[12] , \wRegOut_4_12[17] , 
        \wRegOut_7_32[6] , \wRegInTop_5_0[11] , \wRegOut_6_13[0] , 
        \wRegInTop_7_104[23] , \wRegOut_6_47[17] , \wRegInBot_6_51[2] , 
        \wRegOut_7_84[23] , \wRegOut_6_11[16] , \wRegOut_6_32[27] , 
        \wRegOut_7_49[27] , \wRegEnTop_1_0[0] , \wRegInTop_1_0[7] , 
        \ScanLink53[1] , \wRegOut_6_10[3] , \wRegOut_7_31[5] , 
        \ScanLink210[9] , \ScanLink81[7] , \wRegOut_6_52[23] , 
        \wRegInBot_6_52[1] , \ScanLink89[12] , \wRegOut_6_27[13] , 
        \wRegOut_7_29[23] , \ScanLink111[14] , \wRegInTop_7_0[3] , 
        \ScanLink132[25] , \ScanLink147[15] , \wRegInTop_7_7[15] , 
        \ScanLink164[24] , \wRegInTop_7_81[18] , \ScanLink104[20] , 
        \ScanLink171[10] , \ScanLink152[21] , \wRegEnTop_7_70[0] , 
        \wRegInBot_1_1[1] , \wRegOut_7_108[0] , \wRegInTop_7_122[0] , 
        \wRegInTop_2_2[8] , \wRegOut_3_0[19] , \wRegInTop_6_29[24] , 
        \ScanLink111[5] , \ScanLink127[11] , \ScanLink194[29] , 
        \wRegInTop_7_71[15] , \wRegInBot_6_29[23] , \wRegInBot_6_49[27] , 
        \wRegInTop_6_63[2] , \wRegInTop_7_27[14] , \wRegInTop_7_42[4] , 
        \wRegInTop_7_52[24] , \wRegOut_7_119[23] , \ScanLink194[30] , 
        \wRegInTop_7_47[10] , \wRegInTop_6_49[20] , \wRegInTop_7_32[20] , 
        \wRegInTop_7_11[11] , \wRegInTop_7_64[21] , \wRegOut_3_7[7] , 
        \wRegInBot_4_1[14] , \wRegOut_4_8[10] , \wRegInTop_4_13[6] , 
        \wRegInBot_6_33[8] , \ScanLink32[8] , \wRegOut_5_7[3] , 
        \wRegInTop_7_90[2] , \wRegOut_5_20[8] , \wRegInBot_6_6[10] , 
        \wRegInBot_4_0[9] , \wRegInTop_4_10[5] , \wRegInTop_5_31[3] , 
        \wRegInTop_7_93[1] , \wRegInTop_2_3[14] , \wRegOut_3_4[4] , 
        \wRegEnBot_4_6[0] , \wRegOut_5_4[0] , \wRegOut_7_81[9] , 
        \wRegInBot_5_24[12] , \wRegInTop_5_31[21] , \ScanLink112[6] , 
        \wRegInTop_6_60[1] , \wRegOut_7_0[17] , \wRegInTop_7_41[7] , 
        \ScanLink139[29] , \wRegOut_4_8[23] , \wRegOut_5_7[13] , 
        \wRegInTop_5_12[10] , \ScanLink139[30] , \wRegInBot_5_12[17] , 
        \wRegOut_5_17[18] , \wRegInTop_5_24[15] , \wRegInBot_5_31[26] , 
        \wRegInBot_6_6[23] , \wRegInTop_6_3[29] , \wRegOut_7_29[7] , 
        \ScanLink99[5] , \wRegInTop_2_3[27] , \wRegInBot_4_1[27] , 
        \wRegOut_6_3[2] , \wRegInTop_6_3[30] , \wRegInBot_6_29[10] , 
        \wRegInTop_7_26[0] , \wRegInTop_7_32[13] , \wRegInTop_6_49[13] , 
        \ScanLink224[30] , \wRegInTop_7_47[23] , \ScanLink175[1] , 
        \ScanLink207[18] , \ScanLink19[31] , \ScanLink19[28] , 
        \wRegInTop_7_11[22] , \wRegOut_7_34[8] , \wRegInTop_7_64[12] , 
        \ScanLink224[29] , \ScanLink251[19] , \wRegInTop_7_71[26] , 
        \ScanLink215[4] , \wRegInTop_6_29[17] , \wRegInTop_7_27[27] , 
        \wRegInBot_6_49[14] , \wRegInTop_7_52[17] , \wRegOut_7_119[10] , 
        \wRegOut_7_110[2] , \wRegOut_5_7[20] , \wRegInBot_5_12[24] , 
        \ScanLink48[0] , \wRegInTop_5_24[26] , \wRegInBot_5_31[15] , 
        \wRegInTop_7_25[3] , \ScanLink176[2] , \wRegInBot_5_24[21] , 
        \ScanLink87[9] , \wRegInTop_5_12[23] , \wRegInBot_5_18[2] , 
        \wRegOut_7_113[1] , \wRegInTop_5_31[12] , \ScanLink216[7] , 
        \ScanLink97[19] , \wRegInBot_1_1[24] , \wRegOut_2_0[27] , 
        \wRegOut_3_4[31] , \wRegInBot_4_5[16] , \wRegOut_5_3[11] , 
        \wRegOut_6_0[1] , \wRegOut_6_39[18] , \wRegOut_7_0[24] , 
        \wRegOut_7_42[18] , \wRegOut_7_61[30] , \wRegInBot_6_49[0] , 
        \wRegOut_7_14[19] , \wRegOut_7_37[28] , \wRegOut_7_61[29] , 
        \wRegOut_7_37[31] , \ScanLink232[1] , \wRegOut_5_13[30] , 
        \wRegInTop_5_16[12] , \wRegInBot_5_16[15] , \wRegInTop_5_20[17] , 
        \wRegInBot_5_20[10] , \wRegInTop_6_20[3] , \ScanLink93[31] , 
        \ScanLink152[4] , \ScanLink93[28] , \wRegEnTop_7_117[0] , 
        \wRegInBot_5_22[8] , \ScanLink71[9] , \wRegOut_7_4[15] , 
        \wRegOut_6_48[19] , \wRegOut_7_10[31] , \wRegOut_7_33[19] , 
        \ScanLink180[2] , \wRegInTop_7_100[8] , \wRegOut_7_10[28] , 
        \wRegOut_7_46[29] , \wRegOut_7_46[30] , \wRegOut_7_65[18] , 
        \wRegInBot_6_2[12] , \wRegOut_5_13[29] , \wRegOut_5_30[18] , 
        \wRegInTop_6_7[18] , \wRegOut_6_31[8] , \wRegInTop_6_38[12] , 
        \wRegInBot_6_58[11] , \wRegInTop_7_43[12] , \ScanLink183[1] , 
        \wRegOut_7_108[15] , \ScanLink255[31] , \wRegInTop_7_36[22] , 
        \wRegInTop_7_60[23] , \ScanLink203[29] , \ScanLink231[2] , 
        \ScanLink255[28] , \wRegInTop_7_15[13] , \wRegOut_5_3[22] , 
        \wRegInTop_5_15[5] , \ScanLink68[30] , \ScanLink68[29] , 
        \wRegInTop_7_75[17] , \ScanLink203[30] , \ScanLink220[18] , 
        \wRegInTop_6_8[4] , \ScanLink151[7] , \wRegInBot_6_9[2] , 
        \wRegInTop_6_23[0] , \wRegInTop_6_58[16] , \wRegInTop_7_56[26] , 
        \wRegInTop_7_23[16] , \wRegInBot_6_38[15] , \wRegInTop_5_16[21] , 
        \wRegInBot_5_20[23] , \wRegEnBot_6_47[0] , \wRegInTop_6_59[8] , 
        \wRegOut_7_4[26] , \wRegInTop_7_8[31] , \ScanLink148[28] , 
        \wRegInTop_7_8[28] , \ScanLink148[31] , \wRegOut_7_77[9] , 
        \wRegInBot_5_16[26] , \wRegOut_5_19[1] , \wRegInTop_5_20[24] , 
        \wRegInTop_6_44[7] , \ScanLink136[0] , \wRegInTop_7_65[1] , 
        \ScanLink190[18] , \ScanLink255[6] , \wRegInTop_7_75[24] , 
        \wRegInBot_6_38[26] , \wRegInTop_6_58[25] , \wRegEnTop_7_28[0] , 
        \wRegInTop_7_23[25] , \wRegInTop_7_36[11] , \wRegInTop_7_56[15] , 
        \wRegInTop_7_66[2] , \wRegOut_3_4[28] , \wRegInBot_4_5[25] , 
        \wRegInTop_6_38[21] , \wRegInTop_6_47[4] , \wRegInBot_6_58[22] , 
        \ScanLink135[3] , \wRegInTop_7_43[21] , \wRegOut_7_108[26] , 
        \wRegInTop_5_4[20] , \wRegInTop_5_16[6] , \wRegInBot_6_2[21] , 
        \wRegOut_6_48[3] , \wRegInTop_7_15[20] , \wRegInTop_7_60[10] , 
        \wRegOut_7_69[5] , \ScanLink248[9] , \wRegOut_6_36[16] , 
        \wRegEnTop_7_86[0] , \wRegOut_7_38[26] , \wRegOut_6_15[27] , 
        \wRegOut_6_34[5] , \wRegOut_6_43[26] , \wRegOut_7_15[3] , 
        \wRegOut_6_60[17] , \ScanLink4[31] , \ScanLink4[28] , 
        \wRegOut_6_23[22] , \wRegOut_6_56[12] , \wRegOut_7_58[22] , 
        \ScanLink16[26] , \wRegInBot_5_27[5] , \ScanLink77[7] , 
        \ScanLink136[14] , \ScanLink143[24] , \wRegInTop_7_85[30] , 
        \ScanLink63[16] , \ScanLink98[17] , \ScanLink115[25] , 
        \wRegInTop_7_106[6] , \wRegInTop_7_3[24] , \ScanLink160[15] , 
        \wRegInTop_7_85[29] , \ScanLink229[0] , \ScanLink100[11] , 
        \wRegInTop_6_53[30] , \ScanLink123[20] , \ScanLink149[5] , 
        \ScanLink175[21] , \ScanLink156[10] , \wRegInTop_7_28[30] , 
        \ScanLink35[17] , \ScanLink40[27] , \ScanLink74[4] , 
        \wRegInTop_6_53[29] , \wRegInTop_7_28[29] , \wRegInBot_5_24[6] , 
        \wRegInTop_6_26[19] , \wRegInTop_7_105[5] , \ScanLink55[13] , 
        \wRegInTop_6_38[1] , \wRegInTop_7_19[7] , \wEnable_2[0] , 
        \ScanLink208[16] , \ScanLink13[3] , \wRegInBot_3_6[20] , 
        \ScanLink20[23] , \wRegOut_6_0[29] , \wRegOut_5_18[16] , 
        \wRegOut_6_0[30] , \ScanLink76[22] , \wRegOut_6_37[6] , 
        \wRegOut_7_8[6] , \wRegOut_7_16[0] , \wRegOut_7_95[26] , 
        \wRegInTop_7_115[26] , \ScanLink157[9] , \ScanLink198[0] , 
        \wRegInTop_7_123[23] , \wRegInTop_7_100[12] , \wRegInBot_4_13[29] , 
        \wRegOut_7_80[12] , \ScanLink100[22] , \ScanLink175[12] , 
        \wRegInBot_0_0[23] , \ScanLink1[20] , \ScanLink1[13] , \ScanLink2[7] , 
        \wRegInBot_1_1[17] , \wRegOut_2_0[14] , \wRegInBot_4_13[30] , 
        \wRegInTop_5_9[8] , \ScanLink98[24] , \ScanLink123[13] , 
        \ScanLink156[23] , \wRegInTop_7_3[17] , \ScanLink136[27] , 
        \ScanLink143[17] , \ScanLink160[26] , \wRegOut_6_50[1] , 
        \ScanLink115[16] , \wRegOut_7_71[7] , \wRegInTop_3_3[19] , 
        \wRegInBot_3_6[13] , \wRegInBot_5_1[19] , \wRegInTop_5_4[13] , 
        \wRegInBot_6_12[3] , \wRegOut_6_23[11] , \wRegOut_6_56[21] , 
        \wRegInTop_6_42[9] , \wRegOut_6_43[15] , \wRegOut_7_38[15] , 
        \wRegOut_7_58[11] , \wRegOut_6_15[14] , \wRegOut_6_36[25] , 
        \wRegOut_6_60[24] , \wRegInTop_7_123[10] , \wRegOut_5_18[25] , 
        \wRegOut_6_53[2] , \wRegOut_7_72[4] , \ScanLink253[8] , 
        \wRegOut_7_80[21] , \wRegInTop_7_100[21] , \wRegInBot_6_11[0] , 
        \wRegOut_7_95[15] , \wRegInTop_7_115[15] , \ScanLink20[10] , 
        \wRegOut_7_103[19] , \wRegOut_7_120[31] , \wRegOut_2_1[6] , 
        \wRegInBot_2_3[25] , \wRegInBot_3_0[2] , \ScanLink10[0] , 
        \ScanLink16[15] , \wRegInTop_5_10[8] , \ScanLink55[20] , 
        \ScanLink76[11] , \ScanLink208[25] , \wRegOut_7_120[28] , 
        \wRegInBot_6_46[30] , \wRegInBot_5_0[6] , \wRegInTop_5_1[0] , 
        \ScanLink35[24] , \ScanLink63[25] , \wRegInBot_6_10[28] , 
        \wRegInBot_6_46[29] , \ScanLink40[14] , \wRegInBot_6_10[31] , 
        \wRegOut_5_14[4] , \wRegOut_5_24[15] , \wRegInBot_6_33[19] , 
        \wRegInTop_6_6[21] , \wRegOut_6_58[9] , \wRegInTop_3_1[4] , 
        \wRegOut_5_12[10] , \wRegOut_3_5[22] , \wRegInTop_4_1[25] , 
        \wRegOut_5_31[21] , \ScanLink138[6] , \ScanLink217[24] , 
        \ScanLink69[10] , \wRegOut_6_45[6] , \ScanLink191[12] , 
        \wRegOut_7_64[0] , \ScanLink234[15] , \ScanLink241[25] , 
        \ScanLink18[8] , \wRegInBot_5_21[30] , \wRegInBot_6_59[31] , 
        \ScanLink184[26] , \ScanLink221[21] , \wRegInBot_6_59[28] , 
        \ScanLink125[9] , \wRegInTop_7_76[8] , \ScanLink254[11] , 
        \ScanLink202[10] , \wRegInBot_5_21[29] , \ScanLink92[11] , 
        \wRegOut_6_46[5] , \wRegOut_7_67[3] , \wRegInTop_7_9[22] , 
        \wRegOut_5_2[31] , \ScanLink129[26] , \ScanLink149[22] , 
        \wRegInTop_5_18[0] , \ScanLink87[25] , \wRegInBot_2_3[16] , 
        \wRegInTop_3_2[7] , \wRegInBot_3_3[1] , \wRegOut_5_2[28] , 
        \wRegInTop_5_2[3] , \wRegOut_7_64[21] , \wRegInBot_5_3[5] , 
        \wRegOut_5_17[7] , \wRegInBot_6_19[8] , \wRegOut_7_11[11] , 
        \wRegOut_7_47[10] , \wRegOut_6_29[24] , \wRegOut_6_49[20] , 
        \wRegOut_7_32[20] , \wRegInTop_6_49[2] , \wRegOut_7_52[24] , 
        \wRegInTop_7_68[4] , \wRegOut_7_27[14] , \wRegOut_7_71[15] , 
        \wRegOut_3_5[11] , \wRegOut_6_21[2] , \wRegInTop_7_61[29] , 
        \wRegInBot_6_63[0] , \wRegInTop_7_37[31] , \ScanLink221[8] , 
        \ScanLink254[22] , \wRegInTop_4_1[16] , \wRegInTop_6_39[18] , 
        \wRegInTop_7_14[19] , \wRegInTop_7_42[18] , \ScanLink184[15] , 
        \ScanLink221[12] , \wRegInTop_7_61[30] , \wRegInTop_7_37[28] , 
        \ScanLink202[23] , \wRegInBot_4_10[7] , \wRegInBot_4_13[4] , 
        \wRegOut_5_12[23] , \ScanLink69[23] , \ScanLink191[21] , 
        \ScanLink217[17] , \ScanLink241[16] , \ScanLink234[26] , 
        \ScanLink62[0] , \wRegInBot_6_3[18] , \wRegOut_5_24[26] , 
        \wRegOut_5_31[12] , \wRegInTop_7_113[1] , \wRegInTop_6_5[1] , 
        \ScanLink61[3] , \wRegInBot_6_4[7] , \wRegInTop_6_6[12] , 
        \wRegOut_7_27[27] , \wRegInBot_5_31[1] , \wRegOut_6_29[17] , 
        \wRegOut_7_52[17] , \wRegInTop_7_110[2] , \wRegInTop_6_6[2] , 
        \wRegOut_6_49[13] , \wRegOut_7_11[22] , \wRegOut_7_71[26] , 
        \wRegOut_7_32[13] , \wRegOut_7_64[12] , \ScanLink190[8] , 
        \wRegInBot_6_7[4] , \wRegOut_7_47[23] , \ScanLink129[15] , 
        \wRegEnTop_4_13[0] , \wRegOut_6_22[1] , \ScanLink87[16] , 
        \wRegInBot_5_6[8] , \wRegInTop_5_17[18] , \wRegInBot_6_60[3] , 
        \wRegInTop_6_11[25] , \ScanLink92[22] , \wRegInTop_6_30[9] , 
        \wRegInTop_7_9[11] , \ScanLink149[11] , \wRegOut_7_121[22] , 
        \ScanLink5[22] , \ScanLink5[11] , \wRegEnTop_3_2[0] , \wRegOut_4_1[2] , 
        \wRegOut_6_1[10] , \wRegInTop_6_27[20] , \wRegInBot_6_27[27] , 
        \wRegInTop_6_32[14] , \wRegInBot_6_52[17] , \wRegInTop_7_49[14] , 
        \wRegOut_7_102[13] , \wRegInTop_6_47[24] , \wRegInBot_6_32[13] , 
        \wRegInBot_6_47[23] , \wRegOut_7_117[27] , \wRegInTop_6_52[10] , 
        \wRegInTop_7_29[10] , \wRegInTop_3_2[13] , \wRegInBot_3_7[19] , 
        \wRegOut_4_6[14] , \wRegInBot_6_11[22] , \wRegOut_6_43[8] , 
        \ScanLink243[2] , \wRegInBot_6_8[14] , \wRegInTop_6_51[0] , 
        \wRegInTop_7_70[6] , \ScanLink123[7] , \wRegOut_2_2[5] , 
        \wRegInBot_4_12[23] , \wRegInBot_5_0[13] , \ScanLink240[1] , 
        \wRegInTop_5_5[19] , \ScanLink120[4] , \wRegInTop_7_73[5] , 
        \wRegOut_5_11[9] , \wRegInTop_6_52[3] , \ScanLink101[31] , 
        \ScanLink122[19] , \ScanLink157[29] , \wRegOut_5_9[17] , 
        \ScanLink157[30] , \ScanLink174[18] , \wRegInTop_7_91[24] , 
        \wRegInTop_3_2[20] , \wRegInTop_3_4[9] , \wRegOut_4_2[1] , 
        \ScanLink101[28] , \wRegInTop_4_12[24] , \ScanLink79[1] , 
        \wRegInTop_7_84[10] , \ScanLink21[30] , \wRegOut_4_6[27] , 
        \wRegInBot_5_29[3] , \ScanLink227[6] , \wRegInTop_7_108[0] , 
        \wRegOut_7_122[0] , \wRegInTop_7_122[30] , \wRegInBot_6_8[27] , 
        \ScanLink147[3] , \wRegOut_7_81[18] , \wRegInTop_7_101[18] , 
        \wRegInBot_6_11[11] , \wRegInTop_6_27[13] , \wRegInBot_6_32[20] , 
        \wRegInTop_6_35[4] , \wRegInTop_6_52[23] , \wRegOut_7_5[3] , 
        \wRegInTop_7_14[2] , \wRegInTop_7_122[29] , \wRegInTop_7_29[23] , 
        \wRegInBot_6_47[10] , \wRegOut_7_117[14] , \ScanLink77[28] , 
        \ScanLink21[29] , \ScanLink54[19] , \wRegInTop_6_11[16] , 
        \wRegOut_7_121[11] , \ScanLink77[31] , \wRegInBot_6_27[14] , 
        \wRegInTop_6_47[17] , \ScanLink195[5] , \wRegInTop_7_49[27] , 
        \wRegOut_7_102[20] , \wRegInTop_4_12[17] , \wRegOut_6_1[23] , 
        \wRegInBot_6_2[9] , \wRegInTop_6_32[27] , \wRegInBot_6_52[24] , 
        \wRegInBot_4_12[10] , \wRegEnBot_6_4[0] , \wRegOut_6_39[0] , 
        \wRegOut_7_6[0] , \wRegOut_7_18[6] , \wRegInTop_7_84[23] , 
        \ScanLink196[6] , \wRegEnBot_6_35[0] , \wRegInTop_7_91[17] , 
        \wRegInBot_5_0[20] , \wRegOut_5_9[24] , \wRegOut_6_22[31] , 
        \wRegOut_6_22[28] , \wRegInTop_6_36[7] , \ScanLink224[5] , 
        \wRegOut_7_121[3] , \wRegOut_6_57[18] , \ScanLink144[0] , 
        \wRegInTop_7_17[1] , \wRegOut_7_59[28] , \wRegOut_7_59[31] , 
        \wRegInBot_5_13[9] , \wRegInTop_5_18[16] , \wRegInTop_7_80[12] , 
        \ScanLink88[18] , \wRegInBot_5_18[11] , \wRegInTop_7_95[26] , 
        \wRegInTop_6_12[1] , \ScanLink160[6] , \wRegInTop_7_33[7] , 
        \wRegOut_6_26[19] , \wRegOut_6_53[29] , \wRegOut_7_28[29] , 
        \wRegOut_7_105[5] , \wRegOut_6_53[30] , \ScanLink1[4] , 
        \wRegInTop_1_1[15] , \wRegInTop_3_6[11] , \wRegInBot_5_4[11] , 
        \wRegOut_7_28[30] , \ScanLink200[3] , \wRegInTop_6_11[2] , 
        \wRegInTop_7_30[4] , \ScanLink163[5] , \wRegOut_4_2[16] , 
        \wRegInTop_7_105[29] , \wRegOut_6_8[9] , \wRegInBot_6_41[8] , 
        \ScanLink203[0] , \wRegOut_7_85[29] , \wRegOut_7_85[30] , 
        \wRegInTop_7_105[30] , \wRegInTop_7_126[18] , \wRegOut_7_106[6] , 
        \wRegInTop_6_23[22] , \wRegInBot_6_36[11] , \wRegInBot_6_43[21] , 
        \wRegInTop_7_58[22] , \wRegOut_7_113[25] , \wRegInTop_6_56[12] , 
        \ScanLink218[19] , \wRegInBot_6_60[10] , \ScanLink50[31] , 
        \wRegInTop_6_15[27] , \wRegInBot_6_15[20] , \wRegOut_7_125[20] , 
        \ScanLink73[19] , \ScanLink25[18] , \wRegOut_6_5[12] , 
        \wRegInBot_6_56[15] , \wRegInTop_6_60[17] , \wRegInBot_5_4[22] , 
        \ScanLink40[8] , \wRegOut_7_106[11] , \ScanLink50[28] , 
        \wRegInTop_6_36[16] , \wRegInTop_7_38[26] , \wRegEnBot_5_24[0] , 
        \wRegInBot_6_23[25] , \ScanLink104[2] , \wRegInTop_6_43[26] , 
        \wRegInTop_7_57[3] , \wRegInTop_1_1[26] , \wRegInBot_4_8[1] , 
        \wRegInTop_4_9[7] , \wRegOut_4_14[9] , \wRegInTop_5_1[31] , 
        \wRegInTop_5_1[28] , \wRegOut_5_28[0] , \wRegInTop_5_18[25] , 
        \wRegInBot_5_18[22] , \wRegInTop_5_27[7] , \ScanLink126[28] , 
        \wRegInTop_7_85[5] , \ScanLink153[18] , \ScanLink170[30] , 
        \ScanLink105[19] , \wRegInTop_7_95[15] , \ScanLink126[31] , 
        \ScanLink170[29] , \wRegOut_7_58[4] , \wRegInTop_7_80[21] , 
        \wRegInTop_5_24[4] , \wRegOut_6_5[21] , \wRegInTop_6_15[14] , 
        \wRegInTop_6_60[24] , \wRegOut_7_125[13] , \wRegInBot_6_23[16] , 
        \wRegInTop_6_43[15] , \wRegInTop_7_38[15] , \wRegInTop_7_86[6] , 
        \wRegInBot_6_56[26] , \wRegOut_7_106[22] , \wRegInBot_6_15[13] , 
        \wRegInTop_6_23[11] , \wRegInTop_6_36[25] , \wRegInBot_6_36[22] , 
        \wRegInTop_6_56[21] , \wRegInBot_6_43[12] , \wRegInTop_7_58[11] , 
        \wRegOut_7_113[16] , \wRegInBot_3_3[31] , \wRegInBot_3_3[28] , 
        \wRegInBot_6_38[3] , \wRegInBot_6_60[23] , \wRegOut_4_2[25] , 
        \ScanLink107[1] , \wRegInTop_7_54[0] , \wRegInTop_3_6[22] , 
        \ScanLink39[3] , \wRegInTop_7_28[6] , \wRegOut_7_46[8] , 
        \wRegOut_7_89[1] , \wRegOut_7_56[26] , \wRegInBot_0_0[19] , 
        \wRegInBot_0_0[10] , \ScanLink4[9] , \wRegOut_6_58[16] , 
        \wRegOut_7_15[13] , \wRegOut_7_23[16] , \wRegOut_7_60[23] , 
        \wRegOut_7_75[17] , \wRegOut_3_1[20] , \wRegInTop_5_13[30] , 
        \wRegInTop_5_13[29] , \ScanLink45[5] , \wRegInBot_5_15[7] , 
        \wRegOut_6_38[12] , \wRegOut_7_43[12] , \wRegOut_7_36[22] , 
        \wRegEnTop_5_16[0] , \ScanLink83[27] , \ScanLink158[14] , 
        \wRegInTop_7_35[9] , \ScanLink166[8] , \ScanLink96[13] , 
        \wRegInBot_6_44[5] , \wRegOut_7_27[1] , \wRegInTop_5_30[18] , 
        \ScanLink97[3] , \ScanLink138[10] , \wRegInTop_7_10[28] , 
        \ScanLink18[22] , \wRegInTop_4_5[27] , \ScanLink78[26] , 
        \ScanLink94[0] , \wRegInTop_6_48[19] , \wRegInTop_7_10[31] , 
        \wRegInTop_7_46[30] , \ScanLink180[24] , \ScanLink225[23] , 
        \wRegInTop_7_65[18] , \ScanLink250[13] , \wRegInTop_7_33[19] , 
        \ScanLink206[12] , \wRegInTop_7_46[29] , \ScanLink213[26] , 
        \wRegOut_7_100[8] , \wRegOut_7_24[2] , \ScanLink195[10] , 
        \ScanLink230[17] , \ScanLink245[27] , \wRegOut_4_9[30] , 
        \wRegOut_4_9[29] , \wRegOut_5_16[12] , \wRegInBot_6_7[30] , 
        \wRegInBot_6_47[6] , \wRegInBot_6_7[29] , \ScanLink178[4] , 
        \wRegOut_5_6[19] , \wRegOut_5_9[5] , \ScanLink46[6] , 
        \wRegOut_5_20[17] , \wRegInBot_5_16[4] , \wRegInTop_6_2[23] , 
        \ScanLink218[1] , \ScanLink96[20] , \wRegInBot_5_25[18] , 
        \ScanLink138[23] , \ScanLink158[27] , \wRegInTop_5_21[9] , 
        \ScanLink83[14] , \wRegOut_6_62[3] , \wRegInBot_6_20[1] , 
        \wRegOut_7_43[5] , \wRegOut_7_15[20] , \wRegOut_6_38[21] , 
        \wRegOut_7_36[11] , \wRegOut_7_60[10] , \wRegOut_7_43[21] , 
        \wRegOut_6_58[25] , \wRegOut_1_0[3] , \wRegInBot_1_0[27] , 
        \wRegOut_3_1[13] , \ScanLink18[11] , \wRegInTop_4_5[14] , 
        \ScanLink21[1] , \wRegOut_4_12[7] , \wRegOut_7_23[25] , 
        \ScanLink22[2] , \wRegOut_5_16[21] , \wRegOut_5_20[24] , 
        \wRegOut_7_56[15] , \wRegOut_7_75[24] , \wRegOut_7_91[3] , 
        \wRegInTop_7_80[8] , \wRegInTop_6_2[10] , \wRegOut_7_92[0] , 
        \wRegOut_4_11[4] , \wRegOut_5_30[2] , \wRegOut_7_118[29] , 
        \ScanLink213[15] , \ScanLink245[14] , \wRegOut_7_118[30] , 
        \wRegEnTop_4_9[0] , \wRegInBot_6_23[2] , \wRegOut_6_61[0] , 
        \ScanLink195[23] , \ScanLink230[24] , \wRegOut_7_40[6] , 
        \ScanLink250[20] , \wRegInTop_3_2[30] , \wRegInTop_3_2[29] , 
        \wRegInBot_3_7[23] , \wRegOut_5_19[15] , \ScanLink78[15] , 
        \wRegInBot_6_28[30] , \wRegInBot_6_28[29] , \ScanLink180[17] , 
        \ScanLink225[10] , \ScanLink206[21] , \wRegInTop_7_101[11] , 
        \ScanLink79[8] , \ScanLink188[3] , \wRegOut_7_81[11] , 
        \wRegInTop_7_122[20] , \wRegEnTop_7_95[0] , \wRegInTop_7_108[9] , 
        \wRegOut_7_122[9] , \ScanLink54[10] , \ScanLink77[21] , 
        \wRegOut_6_27[5] , \wRegOut_7_94[25] , \wRegInTop_7_114[25] , 
        \wRegOut_7_102[30] , \wRegOut_7_121[18] , \wRegInTop_6_3[6] , 
        \wRegInTop_6_28[2] , \ScanLink209[15] , \wRegInBot_1_0[14] , 
        \wRegOut_2_1[24] , \ScanLink17[25] , \ScanLink21[20] , 
        \wRegOut_7_102[29] , \wRegInBot_4_15[3] , \ScanLink41[24] , 
        \ScanLink64[7] , \wRegInBot_6_2[0] , \wRegInBot_6_32[29] , 
        \ScanLink34[14] , \wRegInTop_7_115[6] , \ScanLink62[15] , 
        \wRegInBot_6_47[19] , \wRegInBot_6_11[18] , \wRegInBot_6_32[30] , 
        \wRegInBot_4_12[19] , \wRegInTop_6_0[5] , \ScanLink122[23] , 
        \ScanLink159[6] , \wRegInBot_6_1[3] , \ScanLink101[12] , 
        \ScanLink157[13] , \wRegInBot_5_0[30] , \ScanLink67[4] , 
        \ScanLink99[14] , \wRegOut_6_39[9] , \ScanLink114[26] , 
        \ScanLink174[22] , \ScanLink239[3] , \wRegInTop_7_2[27] , 
        \ScanLink161[16] , \wRegOut_7_6[9] , \ScanLink137[17] , 
        \ScanLink142[27] , \wRegInTop_7_17[8] , \wRegInTop_7_116[5] , 
        \wRegInBot_5_0[29] , \wRegOut_6_22[21] , \wRegOut_6_57[11] , 
        \ScanLink144[9] , \wRegOut_7_59[21] , \wRegInBot_3_6[5] , 
        \ScanLink34[27] , \wRegInTop_5_5[23] , \wRegOut_6_14[24] , 
        \wRegOut_6_24[6] , \wRegOut_6_37[15] , \wRegOut_6_61[14] , 
        \wRegOut_6_42[25] , \wRegOut_7_39[25] , \wRegInTop_6_27[29] , 
        \ScanLink41[17] , \wRegInTop_6_52[19] , \wRegInTop_7_29[19] , 
        \wRegInTop_3_7[3] , \ScanLink17[16] , \wRegInTop_6_27[30] , 
        \ScanLink21[13] , \wRegInBot_5_6[1] , \wRegInTop_5_7[7] , 
        \ScanLink62[26] , \ScanLink77[12] , \wRegOut_5_12[3] , 
        \wRegOut_6_1[19] , \wRegOut_2_1[17] , \ScanLink5[18] , 
        \wRegInBot_3_7[10] , \ScanLink54[23] , \wRegInTop_6_51[9] , 
        \ScanLink209[26] , \wRegOut_7_62[7] , \wRegOut_7_94[16] , 
        \wRegInTop_7_114[16] , \wRegInTop_5_5[10] , \wRegOut_5_19[26] , 
        \wRegOut_6_43[1] , \wRegOut_7_81[22] , \wRegInTop_7_101[22] , 
        \wRegOut_6_14[17] , \wRegOut_6_61[27] , \wRegInTop_7_122[13] , 
        \wRegOut_7_39[16] , \wRegOut_6_22[12] , \wRegOut_6_37[26] , 
        \wRegOut_6_42[16] , \wRegOut_6_57[22] , \wRegOut_7_59[12] , 
        \wRegOut_6_40[2] , \wRegOut_7_61[4] , \ScanLink240[8] , 
        \wRegInTop_3_4[0] , \wRegInBot_3_5[6] , \wRegOut_4_2[8] , 
        \ScanLink161[25] , \ScanLink99[27] , \wRegInTop_7_2[14] , 
        \wRegOut_3_5[18] , \wRegInTop_5_4[4] , \wRegOut_5_11[0] , 
        \ScanLink114[15] , \ScanLink137[24] , \ScanLink142[14] , 
        \wRegInTop_7_84[19] , \ScanLink157[20] , \ScanLink122[10] , 
        \wRegInBot_5_5[2] , \ScanLink174[11] , \wRegInTop_6_33[3] , 
        \ScanLink101[21] , \ScanLink141[4] , \wRegInBot_6_39[16] , 
        \wRegInTop_6_59[15] , \wRegInTop_7_12[5] , \wRegInTop_7_57[25] , 
        \ScanLink191[31] , \wRegInTop_7_22[15] , \wRegInTop_7_61[20] , 
        \ScanLink191[28] , \wRegInTop_7_74[14] , \wRegEnTop_7_104[0] , 
        \ScanLink221[1] , \wRegInBot_4_4[15] , \ScanLink62[9] , 
        \wRegInTop_6_5[8] , \wRegInTop_6_39[11] , \wRegInBot_6_59[12] , 
        \wRegInBot_6_63[9] , \wRegInTop_7_14[10] , \wRegInTop_7_42[11] , 
        \wRegOut_7_109[16] , \wRegInTop_7_37[21] , \wRegOut_7_124[7] , 
        \wRegOut_7_3[4] , \ScanLink193[2] , \wRegInBot_6_3[11] , 
        \wRegInTop_7_113[8] , \ScanLink190[1] , \wRegInTop_2_2[17] , 
        \wRegInBot_3_3[8] , \ScanLink18[1] , \wRegInBot_4_4[26] , 
        \wRegOut_4_7[5] , \wRegOut_5_2[12] , \wRegInTop_5_17[11] , 
        \wRegInBot_5_31[8] , \wRegOut_7_0[7] , \wRegOut_7_5[16] , 
        \wRegInTop_7_9[18] , \wRegInTop_5_21[14] , \wRegInBot_5_21[13] , 
        \wRegInTop_6_30[0] , \wRegInTop_7_11[6] , \ScanLink142[7] , 
        \ScanLink149[18] , \ScanLink222[2] , \wRegOut_7_127[4] , 
        \wRegInBot_5_17[16] , \wRegOut_6_22[8] , \wRegInTop_5_1[9] , 
        \wRegOut_5_12[19] , \wRegOut_5_31[31] , \wRegOut_5_31[28] , 
        \wRegInBot_6_3[22] , \wRegEnBot_6_54[0] , \wRegInTop_6_6[31] , 
        \wRegOut_7_79[6] , \wRegInTop_6_6[28] , \wRegOut_6_58[0] , 
        \wRegInTop_7_14[23] , \wRegOut_5_2[21] , \wRegInBot_5_17[25] , 
        \wRegInTop_5_18[9] , \wRegInTop_5_21[27] , \ScanLink69[19] , 
        \wRegInTop_6_39[22] , \wRegInTop_6_57[7] , \wRegInTop_7_37[12] , 
        \wRegInTop_7_61[13] , \ScanLink221[28] , \wRegInTop_7_76[1] , 
        \ScanLink254[18] , \wRegInBot_6_59[21] , \ScanLink125[0] , 
        \ScanLink202[19] , \ScanLink221[31] , \wRegInTop_7_42[22] , 
        \wRegOut_7_109[25] , \wRegInBot_6_39[25] , \wRegInTop_6_59[26] , 
        \wRegInTop_7_22[26] , \wRegInTop_7_57[16] , \wRegOut_7_64[9] , 
        \ScanLink245[5] , \wRegInTop_6_54[4] , \ScanLink126[3] , 
        \wRegInTop_7_74[27] , \wRegInTop_7_75[2] , \wRegInTop_5_17[22] , 
        \ScanLink92[18] , \ScanLink246[6] , \wRegInBot_5_21[20] , 
        \wRegOut_7_5[25] , \wRegOut_4_4[6] , \wRegOut_5_6[10] , 
        \wRegEnTop_5_7[0] , \wRegInTop_5_25[16] , \wRegInBot_6_19[1] , 
        \wRegOut_7_11[18] , \wRegOut_7_64[28] , \wRegOut_6_49[30] , 
        \wRegOut_7_32[30] , \wRegOut_6_49[29] , \wRegOut_7_32[29] , 
        \wRegOut_7_47[19] , \wRegOut_7_64[31] , \wRegInBot_5_30[25] , 
        \wRegInTop_5_13[13] , \wRegInBot_5_13[14] , \wRegInBot_6_20[8] , 
        \wRegInBot_5_25[11] , \wRegInTop_5_30[22] , \ScanLink96[29] , 
        \ScanLink102[5] , \wRegInTop_7_51[4] , \ScanLink96[30] , 
        \wRegOut_7_1[14] , \ScanLink4[0] , \wRegInBot_4_0[17] , 
        \ScanLink21[8] , \wRegOut_4_9[13] , \wRegInTop_5_21[0] , 
        \wRegOut_6_38[31] , \wRegOut_7_15[29] , \wRegOut_7_43[31] , 
        \wRegOut_7_60[19] , \wRegOut_6_38[28] , \wRegOut_7_15[30] , 
        \wRegOut_7_36[18] , \wRegOut_7_43[28] , \wRegInTop_7_83[2] , 
        \wRegOut_5_16[31] , \wRegOut_5_16[28] , \wRegOut_7_92[9] , 
        \wRegInBot_6_7[13] , \wRegInTop_5_22[3] , \wRegInTop_7_80[1] , 
        \wRegInTop_6_2[19] , \wRegOut_6_61[9] , \wRegInTop_7_65[22] , 
        \ScanLink250[29] , \ScanLink18[18] , \wRegInTop_6_28[27] , 
        \wRegInBot_6_28[20] , \wRegInTop_7_10[12] , \wRegInTop_7_46[13] , 
        \ScanLink206[31] , \ScanLink225[19] , \ScanLink250[30] , 
        \ScanLink101[6] , \wRegInTop_6_48[23] , \wRegInTop_7_33[23] , 
        \ScanLink206[28] , \wRegInBot_6_48[24] , \wRegInTop_7_26[17] , 
        \wRegInTop_7_52[7] , \wRegInTop_7_53[27] , \wRegOut_7_118[20] , 
        \wRegInTop_7_70[16] , \wRegInBot_6_59[3] , \ScanLink1[30] , 
        \wRegInTop_2_2[24] , \wRegInTop_5_13[20] , \wRegOut_7_1[27] , 
        \wRegOut_7_27[8] , \ScanLink206[4] , \wRegInBot_5_25[22] , 
        \ScanLink58[3] , \ScanLink138[19] , \ScanLink7[3] , \wRegOut_3_1[30] , 
        \wRegOut_3_1[29] , \wRegInBot_4_0[24] , \wRegOut_5_6[23] , 
        \wRegInBot_5_13[27] , \wRegInTop_5_25[25] , \wRegInTop_5_30[11] , 
        \wRegOut_7_103[2] , \wRegInBot_5_30[16] , \wRegInTop_7_35[0] , 
        \ScanLink166[1] , \wRegInTop_6_14[6] , \wRegInTop_6_28[14] , 
        \ScanLink94[9] , \wRegInTop_7_26[24] , \wRegInBot_6_48[17] , 
        \wRegInTop_7_53[14] , \wRegOut_7_100[1] , \wRegOut_7_118[13] , 
        \wRegInTop_7_10[21] , \ScanLink195[19] , \wRegInTop_7_70[25] , 
        \ScanLink205[7] , \wRegInTop_6_17[5] , \wRegInTop_7_33[10] , 
        \wRegInTop_7_65[11] , \wRegInTop_7_36[3] , \wRegInBot_6_28[13] , 
        \wRegOut_6_18[2] , \ScanLink89[6] , \wRegInTop_6_48[10] , 
        \wRegInTop_7_8[2] , \ScanLink165[2] , \wRegInTop_7_46[20] , 
        \wRegOut_7_39[4] , \ScanLink218[8] , \wRegInBot_4_8[8] , 
        \wRegOut_4_9[20] , \wRegInBot_6_7[20] , \wRegOut_7_45[2] , 
        \wRegInTop_5_1[21] , \wRegOut_5_28[9] , \wRegOut_6_10[26] , 
        \wRegInBot_6_26[6] , \wRegOut_7_48[17] , \wRegOut_6_33[17] , 
        \wRegOut_6_46[27] , \wRegOut_6_26[23] , \wRegOut_6_53[13] , 
        \wRegInTop_7_98[3] , \ScanLink1[29] , \wRegOut_7_28[13] , 
        \wRegInTop_1_0[16] , \wRegInBot_2_0[4] , \wRegInTop_2_1[2] , 
        \wRegOut_3_0[23] , \wRegInBot_3_3[21] , \ScanLink13[27] , 
        \ScanLink24[5] , \ScanLink27[6] , \wRegOut_4_14[0] , \ScanLink110[24] , 
        \ScanLink133[15] , \wRegInTop_7_6[25] , \ScanLink165[14] , 
        \wRegInTop_7_80[28] , \wRegOut_7_97[4] , \wRegInTop_7_80[31] , 
        \ScanLink88[22] , \ScanLink105[10] , \ScanLink119[4] , 
        \ScanLink126[21] , \ScanLink146[25] , \ScanLink153[11] , 
        \ScanLink170[20] , \ScanLink218[23] , \ScanLink30[16] , 
        \ScanLink45[26] , \wRegInTop_6_56[28] , \wRegInTop_6_23[18] , 
        \wRegInTop_7_58[18] , \ScanLink66[17] , \wRegInTop_6_56[31] , 
        \wRegOut_7_94[7] , \ScanLink25[22] , \ScanLink50[12] , 
        \wRegOut_6_5[31] , \ScanLink73[23] , \wRegOut_6_5[28] , 
        \wRegInTop_7_49[6] , \wRegOut_4_13[27] , \wRegInTop_6_9[26] , 
        \wRegInBot_6_25[5] , \wRegOut_7_46[1] , \wRegOut_7_89[8] , 
        \wRegOut_7_90[27] , \wRegInTop_7_110[27] , \wRegInTop_7_105[13] , 
        \wRegInBot_3_3[12] , \wRegInTop_5_1[12] , \wRegInBot_5_4[18] , 
        \ScanLink43[2] , \ScanLink107[8] , \wRegOut_7_85[13] , 
        \wRegInTop_7_54[9] , \wRegInTop_7_126[22] , \wRegInBot_5_13[0] , 
        \ScanLink153[22] , \wRegOut_7_118[3] , \wRegInBot_5_18[18] , 
        \ScanLink88[11] , \ScanLink126[12] , \ScanLink170[13] , 
        \wRegOut_6_26[10] , \ScanLink91[4] , \ScanLink105[23] , 
        \ScanLink110[17] , \wRegInTop_7_6[16] , \ScanLink165[27] , 
        \wRegOut_6_53[20] , \ScanLink133[26] , \ScanLink146[16] , 
        \wRegOut_7_28[20] , \wRegInBot_6_42[2] , \wRegOut_7_21[6] , 
        \wRegOut_6_10[15] , \wRegInTop_6_12[8] , \wRegOut_6_33[24] , 
        \wRegOut_6_46[14] , \wRegOut_7_48[24] , \wRegOut_7_22[5] , 
        \ScanLink203[9] , \ScanLink13[14] , \wRegInTop_3_6[18] , 
        \wRegOut_4_13[14] , \wRegOut_6_8[0] , \ScanLink92[7] , 
        \wRegInBot_6_41[1] , \wRegOut_7_85[20] , \wRegInTop_7_105[20] , 
        \wRegInTop_7_126[11] , \ScanLink25[11] , \wRegInTop_6_9[15] , 
        \wRegOut_7_90[14] , \ScanLink73[10] , \wRegInTop_7_110[14] , 
        \wRegOut_7_125[29] , \ScanLink30[25] , \ScanLink40[1] , 
        \wRegEnTop_7_63[0] , \wRegOut_7_106[18] , \wRegOut_7_125[30] , 
        \wRegInBot_5_10[3] , \ScanLink50[21] , \wRegInBot_6_43[28] , 
        \ScanLink45[15] , \ScanLink218[10] , \wRegInBot_6_15[30] , 
        \wRegInBot_6_36[18] , \ScanLink19[21] , \wRegOut_5_17[11] , 
        \wRegOut_5_21[14] , \ScanLink66[24] , \wRegInBot_6_15[29] , 
        \wRegInBot_6_43[31] , \wRegInBot_6_60[19] , \wRegInTop_6_3[20] , 
        \ScanLink208[2] , \ScanLink56[5] , \wRegInTop_7_5[7] , 
        \ScanLink168[7] , \wRegInTop_7_127[4] , \wRegOut_6_15[7] , 
        \wRegOut_7_34[1] , \ScanLink194[13] , \ScanLink231[14] , 
        \ScanLink244[24] , \wRegInTop_4_4[24] , \ScanLink84[3] , 
        \wRegInBot_6_57[5] , \ScanLink212[25] , \wRegOut_7_119[19] , 
        \wRegInBot_6_29[19] , \wRegInTop_7_26[9] , \ScanLink175[8] , 
        \ScanLink207[11] , \wRegOut_3_0[10] , \ScanLink9[5] , \ScanLink48[9] , 
        \wRegInBot_5_24[28] , \ScanLink79[25] , \ScanLink181[27] , 
        \ScanLink224[20] , \ScanLink251[10] , \ScanLink139[13] , 
        \wRegInBot_5_24[31] , \ScanLink87[0] , \wRegOut_7_113[8] , 
        \wRegOut_6_16[4] , \wRegOut_7_37[2] , \wRegOut_5_7[30] , 
        \wRegOut_5_7[29] , \ScanLink82[24] , \ScanLink97[10] , 
        \wRegInBot_6_54[6] , \ScanLink55[6] , \ScanLink159[17] , 
        \wRegOut_6_0[8] , \wRegOut_6_39[11] , \wRegOut_7_42[11] , 
        \wRegOut_7_37[21] , \wRegInTop_7_124[7] , \wRegInTop_6_19[3] , 
        \wRegInBot_6_49[9] , \wRegOut_7_61[20] , \wRegOut_7_14[10] , 
        \wRegInTop_7_38[5] , \wRegOut_7_57[25] , \wRegOut_7_74[14] , 
        \wRegInBot_6_33[1] , \wRegInTop_6_49[29] , \wRegOut_6_59[15] , 
        \wRegInTop_7_6[4] , \wRegOut_7_22[15] , \wRegInTop_7_32[29] , 
        \wRegInTop_7_47[19] , \wRegInTop_7_64[31] , \wRegOut_7_50[5] , 
        \wRegInTop_7_64[28] , \ScanLink207[22] , \ScanLink251[23] , 
        \wRegInTop_7_11[18] , \wRegInTop_7_32[30] , \wRegInBot_4_0[0] , 
        \ScanLink19[12] , \ScanLink79[16] , \wRegInTop_6_49[30] , 
        \ScanLink181[14] , \ScanLink224[13] , \ScanLink244[17] , 
        \wRegInTop_4_4[17] , \ScanLink194[20] , \ScanLink231[27] , 
        \ScanLink32[1] , \ScanLink212[16] , \wRegOut_5_20[1] , 
        \wRegEnTop_7_11[0] , \wRegInBot_6_6[19] , \wRegInTop_4_1[6] , 
        \wRegOut_4_8[19] , \wRegOut_7_82[3] , \wRegOut_5_17[22] , 
        \wRegInTop_6_3[13] , \wRegInTop_2_2[1] , \wRegInTop_4_2[5] , 
        \wRegInBot_4_3[3] , \wRegOut_5_21[27] , \wRegOut_7_81[0] , 
        \ScanLink31[2] , \wRegOut_5_23[2] , \wRegOut_7_74[27] , 
        \wRegOut_6_59[26] , \wRegOut_7_22[26] , \wRegOut_6_39[22] , 
        \wRegOut_7_37[12] , \wRegOut_7_57[16] , \wRegOut_7_42[22] , 
        \wRegInTop_7_93[8] , \wRegOut_7_14[23] , \wRegInBot_2_3[7] , 
        \wRegOut_5_4[9] , \wRegInTop_5_12[19] , \wRegInTop_5_31[28] , 
        \ScanLink82[17] , \wRegOut_7_61[13] , \wRegInBot_6_30[2] , 
        \wRegOut_7_53[6] , \wRegInTop_6_60[8] , \ScanLink159[24] , 
        \ScanLink97[23] , \ScanLink139[20] , \wRegInTop_5_31[31] , 
        \wRegOut_6_4[11] , \wRegInBot_6_57[16] , \wRegOut_6_5[5] , 
        \wRegInBot_6_22[26] , \wRegInTop_6_37[15] , \wRegOut_7_107[12] , 
        \wRegInTop_7_39[25] , \wRegInTop_6_42[25] , \wRegInTop_6_14[24] , 
        \wRegOut_7_124[23] , \wRegInBot_6_14[23] , \wRegInTop_6_61[14] , 
        \wRegInBot_6_61[13] , \wRegInBot_3_2[18] , \wRegOut_4_3[15] , 
        \wRegOut_6_13[9] , \wRegInTop_6_22[21] , \wRegInBot_6_37[12] , 
        \wRegInBot_6_42[22] , \wRegInTop_7_59[21] , \wRegOut_7_112[26] , 
        \wRegInTop_6_57[11] , \wRegInTop_7_3[9] , \wRegOut_7_116[5] , 
        \ScanLink213[3] , \ScanLink0[10] , \wRegInTop_3_7[12] , 
        \wRegInTop_7_20[7] , \ScanLink173[6] , \wRegInBot_1_1[8] , 
        \wRegInTop_5_0[18] , \wRegInBot_5_5[12] , \ScanLink210[0] , 
        \wRegInBot_6_52[8] , \wRegInTop_7_23[4] , \ScanLink170[5] , 
        \wRegOut_7_115[6] , \wRegInBot_5_19[12] , \ScanLink104[29] , 
        \ScanLink152[31] , \ScanLink171[19] , \wRegInTop_7_94[25] , 
        \ScanLink53[8] , \wRegOut_6_6[6] , \ScanLink152[28] , 
        \wRegInTop_5_19[15] , \ScanLink104[30] , \ScanLink127[18] , 
        \wRegOut_7_108[9] , \wRegInTop_7_122[9] , \wRegEnTop_7_5[0] , 
        \wRegInTop_7_81[11] , \wRegInBot_0_0[27] , \ScanLink0[23] , 
        \wRegInTop_1_0[25] , \wRegOut_3_1[0] , \wRegInTop_3_7[21] , 
        \ScanLink29[0] , \wRegOut_7_99[2] , \wRegOut_4_3[26] , 
        \wRegInTop_5_29[8] , \ScanLink117[2] , \wRegInTop_7_44[3] , 
        \wRegInTop_7_127[28] , \wRegOut_7_84[19] , \wRegInTop_7_104[19] , 
        \wRegInTop_7_127[31] , \ScanLink219[30] , \wRegEnBot_2_3[0] , 
        \wRegInTop_4_7[8] , \wRegInBot_6_14[10] , \wRegInBot_6_28[0] , 
        \ScanLink24[28] , \ScanLink51[18] , \ScanLink72[30] , 
        \wRegInTop_6_22[12] , \wRegInBot_6_37[21] , \wRegInTop_6_57[22] , 
        \wRegInBot_6_61[20] , \ScanLink219[29] , \wRegInBot_6_42[11] , 
        \wRegInTop_7_59[12] , \wRegOut_7_112[15] , \wRegInBot_6_22[15] , 
        \wRegInTop_7_39[16] , \wRegInTop_7_96[5] , \wRegInTop_6_42[16] , 
        \wRegInTop_4_15[1] , \wRegOut_6_4[22] , \wRegInBot_6_57[25] , 
        \wRegOut_7_107[21] , \ScanLink72[29] , \wRegInTop_6_37[26] , 
        \wRegInTop_6_61[27] , \wRegOut_3_2[3] , \ScanLink24[31] , 
        \wRegOut_5_1[4] , \wRegInTop_6_14[17] , \wRegOut_7_124[10] , 
        \wRegOut_7_48[7] , \wRegInTop_7_81[22] , \wRegOut_5_2[7] , 
        \wRegInTop_5_19[26] , \wRegInBot_5_19[21] , \wRegInTop_7_94[16] , 
        \ScanLink89[28] , \wRegInBot_5_5[21] , \ScanLink89[31] , 
        \wRegInTop_7_95[6] , \wRegOut_6_27[30] , \wRegOut_7_55[8] , 
        \ScanLink4[21] , \ScanLink4[12] , \wRegInTop_4_13[27] , 
        \wRegInTop_5_13[2] , \wRegOut_6_27[29] , \ScanLink114[1] , 
        \wRegInTop_7_47[0] , \wRegOut_6_52[19] , \wRegInTop_7_88[9] , 
        \wRegOut_7_29[19] , \wRegInBot_4_13[20] , \wRegInTop_7_85[13] , 
        \wRegOut_5_8[14] , \wRegInTop_6_42[0] , \ScanLink130[7] , 
        \wRegInTop_7_90[27] , \wRegInTop_7_63[6] , \wRegOut_6_56[31] , 
        \ScanLink10[9] , \wRegInTop_3_3[10] , \wRegInBot_5_1[10] , 
        \wRegInTop_5_9[1] , \wRegOut_6_50[8] , \ScanLink250[2] , 
        \wRegInBot_5_8[7] , \wRegOut_6_23[18] , \wRegOut_6_56[28] , 
        \wRegInTop_6_41[3] , \wRegOut_7_58[18] , \wRegInTop_7_60[5] , 
        \ScanLink133[4] , \ScanLink20[19] , \wRegOut_4_7[17] , 
        \wRegInBot_6_9[17] , \wRegOut_7_80[31] , \wRegInTop_7_100[31] , 
        \wRegInTop_7_123[19] , \wRegInTop_7_100[28] , \ScanLink253[1] , 
        \wRegInTop_5_10[1] , \wRegInBot_6_11[9] , \wRegOut_7_80[28] , 
        \wRegOut_6_0[13] , \wRegInBot_6_10[21] , \wRegInTop_6_26[23] , 
        \wRegInBot_6_33[10] , \wRegInBot_6_46[20] , \wRegOut_7_116[24] , 
        \wRegInTop_6_53[13] , \wRegInTop_7_28[13] , \wRegInBot_6_53[14] , 
        \wRegInTop_7_48[17] , \wRegOut_7_103[10] , \wRegInTop_6_33[17] , 
        \wRegInBot_5_1[23] , \ScanLink55[30] , \ScanLink55[29] , 
        \wRegInTop_6_10[26] , \wRegInBot_6_26[24] , \wRegInTop_6_46[27] , 
        \wRegOut_7_120[21] , \ScanLink76[18] , \wRegInTop_2_2[30] , 
        \wRegInTop_2_2[29] , \wRegInBot_2_2[26] , \wRegInTop_3_3[23] , 
        \wRegInBot_3_6[30] , \wRegInTop_4_13[14] , \wRegInBot_4_13[13] , 
        \wRegInTop_5_4[30] , \wRegInTop_5_4[29] , \wRegInTop_6_26[4] , 
        \ScanLink154[3] , \wRegEnTop_7_49[0] , \ScanLink234[6] , 
        \ScanLink100[18] , \wRegInTop_7_90[14] , \ScanLink123[30] , 
        \wRegOut_5_8[27] , \ScanLink123[29] , \ScanLink175[28] , 
        \ScanLink186[5] , \ScanLink156[19] , \ScanLink175[31] , 
        \wRegOut_6_0[20] , \wRegInBot_6_26[17] , \wRegOut_6_29[3] , 
        \wRegInTop_7_85[20] , \ScanLink229[9] , \wRegInTop_6_38[8] , 
        \ScanLink185[6] , \wRegInTop_6_46[14] , \wRegInTop_7_48[24] , 
        \wRegOut_7_103[23] , \wRegInBot_6_9[24] , \wRegInTop_6_10[15] , 
        \wRegEnBot_6_26[0] , \wRegInTop_6_33[24] , \wRegInBot_6_53[27] , 
        \wRegOut_7_120[12] , \wRegInBot_6_10[12] , \wRegInTop_6_26[10] , 
        \wRegInBot_6_33[23] , \wRegInTop_6_53[20] , \wRegInTop_7_28[20] , 
        \wRegInBot_6_46[13] , \ScanLink157[0] , \wRegOut_7_116[17] , 
        \wRegInTop_6_25[7] , \ScanLink198[9] , \wRegInBot_3_6[29] , 
        \wRegOut_4_7[24] , \ScanLink69[2] , \wRegOut_7_16[9] , 
        \ScanLink237[5] , \ScanLink15[4] , \wRegOut_6_28[27] , 
        \wRegOut_7_70[16] , \wRegInTop_7_118[3] , \wRegInTop_6_59[1] , 
        \wRegOut_7_53[27] , \wRegInTop_7_78[7] , \wRegOut_7_26[17] , 
        \wRegOut_4_9[3] , \wRegOut_6_48[23] , \wRegOut_7_33[23] , 
        \wRegOut_7_46[13] , \wRegOut_7_10[12] , \wRegOut_7_65[22] , 
        \ScanLink86[26] , \wRegInBot_2_2[15] , \wRegOut_3_4[21] , 
        \wRegInTop_5_16[31] , \ScanLink128[25] , \ScanLink136[9] , 
        \wRegInTop_7_65[8] , \ScanLink148[21] , \wRegInTop_5_16[28] , 
        \wRegInBot_6_14[4] , \wRegOut_6_56[6] , \wRegOut_7_77[0] , 
        \ScanLink93[12] , \wRegInTop_6_38[28] , \wRegInTop_7_8[21] , 
        \wRegInTop_7_15[30] , \wRegInTop_7_36[18] , \wRegInTop_7_43[28] , 
        \ScanLink203[13] , \wRegInTop_4_0[26] , \wRegEnBot_5_8[0] , 
        \ScanLink68[13] , \wRegInTop_6_38[31] , \wRegInTop_7_15[29] , 
        \wRegInTop_7_43[31] , \ScanLink185[25] , \ScanLink220[22] , 
        \wRegInTop_7_60[19] , \wRegOut_6_55[5] , \ScanLink190[11] , 
        \wRegOut_7_74[3] , \ScanLink235[16] , \ScanLink255[12] , 
        \wRegOut_5_19[8] , \wRegInBot_6_17[7] , \ScanLink240[26] , 
        \ScanLink216[27] , \ScanLink16[7] , \wRegOut_5_13[13] , 
        \wRegOut_5_30[22] , \wRegInBot_6_2[28] , \ScanLink128[5] , 
        \wRegInBot_6_2[31] , \wRegOut_5_25[16] , \wRegInTop_6_7[22] , 
        \ScanLink248[0] , \wRegOut_5_3[18] , \wRegInBot_5_20[19] , 
        \wRegEnTop_6_14[0] , \ScanLink148[12] , \ScanLink93[21] , 
        \wRegOut_6_32[2] , \wRegInTop_7_8[12] , \wRegOut_3_1[24] , 
        \wRegOut_3_4[12] , \wRegInTop_4_0[15] , \wRegOut_5_13[20] , 
        \wRegInBot_5_21[2] , \ScanLink71[0] , \ScanLink86[15] , 
        \wRegOut_7_13[4] , \wRegOut_6_48[10] , \ScanLink128[16] , 
        \ScanLink232[8] , \wRegOut_7_33[10] , \wRegOut_7_10[21] , 
        \wRegOut_7_46[20] , \wRegOut_7_26[24] , \wRegOut_7_65[11] , 
        \wRegOut_7_70[25] , \wRegOut_6_28[14] , \wRegInBot_5_22[1] , 
        \wRegOut_5_25[25] , \wRegInTop_6_7[11] , \wRegOut_7_53[14] , 
        \wRegInTop_7_100[1] , \ScanLink183[8] , \ScanLink72[3] , 
        \wRegOut_5_30[11] , \wRegInTop_7_103[2] , \ScanLink68[20] , 
        \ScanLink190[22] , \ScanLink235[25] , \ScanLink240[15] , 
        \wRegInTop_6_23[9] , \wRegOut_6_31[1] , \wRegInBot_6_58[18] , 
        \ScanLink216[14] , \ScanLink203[20] , \wRegOut_7_10[7] , 
        \ScanLink255[21] , \wRegInBot_4_0[30] , \ScanLink18[26] , 
        \ScanLink46[2] , \wRegOut_5_20[13] , \wRegInTop_6_2[27] , 
        \wRegOut_7_39[9] , \ScanLink185[16] , \ScanLink220[11] , 
        \ScanLink218[5] , \wRegOut_5_16[16] , \wRegInBot_5_16[0] , 
        \ScanLink178[0] , \wRegOut_7_24[6] , \ScanLink195[14] , 
        \ScanLink230[13] , \wRegInTop_7_26[30] , \wRegInTop_7_70[28] , 
        \ScanLink245[23] , \wRegInTop_4_5[23] , \wRegInTop_6_28[19] , 
        \ScanLink94[4] , \wRegInBot_6_47[2] , \wRegInTop_7_26[29] , 
        \ScanLink213[22] , \wRegInTop_7_70[31] , \wRegInTop_7_53[19] , 
        \wRegInBot_4_0[29] , \ScanLink78[22] , \wRegInTop_6_17[8] , 
        \ScanLink206[16] , \ScanLink97[7] , \ScanLink138[14] , 
        \ScanLink180[20] , \ScanLink225[27] , \ScanLink250[17] , 
        \wRegOut_7_27[5] , \ScanLink206[9] , \ScanLink45[1] , 
        \wRegInTop_5_25[31] , \ScanLink83[23] , \ScanLink96[17] , 
        \wRegInBot_6_44[1] , \wRegInTop_5_25[28] , \ScanLink158[10] , 
        \wRegEnTop_7_66[0] , \wRegInBot_5_15[3] , \wRegOut_6_38[16] , 
        \wRegOut_7_43[16] , \wRegOut_7_36[26] , \wRegOut_7_15[17] , 
        \wRegOut_7_60[27] , \wRegInTop_7_28[2] , \wRegOut_7_75[13] , 
        \wRegOut_7_56[22] , \wRegInBot_0_0[14] , \wRegOut_3_1[17] , 
        \ScanLink78[11] , \wRegInBot_6_23[6] , \wRegOut_6_58[12] , 
        \wRegOut_6_61[4] , \wRegOut_7_23[12] , \ScanLink206[25] , 
        \wRegOut_7_40[2] , \ScanLink250[24] , \ScanLink18[15] , 
        \wRegInBot_6_48[30] , \ScanLink180[13] , \ScanLink225[14] , 
        \ScanLink245[10] , \wRegInTop_4_5[10] , \ScanLink195[27] , 
        \ScanLink230[20] , \ScanLink22[6] , \wRegInBot_6_48[29] , 
        \ScanLink213[11] , \wRegOut_4_11[0] , \wRegOut_5_30[6] , 
        \wRegOut_4_12[3] , \wRegOut_5_16[25] , \wRegOut_7_92[4] , 
        \wRegOut_5_20[20] , \wRegInTop_6_2[14] , \wRegOut_6_58[21] , 
        \wRegOut_7_75[20] , \wRegOut_7_91[7] , \wRegOut_7_1[19] , 
        \ScanLink1[24] , \ScanLink1[17] , \ScanLink1[0] , \ScanLink21[5] , 
        \wRegOut_7_23[21] , \wRegOut_5_9[1] , \wRegInBot_5_13[19] , 
        \wRegInBot_5_30[31] , \ScanLink83[10] , \wRegOut_6_38[25] , 
        \wRegOut_7_36[15] , \wRegOut_7_56[11] , \wRegOut_7_43[25] , 
        \wRegOut_6_62[7] , \wRegOut_7_15[24] , \wRegOut_7_60[14] , 
        \wRegOut_7_43[1] , \wRegInBot_6_20[5] , \wRegInBot_5_30[28] , 
        \ScanLink158[23] , \ScanLink96[24] , \ScanLink102[8] , 
        \wRegInTop_7_51[9] , \ScanLink138[27] , \wRegOut_6_5[16] , 
        \wRegInTop_6_15[23] , \wRegInBot_6_23[21] , \wRegInTop_6_36[12] , 
        \wRegInBot_6_56[11] , \wRegOut_7_106[15] , \wRegInTop_7_38[22] , 
        \wRegInTop_6_43[22] , \wRegOut_7_125[24] , \wRegInTop_1_1[11] , 
        \ScanLink13[19] , \ScanLink30[31] , \wRegInTop_6_60[13] , 
        \wRegInBot_6_60[14] , \ScanLink66[29] , \wRegInBot_6_15[24] , 
        \wRegInTop_3_6[15] , \wRegOut_4_2[12] , \wRegOut_4_13[19] , 
        \ScanLink30[28] , \wRegInTop_6_23[26] , \wRegInTop_7_58[26] , 
        \ScanLink45[18] , \ScanLink66[30] , \wRegInBot_6_36[15] , 
        \wRegInBot_6_43[25] , \wRegOut_7_113[21] , \wRegInTop_6_56[16] , 
        \wRegOut_7_106[2] , \ScanLink203[4] , \wRegInTop_6_9[18] , 
        \wRegOut_7_22[8] , \wRegOut_7_90[19] , \wRegInTop_6_11[6] , 
        \wRegInTop_7_30[0] , \wRegInTop_7_110[19] , \ScanLink163[1] , 
        \ScanLink2[3] , \wRegInBot_5_4[15] , \ScanLink200[7] , 
        \wRegOut_6_10[18] , \wRegInTop_6_12[5] , \ScanLink91[9] , 
        \wRegOut_6_46[19] , \ScanLink160[2] , \wRegOut_7_105[1] , 
        \wRegInTop_7_33[3] , \wRegOut_6_33[30] , \wRegOut_6_33[29] , 
        \wRegOut_7_48[29] , \wRegOut_7_48[30] , \wRegInTop_1_1[22] , 
        \wRegInTop_3_6[26] , \ScanLink39[7] , \wRegInTop_5_18[12] , 
        \wRegInBot_5_18[15] , \wRegInTop_7_95[22] , \wRegInBot_6_25[8] , 
        \wRegInTop_7_80[16] , \wRegOut_7_89[5] , \wRegOut_4_2[21] , 
        \ScanLink107[5] , \wRegInTop_7_54[4] , \wRegInBot_4_8[5] , 
        \ScanLink24[8] , \wRegInBot_6_15[17] , \wRegInBot_6_38[7] , 
        \wRegInBot_6_60[27] , \wRegInTop_5_18[21] , \wRegInTop_5_24[0] , 
        \wRegOut_6_5[25] , \wRegInTop_6_23[15] , \wRegInBot_6_36[26] , 
        \wRegInTop_6_56[25] , \wRegInBot_6_23[12] , \wRegInBot_6_43[16] , 
        \wRegInTop_7_58[15] , \wRegOut_7_113[12] , \wRegInTop_6_43[11] , 
        \wRegInTop_7_38[11] , \wRegInTop_7_86[2] , \wRegOut_7_106[26] , 
        \wRegInTop_6_36[21] , \wRegInBot_6_56[22] , \wRegInTop_6_15[10] , 
        \wRegInTop_6_60[20] , \wRegOut_7_125[17] , \ScanLink110[30] , 
        \ScanLink133[18] , \ScanLink110[29] , \wRegInTop_7_6[31] , 
        \ScanLink146[28] , \wRegInTop_7_6[28] , \ScanLink146[31] , 
        \ScanLink165[19] , \wRegOut_7_58[0] , \wRegInTop_7_80[25] , 
        \wRegOut_7_97[9] , \wRegInBot_5_18[26] , \wRegInTop_5_27[3] , 
        \wRegInTop_7_95[11] , \wRegOut_5_28[4] , \ScanLink119[9] , 
        \wRegInTop_7_85[1] , \wRegInTop_4_9[3] , \wRegInBot_5_4[26] , 
        \wRegInBot_1_0[19] , \ScanLink5[15] , \wRegOut_2_2[1] , 
        \wRegOut_4_2[5] , \ScanLink104[6] , \wRegInTop_7_57[7] , 
        \wRegInTop_7_2[19] , \ScanLink137[29] , \ScanLink142[19] , 
        \ScanLink161[31] , \ScanLink161[28] , \wRegInTop_4_12[20] , 
        \ScanLink114[18] , \wRegInBot_4_12[27] , \wRegOut_5_9[13] , 
        \wRegEnBot_6_51[0] , \ScanLink137[30] , \wRegInTop_7_84[14] , 
        \wRegInTop_5_4[9] , \wRegInTop_7_91[20] , \wRegInTop_6_52[7] , 
        \ScanLink120[0] , \wRegInTop_7_73[1] , \wRegInTop_3_2[17] , 
        \wRegInBot_5_0[17] , \wRegOut_7_61[9] , \ScanLink240[5] , 
        \wRegInTop_6_51[4] , \wRegInTop_7_70[2] , \ScanLink123[3] , 
        \wRegInBot_3_6[8] , \wRegOut_4_6[10] , \wRegInBot_6_8[10] , 
        \ScanLink243[6] , \wRegOut_4_1[6] , \wRegOut_6_1[14] , 
        \wRegInBot_6_11[26] , \wRegInTop_6_27[24] , \wRegInBot_6_32[17] , 
        \wRegInBot_6_47[27] , \wRegOut_7_117[23] , \wRegInTop_6_52[14] , 
        \wRegInBot_6_52[13] , \wRegInTop_7_29[14] , \wRegInBot_1_1[20] , 
        \wRegOut_2_1[30] , \wRegOut_2_1[29] , \wRegOut_2_1[2] , 
        \wRegEnTop_5_2[0] , \wRegInBot_6_27[23] , \wRegInTop_6_32[10] , 
        \wRegInTop_7_49[10] , \wRegOut_7_102[17] , \wRegInTop_6_47[20] , 
        \wRegOut_7_121[26] , \wRegInTop_6_11[21] , \wRegInBot_5_0[24] , 
        \ScanLink5[26] , \wRegEnTop_7_101[0] , \wRegInTop_6_36[3] , 
        \wRegInBot_2_3[21] , \wRegInTop_3_2[24] , \ScanLink17[31] , 
        \ScanLink17[28] , \wRegInTop_4_12[13] , \wRegInBot_4_12[14] , 
        \wRegOut_5_9[20] , \wRegOut_6_14[30] , \ScanLink144[4] , 
        \wRegInTop_7_17[5] , \wRegOut_6_14[29] , \wRegOut_6_37[18] , 
        \wRegOut_6_42[28] , \wRegOut_7_39[28] , \ScanLink224[1] , 
        \wRegOut_7_121[7] , \wRegOut_6_42[31] , \wRegOut_7_39[31] , 
        \wRegOut_6_61[19] , \wRegInTop_7_91[13] , \wRegInTop_6_0[8] , 
        \ScanLink196[2] , \ScanLink67[9] , \wRegOut_6_39[4] , \wRegOut_7_6[4] , 
        \wRegInTop_7_116[8] , \ScanLink41[30] , \wRegOut_6_1[27] , 
        \wRegInBot_6_27[10] , \ScanLink99[19] , \wRegOut_7_18[2] , 
        \wRegInTop_7_84[27] , \wRegInTop_6_47[13] , \ScanLink195[1] , 
        \ScanLink209[18] , \wRegInBot_6_52[20] , \wRegInTop_7_49[23] , 
        \wRegOut_7_102[24] , \wRegInTop_6_11[12] , \wRegInTop_6_32[23] , 
        \wRegOut_7_121[15] , \wRegInBot_6_11[15] , \ScanLink62[18] , 
        \ScanLink41[29] , \wRegInTop_6_52[27] , \wRegOut_7_5[7] , 
        \wRegInTop_7_29[27] , \wRegInTop_6_27[17] , \wRegInBot_6_32[24] , 
        \wRegInBot_6_47[14] , \wRegOut_4_6[23] , \ScanLink34[19] , 
        \wRegOut_7_117[10] , \wRegOut_5_19[18] , \wRegInBot_6_8[23] , 
        \ScanLink147[7] , \wRegInTop_6_35[0] , \wRegInTop_7_14[6] , 
        \ScanLink79[5] , \wRegOut_6_27[8] , \ScanLink227[2] , 
        \wRegOut_7_94[28] , \wRegInTop_7_114[28] , \wRegInTop_3_2[3] , 
        \wRegInBot_3_3[5] , \wRegInBot_5_29[7] , \wRegOut_7_94[31] , 
        \wRegInTop_7_108[4] , \wRegInTop_7_114[31] , \wRegOut_7_122[4] , 
        \wRegOut_7_5[31] , \wRegOut_7_71[11] , \wRegInTop_5_2[7] , 
        \wRegOut_5_17[3] , \wRegOut_6_29[20] , \wRegInTop_6_49[6] , 
        \wRegOut_7_52[20] , \wRegInTop_7_68[0] , \wRegOut_7_5[28] , 
        \wRegOut_7_27[10] , \wRegOut_7_47[14] , \wRegOut_6_49[24] , 
        \wRegOut_7_32[24] , \wRegOut_7_64[25] , \wRegInBot_5_3[1] , 
        \wRegInBot_5_17[28] , \wRegOut_7_11[15] , \wRegInTop_5_18[4] , 
        \ScanLink87[21] , \wRegInBot_2_3[12] , \wRegInBot_3_0[6] , 
        \wRegOut_3_5[26] , \wRegInBot_5_17[31] , \wRegInTop_6_54[9] , 
        \ScanLink92[15] , \wRegOut_6_46[1] , \ScanLink129[22] , 
        \ScanLink149[26] , \wRegOut_7_67[7] , \wRegInTop_7_9[26] , 
        \ScanLink202[14] , \wRegOut_7_109[28] , \wRegInTop_4_1[21] , 
        \ScanLink69[14] , \wRegInBot_6_39[31] , \wRegOut_6_45[2] , 
        \ScanLink184[22] , \ScanLink221[25] , \ScanLink191[16] , 
        \wRegOut_7_109[31] , \ScanLink245[8] , \ScanLink254[15] , 
        \wRegOut_7_64[4] , \ScanLink234[11] , \wRegInBot_6_39[28] , 
        \ScanLink217[20] , \ScanLink241[21] , \wRegOut_4_7[8] , 
        \wRegEnBot_5_18[0] , \wRegOut_5_31[25] , \ScanLink138[2] , 
        \wRegInTop_3_1[0] , \wRegOut_5_12[14] , \wRegInBot_5_0[2] , 
        \wRegInTop_5_1[4] , \wRegInTop_6_6[25] , \wRegOut_5_14[0] , 
        \wRegOut_5_24[11] , \wRegOut_6_22[5] , \ScanLink92[26] , 
        \ScanLink149[15] , \wRegInTop_7_9[15] , \wRegOut_3_5[15] , 
        \wRegInTop_4_1[12] , \wRegInBot_4_10[3] , \wRegInTop_5_21[19] , 
        \ScanLink87[12] , \wRegInBot_6_60[7] , \ScanLink61[7] , 
        \wRegInTop_6_6[6] , \ScanLink129[11] , \wRegEnTop_7_90[0] , 
        \wRegOut_7_32[17] , \wRegOut_7_127[9] , \wRegInBot_6_7[0] , 
        \wRegOut_6_49[17] , \wRegOut_7_47[27] , \wRegEnTop_6_63[0] , 
        \wRegOut_7_11[26] , \wRegOut_7_64[16] , \wRegOut_7_71[22] , 
        \wRegOut_7_27[23] , \wRegInBot_5_31[5] , \wRegOut_6_29[13] , 
        \wRegInBot_4_13[0] , \wRegOut_5_24[22] , \wRegInTop_6_5[5] , 
        \wRegInTop_6_6[16] , \wRegOut_7_52[13] , \wRegInTop_7_110[6] , 
        \ScanLink62[4] , \wRegInBot_6_4[3] , \wRegOut_7_3[9] , 
        \wRegInTop_7_113[5] , \wRegOut_5_12[27] , \wRegOut_5_31[16] , 
        \ScanLink69[27] , \wRegInTop_7_57[31] , \ScanLink241[12] , 
        \ScanLink191[25] , \wRegInTop_7_74[19] , \ScanLink234[22] , 
        \ScanLink141[9] , \wRegInTop_7_57[28] , \wRegOut_6_21[6] , 
        \wRegInTop_6_59[18] , \wRegInTop_7_12[8] , \ScanLink217[13] , 
        \wRegInTop_7_22[18] , \ScanLink202[27] , \wRegInBot_6_63[4] , 
        \ScanLink254[26] , \wRegInBot_3_6[24] , \wRegInBot_4_4[18] , 
        \wRegOut_5_18[12] , \wRegInBot_6_9[30] , \ScanLink184[11] , 
        \ScanLink221[16] , \wRegInTop_7_100[16] , \wRegOut_4_7[30] , 
        \wRegOut_4_7[29] , \wRegInBot_6_9[29] , \wRegOut_7_80[16] , 
        \ScanLink198[4] , \wRegInTop_7_123[27] , \ScanLink55[17] , 
        \wRegInTop_6_10[18] , \ScanLink76[26] , \wRegOut_6_37[2] , 
        \wRegOut_7_8[2] , \wRegOut_7_16[4] , \wRegOut_7_95[22] , 
        \ScanLink237[8] , \wRegInTop_7_115[22] , \wRegInTop_7_48[30] , 
        \wRegInTop_6_33[30] , \wRegInTop_6_38[5] , \wRegInTop_6_46[19] , 
        \wRegInTop_7_19[3] , \ScanLink208[12] , \wRegInBot_1_1[13] , 
        \wRegOut_2_0[23] , \ScanLink16[22] , \ScanLink20[27] , 
        \wRegInTop_7_48[29] , \ScanLink35[13] , \ScanLink40[23] , 
        \ScanLink74[0] , \wRegInTop_6_33[29] , \wRegInBot_5_24[2] , 
        \wRegInTop_7_105[1] , \ScanLink63[12] , \wRegInTop_4_13[19] , 
        \ScanLink100[15] , \ScanLink123[24] , \ScanLink186[8] , 
        \ScanLink149[1] , \ScanLink156[14] , \wRegInTop_7_90[19] , 
        \ScanLink115[21] , \ScanLink175[25] , \ScanLink229[4] , 
        \wRegInBot_5_27[1] , \ScanLink77[3] , \ScanLink98[13] , 
        \wRegInTop_7_3[20] , \ScanLink160[11] , \ScanLink136[10] , 
        \ScanLink143[20] , \wRegOut_6_23[26] , \wRegInTop_7_106[2] , 
        \wRegInTop_6_26[9] , \wRegOut_6_56[16] , \wRegOut_7_58[26] , 
        \ScanLink16[11] , \ScanLink35[20] , \wRegInTop_5_4[24] , 
        \wRegOut_6_15[23] , \wRegOut_6_34[1] , \wRegOut_7_15[7] , 
        \wRegOut_6_36[12] , \wRegOut_6_60[13] , \wRegOut_6_43[22] , 
        \wRegOut_7_38[22] , \wRegOut_7_116[29] , \ScanLink40[10] , 
        \ScanLink20[14] , \ScanLink63[21] , \wRegOut_7_116[30] , 
        \ScanLink76[15] , \wRegInBot_6_26[30] , \wRegOut_2_0[10] , 
        \ScanLink10[4] , \wRegInBot_6_53[19] , \wRegInBot_3_6[17] , 
        \ScanLink55[24] , \wRegInBot_6_26[29] , \ScanLink133[9] , 
        \wRegInTop_7_60[8] , \ScanLink208[21] , \wRegOut_7_72[0] , 
        \wRegOut_7_95[11] , \wRegInTop_7_115[11] , \wRegInTop_5_4[17] , 
        \wRegOut_5_18[21] , \wRegOut_6_53[6] , \wRegOut_7_80[25] , 
        \wRegInTop_7_100[25] , \wRegInBot_6_11[4] , \wRegOut_6_15[10] , 
        \wRegOut_6_60[20] , \wRegInTop_7_123[14] , \wRegOut_7_38[11] , 
        \wRegInBot_6_12[7] , \wRegOut_6_23[15] , \wRegOut_6_36[21] , 
        \wRegOut_6_43[11] , \wRegOut_6_56[25] , \wRegOut_6_50[5] , 
        \wRegOut_7_58[15] , \wRegOut_7_71[3] , \ScanLink13[7] , 
        \ScanLink98[20] , \wRegInTop_7_3[13] , \ScanLink160[22] , 
        \ScanLink115[12] , \ScanLink136[23] , \ScanLink143[13] , 
        \wRegOut_0_0[1] , \wRegInBot_2_0[9] , \wRegInBot_2_2[18] , 
        \wRegInTop_4_0[18] , \wRegOut_5_8[19] , \wRegEnTop_6_11[0] , 
        \ScanLink123[17] , \ScanLink156[27] , \wRegInTop_6_8[0] , 
        \ScanLink100[26] , \ScanLink175[16] , \ScanLink151[3] , 
        \wRegInTop_6_23[4] , \wRegInBot_4_5[12] , \wRegInBot_6_9[6] , 
        \wRegInTop_6_58[12] , \wRegInTop_7_56[22] , \ScanLink235[31] , 
        \wRegInTop_7_23[12] , \ScanLink216[19] , \wRegInBot_6_38[11] , 
        \wRegInTop_7_60[27] , \wRegInTop_7_75[13] , \ScanLink240[18] , 
        \ScanLink235[28] , \ScanLink231[6] , \wRegOut_5_3[15] , 
        \wRegInTop_5_16[16] , \wRegOut_5_25[31] , \wRegOut_5_25[28] , 
        \wRegInTop_6_38[16] , \wRegInBot_6_58[15] , \wRegInTop_7_15[17] , 
        \wRegInTop_7_43[16] , \wRegOut_7_108[11] , \wRegInTop_7_36[26] , 
        \ScanLink183[5] , \wRegInBot_6_2[16] , \wRegEnBot_6_23[0] , 
        \wRegOut_6_28[19] , \wRegOut_7_4[11] , \ScanLink180[6] , 
        \wRegOut_7_26[29] , \wRegOut_7_26[30] , \wRegOut_7_53[19] , 
        \wRegOut_7_70[31] , \wRegOut_7_70[28] , \wRegInTop_5_20[13] , 
        \wRegInBot_5_20[14] , \wRegInTop_6_20[7] , \ScanLink152[0] , 
        \ScanLink86[18] , \wRegOut_7_13[9] , \ScanLink232[5] , 
        \wRegInTop_2_3[10] , \ScanLink15[9] , \wRegInBot_4_5[21] , 
        \wRegInTop_5_16[2] , \wRegInBot_5_16[11] , \wRegInBot_6_2[25] , 
        \wRegOut_6_48[7] , \ScanLink128[8] , \wRegOut_7_69[1] , 
        \wRegInTop_7_15[24] , \wRegOut_5_3[26] , \wRegInBot_5_16[22] , 
        \wRegOut_5_19[5] , \wRegInTop_6_38[25] , \wRegInTop_6_47[0] , 
        \wRegInTop_7_36[15] , \ScanLink185[28] , \wRegInTop_7_60[14] , 
        \wRegInTop_7_66[6] , \wRegInBot_6_58[26] , \ScanLink135[7] , 
        \ScanLink185[31] , \wRegInTop_7_43[25] , \wRegOut_7_108[22] , 
        \wRegInTop_6_58[21] , \wRegInTop_5_20[20] , \wRegInBot_6_38[22] , 
        \wRegInTop_6_44[3] , \wRegOut_6_55[8] , \wRegInTop_7_23[21] , 
        \wRegInTop_7_56[11] , \ScanLink128[28] , \ScanLink136[4] , 
        \wRegInTop_7_75[20] , \ScanLink255[2] , \wRegInTop_7_65[5] , 
        \ScanLink128[31] , \wRegInTop_5_15[1] , \wRegInTop_5_16[25] , 
        \wRegInBot_6_14[9] , \wRegInBot_5_20[27] , \wRegOut_7_4[22] , 
        \wRegOut_5_7[17] , \wRegInTop_5_24[11] , \wRegInBot_5_31[22] , 
        \ScanLink159[29] , \wRegInTop_5_12[14] , \wRegInBot_5_12[13] , 
        \ScanLink159[30] , \wRegInBot_5_24[16] , \wRegInTop_5_31[25] , 
        \wRegInTop_6_60[5] , \wRegInTop_7_41[3] , \ScanLink112[2] , 
        \wRegOut_3_4[0] , \wRegOut_7_0[13] , \wRegOut_3_7[3] , 
        \wRegInTop_4_2[8] , \wRegOut_4_8[14] , \wRegInTop_4_10[1] , 
        \wRegInTop_5_31[7] , \wRegOut_5_4[4] , \wRegInTop_7_93[5] , 
        \wRegInTop_4_13[2] , \wRegInBot_6_6[14] , \wRegInTop_7_90[6] , 
        \wRegOut_5_7[7] , \wRegInBot_4_1[10] , \wRegOut_7_50[8] , 
        \wRegInTop_7_64[25] , \wRegOut_6_0[5] , \wRegInTop_6_29[20] , 
        \wRegInBot_6_29[27] , \wRegInTop_7_11[15] , \wRegInTop_7_47[14] , 
        \ScanLink181[19] , \ScanLink111[1] , \wRegInTop_6_49[24] , 
        \wRegInTop_7_32[24] , \wRegInBot_6_49[23] , \wRegInBot_6_49[4] , 
        \wRegInTop_6_63[6] , \wRegInTop_7_27[10] , \wRegInTop_7_42[0] , 
        \wRegInTop_7_52[20] , \wRegOut_7_119[27] , \wRegInTop_7_71[11] , 
        \wRegInTop_1_0[31] , \wRegInTop_2_3[23] , \ScanLink9[8] , 
        \wRegOut_6_16[9] , \wRegOut_6_59[18] , \wRegInTop_7_6[9] , 
        \wRegInTop_7_38[8] , \wRegOut_7_57[28] , \wRegOut_7_0[20] , 
        \wRegOut_7_22[18] , \wRegOut_7_57[31] , \wRegOut_7_74[19] , 
        \ScanLink216[3] , \wRegInTop_5_12[27] , \ScanLink48[4] , 
        \wRegInBot_5_24[25] , \wRegInBot_4_1[23] , \wRegInTop_4_4[30] , 
        \wRegInTop_4_4[29] , \wRegOut_5_7[24] , \wRegInBot_5_12[20] , 
        \wRegInBot_5_18[6] , \wRegOut_7_113[5] , \wRegInTop_5_24[22] , 
        \wRegInTop_5_31[16] , \wRegInBot_5_31[11] , \ScanLink176[6] , 
        \wRegInTop_7_25[7] , \ScanLink82[30] , \ScanLink82[29] , 
        \wRegInTop_6_29[13] , \wRegEnTop_6_49[0] , \ScanLink212[28] , 
        \wRegInTop_7_27[23] , \ScanLink244[30] , \wRegInTop_7_52[13] , 
        \wRegOut_7_110[6] , \wRegInBot_6_49[10] , \wRegOut_7_119[14] , 
        \ScanLink212[31] , \ScanLink215[0] , \ScanLink231[19] , 
        \ScanLink244[29] , \wRegInBot_6_57[8] , \wRegInTop_7_11[26] , 
        \wRegInTop_7_71[22] , \wRegInTop_4_4[6] , \wRegInBot_4_5[0] , 
        \wRegOut_4_8[27] , \wRegOut_5_21[19] , \ScanLink79[31] , 
        \ScanLink79[28] , \wRegInBot_6_29[14] , \wRegInTop_7_26[4] , 
        \wRegInTop_7_64[16] , \wRegInTop_7_32[17] , \ScanLink99[1] , 
        \wRegInTop_6_49[17] , \wRegInTop_7_47[27] , \ScanLink175[5] , 
        \ScanLink56[8] , \wRegOut_6_3[6] , \wRegOut_7_29[3] , 
        \wRegInTop_7_127[9] , \wRegInTop_5_0[26] , \wRegInBot_6_6[27] , 
        \wRegOut_6_11[21] , \wRegEnTop_7_0[0] , \wRegOut_7_55[5] , 
        \wRegOut_6_32[10] , \wRegInBot_6_36[1] , \wRegOut_7_49[10] , 
        \wRegOut_6_47[20] , \wRegOut_6_27[24] , \ScanLink111[23] , 
        \wRegOut_6_52[14] , \wRegInTop_7_88[4] , \wRegOut_7_29[14] , 
        \wRegOut_7_87[3] , \ScanLink34[2] , \ScanLink37[1] , \wRegOut_5_25[1] , 
        \wRegInTop_7_7[22] , \ScanLink164[13] , \ScanLink132[12] , 
        \ScanLink89[25] , \ScanLink104[17] , \ScanLink109[3] , 
        \wRegEnTop_7_14[0] , \ScanLink147[22] , \ScanLink127[26] , 
        \ScanLink152[16] , \ScanLink171[27] , \ScanLink219[24] , 
        \wRegOut_5_26[2] , \wRegInTop_1_0[28] , \wRegInBot_4_6[3] , 
        \ScanLink31[11] , \ScanLink44[21] , \wRegOut_7_112[18] , 
        \ScanLink67[10] , \wRegOut_7_84[0] , \wRegInTop_1_0[3] , 
        \wRegInBot_3_2[26] , \ScanLink12[20] , \wRegInTop_4_7[5] , 
        \ScanLink24[25] , \wRegOut_5_1[9] , \ScanLink72[24] , 
        \wRegInBot_6_57[31] , \ScanLink51[15] , \wRegInBot_6_22[18] , 
        \wRegInTop_7_96[8] , \wRegInBot_6_57[28] , \wRegInTop_7_59[1] , 
        \wRegOut_4_12[20] , \wRegInTop_5_29[5] , \wRegInTop_6_8[21] , 
        \wRegInBot_6_35[2] , \wRegOut_7_56[6] , \wRegOut_7_91[20] , 
        \wRegInTop_7_111[20] , \wRegInTop_7_104[14] , \ScanLink53[5] , 
        \wRegOut_7_84[14] , \wRegInTop_7_127[25] , \ScanLink152[25] , 
        \wRegInBot_1_1[5] , \wRegOut_7_108[4] , \wRegInTop_7_122[4] , 
        \wRegInBot_3_2[15] , \wRegOut_4_3[18] , \wRegInTop_5_0[15] , 
        \wRegInTop_5_19[18] , \ScanLink89[16] , \ScanLink127[15] , 
        \wRegInTop_7_94[31] , \ScanLink104[24] , \ScanLink171[14] , 
        \wRegInTop_7_94[28] , \ScanLink164[20] , \wRegOut_6_10[7] , 
        \ScanLink81[3] , \ScanLink111[10] , \wRegInTop_7_7[11] , 
        \wRegOut_6_52[27] , \wRegInTop_7_0[7] , \ScanLink132[21] , 
        \ScanLink147[11] , \wRegOut_6_27[17] , \wRegOut_7_29[27] , 
        \wRegOut_7_31[1] , \wRegOut_6_11[12] , \wRegInBot_6_52[5] , 
        \ScanLink170[8] , \wRegOut_6_32[23] , \wRegOut_6_47[13] , 
        \wRegInTop_7_23[9] , \wRegOut_7_49[23] , \wRegOut_7_32[2] , 
        \wRegOut_4_12[13] , \wRegOut_6_13[4] , \wRegInTop_7_104[27] , 
        \ScanLink82[0] , \wRegInBot_6_51[6] , \wRegOut_7_84[27] , 
        \wRegOut_7_116[8] , \wRegInTop_7_127[16] , \wRegInTop_6_8[12] , 
        \wRegOut_7_91[13] , \wRegInTop_7_111[13] , \ScanLink0[14] , 
        \wRegInBot_1_1[30] , \wRegOut_2_0[19] , \ScanLink4[16] , 
        \wRegInBot_2_2[22] , \wRegOut_3_4[25] , \ScanLink12[13] , 
        \ScanLink24[16] , \ScanLink72[17] , \wRegInTop_6_14[29] , 
        \wRegInTop_6_42[31] , \wRegInTop_6_61[19] , \wRegInTop_7_39[31] , 
        \ScanLink31[22] , \ScanLink50[6] , \ScanLink51[26] , 
        \wRegInTop_6_14[30] , \wRegInTop_6_37[18] , \wRegInTop_7_39[28] , 
        \wRegOut_6_5[8] , \wRegInTop_6_42[28] , \wRegInTop_7_121[7] , 
        \ScanLink44[12] , \ScanLink219[17] , \wRegInTop_7_3[4] , 
        \wRegInTop_4_0[22] , \ScanLink16[3] , \wRegOut_5_25[12] , 
        \ScanLink67[23] , \wRegOut_5_13[17] , \wRegInTop_6_7[26] , 
        \wRegOut_7_69[8] , \ScanLink248[4] , \wRegOut_5_30[26] , 
        \wRegInTop_6_58[28] , \ScanLink128[1] , \wRegInTop_7_23[28] , 
        \ScanLink216[23] , \wRegInTop_7_56[18] , \wRegInTop_7_75[30] , 
        \wRegInBot_4_5[28] , \ScanLink68[17] , \wRegOut_6_55[1] , 
        \wRegInTop_6_58[31] , \ScanLink190[15] , \wRegOut_7_74[7] , 
        \ScanLink235[12] , \wRegInTop_7_23[31] , \wRegInBot_6_17[3] , 
        \wRegInTop_7_75[29] , \ScanLink240[22] , \wRegInBot_4_5[31] , 
        \wRegInTop_6_47[9] , \ScanLink185[21] , \ScanLink220[26] , 
        \ScanLink255[16] , \wRegOut_4_9[7] , \wRegInTop_5_20[29] , 
        \wRegInBot_6_14[0] , \wRegOut_6_56[2] , \ScanLink203[17] , 
        \wRegOut_7_77[4] , \ScanLink93[16] , \ScanLink128[21] , 
        \wRegInTop_7_8[25] , \ScanLink148[25] , \wRegInTop_5_20[30] , 
        \ScanLink86[22] , \wRegInBot_2_2[11] , \wRegOut_3_4[16] , 
        \ScanLink15[0] , \wRegOut_7_10[16] , \wRegOut_7_65[26] , 
        \wRegInTop_5_15[8] , \wRegOut_6_28[23] , \wRegOut_6_48[27] , 
        \wRegOut_7_33[27] , \wRegOut_7_46[17] , \wRegInTop_6_59[5] , 
        \wRegOut_7_53[23] , \wRegInTop_7_78[3] , \wRegOut_7_26[13] , 
        \wRegOut_6_31[5] , \wRegOut_7_70[12] , \wRegOut_7_10[3] , 
        \ScanLink255[25] , \wRegInTop_4_0[11] , \wRegInTop_6_8[9] , 
        \ScanLink185[12] , \ScanLink203[24] , \wRegEnTop_7_83[0] , 
        \ScanLink220[15] , \wRegOut_7_108[18] , \wRegOut_5_13[24] , 
        \ScanLink68[24] , \wRegInBot_6_38[18] , \ScanLink216[10] , 
        \ScanLink190[26] , \ScanLink235[21] , \ScanLink240[11] , 
        \wRegInBot_5_21[6] , \wRegInBot_5_22[5] , \ScanLink72[7] , 
        \wRegOut_5_25[21] , \wRegOut_5_30[15] , \wRegInTop_7_103[6] , 
        \wRegInTop_6_7[15] , \ScanLink71[4] , \wRegOut_7_4[18] , 
        \wRegOut_7_26[20] , \wRegOut_6_28[10] , \wRegOut_6_48[14] , 
        \wRegOut_7_10[25] , \wRegOut_7_53[10] , \wRegOut_7_70[21] , 
        \wRegInTop_7_100[5] , \wRegOut_7_33[14] , \wRegOut_7_65[15] , 
        \ScanLink128[12] , \wRegOut_7_46[24] , \wRegInTop_3_3[14] , 
        \ScanLink16[18] , \ScanLink35[30] , \ScanLink35[29] , 
        \wRegInBot_5_16[18] , \ScanLink86[11] , \wRegOut_6_32[6] , 
        \wRegOut_7_13[0] , \wRegOut_6_0[17] , \wRegInTop_6_10[22] , 
        \ScanLink93[25] , \wRegInTop_7_8[16] , \ScanLink148[16] , 
        \ScanLink152[9] , \wRegOut_7_120[25] , \wRegInBot_6_53[10] , 
        \ScanLink208[31] , \wRegInTop_6_26[27] , \wRegInBot_6_26[20] , 
        \wRegInTop_6_33[13] , \wRegInTop_7_48[13] , \wRegOut_7_103[14] , 
        \wRegInTop_6_46[23] , \ScanLink208[28] , \wRegOut_7_116[20] , 
        \ScanLink40[19] , \ScanLink63[31] , \wRegInBot_6_46[24] , 
        \wRegInTop_6_53[17] , \wRegInBot_6_33[14] , \wRegInTop_7_28[17] , 
        \wRegInTop_5_10[5] , \wRegOut_4_7[13] , \ScanLink63[28] , 
        \wRegEnBot_6_42[0] , \wRegInBot_6_10[25] , \wRegOut_7_72[9] , 
        \wRegOut_5_18[31] , \wRegOut_5_18[28] , \ScanLink253[5] , 
        \wRegInBot_6_9[13] , \wRegInTop_6_41[7] , \wRegInTop_7_60[1] , 
        \ScanLink133[0] , \wRegOut_7_95[18] , \wRegInTop_7_115[18] , 
        \wRegInBot_5_8[3] , \wRegInTop_5_9[5] , \ScanLink250[6] , 
        \wRegInTop_3_3[27] , \wRegInTop_4_13[23] , \wRegInBot_4_13[24] , 
        \wRegInBot_5_1[14] , \wRegOut_5_8[10] , \wRegOut_6_15[19] , 
        \wRegOut_6_36[31] , \wRegOut_6_60[29] , \wRegOut_6_36[28] , 
        \wRegInTop_6_42[4] , \wRegOut_6_60[30] , \ScanLink130[3] , 
        \wRegOut_7_38[18] , \wRegInTop_7_63[2] , \wRegOut_6_43[18] , 
        \wRegInTop_5_13[6] , \ScanLink98[29] , \wRegInTop_7_90[23] , 
        \ScanLink69[6] , \ScanLink98[30] , \wRegInTop_7_85[17] , 
        \wRegOut_4_7[20] , \ScanLink237[1] , \wRegInTop_7_118[7] , 
        \wRegEnTop_7_112[0] , \wRegInBot_6_9[20] , \ScanLink157[4] , 
        \wRegInBot_6_10[16] , \ScanLink74[9] , \wRegInTop_6_25[3] , 
        \wRegInTop_6_53[24] , \wRegInTop_6_26[14] , \wRegInBot_6_33[27] , 
        \wRegInTop_7_28[24] , \wRegInTop_7_105[8] , \wRegInBot_6_46[17] , 
        \wRegOut_7_116[13] , \wRegInBot_1_1[29] , \wRegInTop_6_10[11] , 
        \wRegOut_7_120[16] , \wRegInBot_6_26[13] , \wRegInTop_6_46[10] , 
        \ScanLink185[2] , \wRegInBot_6_53[23] , \wRegInTop_7_48[20] , 
        \wRegOut_7_103[27] , \ScanLink4[25] , \wRegInTop_4_13[10] , 
        \wRegOut_6_0[24] , \wRegOut_6_29[7] , \wRegInTop_6_33[20] , 
        \wRegInBot_4_13[17] , \wRegOut_5_8[23] , \wRegInBot_5_27[8] , 
        \ScanLink115[31] , \ScanLink115[28] , \wRegInTop_7_3[29] , 
        \ScanLink143[30] , \ScanLink160[18] , \wRegInTop_7_85[24] , 
        \ScanLink136[19] , \ScanLink143[29] , \wRegInTop_7_3[30] , 
        \ScanLink149[8] , \ScanLink186[1] , \wRegInTop_7_90[10] , 
        \wRegInBot_5_1[27] , \wRegInTop_6_26[0] , \wRegOut_6_34[8] , 
        \ScanLink234[2] , \ScanLink154[7] , \wRegInTop_5_19[11] , 
        \wRegInTop_7_7[18] , \ScanLink164[29] , \wRegInBot_5_19[16] , 
        \wRegOut_6_6[2] , \ScanLink111[19] , \ScanLink132[31] , 
        \ScanLink132[28] , \ScanLink147[18] , \wRegInTop_7_81[15] , 
        \ScanLink164[30] , \wRegInTop_7_94[21] , \wRegInTop_7_23[0] , 
        \ScanLink170[1] , \wRegOut_7_115[2] , \wRegInTop_3_7[16] , 
        \wRegInBot_5_5[16] , \wRegOut_7_31[8] , \ScanLink210[4] , 
        \wRegInTop_7_20[3] , \ScanLink173[2] , \ScanLink0[27] , 
        \wRegInTop_1_0[12] , \wRegOut_4_3[11] , \ScanLink213[7] , 
        \ScanLink82[9] , \wRegInTop_6_22[25] , \wRegOut_7_116[1] , 
        \wRegInBot_6_37[16] , \wRegInBot_6_42[26] , \wRegInTop_7_59[25] , 
        \wRegOut_7_112[22] , \wRegInTop_6_57[15] , \wRegInBot_6_61[17] , 
        \wRegInBot_5_5[25] , \wRegOut_6_4[15] , \wRegInTop_6_14[20] , 
        \wRegInBot_6_14[27] , \wRegOut_7_124[27] , \wRegInTop_6_61[10] , 
        \wRegOut_6_5[1] , \wRegInBot_6_22[22] , \wRegInTop_6_37[11] , 
        \wRegInBot_6_57[12] , \wRegOut_7_107[16] , \wRegInTop_7_39[21] , 
        \wRegInTop_6_42[21] , \ScanLink114[5] , \wRegInTop_7_47[4] , 
        \wRegInTop_1_0[21] , \wRegOut_3_1[4] , \wRegOut_3_2[7] , 
        \wRegOut_5_2[3] , \wRegInBot_5_19[25] , \wRegOut_6_11[31] , 
        \wRegOut_6_11[28] , \wRegEnTop_6_28[0] , \wRegInBot_6_36[8] , 
        \wRegOut_6_47[30] , \wRegOut_7_49[19] , \wRegOut_6_32[19] , 
        \wRegOut_6_47[29] , \wRegInTop_7_94[12] , \wRegInTop_7_95[2] , 
        \wRegOut_7_48[3] , \wRegInTop_7_81[26] , \ScanLink12[30] , 
        \wRegInBot_4_5[9] , \wRegInTop_4_15[5] , \ScanLink37[8] , 
        \wRegInTop_5_19[22] , \wRegOut_5_25[8] , \wRegInTop_6_61[23] , 
        \wRegOut_5_1[0] , \wRegOut_7_124[14] , \ScanLink44[28] , 
        \wRegOut_6_4[26] , \wRegInTop_6_14[13] , \wRegInBot_6_22[11] , 
        \wRegInTop_6_42[12] , \wRegInTop_7_39[12] , \wRegInTop_7_96[1] , 
        \wRegInTop_7_59[8] , \wRegOut_7_107[25] , \wRegInTop_6_37[22] , 
        \wRegInBot_6_57[21] , \wRegInTop_6_57[26] , \wRegInTop_6_22[16] , 
        \wRegInBot_6_37[25] , \ScanLink31[18] , \wRegInBot_6_42[15] , 
        \wRegInTop_7_59[16] , \wRegOut_7_84[9] , \wRegOut_7_112[11] , 
        \wRegEnBot_4_3[0] , \ScanLink44[31] , \wRegInBot_6_14[14] , 
        \ScanLink12[29] , \ScanLink67[19] , \wRegInBot_6_28[4] , 
        \wRegInTop_3_7[25] , \wRegOut_4_3[22] , \wRegInBot_6_61[24] , 
        \wRegOut_4_12[30] , \wRegOut_4_12[29] , \ScanLink117[6] , 
        \wRegInTop_7_44[7] , \ScanLink29[4] , \wRegInTop_6_8[31] , 
        \wRegOut_7_91[30] , \wRegInTop_7_111[30] , \wRegOut_0_0[8] , 
        \wRegInTop_6_8[28] , \wRegOut_7_91[29] , \wRegOut_7_99[6] , 
        \wRegInTop_6_19[7] , \wRegInTop_7_38[1] , \wRegInTop_7_111[29] , 
        \wRegOut_7_57[21] , \ScanLink1[9] , \wRegInTop_1_1[18] , 
        \wRegInBot_2_0[0] , \wRegInTop_2_1[6] , \wRegInTop_2_2[5] , 
        \wRegInTop_2_3[19] , \wRegOut_3_0[27] , \ScanLink9[1] , 
        \wRegInBot_5_12[30] , \ScanLink55[2] , \wRegOut_6_59[11] , 
        \wRegOut_7_0[29] , \wRegOut_7_0[30] , \wRegInTop_7_6[0] , 
        \wRegOut_7_22[11] , \wRegOut_7_74[10] , \wRegOut_7_14[14] , 
        \wRegOut_7_61[24] , \wRegOut_6_39[15] , \wRegOut_7_42[15] , 
        \wRegOut_7_37[25] , \wRegInTop_7_124[3] , \wRegInBot_5_12[29] , 
        \wRegInBot_5_31[18] , \ScanLink159[13] , \wRegOut_6_16[0] , 
        \ScanLink82[20] , \wRegOut_7_37[6] , \ScanLink79[21] , \ScanLink87[4] , 
        \ScanLink97[14] , \wRegInBot_6_54[2] , \ScanLink139[17] , 
        \ScanLink19[25] , \wRegInTop_4_4[20] , \ScanLink84[7] , 
        \ScanLink181[23] , \ScanLink207[15] , \ScanLink224[24] , 
        \ScanLink251[14] , \wRegInBot_6_49[19] , \ScanLink212[21] , 
        \wRegOut_6_15[3] , \wRegOut_7_34[5] , \ScanLink231[10] , 
        \ScanLink194[17] , \ScanLink215[9] , \ScanLink244[20] , 
        \wRegOut_5_17[15] , \wRegInBot_6_57[1] , \wRegOut_5_21[10] , 
        \wRegInTop_7_5[3] , \ScanLink168[3] , \ScanLink56[1] , \ScanLink99[8] , 
        \wRegInTop_6_3[24] , \wRegEnTop_7_75[0] , \ScanLink208[6] , 
        \wRegInTop_7_127[0] , \ScanLink97[27] , \ScanLink139[24] , 
        \wRegInTop_4_10[8] , \wRegInTop_5_24[18] , \ScanLink82[13] , 
        \ScanLink159[20] , \wRegOut_7_53[2] , \wRegInBot_6_30[6] , 
        \wRegOut_7_14[27] , \wRegInBot_2_3[3] , \wRegOut_3_4[9] , 
        \wRegInBot_4_3[7] , \ScanLink31[6] , \wRegOut_5_23[6] , 
        \wRegOut_6_39[26] , \wRegOut_7_37[16] , \wRegOut_7_61[17] , 
        \wRegOut_7_42[26] , \wRegOut_6_59[22] , \wRegOut_7_22[22] , 
        \wRegOut_7_57[12] , \wRegInTop_4_2[1] , \wRegOut_7_81[4] , 
        \wRegOut_5_21[23] , \wRegOut_7_74[23] , \wRegInTop_6_3[17] , 
        \wRegOut_3_0[14] , \wRegInBot_4_0[4] , \wRegInTop_4_1[2] , 
        \wRegOut_7_82[7] , \ScanLink19[16] , \wRegInTop_4_4[13] , 
        \ScanLink32[5] , \wRegOut_5_17[26] , \wRegOut_5_20[5] , 
        \wRegInTop_6_29[29] , \ScanLink111[8] , \wRegInTop_7_42[9] , 
        \wRegInTop_6_29[30] , \wRegInTop_7_27[19] , \wRegInTop_7_52[29] , 
        \ScanLink212[12] , \wRegInTop_7_52[30] , \ScanLink244[13] , 
        \wRegInTop_7_71[18] , \ScanLink79[12] , \wRegInBot_6_33[5] , 
        \wRegOut_7_50[1] , \ScanLink194[24] , \ScanLink231[23] , 
        \ScanLink251[27] , \wRegInBot_3_3[25] , \wRegInBot_4_1[19] , 
        \wRegOut_4_2[31] , \ScanLink181[10] , \ScanLink207[26] , 
        \ScanLink224[17] , \wRegOut_4_13[23] , \wRegInTop_7_105[17] , 
        \wRegInTop_7_126[26] , \ScanLink13[23] , \wRegOut_4_2[28] , 
        \ScanLink25[26] , \ScanLink50[16] , \wRegInTop_6_9[22] , 
        \wRegInBot_6_25[1] , \wRegOut_7_46[5] , \wRegOut_7_85[17] , 
        \wRegOut_7_90[23] , \wRegInTop_7_110[23] , \wRegInTop_7_38[18] , 
        \wRegInTop_6_43[18] , \wRegInTop_6_60[30] , \wRegInTop_7_49[2] , 
        \wRegInTop_5_24[9] , \ScanLink73[27] , \wRegInTop_6_36[28] , 
        \wRegInTop_6_60[29] , \ScanLink66[13] , \wRegInTop_6_15[19] , 
        \wRegInTop_6_36[31] , \wRegOut_7_94[3] , \ScanLink13[10] , 
        \ScanLink24[1] , \ScanLink218[27] , \ScanLink27[2] , \wRegOut_4_14[4] , 
        \ScanLink30[12] , \ScanLink45[22] , \ScanLink88[26] , 
        \ScanLink105[14] , \wRegInTop_7_95[18] , \ScanLink119[0] , 
        \ScanLink170[24] , \ScanLink126[25] , \wRegInTop_7_85[8] , 
        \ScanLink153[15] , \ScanLink133[11] , \wRegInTop_5_1[25] , 
        \wRegInTop_5_18[31] , \ScanLink146[21] , \wRegInTop_5_18[28] , 
        \ScanLink110[20] , \wRegOut_7_58[9] , \ScanLink165[10] , 
        \wRegOut_7_97[0] , \wRegOut_6_26[27] , \wRegInTop_7_6[21] , 
        \wRegOut_6_33[13] , \wRegOut_6_53[17] , \wRegInTop_7_98[7] , 
        \wRegOut_7_28[17] , \wRegOut_7_48[13] , \wRegOut_6_10[22] , 
        \wRegOut_6_46[23] , \wRegOut_7_45[6] , \wRegInBot_6_26[2] , 
        \wRegOut_7_113[31] , \ScanLink25[15] , \ScanLink30[21] , 
        \ScanLink66[20] , \ScanLink45[11] , \ScanLink218[14] , 
        \wRegOut_7_113[28] , \ScanLink40[5] , \wRegInBot_6_56[18] , 
        \wRegInBot_5_10[7] , \ScanLink50[25] , \wRegInBot_6_23[28] , 
        \ScanLink73[14] , \wRegInBot_6_23[31] , \ScanLink4[4] , 
        \wRegInTop_2_2[20] , \wRegInTop_2_2[13] , \wRegInBot_3_3[16] , 
        \wRegOut_6_8[4] , \wRegInTop_6_9[11] , \wRegOut_7_90[10] , 
        \wRegInTop_7_110[10] , \ScanLink92[3] , \wRegInTop_7_30[9] , 
        \ScanLink163[8] , \wRegInTop_7_126[15] , \wRegInBot_4_0[13] , 
        \wRegInTop_4_5[19] , \wRegOut_4_13[10] , \wRegOut_7_22[1] , 
        \wRegInTop_7_105[24] , \wRegInTop_5_1[16] , \wRegEnTop_5_13[0] , 
        \wRegInBot_6_41[5] , \wRegOut_7_85[24] , \wRegOut_6_46[10] , 
        \ScanLink43[6] , \wRegOut_6_10[11] , \wRegOut_6_33[20] , 
        \wRegOut_7_48[20] , \ScanLink88[15] , \wRegOut_6_26[14] , 
        \ScanLink91[0] , \wRegInBot_6_42[6] , \wRegOut_7_21[2] , 
        \wRegOut_6_53[24] , \wRegOut_7_28[24] , \ScanLink110[13] , 
        \ScanLink133[22] , \ScanLink146[12] , \wRegOut_7_105[8] , 
        \wRegInTop_7_6[12] , \ScanLink165[23] , \ScanLink105[27] , 
        \ScanLink170[17] , \wRegInBot_5_13[4] , \ScanLink153[26] , 
        \wRegOut_7_118[7] , \wRegInTop_6_28[23] , \ScanLink101[2] , 
        \ScanLink126[16] , \wRegInTop_7_70[12] , \ScanLink245[19] , 
        \ScanLink230[29] , \wRegInBot_6_48[20] , \wRegInTop_7_53[23] , 
        \wRegEnBot_5_21[0] , \wRegInTop_7_52[3] , \ScanLink213[18] , 
        \ScanLink230[30] , \wRegOut_7_118[24] , \wRegInBot_6_28[24] , 
        \wRegInTop_7_26[13] , \wRegInTop_7_46[17] , \wRegInTop_6_48[27] , 
        \wRegInTop_7_33[27] , \wRegInTop_7_10[16] , \wRegInTop_7_65[26] , 
        \wRegOut_4_9[17] , \wRegOut_4_11[9] , \wRegOut_5_20[30] , 
        \wRegInTop_5_22[7] , \ScanLink78[18] , \wRegOut_5_20[29] , 
        \wRegInTop_7_80[5] , \wRegInBot_6_7[17] , \wRegInTop_5_21[4] , 
        \wRegInTop_7_83[6] , \wRegInBot_5_25[15] , \wRegInTop_5_30[26] , 
        \wRegOut_6_58[31] , \wRegOut_6_58[28] , \wRegOut_7_1[10] , 
        \wRegOut_7_23[31] , \wRegOut_7_75[29] , \wRegOut_7_23[28] , 
        \wRegInTop_7_51[0] , \wRegOut_7_56[18] , \wRegOut_7_75[30] , 
        \ScanLink102[1] , \ScanLink7[7] , \wRegOut_4_9[24] , \wRegOut_5_6[14] , 
        \wRegOut_5_9[8] , \wRegInTop_5_13[17] , \ScanLink83[19] , 
        \wRegOut_7_43[8] , \wRegInBot_5_13[10] , \wRegInTop_5_25[12] , 
        \wRegInBot_5_30[21] , \wRegInBot_6_7[24] , \ScanLink178[9] , 
        \wRegOut_6_18[6] , \wRegOut_7_39[0] , \wRegInBot_4_0[20] , 
        \wRegInBot_5_16[9] , \ScanLink89[2] , \wRegInTop_6_17[1] , 
        \wRegInTop_7_33[14] , \wRegInTop_7_36[7] , \wRegInBot_6_28[17] , 
        \wRegInTop_6_48[14] , \ScanLink180[30] , \wRegInTop_7_8[6] , 
        \ScanLink165[6] , \wRegInTop_7_46[24] , \wRegOut_5_6[27] , 
        \wRegInBot_5_13[23] , \wRegInTop_6_28[10] , \wRegInTop_7_10[25] , 
        \wRegInTop_7_26[20] , \ScanLink180[29] , \wRegInTop_7_65[15] , 
        \wRegInTop_7_70[21] , \ScanLink205[3] , \wRegInBot_6_48[13] , 
        \wRegInTop_7_53[10] , \wRegOut_7_100[5] , \wRegOut_7_118[17] , 
        \wRegInTop_5_25[21] , \wRegInBot_5_30[12] , \ScanLink166[5] , 
        \wRegInTop_6_14[2] , \wRegInTop_7_35[4] , \wRegInBot_5_25[26] , 
        \ScanLink58[7] , \ScanLink158[19] , \wRegInTop_5_13[24] , 
        \wRegInTop_5_30[15] , \wRegOut_7_103[6] , \wRegInBot_6_44[8] , 
        \ScanLink206[0] , \ScanLink45[8] , \wRegOut_7_1[23] , 
        \wRegInBot_6_59[7] , \wRegOut_1_0[7] , \wRegOut_5_2[16] , 
        \ScanLink222[6] , \wRegInTop_5_17[15] , \wRegInBot_5_17[12] , 
        \wRegInTop_5_21[10] , \wRegInBot_5_21[17] , \wRegInTop_6_30[4] , 
        \ScanLink129[18] , \wRegOut_7_127[0] , \wRegInTop_7_11[2] , 
        \ScanLink142[3] , \wRegInBot_6_7[9] , \wRegOut_7_0[3] , 
        \wRegOut_7_5[12] , \ScanLink190[5] , \wRegInBot_1_0[23] , 
        \wRegOut_2_1[20] , \wRegInBot_2_3[31] , \wRegInBot_2_3[28] , 
        \wRegEnTop_3_7[0] , \wRegOut_4_4[2] , \wRegInBot_4_4[11] , 
        \wRegInBot_4_13[9] , \wRegOut_7_3[0] , \wRegEnBot_6_1[0] , 
        \wRegInBot_6_3[15] , \wRegEnBot_6_30[0] , \ScanLink193[6] , 
        \wRegInTop_6_39[15] , \wRegInBot_6_59[16] , \wRegInTop_7_42[15] , 
        \wRegOut_7_109[12] , \wRegInTop_7_14[14] , \wRegInTop_7_37[25] , 
        \wRegOut_7_124[3] , \wRegInTop_7_61[24] , \ScanLink221[5] , 
        \wRegInBot_5_3[8] , \wRegInTop_6_33[7] , \ScanLink141[0] , 
        \ScanLink184[18] , \wRegInTop_7_74[10] , \wRegInBot_6_39[12] , 
        \wRegInTop_6_59[11] , \wRegInTop_7_12[1] , \wRegInTop_7_57[21] , 
        \wRegInTop_7_22[11] , \wRegInBot_6_19[5] , \wRegOut_6_29[30] , 
        \wRegOut_7_71[18] , \wRegOut_7_52[30] , \ScanLink18[5] , 
        \wRegOut_6_29[29] , \wRegOut_7_5[21] , \wRegOut_7_52[29] , 
        \wRegInTop_7_68[9] , \wRegOut_7_27[19] , \wRegInTop_5_17[26] , 
        \wRegInBot_5_21[24] , \wRegOut_6_46[8] , \ScanLink246[2] , 
        \wRegInBot_5_17[21] , \wRegOut_5_2[25] , \ScanLink87[28] , 
        \wRegInTop_6_54[0] , \ScanLink126[7] , \wRegInTop_7_75[6] , 
        \wRegInTop_3_1[9] , \wRegInTop_4_1[31] , \wRegInTop_5_21[23] , 
        \ScanLink87[31] , \ScanLink217[30] , \ScanLink234[18] , 
        \ScanLink241[28] , \ScanLink245[1] , \wRegInTop_4_1[28] , 
        \wRegInBot_6_39[21] , \wRegInTop_6_59[22] , \wRegInTop_7_74[23] , 
        \ScanLink217[29] , \wRegInTop_7_22[22] , \ScanLink241[31] , 
        \wRegInBot_4_4[22] , \wRegInTop_6_39[26] , \wRegInTop_6_57[3] , 
        \wRegInTop_7_37[16] , \wRegInTop_7_57[12] , \wRegInTop_7_76[5] , 
        \wRegInBot_6_59[25] , \ScanLink125[4] , \wRegInTop_7_42[26] , 
        \wRegOut_7_109[21] , \wRegOut_4_7[1] , \wRegOut_5_14[9] , 
        \wRegOut_6_58[4] , \wRegInTop_7_14[27] , \wRegInTop_7_61[17] , 
        \wRegOut_7_79[2] , \wRegOut_5_24[18] , \wRegInBot_6_3[26] , 
        \wRegInTop_5_5[27] , \wRegOut_6_37[11] , \wRegOut_7_39[21] , 
        \wRegOut_6_14[20] , \wRegOut_6_24[2] , \wRegOut_6_42[21] , 
        \ScanLink224[8] , \wRegOut_6_61[10] , \ScanLink17[21] , 
        \wRegOut_5_9[30] , \wRegOut_5_9[29] , \ScanLink67[0] , 
        \wRegOut_6_22[25] , \wRegOut_6_57[15] , \wRegOut_7_59[25] , 
        \ScanLink137[13] , \ScanLink99[10] , \ScanLink114[22] , 
        \ScanLink142[23] , \ScanLink239[7] , \wRegInTop_7_116[1] , 
        \wRegInTop_7_2[23] , \ScanLink161[12] , \ScanLink101[16] , 
        \wRegInTop_6_0[1] , \ScanLink122[27] , \ScanLink174[26] , 
        \ScanLink159[2] , \ScanLink62[11] , \wRegInBot_6_1[7] , 
        \ScanLink157[17] , \wRegInBot_4_15[7] , \ScanLink41[20] , 
        \ScanLink64[3] , \wRegInTop_7_115[2] , \ScanLink34[10] , 
        \wRegOut_7_117[19] , \ScanLink54[14] , \wRegInTop_6_3[2] , 
        \wRegInBot_6_27[19] , \wRegInTop_6_28[6] , \ScanLink195[8] , 
        \ScanLink209[11] , \wRegInBot_1_0[10] , \wRegOut_2_1[13] , 
        \wRegOut_2_2[8] , \wRegInBot_3_7[27] , \ScanLink21[24] , 
        \wRegInBot_6_52[29] , \wRegOut_5_19[11] , \wRegInBot_6_2[4] , 
        \ScanLink77[25] , \wRegOut_6_27[1] , \wRegInBot_6_52[30] , 
        \wRegInTop_6_35[9] , \ScanLink188[7] , \wRegOut_7_94[21] , 
        \wRegInTop_7_114[21] , \wRegInTop_7_122[24] , \wRegInTop_7_101[15] , 
        \wRegInTop_5_4[0] , \wRegOut_7_81[15] , \ScanLink174[15] , 
        \wRegInTop_3_4[4] , \wRegInBot_3_5[2] , \wRegInTop_4_12[30] , 
        \wRegInBot_5_5[6] , \wRegOut_5_11[4] , \ScanLink101[25] , 
        \wRegInTop_7_91[29] , \ScanLink157[24] , \ScanLink122[14] , 
        \wRegInTop_7_91[30] , \ScanLink142[10] , \ScanLink137[20] , 
        \ScanLink161[21] , \wRegInTop_4_12[29] , \ScanLink99[23] , 
        \wRegInTop_7_2[10] , \wRegOut_6_40[6] , \ScanLink114[11] , 
        \wRegOut_7_61[0] , \wRegInBot_3_7[14] , \wRegOut_4_6[19] , 
        \wRegInTop_5_5[14] , \wRegOut_6_22[16] , \wRegOut_6_57[26] , 
        \wRegOut_6_42[12] , \ScanLink120[9] , \wRegOut_7_59[16] , 
        \wRegOut_7_39[12] , \wRegInBot_6_8[19] , \wRegOut_6_14[13] , 
        \wRegOut_6_37[22] , \wRegInTop_7_73[8] , \wRegOut_6_61[23] , 
        \wRegInTop_7_122[17] , \ScanLink21[17] , \wRegOut_5_19[22] , 
        \wRegOut_6_43[5] , \wRegOut_7_62[3] , \wRegOut_7_81[26] , 
        \wRegInTop_7_101[26] , \wRegInTop_7_49[19] , \wRegOut_7_94[12] , 
        \wRegInTop_7_114[12] , \ScanLink2[8] , \wRegInTop_1_1[30] , 
        \wRegInTop_1_1[29] , \ScanLink13[21] , \wRegInBot_3_6[1] , 
        \wRegInBot_5_6[5] , \wRegInTop_5_7[3] , \wRegOut_5_12[7] , 
        \ScanLink54[27] , \wRegInTop_6_11[31] , \wRegInTop_6_32[19] , 
        \wRegInTop_6_47[29] , \ScanLink209[22] , \wRegInTop_6_11[28] , 
        \ScanLink77[16] , \wRegInTop_6_47[30] , \wRegInTop_3_7[7] , 
        \ScanLink17[12] , \wRegInTop_4_9[8] , \wRegInTop_5_1[27] , 
        \ScanLink34[23] , \ScanLink62[22] , \ScanLink41[13] , 
        \wRegOut_6_46[21] , \wRegOut_6_33[11] , \wRegOut_7_48[11] , 
        \ScanLink27[0] , \wRegOut_4_14[6] , \wRegOut_6_10[20] , 
        \wRegInBot_6_26[0] , \wRegOut_7_45[4] , \wRegOut_6_26[25] , 
        \wRegOut_6_53[15] , \wRegOut_7_28[15] , \ScanLink146[23] , 
        \wRegInTop_7_98[5] , \ScanLink133[13] , \wRegInTop_5_27[8] , 
        \ScanLink88[24] , \ScanLink110[22] , \wRegInTop_7_6[23] , 
        \ScanLink165[12] , \wRegOut_7_97[2] , \ScanLink170[26] , 
        \ScanLink105[16] , \ScanLink119[2] , \ScanLink126[27] , 
        \ScanLink153[17] , \wRegOut_7_94[1] , \ScanLink24[3] , 
        \ScanLink30[10] , \ScanLink66[11] , \wRegOut_7_113[19] , 
        \ScanLink45[20] , \ScanLink218[25] , \wRegInBot_3_3[27] , 
        \ScanLink25[24] , \ScanLink50[14] , \wRegInBot_6_23[19] , 
        \wRegInBot_6_56[29] , \wRegInTop_6_9[20] , \ScanLink73[25] , 
        \wRegInBot_6_56[30] , \wRegInTop_7_49[0] , \wRegInTop_7_86[9] , 
        \wRegInBot_6_25[3] , \wRegOut_7_90[21] , \wRegOut_7_46[7] , 
        \wRegInTop_7_110[21] , \wRegInTop_7_126[24] , \wRegOut_4_13[21] , 
        \wRegOut_7_85[15] , \wRegInTop_7_105[15] , \ScanLink4[6] , 
        \wRegInTop_2_2[11] , \wRegInBot_3_3[14] , \wRegOut_4_2[19] , 
        \wRegOut_4_13[12] , \wRegInTop_5_1[14] , \ScanLink43[4] , 
        \wRegInBot_5_13[6] , \ScanLink88[17] , \ScanLink105[25] , 
        \wRegInTop_7_95[29] , \ScanLink170[15] , \wRegInTop_7_95[30] , 
        \ScanLink126[14] , \wRegOut_7_118[5] , \wRegInTop_5_18[19] , 
        \ScanLink110[11] , \ScanLink133[20] , \ScanLink153[24] , 
        \ScanLink146[10] , \wRegInTop_7_6[10] , \ScanLink165[21] , 
        \wRegOut_6_26[16] , \wRegInBot_6_42[4] , \wRegOut_7_21[0] , 
        \ScanLink91[2] , \wRegOut_6_53[26] , \wRegOut_7_28[26] , 
        \wRegOut_6_33[22] , \wRegOut_7_48[22] , \ScanLink160[9] , 
        \wRegInTop_7_33[8] , \wRegOut_6_8[6] , \wRegOut_6_10[13] , 
        \wRegOut_6_46[12] , \wRegOut_7_106[9] , \ScanLink92[1] , 
        \wRegInBot_6_41[7] , \wRegInTop_7_126[17] , \wRegOut_7_22[3] , 
        \wRegInTop_7_105[26] , \ScanLink13[12] , \ScanLink25[17] , 
        \wRegInBot_5_10[5] , \ScanLink50[27] , \wRegInTop_6_9[13] , 
        \wRegOut_7_85[26] , \wRegOut_7_90[12] , \wRegInTop_7_110[12] , 
        \wRegInTop_7_38[29] , \wRegInTop_6_43[29] , \ScanLink40[7] , 
        \wRegInTop_6_15[31] , \wRegEnTop_6_42[0] , \wRegInTop_6_36[19] , 
        \ScanLink66[22] , \ScanLink73[16] , \wRegInTop_7_38[30] , 
        \wRegInTop_6_15[28] , \wRegInTop_6_43[30] , \wRegInTop_6_60[18] , 
        \ScanLink30[23] , \ScanLink45[13] , \ScanLink218[16] , 
        \wRegOut_5_6[16] , \wRegInBot_5_13[12] , \wRegInTop_5_25[10] , 
        \wRegInBot_5_30[23] , \ScanLink158[31] , \wRegInBot_5_25[17] , 
        \ScanLink158[28] , \wRegInBot_4_0[11] , \wRegOut_4_9[15] , 
        \wRegOut_4_12[8] , \wRegInTop_5_13[15] , \wRegInTop_5_30[24] , 
        \ScanLink102[3] , \wRegInTop_7_51[2] , \wRegOut_7_1[12] , 
        \wRegInTop_5_21[6] , \wRegInTop_7_83[4] , \wRegInBot_6_7[15] , 
        \wRegInTop_5_22[5] , \wRegInBot_6_28[26] , \wRegInTop_7_33[25] , 
        \wRegInTop_7_80[7] , \wRegInTop_6_48[25] , \wRegInTop_7_46[15] , 
        \wRegInBot_5_15[8] , \wRegInTop_6_28[21] , \wRegInTop_7_10[14] , 
        \wRegInTop_7_26[11] , \wRegOut_7_40[9] , \ScanLink180[18] , 
        \wRegInTop_7_65[24] , \wRegInTop_7_70[10] , \ScanLink101[0] , 
        \wRegInBot_6_48[22] , \wRegInTop_7_52[1] , \wRegOut_7_118[26] , 
        \wRegInTop_7_53[21] , \wRegInBot_6_59[5] , \wRegOut_1_0[5] , 
        \wRegInTop_2_2[22] , \wRegInBot_5_25[24] , \wRegInTop_5_30[17] , 
        \wRegOut_6_58[19] , \wRegOut_7_1[21] , \wRegOut_7_56[30] , 
        \wRegOut_7_75[18] , \wRegOut_7_23[19] , \wRegInTop_7_28[9] , 
        \wRegOut_7_56[29] , \wRegOut_7_103[4] , \ScanLink58[5] , 
        \ScanLink7[5] , \wRegInBot_4_0[22] , \wRegInTop_4_5[31] , 
        \wRegOut_5_6[25] , \wRegInTop_5_13[26] , \ScanLink83[28] , 
        \ScanLink206[2] , \wRegInBot_5_13[21] , \wRegInTop_5_25[23] , 
        \ScanLink83[31] , \wRegInBot_5_30[10] , \wRegInTop_6_14[0] , 
        \ScanLink166[7] , \wRegInTop_7_35[6] , \wRegInBot_6_47[9] , 
        \wRegInTop_7_70[23] , \ScanLink245[28] , \wRegInTop_4_5[28] , 
        \wRegInTop_6_28[12] , \ScanLink205[1] , \ScanLink230[18] , 
        \ScanLink213[30] , \wRegInBot_6_48[11] , \ScanLink245[31] , 
        \wRegOut_7_118[15] , \ScanLink78[30] , \wRegInTop_7_8[4] , 
        \wRegInTop_7_26[22] , \wRegInTop_7_53[12] , \ScanLink213[29] , 
        \wRegOut_7_100[7] , \wRegInTop_7_46[26] , \ScanLink78[29] , 
        \wRegInTop_6_17[3] , \wRegInBot_6_28[15] , \wRegInTop_6_48[16] , 
        \wRegInTop_7_33[16] , \wRegInTop_7_36[5] , \ScanLink165[4] , 
        \wRegInTop_7_65[17] , \wRegInTop_7_10[27] , \wRegEnTop_7_120[0] , 
        \wRegInTop_4_1[19] , \wRegOut_4_9[26] , \ScanLink46[9] , 
        \wRegOut_5_20[18] , \wRegOut_6_18[4] , \wRegOut_7_39[2] , 
        \ScanLink89[0] , \wRegInBot_6_7[26] , \wRegInBot_6_39[10] , 
        \wRegInTop_6_59[13] , \wRegInTop_7_74[12] , \ScanLink234[29] , 
        \ScanLink241[19] , \ScanLink217[18] , \ScanLink234[30] , 
        \wRegInTop_7_12[3] , \ScanLink141[2] , \wRegInTop_7_22[13] , 
        \wRegInTop_7_57[23] , \wRegInBot_4_4[13] , \wRegInTop_6_33[5] , 
        \wRegInTop_6_39[17] , \wRegInBot_6_59[14] , \wRegInTop_7_37[27] , 
        \wRegOut_7_124[1] , \wRegInTop_7_42[17] , \wRegOut_7_109[10] , 
        \wRegOut_5_24[30] , \wRegInTop_7_14[16] , \wRegInTop_7_61[26] , 
        \ScanLink221[7] , \wRegOut_5_24[29] , \wRegInBot_6_3[17] , 
        \wRegInBot_6_4[8] , \ScanLink193[4] , \wRegOut_7_3[2] , 
        \wRegInTop_1_0[10] , \wRegInBot_1_0[21] , \wRegInBot_2_3[19] , 
        \wRegInBot_4_10[8] , \wRegOut_6_29[18] , \wRegOut_7_27[31] , 
        \ScanLink190[7] , \wRegOut_7_71[29] , \wRegOut_7_52[18] , 
        \wRegOut_7_71[30] , \wRegOut_5_2[14] , \wRegInTop_5_17[17] , 
        \wRegInBot_5_21[15] , \wRegOut_7_0[1] , \wRegOut_7_5[10] , 
        \wRegOut_7_27[28] , \wRegInTop_6_30[6] , \wRegInTop_7_11[0] , 
        \ScanLink142[1] , \wRegInBot_5_17[10] , \wRegInTop_3_2[8] , 
        \ScanLink18[7] , \wRegInBot_4_4[20] , \wRegOut_4_7[3] , 
        \wRegInTop_5_21[12] , \ScanLink87[19] , \ScanLink222[4] , 
        \wRegOut_7_127[2] , \wRegInBot_6_3[24] , \ScanLink138[9] , 
        \wRegInBot_5_0[9] , \wRegInTop_6_39[24] , \wRegOut_6_58[6] , 
        \wRegInBot_6_59[27] , \wRegInTop_7_42[24] , \wRegOut_7_79[0] , 
        \wRegOut_7_109[23] , \wRegInTop_6_57[1] , \ScanLink125[6] , 
        \wRegInTop_7_37[14] , \wRegInTop_7_76[7] , \wRegInTop_7_14[25] , 
        \ScanLink184[30] , \wRegInTop_7_61[15] , \wRegOut_5_2[27] , 
        \wRegInBot_6_39[23] , \wRegOut_6_45[9] , \ScanLink184[29] , 
        \wRegInTop_7_74[21] , \ScanLink245[3] , \wRegInTop_6_59[20] , 
        \wRegInTop_7_57[10] , \wRegInTop_7_22[20] , \wRegInBot_5_17[23] , 
        \wRegInTop_5_21[21] , \ScanLink129[30] , \wRegInBot_5_21[26] , 
        \wRegInTop_6_54[2] , \ScanLink126[5] , \ScanLink129[29] , 
        \wRegInTop_7_75[4] , \wRegInTop_5_17[24] , \ScanLink246[0] , 
        \wRegInBot_3_7[25] , \wRegOut_4_4[0] , \wRegOut_4_6[31] , 
        \wRegEnBot_5_6[0] , \wRegOut_5_17[8] , \wRegOut_7_5[23] , 
        \wRegInBot_6_19[7] , \wRegInBot_6_8[28] , \wRegInTop_7_122[26] , 
        \ScanLink188[5] , \ScanLink21[26] , \wRegOut_4_6[28] , 
        \wRegOut_5_19[13] , \wRegInBot_6_8[31] , \wRegOut_7_81[17] , 
        \wRegInTop_7_101[17] , \wRegOut_6_27[3] , \wRegOut_7_94[23] , 
        \ScanLink227[9] , \wRegInTop_7_114[23] , \wRegInTop_7_49[28] , 
        \wRegInBot_1_0[12] , \wRegOut_2_1[22] , \ScanLink17[23] , 
        \ScanLink54[16] , \wRegInBot_6_2[6] , \wRegInTop_6_32[28] , 
        \wRegInTop_6_3[0] , \wRegInTop_6_11[19] , \wRegInTop_6_28[4] , 
        \ScanLink209[13] , \wRegInTop_6_32[31] , \wRegInTop_6_47[18] , 
        \wRegInTop_7_49[31] , \ScanLink77[27] , \wRegInTop_4_12[18] , 
        \wRegInBot_4_15[5] , \ScanLink62[13] , \ScanLink34[12] , 
        \wRegInTop_7_115[0] , \ScanLink41[22] , \ScanLink64[1] , 
        \wRegEnTop_7_47[0] , \wRegInTop_6_0[3] , \wRegInBot_6_1[5] , 
        \ScanLink101[14] , \ScanLink174[24] , \wRegInTop_7_91[18] , 
        \ScanLink157[15] , \ScanLink196[9] , \ScanLink67[2] , 
        \ScanLink122[25] , \ScanLink159[0] , \ScanLink137[11] , 
        \ScanLink142[21] , \wRegInTop_7_116[3] , \ScanLink99[12] , 
        \ScanLink161[10] , \wRegInTop_7_2[21] , \wRegEnBot_6_28[0] , 
        \ScanLink114[20] , \wRegOut_7_18[9] , \ScanLink239[5] , 
        \wRegInBot_3_6[3] , \wRegInTop_3_7[5] , \wRegInTop_5_5[25] , 
        \wRegOut_6_22[27] , \wRegInTop_6_36[8] , \wRegOut_6_57[17] , 
        \wRegOut_6_42[23] , \wRegOut_7_39[23] , \wRegOut_7_59[27] , 
        \ScanLink62[20] , \wRegOut_6_14[22] , \wRegOut_6_24[0] , 
        \wRegOut_6_37[13] , \wRegOut_6_61[12] , \ScanLink17[10] , 
        \wRegOut_7_117[31] , \ScanLink34[21] , \ScanLink41[11] , 
        \wRegOut_7_117[28] , \wRegOut_5_12[5] , \ScanLink54[25] , 
        \wRegInBot_6_27[28] , \wRegInBot_6_52[18] , \ScanLink209[20] , 
        \wRegInBot_1_1[18] , \ScanLink4[14] , \wRegOut_2_1[11] , 
        \wRegOut_2_1[9] , \ScanLink21[15] , \ScanLink77[14] , 
        \wRegInBot_6_27[31] , \wRegInBot_3_7[16] , \wRegInBot_5_6[7] , 
        \wRegInTop_5_7[1] , \wRegOut_5_19[20] , \ScanLink123[8] , 
        \wRegInTop_7_70[9] , \wRegOut_7_94[10] , \wRegInTop_7_114[10] , 
        \wRegInTop_7_122[15] , \wRegOut_6_43[7] , \wRegInTop_7_101[24] , 
        \wRegOut_7_62[1] , \wRegInTop_5_5[16] , \wRegOut_6_37[20] , 
        \wRegOut_7_81[24] , \wRegOut_7_39[10] , \wRegOut_6_14[11] , 
        \wRegOut_6_42[10] , \wRegOut_6_61[21] , \wRegInBot_2_2[20] , 
        \wRegInTop_3_4[6] , \wRegOut_6_22[14] , \wRegOut_6_40[4] , 
        \wRegOut_7_61[2] , \ScanLink114[13] , \wRegOut_6_57[24] , 
        \wRegOut_7_59[14] , \ScanLink137[22] , \ScanLink142[12] , 
        \wRegInBot_3_5[0] , \ScanLink99[21] , \ScanLink161[23] , 
        \wRegInTop_7_2[12] , \ScanLink15[2] , \wRegInTop_5_4[2] , 
        \wRegInBot_5_5[4] , \wRegOut_5_9[18] , \ScanLink101[27] , 
        \ScanLink174[17] , \wRegOut_5_11[6] , \ScanLink122[16] , 
        \wRegOut_6_28[21] , \wRegOut_7_4[29] , \ScanLink157[26] , 
        \wRegOut_7_26[11] , \wRegOut_6_48[25] , \wRegInTop_6_59[7] , 
        \wRegOut_7_4[30] , \wRegOut_7_53[21] , \wRegInTop_7_78[1] , 
        \wRegOut_7_10[14] , \wRegOut_7_70[10] , \wRegOut_7_33[25] , 
        \wRegOut_7_65[24] , \wCtrlOut_2[0] , \wRegOut_7_46[15] , 
        \wRegInBot_5_16[30] , \wRegInTop_6_44[8] , \ScanLink128[23] , 
        \wRegInBot_2_2[13] , \wRegOut_3_4[27] , \wRegOut_4_9[5] , 
        \ScanLink86[20] , \wRegInBot_5_16[29] , \wRegInBot_6_14[2] , 
        \ScanLink93[14] , \wRegInTop_7_8[27] , \wRegOut_6_56[0] , 
        \ScanLink148[27] , \wRegOut_7_77[6] , \wRegOut_7_108[30] , 
        \ScanLink255[14] , \wRegInTop_4_0[20] , \ScanLink185[23] , 
        \ScanLink220[24] , \ScanLink203[15] , \wRegOut_7_108[29] , 
        \ScanLink16[1] , \wRegEnTop_5_9[0] , \ScanLink68[15] , 
        \wRegInBot_6_17[1] , \wRegInBot_6_38[29] , \ScanLink216[21] , 
        \ScanLink240[20] , \wRegOut_6_55[3] , \ScanLink190[17] , 
        \wRegOut_7_74[5] , \ScanLink235[10] , \ScanLink255[9] , 
        \wRegInBot_6_38[30] , \wRegOut_5_13[15] , \wRegInTop_5_16[9] , 
        \wRegOut_5_25[10] , \wRegOut_5_30[24] , \ScanLink128[3] , 
        \wRegInTop_5_20[18] , \wRegInTop_6_7[24] , \wRegEnTop_7_35[0] , 
        \ScanLink93[27] , \wRegInTop_7_8[14] , \ScanLink248[6] , 
        \ScanLink128[10] , \ScanLink148[14] , \ScanLink86[13] , 
        \wRegOut_7_13[2] , \wRegOut_6_32[4] , \wRegOut_3_4[14] , 
        \wRegInTop_4_0[13] , \wRegOut_5_13[26] , \wRegInBot_5_21[4] , 
        \wRegOut_6_28[12] , \wRegOut_6_48[16] , \wRegOut_7_10[27] , 
        \wRegOut_7_65[17] , \wRegOut_7_33[16] , \wRegOut_7_46[26] , 
        \wRegOut_7_53[12] , \wRegInTop_7_100[7] , \wRegOut_5_25[23] , 
        \ScanLink71[6] , \wRegOut_7_26[22] , \wRegOut_7_70[23] , 
        \wRegInTop_6_7[17] , \wRegInBot_5_22[7] , \wRegInTop_7_103[4] , 
        \wRegOut_5_30[17] , \ScanLink72[5] , \wRegInTop_6_58[19] , 
        \wRegInTop_7_23[19] , \ScanLink216[12] , \ScanLink151[8] , 
        \ScanLink68[26] , \wRegInTop_7_56[29] , \ScanLink190[24] , 
        \ScanLink235[23] , \wRegInTop_7_56[30] , \wRegInTop_7_75[18] , 
        \ScanLink240[13] , \wRegInBot_4_5[19] , \wRegInTop_4_13[21] , 
        \wRegEnTop_5_21[0] , \ScanLink185[10] , \ScanLink220[17] , 
        \wRegOut_6_31[7] , \wRegOut_7_10[1] , \ScanLink255[27] , 
        \ScanLink203[26] , \wRegInBot_4_13[26] , \wRegInTop_5_13[4] , 
        \ScanLink115[19] , \ScanLink136[31] , \ScanLink160[29] , 
        \wRegInTop_7_85[15] , \wRegInTop_7_3[18] , \ScanLink136[28] , 
        \ScanLink143[18] , \ScanLink160[30] , \wRegInTop_7_90[21] , 
        \wRegInBot_5_1[16] , \wRegOut_5_8[12] , \wRegInTop_6_42[6] , 
        \ScanLink130[1] , \wRegInTop_7_63[0] , \wRegInBot_5_8[1] , 
        \wRegInTop_3_3[16] , \wRegInTop_5_9[7] , \wRegOut_7_71[8] , 
        \ScanLink250[4] , \wRegEnBot_5_13[0] , \wRegOut_4_7[11] , 
        \wRegInTop_6_41[5] , \ScanLink133[2] , \wRegInTop_7_60[3] , 
        \ScanLink253[7] , \wRegInTop_5_10[7] , \wRegInBot_6_9[11] , 
        \wRegInBot_6_10[27] , \wRegInTop_6_26[25] , \wRegInBot_6_33[16] , 
        \wRegInTop_6_53[15] , \wRegInTop_7_28[15] , \wRegInBot_6_46[26] , 
        \wRegOut_7_116[22] , \wRegOut_6_0[15] , \wRegInTop_6_10[20] , 
        \wRegOut_7_120[27] , \wRegInBot_6_26[22] , \wRegInTop_6_46[21] , 
        \wRegInTop_7_48[11] , \wRegOut_7_103[16] , \wRegOut_2_0[31] , 
        \wRegInTop_6_33[11] , \wRegInBot_6_53[12] , \wRegOut_2_0[28] , 
        \ScanLink4[27] , \wRegInTop_6_26[2] , \ScanLink154[5] , 
        \wRegInBot_5_1[25] , \wRegInTop_3_3[25] , \ScanLink16[30] , 
        \wRegInTop_4_13[12] , \wRegInBot_4_13[15] , \wRegOut_6_15[31] , 
        \wRegOut_6_15[28] , \wRegOut_6_43[30] , \wRegOut_6_60[18] , 
        \wRegOut_7_38[30] , \ScanLink234[0] , \wRegOut_6_36[19] , 
        \wRegOut_6_43[29] , \wRegOut_7_38[29] , \ScanLink186[3] , 
        \wRegOut_5_8[21] , \ScanLink98[18] , \wRegInTop_7_90[12] , 
        \ScanLink35[18] , \wRegInBot_5_24[9] , \wRegOut_6_0[26] , 
        \wRegInTop_6_10[13] , \ScanLink77[8] , \wRegOut_6_29[5] , 
        \wRegInTop_7_85[26] , \wRegInTop_7_106[9] , \wRegOut_7_120[14] , 
        \wRegInTop_6_26[16] , \wRegInBot_6_26[11] , \wRegInTop_6_33[22] , 
        \wRegInBot_6_53[21] , \wRegInTop_7_48[22] , \wRegOut_7_103[25] , 
        \wRegInTop_6_46[12] , \wRegInTop_7_19[8] , \ScanLink208[19] , 
        \ScanLink185[0] , \wRegOut_7_116[11] , \ScanLink16[29] , 
        \ScanLink40[28] , \wRegInBot_6_33[25] , \wRegInBot_6_46[15] , 
        \wRegInTop_6_53[26] , \wRegInTop_7_28[26] , \wRegOut_4_7[22] , 
        \ScanLink40[31] , \ScanLink63[19] , \wRegInBot_6_10[14] , 
        \wRegOut_5_18[19] , \ScanLink69[4] , \wRegInBot_6_9[22] , 
        \wRegInTop_6_25[1] , \ScanLink157[6] , \wRegOut_7_95[30] , 
        \wRegInTop_7_118[5] , \wRegInTop_7_115[30] , \wRegOut_7_8[9] , 
        \ScanLink31[29] , \ScanLink44[19] , \wRegOut_6_4[17] , 
        \wRegOut_6_5[3] , \wRegInTop_6_14[22] , \wRegOut_6_37[9] , 
        \wRegOut_7_95[29] , \wRegInTop_7_115[29] , \wRegInTop_6_61[12] , 
        \ScanLink237[3] , \wRegOut_7_124[25] , \wRegInBot_6_22[20] , 
        \wRegInTop_6_42[23] , \wRegInTop_7_39[23] , \wRegInBot_6_57[10] , 
        \wRegOut_7_107[14] , \wRegInTop_6_37[13] , \wRegInTop_6_57[17] , 
        \ScanLink67[31] , \wRegInTop_6_22[27] , \wRegInBot_6_37[14] , 
        \wRegInBot_6_42[24] , \wRegInBot_6_14[25] , \wRegInTop_7_59[27] , 
        \wRegOut_7_112[20] , \ScanLink12[18] , \ScanLink67[28] , 
        \wRegInTop_3_7[14] , \wRegOut_4_3[13] , \ScanLink31[30] , 
        \wRegInBot_6_61[15] , \wRegOut_4_12[18] , \wRegOut_7_32[9] , 
        \ScanLink213[5] , \wRegOut_7_116[3] , \wRegInTop_7_20[1] , 
        \ScanLink173[0] , \ScanLink0[16] , \wRegInBot_5_5[14] , 
        \wRegInTop_6_8[19] , \wRegOut_7_91[18] , \wRegInTop_7_111[18] , 
        \ScanLink81[8] , \wRegOut_7_115[0] , \wRegInTop_1_0[8] , 
        \wRegOut_6_6[0] , \wRegOut_6_11[19] , \wRegOut_7_49[31] , 
        \ScanLink210[6] , \wRegOut_6_32[31] , \wRegOut_6_32[28] , 
        \wRegOut_7_49[28] , \wRegOut_6_47[18] , \ScanLink170[3] , 
        \wRegInTop_7_23[2] , \wRegInTop_3_7[27] , \ScanLink29[6] , 
        \wRegInTop_5_19[13] , \wRegInBot_5_19[14] , \wRegInTop_7_94[23] , 
        \wRegInTop_7_81[17] , \wRegInBot_6_35[9] , \wRegOut_7_99[4] , 
        \wRegOut_0_0[3] , \ScanLink0[25] , \wRegInTop_1_0[23] , 
        \wRegOut_3_1[6] , \wRegOut_4_3[20] , \ScanLink34[9] , 
        \wRegInTop_6_22[14] , \ScanLink117[4] , \wRegInTop_7_44[5] , 
        \wRegInBot_6_42[17] , \wRegInTop_7_59[14] , \wRegOut_7_112[13] , 
        \wRegInTop_6_57[24] , \wRegOut_5_26[9] , \wRegInBot_6_28[6] , 
        \wRegInBot_6_37[27] , \wRegInBot_6_61[26] , \wRegInBot_4_6[8] , 
        \wRegEnTop_2_2[0] , \wRegInTop_4_15[7] , \wRegOut_5_1[2] , 
        \wRegInTop_6_14[11] , \wRegInBot_6_14[16] , \wRegOut_7_124[16] , 
        \wRegInTop_6_61[21] , \wRegOut_3_2[5] , \wRegInTop_5_19[20] , 
        \wRegOut_6_4[24] , \wRegInBot_6_57[23] , \wRegInBot_6_22[13] , 
        \wRegInTop_6_37[20] , \wRegOut_7_107[27] , \wRegInTop_7_39[10] , 
        \wRegInTop_7_96[3] , \wRegInTop_6_42[10] , \ScanLink147[30] , 
        \ScanLink164[18] , \ScanLink111[28] , \wRegInTop_7_7[29] , 
        \wRegOut_7_48[1] , \wRegOut_5_2[1] , \ScanLink109[8] , 
        \ScanLink111[31] , \wRegInTop_7_7[30] , \ScanLink147[29] , 
        \wRegInTop_7_81[24] , \wRegOut_7_87[8] , \ScanLink132[19] , 
        \wRegInTop_7_95[0] , \wRegInBot_5_19[27] , \wRegInTop_7_94[10] , 
        \ScanLink114[7] , \wRegInTop_7_47[6] , \wRegEnBot_1_1[0] , 
        \wRegInBot_1_1[22] , \wRegOut_2_0[21] , \wRegInBot_2_0[2] , 
        \wRegInTop_2_3[31] , \wRegOut_3_0[25] , \wRegInBot_4_1[28] , 
        \ScanLink19[27] , \wRegInTop_4_4[22] , \wRegInBot_5_5[27] , 
        \wRegOut_5_17[17] , \wRegOut_5_21[12] , \wRegInTop_7_127[2] , 
        \ScanLink56[3] , \wRegInTop_6_3[26] , \wRegOut_7_29[8] , 
        \ScanLink208[4] , \wRegInTop_6_29[18] , \wRegInTop_7_5[1] , 
        \ScanLink168[1] , \wRegInTop_7_52[18] , \ScanLink84[5] , 
        \wRegInTop_7_71[30] , \ScanLink212[23] , \wRegInBot_6_57[3] , 
        \wRegInTop_7_27[28] , \ScanLink244[22] , \wRegOut_6_15[1] , 
        \wRegInTop_7_71[29] , \wRegInTop_7_27[31] , \wRegOut_7_34[7] , 
        \ScanLink194[15] , \ScanLink231[12] , \ScanLink251[16] , 
        \ScanLink9[3] , \wRegInBot_4_1[31] , \ScanLink79[23] , 
        \ScanLink181[21] , \ScanLink224[26] , \wRegInBot_6_54[0] , 
        \ScanLink207[17] , \wRegOut_6_16[2] , \ScanLink97[16] , 
        \wRegInTop_2_3[28] , \ScanLink139[15] , \wRegOut_7_37[4] , 
        \ScanLink216[8] , \wRegOut_3_0[16] , \ScanLink55[0] , 
        \wRegInTop_5_24[30] , \wRegInTop_5_24[29] , \ScanLink87[6] , 
        \ScanLink159[11] , \ScanLink82[22] , \wRegOut_7_14[16] , 
        \wRegOut_7_37[27] , \wRegOut_7_61[26] , \wRegOut_7_42[17] , 
        \wRegInTop_7_124[1] , \wRegInTop_6_19[5] , \wRegOut_6_39[17] , 
        \wRegOut_6_59[13] , \wRegInTop_7_6[2] , \wRegOut_7_22[13] , 
        \wRegInTop_7_38[3] , \wRegOut_7_57[23] , \wRegOut_7_74[12] , 
        \wRegOut_3_7[8] , \wRegInBot_4_0[6] , \wRegInTop_4_1[0] , 
        \ScanLink19[14] , \wRegInTop_4_4[11] , \ScanLink79[10] , 
        \wRegInBot_6_33[7] , \wRegInBot_6_49[28] , \wRegOut_7_50[3] , 
        \ScanLink181[12] , \ScanLink224[15] , \ScanLink207[24] , 
        \ScanLink251[25] , \ScanLink212[10] , \ScanLink194[26] , 
        \ScanLink231[21] , \ScanLink244[11] , \wRegOut_5_17[24] , 
        \wRegInBot_6_49[31] , \wRegOut_7_82[5] , \ScanLink32[7] , 
        \wRegOut_5_20[7] , \wRegEnTop_6_30[0] , \wRegOut_5_21[21] , 
        \wRegInTop_2_1[4] , \wRegInTop_2_2[7] , \wRegInBot_2_3[1] , 
        \wRegInTop_4_2[3] , \wRegInTop_4_13[9] , \wRegInTop_6_3[15] , 
        \ScanLink31[4] , \wRegOut_5_23[4] , \wRegOut_7_0[18] , 
        \wRegOut_7_57[10] , \wRegOut_6_59[20] , \wRegOut_7_22[20] , 
        \wRegInBot_4_3[5] , \wRegOut_7_74[21] , \wRegOut_7_81[6] , 
        \wRegOut_7_61[15] , \wRegOut_7_14[25] , \wRegInTop_5_4[26] , 
        \wRegInBot_5_12[18] , \wRegInBot_5_31[29] , \wRegOut_6_39[24] , 
        \wRegOut_7_42[24] , \wRegOut_7_37[14] , \ScanLink159[22] , 
        \wRegInBot_5_31[30] , \wRegOut_6_15[21] , \ScanLink82[11] , 
        \wRegInBot_6_30[4] , \ScanLink97[25] , \wRegOut_7_53[0] , 
        \wRegOut_6_34[3] , \ScanLink112[9] , \ScanLink139[26] , 
        \wRegInTop_7_41[8] , \wRegOut_6_60[11] , \wRegOut_7_15[5] , 
        \ScanLink234[9] , \wRegOut_7_38[20] , \wRegOut_6_23[24] , 
        \wRegOut_6_36[10] , \wRegOut_6_43[20] , \wRegOut_6_56[14] , 
        \wRegOut_7_58[24] , \ScanLink16[20] , \ScanLink35[11] , 
        \wRegOut_5_8[31] , \wRegInBot_5_27[3] , \ScanLink98[11] , 
        \ScanLink160[13] , \ScanLink115[23] , \wRegInTop_7_3[22] , 
        \ScanLink143[22] , \ScanLink229[6] , \wRegInTop_7_106[0] , 
        \ScanLink77[1] , \ScanLink136[12] , \wRegEnTop_7_54[0] , 
        \wRegOut_5_8[28] , \ScanLink123[26] , \ScanLink149[3] , 
        \ScanLink156[16] , \wRegInBot_5_24[0] , \ScanLink100[17] , 
        \ScanLink175[27] , \wRegInTop_7_105[3] , \wRegOut_7_116[18] , 
        \ScanLink40[21] , \ScanLink74[2] , \ScanLink20[25] , \ScanLink63[10] , 
        \ScanLink76[24] , \wRegInBot_6_53[31] , \wRegInBot_6_53[28] , 
        \wRegInBot_1_1[11] , \wRegOut_2_0[12] , \ScanLink13[5] , 
        \wRegInBot_3_6[26] , \ScanLink55[15] , \wRegInBot_6_26[18] , 
        \wRegOut_6_37[0] , \wRegInTop_6_38[7] , \wRegInTop_7_19[1] , 
        \ScanLink185[9] , \ScanLink208[10] , \wRegOut_7_8[0] , 
        \wRegOut_7_16[6] , \wRegOut_7_95[20] , \wRegInTop_7_115[20] , 
        \wRegOut_5_18[10] , \wRegOut_7_80[14] , \wRegInTop_7_100[14] , 
        \wRegInTop_6_25[8] , \wRegInTop_7_123[25] , \ScanLink123[15] , 
        \ScanLink198[6] , \wRegInTop_7_90[31] , \wRegInTop_4_13[31] , 
        \wRegInTop_4_13[28] , \ScanLink100[24] , \ScanLink156[25] , 
        \wRegInTop_7_90[28] , \ScanLink115[10] , \ScanLink175[14] , 
        \ScanLink98[22] , \ScanLink160[20] , \wRegInTop_7_3[11] , 
        \wRegInBot_5_8[8] , \wRegOut_6_23[17] , \ScanLink136[21] , 
        \ScanLink143[11] , \wRegOut_6_56[27] , \wRegOut_7_58[17] , 
        \wRegInBot_3_6[15] , \wRegOut_4_7[18] , \wRegInTop_5_4[15] , 
        \wRegInBot_6_12[5] , \wRegOut_6_15[12] , \wRegOut_6_50[7] , 
        \wRegOut_7_71[1] , \wRegOut_6_36[23] , \wRegOut_6_60[22] , 
        \wRegOut_6_43[13] , \ScanLink130[8] , \wRegOut_7_38[13] , 
        \wRegInTop_7_63[9] , \wRegOut_5_18[23] , \wRegInBot_6_11[6] , 
        \wRegOut_6_53[4] , \wRegInTop_7_100[27] , \ScanLink55[26] , 
        \wRegInBot_6_9[18] , \wRegOut_7_72[2] , \wRegOut_7_80[27] , 
        \wRegInTop_6_10[29] , \ScanLink76[17] , \wRegOut_7_95[13] , 
        \wRegInTop_7_123[16] , \wRegInTop_7_115[13] , \wRegInTop_6_46[31] , 
        \wRegInTop_6_46[28] , \ScanLink208[23] , \wRegInBot_2_2[30] , 
        \ScanLink10[6] , \ScanLink20[16] , \wRegInTop_6_10[30] , 
        \wRegInTop_7_48[18] , \ScanLink16[13] , \ScanLink35[22] , 
        \ScanLink40[12] , \wRegInTop_6_33[18] , \ScanLink63[23] , 
        \wRegInBot_4_5[10] , \wRegOut_5_3[17] , \wRegInBot_5_16[13] , 
        \wRegInTop_5_20[11] , \ScanLink128[19] , \wRegInTop_5_16[14] , 
        \ScanLink232[7] , \wRegInBot_5_20[16] , \wRegInBot_6_2[14] , 
        \wRegInTop_6_20[5] , \wRegOut_7_4[13] , \ScanLink152[2] , 
        \ScanLink180[4] , \wRegInTop_7_15[15] , \ScanLink183[7] , 
        \wRegInTop_5_15[3] , \wRegInTop_6_8[2] , \wRegInBot_6_9[4] , 
        \wRegInTop_6_38[14] , \wRegInBot_6_58[17] , \wRegOut_7_10[8] , 
        \ScanLink185[19] , \wRegInTop_7_60[25] , \wRegInTop_7_36[24] , 
        \ScanLink231[4] , \wRegInTop_7_43[14] , \wRegOut_7_108[13] , 
        \wRegInBot_6_38[13] , \wRegInTop_6_58[10] , \wRegInTop_7_23[10] , 
        \wRegInTop_6_23[6] , \ScanLink151[1] , \wRegInTop_7_56[20] , 
        \wRegOut_6_28[31] , \wRegOut_6_28[28] , \wRegOut_7_4[20] , 
        \wRegInTop_7_75[11] , \wRegOut_7_26[18] , \wRegOut_7_53[28] , 
        \wRegInTop_7_78[8] , \wRegOut_7_53[31] , \wRegInTop_5_16[27] , 
        \wRegOut_7_70[19] , \wRegInTop_5_20[22] , \wRegInBot_5_20[25] , 
        \wRegOut_6_56[9] , \ScanLink86[30] , \wRegInBot_2_2[29] , 
        \ScanLink86[29] , \wRegInTop_6_44[1] , \ScanLink136[6] , 
        \wRegInTop_7_65[7] , \wRegInTop_2_3[12] , \wRegInBot_2_3[8] , 
        \wRegOut_3_7[1] , \wRegInTop_4_0[30] , \wRegInTop_4_0[29] , 
        \wRegOut_5_3[24] , \wRegInBot_5_16[20] , \wRegInTop_7_56[13] , 
        \ScanLink240[30] , \wRegOut_5_19[7] , \wRegInBot_6_38[20] , 
        \wRegInTop_6_58[23] , \wRegInTop_7_23[23] , \ScanLink216[28] , 
        \wRegInTop_7_75[22] , \ScanLink240[29] , \ScanLink16[8] , 
        \wRegInBot_4_5[23] , \wRegInBot_6_17[8] , \wRegInTop_7_60[16] , 
        \ScanLink216[31] , \ScanLink235[19] , \ScanLink255[0] , 
        \wRegOut_5_25[19] , \wRegInTop_6_38[27] , \wRegInBot_6_58[24] , 
        \wRegInTop_7_15[26] , \wRegInTop_7_43[27] , \wRegOut_7_108[20] , 
        \wRegInTop_6_47[2] , \ScanLink135[5] , \wRegInTop_7_36[17] , 
        \wRegInTop_7_66[4] , \wRegInTop_4_1[9] , \wRegInBot_4_1[12] , 
        \wRegInTop_4_4[18] , \wRegInTop_5_16[0] , \wRegOut_6_48[5] , 
        \wRegOut_7_69[3] , \wRegInBot_6_2[27] , \wRegInTop_6_29[22] , 
        \wRegInTop_7_27[12] , \ScanLink212[19] , \ScanLink231[31] , 
        \ScanLink111[3] , \wRegOut_7_119[25] , \ScanLink79[19] , 
        \wRegInBot_6_49[21] , \wRegInTop_6_63[4] , \wRegInTop_7_42[2] , 
        \wRegInTop_7_52[22] , \wRegInTop_7_71[13] , \ScanLink231[28] , 
        \ScanLink244[18] , \wRegInTop_7_11[17] , \wRegInTop_4_13[0] , 
        \wRegOut_5_7[5] , \wRegOut_5_21[31] , \wRegOut_5_21[28] , 
        \wRegInBot_6_29[25] , \wRegInTop_7_32[26] , \wRegInTop_7_64[27] , 
        \wRegInTop_6_49[26] , \wRegInTop_7_47[16] , \wRegInTop_7_90[4] , 
        \wRegOut_4_8[16] , \wRegOut_5_4[6] , \wRegInBot_6_6[16] , 
        \wRegOut_3_4[2] , \wRegEnTop_4_7[0] , \wRegInTop_4_10[3] , 
        \wRegEnBot_6_63[0] , \wRegInTop_5_31[5] , \wRegOut_6_59[29] , 
        \wRegOut_7_57[19] , \wRegOut_7_74[31] , \wRegInTop_7_93[7] , 
        \wRegOut_7_0[11] , \wRegOut_7_22[29] , \wRegOut_7_74[28] , 
        \wRegOut_6_59[30] , \wRegOut_7_22[30] , \wRegInTop_5_12[16] , 
        \wRegInBot_5_24[14] , \wRegOut_4_8[25] , \wRegOut_5_7[15] , 
        \wRegInBot_5_12[11] , \wRegInTop_5_24[13] , \wRegInTop_5_31[27] , 
        \ScanLink112[0] , \wRegInTop_6_60[7] , \wRegInTop_7_41[1] , 
        \wRegInBot_5_31[20] , \ScanLink82[18] , \wRegOut_7_53[9] , 
        \wRegInBot_6_6[25] , \wRegInTop_7_5[8] , \ScanLink168[8] , 
        \wRegInTop_2_3[21] , \wRegInBot_4_1[21] , \wRegEnTop_5_18[0] , 
        \wRegOut_6_3[4] , \ScanLink99[3] , \wRegOut_7_29[1] , 
        \wRegInTop_7_64[14] , \wRegOut_5_7[26] , \wRegInTop_5_24[20] , 
        \wRegOut_6_15[8] , \wRegInTop_6_29[11] , \wRegInBot_6_29[16] , 
        \wRegInTop_7_11[24] , \wRegInTop_7_47[25] , \ScanLink181[28] , 
        \wRegInTop_6_49[15] , \wRegInTop_7_26[6] , \wRegInTop_7_32[15] , 
        \ScanLink175[7] , \ScanLink181[31] , \wRegInBot_6_49[12] , 
        \wRegInTop_7_27[21] , \wRegInTop_7_52[11] , \wRegOut_7_110[4] , 
        \wRegOut_7_119[16] , \wRegInTop_7_71[20] , \ScanLink215[2] , 
        \wRegInBot_5_31[13] , \wRegInTop_7_25[5] , \ScanLink159[18] , 
        \ScanLink176[4] , \wRegInTop_5_12[25] , \wRegInBot_5_12[22] , 
        \wRegInBot_6_54[9] , \ScanLink48[6] , \wRegInBot_5_18[4] , 
        \ScanLink216[1] , \wRegInBot_5_24[27] , \wRegInTop_5_31[14] , 
        \wRegOut_7_113[7] , \wRegOut_7_0[22] , \wRegInBot_3_2[24] , 
        \ScanLink55[9] , \wRegOut_6_0[7] , \wRegInBot_6_49[6] , 
        \wRegInTop_7_124[8] , \wRegOut_4_3[30] , \wRegOut_4_3[29] , 
        \wRegOut_4_12[22] , \wRegInTop_5_29[7] , \wRegOut_7_84[16] , 
        \wRegInTop_7_104[16] , \wRegInTop_7_127[27] , \wRegInTop_6_8[23] , 
        \wRegInBot_6_35[0] , \wRegOut_7_91[22] , \wRegInTop_7_111[22] , 
        \wRegInBot_0_0[25] , \wRegInTop_1_0[19] , \ScanLink12[22] , 
        \ScanLink24[27] , \ScanLink72[26] , \wRegInTop_6_14[18] , 
        \wRegInTop_6_37[30] , \wRegOut_7_56[4] , \wRegInTop_6_61[28] , 
        \ScanLink31[13] , \ScanLink51[17] , \wRegInTop_6_37[29] , 
        \wRegInTop_6_42[19] , \wRegInTop_6_61[31] , \wRegInTop_7_39[19] , 
        \wRegInTop_7_59[3] , \ScanLink34[0] , \ScanLink44[23] , 
        \ScanLink219[26] , \wRegOut_5_26[0] , \wRegInTop_4_4[4] , 
        \wRegInBot_4_6[1] , \wRegInTop_4_7[7] , \wRegOut_7_84[2] , 
        \wRegOut_5_2[8] , \ScanLink67[12] , \ScanLink89[27] , \ScanLink109[1] , 
        \ScanLink127[24] , \ScanLink152[14] , \wRegInTop_7_95[9] , 
        \ScanLink104[15] , \ScanLink171[25] , \wRegInTop_7_94[19] , 
        \ScanLink164[11] , \wRegInBot_4_5[2] , \wRegInTop_5_19[29] , 
        \wRegInTop_7_7[20] , \ScanLink111[21] , \wRegOut_7_48[8] , 
        \wRegOut_7_87[1] , \ScanLink31[20] , \wRegInTop_5_0[24] , 
        \ScanLink37[3] , \wRegInTop_5_19[30] , \ScanLink147[20] , 
        \wRegOut_5_25[3] , \ScanLink132[10] , \wRegOut_6_11[23] , 
        \wRegOut_6_27[26] , \wRegOut_6_52[16] , \wRegOut_7_29[16] , 
        \wRegInBot_6_36[3] , \wRegInTop_7_88[6] , \wRegOut_7_55[7] , 
        \ScanLink44[10] , \wRegOut_6_32[12] , \wRegOut_6_47[22] , 
        \wRegOut_7_49[12] , \wRegInTop_7_3[6] , \ScanLink219[15] , 
        \ScanLink67[21] , \wRegOut_7_112[29] , \wRegInTop_1_0[1] , 
        \wRegInBot_1_1[7] , \wRegInBot_3_2[17] , \ScanLink12[11] , 
        \wRegOut_7_112[30] , \ScanLink24[14] , \ScanLink51[24] , 
        \ScanLink72[15] , \wRegInBot_6_22[30] , \wRegInBot_6_22[29] , 
        \wRegInBot_6_57[19] , \wRegInTop_7_121[5] , \wRegOut_4_12[11] , 
        \ScanLink50[4] , \wRegInTop_6_8[10] , \wRegInTop_7_20[8] , 
        \ScanLink173[9] , \wRegOut_7_91[11] , \wRegInBot_6_51[4] , 
        \wRegInTop_7_111[11] , \wRegOut_6_13[6] , \wRegInTop_7_104[25] , 
        \wRegInTop_5_0[17] , \wRegOut_6_11[10] , \ScanLink82[2] , 
        \wRegOut_7_32[0] , \wRegOut_7_84[25] , \wRegInTop_7_127[14] , 
        \wRegOut_6_32[21] , \wRegOut_7_49[21] , \wRegOut_6_47[11] , 
        \wRegOut_6_10[5] , \ScanLink81[1] , \wRegOut_6_27[15] , 
        \wRegOut_7_115[9] , \wRegOut_6_52[25] , \wRegOut_7_29[25] , 
        \wRegInBot_6_52[7] , \ScanLink111[12] , \wRegOut_7_31[3] , 
        \wRegInTop_7_0[5] , \wRegInTop_7_7[13] , \ScanLink164[22] , 
        \ScanLink132[23] , \ScanLink147[13] , \ScanLink53[7] , 
        \wRegOut_6_6[9] , \wRegEnTop_6_51[0] , \ScanLink127[17] , 
        \wRegOut_7_108[6] , \wRegInTop_7_122[6] , \ScanLink89[14] , 
        \ScanLink104[26] , \ScanLink152[27] , \wRegOut_6_58[10] , 
        \wRegOut_7_1[31] , \ScanLink171[16] , \wRegOut_7_75[11] , 
        \ScanLink45[3] , \wRegInBot_5_15[1] , \wRegOut_7_1[28] , 
        \wRegOut_7_23[10] , \wRegInTop_7_28[0] , \wRegOut_7_56[20] , 
        \wRegOut_7_36[24] , \wRegOut_7_43[14] , \wRegOut_6_38[14] , 
        \wRegOut_7_15[15] , \wRegInBot_0_0[16] , \wRegInTop_2_2[18] , 
        \wRegOut_3_1[26] , \wRegInBot_5_13[31] , \wRegInBot_5_13[28] , 
        \ScanLink83[21] , \wRegOut_7_60[25] , \wRegInBot_5_30[19] , 
        \ScanLink158[12] , \wRegInTop_6_14[9] , \ScanLink96[15] , 
        \ScanLink97[5] , \ScanLink138[16] , \wRegInBot_6_44[3] , 
        \wRegOut_7_27[7] , \ScanLink206[14] , \ScanLink250[15] , 
        \ScanLink18[24] , \ScanLink78[20] , \wRegInBot_6_47[0] , 
        \ScanLink180[22] , \ScanLink225[25] , \ScanLink245[21] , 
        \wRegInTop_4_5[21] , \wRegOut_7_24[4] , \ScanLink205[8] , 
        \ScanLink230[11] , \ScanLink195[16] , \ScanLink46[0] , 
        \wRegOut_5_16[14] , \ScanLink94[6] , \wRegInBot_6_48[18] , 
        \ScanLink213[20] , \ScanLink178[2] , \wRegInBot_5_16[2] , 
        \wRegInTop_6_2[25] , \ScanLink218[7] , \wRegOut_5_20[11] , 
        \ScanLink89[9] , \ScanLink138[25] , \wRegOut_5_9[3] , 
        \wRegInTop_5_25[19] , \ScanLink83[12] , \wRegInBot_6_20[7] , 
        \ScanLink96[26] , \wRegOut_6_62[5] , \wRegOut_7_43[3] , 
        \wRegOut_6_38[27] , \ScanLink158[21] , \wRegOut_7_43[27] , 
        \wRegOut_7_15[26] , \wRegOut_7_36[17] , \wRegOut_7_60[16] , 
        \wRegOut_7_56[13] , \wRegOut_7_75[22] , \wRegOut_7_91[5] , 
        \ScanLink1[26] , \ScanLink1[15] , \ScanLink2[1] , \wRegOut_3_1[15] , 
        \ScanLink18[17] , \ScanLink21[7] , \wRegOut_4_12[1] , 
        \wRegOut_6_58[23] , \ScanLink22[4] , \wRegOut_5_20[22] , 
        \wRegInTop_6_2[16] , \wRegEnTop_6_23[0] , \wRegOut_7_23[23] , 
        \wRegOut_4_11[2] , \wRegOut_5_16[27] , \wRegOut_5_30[4] , 
        \wRegInTop_6_28[31] , \ScanLink195[25] , \wRegOut_7_92[6] , 
        \ScanLink230[22] , \ScanLink245[12] , \wRegInTop_4_5[12] , 
        \wRegInTop_6_28[28] , \ScanLink101[9] , \wRegInTop_7_26[18] , 
        \wRegInTop_7_53[31] , \wRegInTop_7_70[19] , \ScanLink213[13] , 
        \wRegInTop_7_52[8] , \wRegInTop_7_53[28] , \ScanLink206[27] , 
        \wRegInBot_4_0[18] , \wRegEnBot_4_8[0] , \ScanLink78[13] , 
        \wRegInBot_6_23[4] , \wRegOut_6_61[6] , \wRegOut_7_40[0] , 
        \ScanLink180[11] , \ScanLink225[16] , \ScanLink250[26] , 
        \wRegInTop_5_18[10] , \wRegEnBot_6_11[0] , \ScanLink110[18] , 
        \ScanLink133[30] , \ScanLink133[29] , \ScanLink146[19] , 
        \ScanLink165[31] , \wRegInTop_7_80[14] , \ScanLink165[28] , 
        \wRegInTop_7_6[19] , \wRegInTop_7_95[20] , \wRegInBot_5_4[17] , 
        \wRegInBot_5_18[17] , \wRegInTop_6_12[7] , \ScanLink160[0] , 
        \wRegInTop_7_33[1] , \ScanLink1[2] , \wRegInTop_1_1[13] , 
        \wRegInTop_3_6[17] , \wRegOut_7_21[9] , \ScanLink200[5] , 
        \wRegOut_7_105[3] , \wRegOut_4_2[10] , \wRegInTop_6_11[4] , 
        \ScanLink92[8] , \wRegInTop_7_30[2] , \ScanLink163[3] , 
        \wRegOut_7_106[0] , \ScanLink203[6] , \wRegOut_6_5[14] , 
        \wRegInBot_6_15[26] , \wRegInTop_6_23[24] , \wRegInBot_6_36[17] , 
        \wRegInTop_6_56[14] , \wRegInBot_6_60[16] , \wRegInBot_6_23[23] , 
        \wRegInBot_6_43[27] , \wRegInTop_7_58[24] , \wRegOut_7_113[23] , 
        \wRegInTop_6_43[20] , \wRegInTop_7_38[20] , \wRegInBot_6_56[13] , 
        \wRegOut_7_106[17] , \wRegInTop_6_36[10] , \wRegInTop_6_60[11] , 
        \wRegInTop_6_15[21] , \wRegOut_7_125[26] , \ScanLink0[12] , 
        \wRegInBot_1_0[31] , \wRegInBot_1_0[28] , \wRegInTop_1_1[20] , 
        \ScanLink13[28] , \wRegInBot_4_8[7] , \wRegInTop_4_9[1] , 
        \wRegInBot_5_4[24] , \wRegOut_5_28[6] , \ScanLink104[4] , 
        \wRegInTop_7_57[5] , \wRegOut_6_46[28] , \wRegOut_7_48[18] , 
        \wRegOut_6_10[30] , \wRegOut_6_33[18] , \wRegInBot_6_26[9] , 
        \wRegOut_6_46[31] , \ScanLink27[9] , \wRegInBot_5_18[24] , 
        \wRegInTop_5_27[1] , \wRegOut_6_10[29] , \wRegInTop_7_95[13] , 
        \wRegInTop_7_85[3] , \wRegInTop_5_18[23] , \wRegInTop_5_24[2] , 
        \wRegOut_6_5[27] , \wRegInBot_6_56[20] , \wRegOut_7_58[2] , 
        \wRegInTop_7_80[27] , \wRegInTop_6_15[12] , \wRegInBot_6_23[10] , 
        \wRegInTop_6_36[23] , \wRegOut_7_106[24] , \wRegInTop_7_38[13] , 
        \wRegInTop_7_86[0] , \wRegInTop_6_43[13] , \wRegInTop_7_49[9] , 
        \wRegOut_7_125[15] , \wRegInTop_6_60[22] , \wRegInBot_6_38[5] , 
        \wRegInBot_6_60[25] , \ScanLink66[18] , \wRegOut_7_94[8] , 
        \wRegInBot_6_15[15] , \wRegOut_2_1[18] , \wRegOut_2_1[0] , 
        \ScanLink13[31] , \ScanLink30[19] , \ScanLink45[30] , 
        \wRegInTop_6_23[17] , \wRegInBot_6_43[14] , \wRegInTop_7_58[17] , 
        \wRegOut_7_113[10] , \wRegInTop_3_6[24] , \wRegOut_4_2[23] , 
        \wRegOut_4_13[31] , \ScanLink45[29] , \wRegInBot_6_36[24] , 
        \wRegInTop_6_56[27] , \wRegOut_4_13[28] , \ScanLink107[7] , 
        \wRegInTop_7_54[6] , \ScanLink39[5] , \wRegInTop_6_9[30] , 
        \wRegInTop_6_9[29] , \wRegOut_7_90[28] , \wRegInTop_7_110[28] , 
        \wRegOut_7_89[7] , \wRegOut_7_90[31] , \wRegInTop_7_110[31] , 
        \wRegOut_6_1[16] , \wRegInBot_6_27[21] , \wRegInTop_6_47[22] , 
        \ScanLink209[29] , \wRegInTop_7_49[12] , \wRegOut_7_102[15] , 
        \wRegInTop_6_32[12] , \wRegInBot_6_52[11] , \ScanLink209[30] , 
        \wRegInTop_3_2[15] , \wRegEnBot_3_3[0] , \wRegOut_4_1[4] , 
        \wRegInTop_5_7[8] , \ScanLink62[29] , \wRegInTop_6_11[23] , 
        \wRegOut_7_121[24] , \wRegInBot_6_11[24] , \ScanLink17[19] , 
        \ScanLink34[31] , \wRegOut_4_6[12] , \ScanLink34[28] , 
        \ScanLink41[18] , \wRegInTop_6_52[16] , \ScanLink62[30] , 
        \wRegInBot_6_32[15] , \wRegInTop_7_29[16] , \wRegInTop_6_27[26] , 
        \wRegInBot_6_47[25] , \wRegOut_7_117[21] , \wRegOut_5_19[30] , 
        \wRegInBot_6_8[12] , \wRegOut_5_19[29] , \wRegOut_7_62[8] , 
        \ScanLink243[4] , \wRegOut_7_94[19] , \wRegInTop_7_114[19] , 
        \wRegInTop_6_51[6] , \ScanLink123[1] , \wRegInTop_7_70[0] , 
        \ScanLink5[17] , \wRegInBot_5_0[15] , \wRegOut_2_2[3] , 
        \wRegOut_6_14[18] , \wRegOut_6_37[29] , \ScanLink240[7] , 
        \wRegOut_6_42[19] , \ScanLink120[2] , \wRegOut_7_39[19] , 
        \wRegInTop_6_52[5] , \wRegOut_6_61[31] , \wRegInTop_7_73[3] , 
        \wRegOut_6_37[30] , \wRegOut_6_61[28] , \wRegInTop_3_2[26] , 
        \wRegInBot_3_5[9] , \wRegInTop_4_12[22] , \wRegInBot_4_12[25] , 
        \wRegInTop_7_91[22] , \wRegOut_5_9[11] , \ScanLink99[31] , 
        \wRegInTop_7_84[16] , \wRegOut_4_2[7] , \wRegInBot_5_29[5] , 
        \ScanLink99[28] , \ScanLink227[0] , \wRegInTop_7_108[6] , 
        \wRegOut_7_122[6] , \ScanLink79[7] , \wRegOut_4_6[21] , 
        \wRegInBot_6_8[21] , \wRegInTop_6_35[2] , \wRegInTop_7_14[4] , 
        \ScanLink147[5] , \ScanLink64[8] , \wRegInBot_6_11[17] , 
        \wRegInTop_6_27[15] , \wRegInBot_6_47[16] , \wRegInTop_7_115[9] , 
        \wRegOut_7_117[12] , \wRegOut_7_5[5] , \wRegInBot_6_32[26] , 
        \wRegInTop_6_52[25] , \wRegEnTop_7_88[0] , \wRegInTop_7_29[25] , 
        \wRegOut_6_1[25] , \wRegInTop_6_3[9] , \wRegInBot_6_27[12] , 
        \wRegInTop_6_32[21] , \wRegInBot_6_52[22] , \wRegInTop_7_49[21] , 
        \wRegOut_7_102[26] , \wRegInTop_6_47[11] , \ScanLink195[3] , 
        \wRegOut_7_121[17] , \wRegInBot_2_0[6] , \ScanLink5[24] , 
        \wRegInTop_4_12[11] , \wRegInTop_6_11[10] , \ScanLink114[30] , 
        \wRegInTop_7_2[31] , \ScanLink142[28] , \ScanLink114[29] , 
        \wRegInTop_7_2[28] , \wRegOut_7_6[6] , \ScanLink137[18] , 
        \ScanLink142[31] , \ScanLink161[19] , \wRegOut_7_18[0] , 
        \wRegInBot_4_12[16] , \wRegOut_6_39[6] , \wRegInTop_7_84[25] , 
        \wRegOut_5_9[22] , \wRegEnTop_6_5[0] , \wRegInTop_7_91[11] , 
        \wRegOut_6_24[9] , \ScanLink159[9] , \ScanLink196[0] , 
        \wRegOut_7_121[5] , \ScanLink224[3] , \wRegInTop_2_2[3] , 
        \wRegInBot_2_3[23] , \wRegInBot_3_0[4] , \wRegInTop_3_1[2] , 
        \wRegInBot_5_0[26] , \wRegInBot_5_0[0] , \wRegInTop_6_36[1] , 
        \wRegInTop_7_17[7] , \ScanLink144[6] , \wRegInTop_5_1[6] , 
        \wRegInTop_6_6[27] , \wRegOut_7_79[9] , \wRegOut_5_14[2] , 
        \wRegOut_5_24[13] , \wRegOut_5_31[27] , \ScanLink138[0] , 
        \wRegOut_3_5[24] , \wRegInTop_4_1[23] , \wRegOut_5_12[16] , 
        \ScanLink69[16] , \wRegOut_6_45[0] , \wRegInTop_7_74[28] , 
        \ScanLink241[23] , \wRegInTop_6_59[30] , \ScanLink191[14] , 
        \wRegOut_7_64[6] , \ScanLink234[13] , \wRegInTop_7_22[30] , 
        \wRegInBot_4_4[30] , \wRegInTop_6_59[29] , \wRegInTop_7_57[19] , 
        \wRegInTop_7_74[31] , \ScanLink217[22] , \wRegInTop_7_22[29] , 
        \wRegInBot_4_4[29] , \wRegEnBot_6_49[0] , \wRegInTop_6_57[8] , 
        \ScanLink202[16] , \ScanLink254[17] , \ScanLink92[17] , 
        \wRegInTop_7_9[24] , \ScanLink149[24] , \ScanLink184[20] , 
        \ScanLink221[27] , \wRegOut_6_46[3] , \wRegOut_7_67[5] , 
        \ScanLink246[9] , \wRegInBot_2_3[10] , \wRegInTop_3_2[1] , 
        \wRegInTop_5_2[5] , \wRegInBot_5_3[3] , \wRegOut_5_17[1] , 
        \wRegInTop_5_18[6] , \wRegInTop_5_21[31] , \ScanLink87[23] , 
        \wRegInTop_5_21[28] , \wRegOut_6_49[26] , \ScanLink129[20] , 
        \wRegOut_7_32[26] , \wRegEnTop_7_26[0] , \wRegOut_7_47[16] , 
        \wRegOut_7_11[17] , \wRegOut_7_64[27] , \wRegInBot_3_3[7] , 
        \wRegOut_4_4[9] , \wRegOut_7_71[13] , \wRegOut_3_5[17] , 
        \wRegOut_6_29[22] , \wRegOut_7_27[12] , \wRegInTop_6_49[4] , 
        \wRegOut_7_52[22] , \wRegInTop_7_68[2] , \ScanLink202[25] , 
        \wRegOut_7_124[8] , \wRegOut_7_109[19] , \wRegInTop_4_1[10] , 
        \ScanLink69[25] , \wRegOut_6_21[4] , \wRegInBot_6_63[6] , 
        \ScanLink184[13] , \ScanLink221[14] , \ScanLink254[24] , 
        \ScanLink191[27] , \ScanLink234[20] , \wRegInBot_6_39[19] , 
        \ScanLink217[11] , \ScanLink241[10] , \wRegInBot_4_10[1] , 
        \wRegInBot_4_13[2] , \wRegOut_5_12[25] , \ScanLink62[6] , 
        \wRegOut_5_31[14] , \wRegInTop_7_113[7] , \wRegOut_5_24[20] , 
        \wRegInTop_6_6[14] , \wRegEnTop_7_119[0] , \wRegInBot_6_4[1] , 
        \wRegInTop_6_5[7] , \wRegOut_6_29[11] , \wRegOut_7_71[20] , 
        \wRegOut_7_52[11] , \wRegInTop_7_110[4] , \wRegInBot_5_17[19] , 
        \ScanLink61[5] , \wRegInBot_5_31[7] , \wRegOut_7_0[8] , 
        \wRegOut_7_5[19] , \wRegInTop_6_6[4] , \wRegInBot_6_7[2] , 
        \wRegOut_7_27[21] , \wRegOut_6_49[15] , \wRegOut_7_32[15] , 
        \wRegOut_7_47[25] , \wRegOut_7_11[24] , \wRegOut_7_64[14] , 
        \ScanLink87[10] , \wRegInBot_6_60[5] , \wRegInBot_2_3[5] , 
        \wRegOut_3_0[21] , \ScanLink9[7] , \wRegInTop_5_12[31] , 
        \wRegInBot_5_18[9] , \ScanLink55[4] , \wRegInTop_6_19[1] , 
        \wRegOut_6_22[7] , \ScanLink92[24] , \ScanLink129[13] , 
        \wRegInTop_7_9[17] , \wRegInTop_7_11[9] , \ScanLink149[17] , 
        \ScanLink142[8] , \wRegOut_6_59[17] , \wRegOut_7_74[16] , 
        \wRegInTop_7_6[6] , \wRegOut_7_22[17] , \wRegOut_7_37[23] , 
        \wRegInTop_7_38[7] , \wRegOut_7_57[27] , \wRegOut_7_42[13] , 
        \wRegInTop_7_124[5] , \ScanLink82[26] , \wRegOut_6_39[13] , 
        \wRegOut_7_14[12] , \wRegOut_7_61[22] , \wRegInTop_7_25[8] , 
        \ScanLink159[15] , \ScanLink176[9] , \wRegInTop_5_31[19] , 
        \ScanLink87[2] , \ScanLink139[11] , \wRegInBot_6_54[4] , 
        \wRegInTop_5_12[28] , \ScanLink79[27] , \wRegOut_6_16[6] , 
        \ScanLink97[12] , \wRegInTop_6_49[18] , \wRegInTop_7_11[30] , 
        \wRegInTop_7_32[18] , \wRegOut_7_37[0] , \wRegInTop_7_47[28] , 
        \wRegInTop_7_47[31] , \wRegInTop_7_64[19] , \ScanLink207[13] , 
        \ScanLink251[12] , \wRegInTop_7_11[29] , \ScanLink19[23] , 
        \wRegInBot_6_57[7] , \ScanLink181[25] , \ScanLink224[22] , 
        \ScanLink244[26] , \wRegInTop_4_4[26] , \wRegOut_6_15[5] , 
        \wRegOut_7_34[3] , \ScanLink194[11] , \ScanLink231[16] , 
        \wRegOut_4_8[31] , \ScanLink84[1] , \ScanLink212[27] , 
        \wRegOut_7_110[9] , \wRegOut_4_8[28] , \wRegInBot_6_6[28] , 
        \wRegInTop_7_5[5] , \ScanLink168[5] , \wRegOut_5_7[18] , 
        \wRegOut_5_17[13] , \wRegInBot_6_6[31] , \wRegOut_5_21[16] , 
        \wRegOut_6_3[9] , \wRegInTop_6_3[22] , \ScanLink208[0] , 
        \wRegInTop_7_127[6] , \wRegInBot_5_24[19] , \ScanLink56[7] , 
        \wRegEnTop_6_54[0] , \ScanLink82[15] , \wRegInBot_6_30[0] , 
        \ScanLink97[21] , \ScanLink139[22] , \wRegOut_7_53[4] , 
        \wRegOut_6_39[20] , \ScanLink159[26] , \wRegOut_7_42[20] , 
        \wRegOut_7_37[10] , \wRegOut_7_61[11] , \wRegInTop_5_31[8] , 
        \wRegOut_7_14[21] , \wRegInTop_4_2[7] , \wRegInBot_4_3[1] , 
        \wRegOut_7_74[25] , \wRegOut_7_81[2] , \ScanLink31[0] , 
        \wRegOut_5_23[0] , \wRegOut_6_59[24] , \wRegOut_7_57[14] , 
        \wRegOut_7_22[24] , \wRegInTop_2_1[0] , \wRegOut_5_7[8] , 
        \wRegOut_3_0[12] , \wRegInBot_4_0[2] , \wRegInTop_4_1[4] , 
        \ScanLink32[3] , \wRegOut_5_21[25] , \wRegInTop_6_3[11] , 
        \wRegInTop_7_90[9] , \wRegOut_5_17[20] , \wRegOut_5_20[3] , 
        \wRegOut_7_82[1] , \ScanLink19[10] , \ScanLink194[22] , 
        \ScanLink231[25] , \ScanLink244[15] , \wRegInTop_4_4[15] , 
        \wRegInTop_6_63[9] , \ScanLink212[14] , \wRegOut_7_119[31] , 
        \ScanLink79[14] , \wRegInBot_6_29[28] , \wRegOut_7_119[28] , 
        \ScanLink207[20] , \wRegInBot_5_5[10] , \wRegInTop_5_19[17] , 
        \wRegInBot_6_29[31] , \wRegInBot_6_33[3] , \wRegInTop_7_0[8] , 
        \wRegOut_7_50[7] , \ScanLink181[16] , \ScanLink224[11] , 
        \ScanLink251[21] , \wRegInTop_7_81[13] , \wRegInBot_5_19[10] , 
        \wRegInTop_7_94[27] , \wRegOut_6_6[4] , \ScanLink89[19] , 
        \wRegInTop_7_23[6] , \ScanLink170[7] , \wRegOut_6_10[8] , 
        \wRegOut_6_52[31] , \ScanLink210[2] , \wRegOut_6_27[18] , 
        \wRegOut_7_29[31] , \wRegOut_6_52[28] , \wRegOut_7_115[4] , 
        \wRegOut_7_29[28] , \ScanLink0[21] , \wRegInTop_1_0[14] , 
        \wRegInTop_3_7[10] , \wRegOut_4_3[17] , \wRegInBot_6_51[9] , 
        \wRegInTop_7_20[5] , \ScanLink173[4] , \wRegOut_7_84[31] , 
        \wRegInTop_7_104[31] , \wRegOut_7_116[7] , \wRegInTop_7_127[19] , 
        \ScanLink213[1] , \wRegOut_7_84[28] , \wRegInTop_7_104[28] , 
        \ScanLink24[19] , \ScanLink51[29] , \wRegInBot_6_14[21] , 
        \wRegInTop_6_22[23] , \wRegInBot_6_37[10] , \wRegInTop_6_57[13] , 
        \wRegInBot_6_61[11] , \ScanLink219[18] , \wRegInBot_6_22[24] , 
        \wRegInBot_6_42[20] , \wRegInTop_7_59[23] , \wRegOut_7_112[24] , 
        \wRegOut_6_5[7] , \wRegInTop_7_39[27] , \wRegInTop_7_121[8] , 
        \wRegInTop_6_42[27] , \ScanLink50[9] , \wRegOut_6_4[13] , 
        \wRegOut_7_107[10] , \wRegInTop_6_37[17] , \wRegInBot_6_57[14] , 
        \ScanLink51[30] , \ScanLink72[18] , \wRegInTop_6_14[26] , 
        \wRegInTop_6_61[16] , \wRegOut_7_124[21] , \wRegInTop_1_0[27] , 
        \wRegOut_3_1[2] , \wRegOut_3_2[1] , \wRegInTop_4_4[9] , 
        \wRegInTop_5_0[30] , \wRegInTop_5_0[29] , \wRegInBot_5_5[23] , 
        \ScanLink114[3] , \wRegInTop_7_47[2] , \wRegOut_5_2[5] , 
        \wRegInBot_5_19[23] , \ScanLink104[18] , \ScanLink127[30] , 
        \ScanLink171[28] , \wRegInTop_7_94[14] , \ScanLink127[29] , 
        \ScanLink152[19] , \ScanLink171[31] , \wRegInTop_7_95[4] , 
        \wRegInTop_5_19[24] , \wRegOut_7_48[5] , \wRegEnTop_4_2[0] , 
        \wRegInTop_4_15[3] , \wRegOut_5_1[6] , \wRegOut_6_4[20] , 
        \wRegInTop_7_81[20] , \wRegInBot_6_22[17] , \wRegInTop_6_37[24] , 
        \wRegInBot_6_57[27] , \wRegOut_7_107[23] , \wRegInTop_7_39[14] , 
        \wRegInTop_7_96[7] , \wRegInTop_6_42[14] , \wRegOut_7_124[12] , 
        \wRegInTop_6_14[15] , \wRegInBot_6_28[2] , \wRegInTop_6_61[25] , 
        \wRegInBot_6_61[22] , \wRegInBot_6_14[12] , \wRegInBot_3_2[30] , 
        \wRegInTop_6_22[10] , \wRegInBot_6_37[23] , \wRegInBot_6_42[13] , 
        \wRegInTop_7_59[10] , \wRegOut_7_112[17] , \wRegInTop_6_57[20] , 
        \wRegInBot_3_2[29] , \ScanLink117[0] , \wRegInTop_7_44[1] , 
        \wRegOut_4_3[24] , \wRegOut_7_99[0] , \wRegInBot_0_0[31] , 
        \wRegInBot_0_0[28] , \wRegOut_1_0[1] , \wRegInBot_1_0[25] , 
        \ScanLink4[23] , \ScanLink4[10] , \wRegInTop_3_3[12] , 
        \wRegInBot_3_6[18] , \wRegInTop_3_7[23] , \ScanLink29[2] , 
        \wRegOut_7_56[9] , \wRegOut_4_7[15] , \wRegInTop_5_10[3] , 
        \wRegOut_6_0[11] , \wRegInBot_6_26[26] , \wRegInTop_6_46[25] , 
        \wRegInBot_6_53[16] , \wRegInTop_7_48[15] , \wRegOut_7_103[12] , 
        \wRegInTop_6_10[24] , \wRegInTop_6_33[15] , \wRegOut_7_120[23] , 
        \wRegInBot_6_10[23] , \wRegInBot_6_9[15] , \wRegInTop_6_26[21] , 
        \wRegInBot_6_33[12] , \wRegInTop_6_53[11] , \wRegInTop_7_28[11] , 
        \wRegInBot_6_46[22] , \wRegOut_7_116[26] , \wRegOut_6_53[9] , 
        \ScanLink253[3] , \wRegInBot_5_1[12] , \wRegInBot_5_8[5] , 
        \wRegInTop_6_41[1] , \ScanLink133[6] , \wRegInTop_7_60[7] , 
        \wRegInBot_6_12[8] , \wRegInTop_3_3[21] , \ScanLink13[8] , 
        \wRegInBot_4_13[22] , \wRegInTop_5_4[18] , \wRegInTop_5_9[3] , 
        \ScanLink250[0] , \ScanLink130[5] , \wRegOut_5_8[16] , 
        \ScanLink100[29] , \wRegInTop_6_42[2] , \wRegInTop_7_63[4] , 
        \wRegInTop_7_90[25] , \ScanLink100[30] , \ScanLink156[31] , 
        \ScanLink175[19] , \ScanLink123[18] , \wRegInTop_4_13[25] , 
        \ScanLink156[28] , \wRegInTop_5_13[0] , \wRegInTop_7_85[11] , 
        \ScanLink69[0] , \ScanLink237[7] , \wRegInTop_7_118[1] , 
        \ScanLink20[31] , \ScanLink20[28] , \wRegOut_4_7[26] , 
        \wRegInBot_6_9[26] , \wRegInTop_7_123[28] , \wRegInTop_6_25[5] , 
        \ScanLink157[2] , \wRegInTop_7_100[19] , \wRegOut_6_0[22] , 
        \wRegInBot_6_10[10] , \wRegOut_7_80[19] , \wRegInTop_7_123[31] , 
        \wRegInTop_6_26[12] , \wRegInBot_6_33[21] , \wRegInBot_6_46[11] , 
        \wRegOut_7_116[15] , \wRegInTop_6_53[22] , \wRegInBot_6_53[25] , 
        \wRegInTop_7_28[22] , \wRegOut_7_103[21] , \ScanLink55[18] , 
        \wRegInTop_6_33[26] , \wRegInTop_7_48[26] , \ScanLink76[30] , 
        \wRegInBot_6_26[15] , \wRegInTop_6_46[16] , \ScanLink185[4] , 
        \wRegOut_7_120[10] , \wRegInTop_4_13[16] , \wRegInTop_6_10[17] , 
        \ScanLink76[29] , \wRegOut_6_29[1] , \wRegInBot_4_13[11] , 
        \wRegOut_5_8[25] , \wRegInTop_7_85[22] , \wRegOut_7_15[8] , 
        \ScanLink186[7] , \wRegInTop_7_90[16] , \ScanLink234[4] , 
        \wRegOut_2_1[26] , \ScanLink5[30] , \wRegInBot_2_2[24] , 
        \wRegOut_3_4[23] , \wRegInTop_4_0[24] , \ScanLink16[5] , 
        \wRegInBot_5_1[21] , \wRegOut_5_25[14] , \wRegInTop_6_7[20] , 
        \wRegOut_6_23[30] , \wRegOut_6_23[29] , \wRegOut_6_56[19] , 
        \wRegOut_7_58[30] , \wRegInTop_6_26[6] , \ScanLink154[1] , 
        \wRegOut_7_58[29] , \wRegOut_6_48[8] , \ScanLink248[2] , 
        \wRegOut_5_13[11] , \wRegOut_5_30[20] , \ScanLink128[7] , 
        \ScanLink68[11] , \wRegInBot_6_17[5] , \ScanLink240[24] , 
        \wRegOut_6_55[7] , \ScanLink190[13] , \wRegOut_7_74[1] , 
        \ScanLink235[14] , \wRegInBot_6_58[30] , \wRegInBot_6_58[29] , 
        \ScanLink216[25] , \ScanLink135[8] , \wRegInTop_7_66[9] , 
        \ScanLink203[11] , \ScanLink255[10] , \wRegInBot_5_20[31] , 
        \wRegInBot_5_20[28] , \ScanLink148[23] , \ScanLink185[27] , 
        \ScanLink220[20] , \wRegInBot_6_14[6] , \ScanLink93[10] , 
        \wRegInTop_7_8[23] , \wRegOut_6_56[4] , \wRegOut_7_77[2] , 
        \wRegInBot_2_2[17] , \wRegOut_3_4[10] , \ScanLink15[6] , 
        \wRegOut_4_9[1] , \wRegOut_5_3[29] , \ScanLink86[24] , 
        \wRegOut_5_3[30] , \wRegOut_6_48[21] , \ScanLink128[27] , 
        \wRegOut_7_33[21] , \wRegOut_7_46[11] , \wRegOut_6_28[25] , 
        \wRegOut_7_10[10] , \wRegOut_7_26[15] , \wRegOut_7_65[20] , 
        \wRegOut_7_70[14] , \wRegInTop_6_38[19] , \wRegInTop_6_59[3] , 
        \wRegInTop_7_36[29] , \wRegOut_7_53[25] , \wRegInTop_7_78[5] , 
        \wRegInTop_7_43[19] , \ScanLink203[22] , \wRegInTop_7_60[31] , 
        \wRegInTop_4_0[17] , \ScanLink68[22] , \wRegOut_6_31[3] , 
        \wRegOut_7_10[5] , \wRegInTop_7_15[18] , \wRegInTop_7_36[30] , 
        \ScanLink185[14] , \ScanLink220[13] , \wRegInTop_7_60[28] , 
        \ScanLink255[23] , \ScanLink231[9] , \ScanLink190[20] , 
        \ScanLink235[27] , \wRegInBot_6_9[9] , \ScanLink216[16] , 
        \ScanLink240[17] , \wRegOut_5_13[22] , \wRegInBot_5_22[3] , 
        \wRegInBot_6_2[19] , \wRegInTop_7_103[0] , \wRegOut_5_30[13] , 
        \ScanLink72[1] , \wRegEnTop_7_51[0] , \wRegInBot_5_21[0] , 
        \wRegOut_5_25[27] , \wRegInTop_6_7[13] , \wRegOut_6_28[16] , 
        \wRegOut_7_70[27] , \wRegOut_7_53[16] , \wRegInTop_7_100[3] , 
        \ScanLink71[2] , \ScanLink86[17] , \wRegOut_6_48[12] , 
        \wRegOut_7_26[26] , \wRegOut_7_33[12] , \wRegOut_7_46[22] , 
        \ScanLink180[9] , \wRegOut_7_10[23] , \wRegOut_7_65[13] , 
        \wRegOut_7_13[6] , \wRegInTop_5_5[21] , \wRegInTop_5_16[19] , 
        \wRegInTop_6_20[8] , \wRegOut_6_32[0] , \ScanLink128[14] , 
        \ScanLink93[23] , \wRegInTop_7_8[10] , \ScanLink148[10] , 
        \wRegOut_6_14[26] , \wRegOut_6_24[4] , \wRegOut_6_61[16] , 
        \wRegOut_7_39[27] , \wRegOut_6_37[17] , \wRegOut_6_42[27] , 
        \wRegOut_7_121[8] , \ScanLink5[29] , \wRegOut_6_22[23] , 
        \wRegOut_6_57[13] , \wRegOut_7_59[23] , \ScanLink17[27] , 
        \wRegInBot_4_15[1] , \wRegInTop_6_0[7] , \wRegInBot_6_1[1] , 
        \ScanLink67[6] , \ScanLink99[16] , \ScanLink161[14] , 
        \ScanLink114[24] , \wRegInTop_7_2[25] , \ScanLink239[1] , 
        \ScanLink137[15] , \ScanLink142[25] , \wRegInTop_7_84[28] , 
        \wRegInTop_7_116[7] , \wRegInTop_7_84[31] , \ScanLink157[11] , 
        \ScanLink101[10] , \ScanLink122[21] , \ScanLink159[4] , 
        \ScanLink174[20] , \wRegInTop_7_115[4] , \ScanLink34[16] , 
        \wRegInTop_6_27[18] , \ScanLink41[26] , \ScanLink64[5] , 
        \wRegInTop_6_52[28] , \wRegOut_7_5[8] , \wRegInTop_7_29[28] , 
        \ScanLink21[22] , \ScanLink62[17] , \wRegInTop_6_52[31] , 
        \wRegInTop_7_29[31] , \wRegOut_6_1[31] , \ScanLink77[23] , 
        \wRegInBot_1_0[16] , \wRegOut_2_1[15] , \wRegInTop_3_4[2] , 
        \wRegInBot_3_7[21] , \ScanLink54[12] , \wRegOut_6_1[28] , 
        \wRegInBot_6_2[2] , \wRegInTop_6_3[4] , \wRegInBot_5_29[8] , 
        \wRegInTop_6_28[0] , \ScanLink209[17] , \wRegOut_6_27[7] , 
        \wRegOut_7_94[27] , \wRegInTop_7_114[27] , \wRegInBot_4_12[31] , 
        \wRegOut_5_19[17] , \wRegOut_7_81[13] , \wRegInTop_7_101[13] , 
        \ScanLink122[12] , \wRegInTop_7_14[9] , \ScanLink147[8] , 
        \wRegInTop_7_122[22] , \ScanLink188[1] , \wRegInBot_4_12[28] , 
        \wRegInBot_5_5[0] , \wRegOut_5_11[2] , \ScanLink157[22] , 
        \ScanLink101[23] , \wRegInTop_5_4[6] , \ScanLink174[13] , 
        \ScanLink114[17] , \wRegInBot_3_5[4] , \ScanLink99[25] , 
        \ScanLink161[27] , \wRegInTop_7_2[16] , \wRegOut_6_22[10] , 
        \ScanLink137[26] , \ScanLink142[16] , \wRegOut_6_57[20] , 
        \wRegOut_7_59[10] , \wRegInTop_3_2[18] , \wRegInBot_3_7[12] , 
        \wRegInBot_5_0[18] , \wRegInTop_5_5[12] , \wRegOut_6_14[15] , 
        \wRegOut_6_40[0] , \wRegOut_7_61[6] , \wRegOut_6_37[24] , 
        \wRegOut_6_61[25] , \wRegOut_6_42[14] , \wRegInTop_6_52[8] , 
        \wRegOut_7_39[14] , \wRegOut_5_19[24] , \wRegOut_6_43[3] , 
        \wRegInTop_7_101[20] , \ScanLink243[9] , \wRegOut_7_62[5] , 
        \wRegOut_7_81[20] , \wRegInTop_7_122[11] , \wRegInBot_5_6[3] , 
        \ScanLink77[10] , \wRegOut_7_94[14] , \wRegInTop_7_114[14] , 
        \wRegInTop_5_7[5] , \wRegOut_7_121[29] , \ScanLink54[21] , 
        \ScanLink209[24] , \wRegInBot_3_6[7] , \wRegInTop_3_7[1] , 
        \ScanLink21[11] , \wRegOut_5_12[1] , \wRegOut_7_102[18] , 
        \wRegOut_7_121[30] , \ScanLink34[25] , \ScanLink41[15] , 
        \wRegInBot_6_32[18] , \wRegEnTop_7_23[0] , \wRegInBot_6_11[30] , 
        \ScanLink62[24] , \wRegInBot_6_47[28] , \wRegOut_4_1[9] , 
        \wRegInBot_6_11[29] , \ScanLink17[14] , \wRegOut_5_2[10] , 
        \wRegInBot_5_17[14] , \wRegInTop_5_21[16] , \wRegInBot_6_47[31] , 
        \wRegOut_7_127[6] , \wRegInBot_6_60[8] , \wRegInTop_5_17[13] , 
        \ScanLink222[0] , \wRegInBot_5_21[11] , \ScanLink92[29] , 
        \ScanLink61[8] , \ScanLink92[30] , \wRegInTop_6_30[2] , 
        \wRegInTop_7_11[4] , \wRegOut_7_5[14] , \ScanLink142[5] , 
        \wRegInTop_7_110[9] , \wRegOut_7_0[5] , \wRegOut_7_11[29] , 
        \wRegOut_7_47[31] , \wRegOut_7_64[19] , \wRegOut_7_47[28] , 
        \wRegInTop_2_2[26] , \wRegInTop_2_2[15] , \wRegInBot_3_0[9] , 
        \wRegOut_3_5[30] , \wRegOut_3_5[29] , \wRegEnBot_3_6[0] , 
        \wRegInBot_4_4[17] , \wRegOut_5_12[31] , \wRegOut_5_12[28] , 
        \wRegInTop_6_6[9] , \wRegOut_6_49[18] , \wRegOut_7_11[30] , 
        \wRegOut_7_32[18] , \ScanLink190[3] , \wRegOut_5_31[19] , 
        \wRegInBot_6_3[13] , \wRegEnTop_6_0[0] , \wRegOut_7_3[6] , 
        \wRegInTop_6_6[19] , \ScanLink193[0] , \wRegInTop_7_14[12] , 
        \wRegInTop_5_2[8] , \ScanLink69[31] , \wRegOut_6_21[9] , 
        \wRegInTop_7_61[22] , \ScanLink202[31] , \ScanLink221[19] , 
        \wRegInTop_6_39[13] , \wRegInBot_6_59[10] , \wRegInTop_7_37[23] , 
        \ScanLink221[3] , \ScanLink254[29] , \ScanLink202[28] , 
        \wRegOut_7_124[5] , \wRegInTop_7_42[13] , \wRegOut_7_109[14] , 
        \wRegInTop_6_59[17] , \ScanLink254[30] , \ScanLink69[28] , 
        \wRegInTop_6_33[1] , \wRegInBot_6_39[14] , \wRegInTop_7_12[7] , 
        \ScanLink141[6] , \wRegInTop_7_22[17] , \wRegInTop_7_57[27] , 
        \wRegInBot_6_19[3] , \wRegInTop_7_74[16] , \wRegInTop_6_49[9] , 
        \wRegOut_7_5[27] , \ScanLink18[3] , \wRegOut_4_4[4] , 
        \wRegInTop_5_17[20] , \ScanLink149[30] , \wRegInBot_5_21[22] , 
        \wRegInTop_7_9[30] , \wRegInTop_7_9[29] , \ScanLink149[29] , 
        \wRegOut_7_67[8] , \ScanLink246[4] , \wRegInBot_4_4[24] , 
        \wRegOut_5_2[23] , \wRegInTop_5_21[25] , \wRegInTop_6_54[6] , 
        \ScanLink126[1] , \wRegInTop_7_75[0] , \wRegInBot_5_17[27] , 
        \wRegInBot_6_39[27] , \wRegInTop_6_59[24] , \wRegInTop_7_57[14] , 
        \wRegInTop_7_22[24] , \wRegInTop_7_61[11] , \ScanLink191[19] , 
        \wRegInTop_7_74[25] , \ScanLink245[7] , \wRegInTop_6_39[20] , 
        \wRegInBot_6_59[23] , \wRegInTop_7_14[21] , \wRegInTop_7_42[20] , 
        \wRegOut_7_109[27] , \wRegInTop_6_57[5] , \wRegOut_6_58[2] , 
        \ScanLink125[2] , \wRegInTop_7_37[10] , \wRegInTop_7_76[3] , 
        \wRegOut_7_79[4] , \wRegOut_3_1[18] , \wRegOut_4_7[7] , 
        \wRegInBot_6_3[20] , \wRegInBot_6_23[9] , \wRegInTop_6_28[25] , 
        \wRegInTop_7_26[15] , \ScanLink195[31] , \ScanLink101[4] , 
        \wRegInBot_6_48[26] , \wRegInTop_7_52[5] , \wRegInTop_7_53[25] , 
        \wRegOut_7_118[22] , \ScanLink195[28] , \wRegInTop_7_70[14] , 
        \wRegInTop_7_10[10] , \wRegInBot_4_0[15] , \ScanLink22[9] , 
        \wRegOut_4_9[11] , \wRegInTop_5_22[1] , \wRegInBot_6_28[22] , 
        \wRegInTop_7_33[21] , \wRegInTop_7_65[20] , \wRegInTop_6_48[21] , 
        \wRegInTop_7_46[11] , \wRegInTop_7_80[3] , \wRegInBot_6_7[11] , 
        \wRegInTop_5_13[11] , \wRegInTop_5_21[2] , \wRegOut_5_30[9] , 
        \wRegOut_7_1[16] , \wRegInTop_7_83[0] , \ScanLink138[31] , 
        \wRegOut_7_91[8] , \wRegInBot_5_25[13] , \ScanLink138[28] , 
        \ScanLink7[1] , \wRegOut_4_9[22] , \wRegOut_5_6[12] , 
        \wRegInBot_5_13[16] , \wRegInTop_5_25[14] , \wRegInTop_5_30[20] , 
        \wRegInTop_7_51[6] , \wRegInBot_5_30[27] , \ScanLink102[7] , 
        \wRegOut_6_62[8] , \wRegOut_5_16[19] , \wRegEnBot_6_14[0] , 
        \wRegInTop_6_2[31] , \wRegInBot_6_7[22] , \wRegInTop_6_2[28] , 
        \ScanLink89[4] , \wRegInBot_4_0[26] , \wRegOut_6_18[0] , 
        \wRegOut_7_39[6] , \wRegInTop_7_65[13] , \ScanLink250[18] , 
        \ScanLink18[30] , \wRegInTop_6_17[7] , \wRegInBot_6_28[11] , 
        \wRegInTop_7_8[0] , \wRegInTop_7_10[23] , \wRegInTop_7_46[22] , 
        \ScanLink225[28] , \wRegInTop_6_28[16] , \wRegInTop_6_48[12] , 
        \wRegInTop_7_33[12] , \wRegInTop_7_36[1] , \ScanLink165[0] , 
        \ScanLink206[19] , \ScanLink225[31] , \ScanLink18[29] , 
        \wRegInBot_6_48[15] , \wRegInTop_7_26[26] , \wRegInTop_7_53[16] , 
        \wRegOut_7_100[3] , \wRegOut_7_118[11] , \wRegOut_5_6[21] , 
        \wRegInTop_5_25[27] , \wRegOut_7_24[9] , \wRegInTop_7_70[27] , 
        \ScanLink205[5] , \wRegInBot_5_30[14] , \wRegInTop_6_14[4] , 
        \ScanLink166[3] , \wRegInTop_7_35[2] , \wRegInTop_5_13[22] , 
        \wRegInBot_5_13[25] , \ScanLink96[18] , \wRegInBot_5_25[20] , 
        \wRegInTop_5_30[13] , \ScanLink206[6] , \wRegOut_7_103[0] , 
        \ScanLink58[1] , \ScanLink97[8] , \wRegOut_7_1[25] , \ScanLink4[2] , 
        \wRegInBot_6_59[1] , \wRegOut_7_15[18] , \wRegOut_7_36[30] , 
        \wRegOut_0_0[7] , \wRegInBot_0_0[21] , \ScanLink1[22] , 
        \ScanLink1[18] , \wRegInBot_3_3[23] , \wRegOut_6_38[19] , 
        \wRegOut_7_36[29] , \wRegOut_7_60[28] , \wRegOut_7_43[19] , 
        \wRegOut_7_60[31] , \wRegInBot_3_3[10] , \ScanLink13[25] , 
        \wRegInTop_3_6[30] , \wRegInTop_3_6[29] , \wRegOut_4_13[25] , 
        \wRegInTop_7_105[11] , \ScanLink39[8] , \wRegOut_7_85[11] , 
        \wRegInTop_7_126[20] , \wRegInTop_6_9[24] , \wRegInBot_6_25[7] , 
        \wRegOut_7_90[25] , \wRegInTop_7_110[25] , \wRegOut_7_46[3] , 
        \ScanLink24[7] , \ScanLink25[20] , \ScanLink73[21] , 
        \wRegOut_7_106[30] , \wRegOut_7_125[18] , \ScanLink30[14] , 
        \ScanLink50[10] , \wRegOut_7_106[29] , \wRegInBot_6_43[19] , 
        \wRegInTop_7_49[4] , \wRegInBot_6_60[31] , \ScanLink45[24] , 
        \wRegEnTop_6_26[0] , \ScanLink218[21] , \wRegInBot_6_36[29] , 
        \wRegInBot_6_38[8] , \ScanLink13[16] , \ScanLink27[4] , 
        \wRegOut_4_14[2] , \wRegInBot_5_18[30] , \ScanLink66[15] , 
        \wRegInBot_6_15[18] , \wRegInBot_6_60[28] , \wRegOut_7_94[5] , 
        \wRegInBot_6_36[30] , \ScanLink153[13] , \wRegInBot_5_18[29] , 
        \ScanLink88[20] , \ScanLink119[6] , \ScanLink126[23] , 
        \ScanLink170[22] , \ScanLink105[12] , \ScanLink110[26] , 
        \wRegInTop_7_6[27] , \ScanLink165[16] , \ScanLink133[17] , 
        \ScanLink146[27] , \wRegOut_7_97[6] , \ScanLink30[27] , 
        \wRegInTop_5_1[23] , \wRegInBot_5_4[30] , \wRegOut_6_26[21] , 
        \wRegOut_6_53[11] , \wRegOut_7_28[11] , \wRegInTop_7_57[8] , 
        \wRegInBot_5_4[29] , \ScanLink104[9] , \wRegInTop_7_98[1] , 
        \wRegOut_6_10[24] , \wRegInBot_6_26[4] , \wRegOut_7_45[0] , 
        \ScanLink45[17] , \wRegOut_6_33[15] , \wRegOut_6_46[25] , 
        \wRegOut_7_48[15] , \wRegInTop_6_56[19] , \ScanLink218[12] , 
        \wRegInTop_6_23[29] , \ScanLink66[26] , \wRegInTop_7_58[29] , 
        \wRegInTop_6_23[30] , \wRegInTop_7_58[30] , \ScanLink25[13] , 
        \wRegInBot_5_10[1] , \ScanLink50[23] , \ScanLink73[12] , 
        \wRegOut_6_5[19] , \wRegOut_4_13[16] , \ScanLink40[3] , 
        \wRegInTop_6_9[17] , \wRegInTop_6_11[9] , \wRegOut_7_90[16] , 
        \wRegInTop_7_110[16] , \wRegInBot_6_41[3] , \wRegInTop_7_105[22] , 
        \wRegInTop_5_1[10] , \wRegOut_6_8[2] , \wRegOut_7_22[7] , 
        \wRegOut_7_85[22] , \wRegOut_6_10[17] , \ScanLink92[5] , 
        \wRegInTop_7_126[13] , \wRegOut_6_33[26] , \wRegOut_7_48[26] , 
        \wRegOut_6_46[16] , \wRegOut_6_26[12] , \ScanLink91[6] , 
        \wRegOut_6_53[22] , \wRegOut_7_28[22] , \wRegInBot_6_42[0] , 
        \ScanLink1[11] , \ScanLink1[6] , \wRegOut_1_0[8] , \wRegInBot_2_3[27] , 
        \wRegInTop_3_2[5] , \ScanLink43[0] , \wRegInBot_5_13[2] , 
        \ScanLink110[15] , \wRegOut_7_21[4] , \ScanLink200[8] , 
        \ScanLink133[24] , \wRegInTop_7_6[14] , \ScanLink165[25] , 
        \wRegInTop_7_80[19] , \ScanLink146[14] , \ScanLink126[10] , 
        \wRegOut_7_118[1] , \ScanLink88[13] , \ScanLink105[21] , 
        \ScanLink153[20] , \wRegOut_6_29[26] , \wRegOut_7_27[16] , 
        \ScanLink170[11] , \wRegInTop_6_49[0] , \wRegOut_7_52[26] , 
        \wRegInTop_7_68[6] , \wRegInBot_3_3[3] , \wRegOut_7_71[17] , 
        \wRegInTop_5_2[1] , \wRegInBot_5_3[7] , \wRegOut_7_11[13] , 
        \wRegOut_7_64[23] , \wRegOut_5_17[5] , \wRegOut_6_49[22] , 
        \wRegOut_7_32[22] , \wRegOut_7_47[12] , \ScanLink126[8] , 
        \ScanLink129[24] , \wRegInTop_7_75[9] , \wRegInBot_2_3[14] , 
        \wRegInBot_3_0[0] , \wRegInTop_3_1[6] , \wRegOut_3_5[20] , 
        \wRegInTop_5_17[30] , \wRegInTop_5_17[29] , \wRegInTop_5_18[2] , 
        \ScanLink87[27] , \ScanLink92[13] , \wRegInTop_7_9[20] , 
        \wRegOut_6_46[7] , \ScanLink149[20] , \wRegOut_7_67[1] , 
        \wRegInTop_6_39[30] , \wRegInTop_7_42[30] , \wRegInTop_7_61[18] , 
        \ScanLink254[13] , \wRegInTop_4_1[27] , \wRegInTop_6_39[29] , 
        \wRegInTop_7_14[28] , \wRegInTop_7_42[29] , \ScanLink184[24] , 
        \ScanLink221[23] , \wRegInTop_7_14[31] , \wRegInTop_7_37[19] , 
        \ScanLink202[12] , \ScanLink69[12] , \wRegOut_6_45[4] , 
        \ScanLink217[26] , \ScanLink241[27] , \ScanLink191[10] , 
        \wRegOut_7_64[2] , \ScanLink234[17] , \wRegInBot_6_3[30] , 
        \wRegInBot_5_0[4] , \wRegOut_5_12[12] , \wRegOut_5_14[6] , 
        \wRegOut_5_31[23] , \wRegInBot_6_3[29] , \ScanLink138[4] , 
        \wRegOut_5_24[17] , \wRegInTop_5_1[2] , \wRegInTop_6_6[23] , 
        \wRegOut_5_2[19] , \wRegInBot_5_21[18] , \ScanLink92[20] , 
        \wRegInTop_7_9[13] , \wRegOut_6_22[3] , \ScanLink87[14] , 
        \wRegInBot_6_60[1] , \ScanLink129[17] , \ScanLink149[13] , 
        \ScanLink222[9] , \wRegOut_7_11[20] , \wRegOut_7_64[10] , 
        \wRegOut_2_1[4] , \ScanLink5[13] , \wRegOut_2_2[7] , \wRegOut_3_5[13] , 
        \wRegInTop_4_1[14] , \wRegInBot_4_10[5] , \wRegInTop_6_6[0] , 
        \wRegInBot_6_7[6] , \wRegOut_7_32[11] , \wRegOut_7_47[21] , 
        \wRegOut_6_29[15] , \wRegOut_6_49[11] , \wRegInBot_4_13[6] , 
        \wRegOut_5_12[21] , \wRegOut_5_24[24] , \ScanLink61[1] , 
        \wRegInBot_5_31[3] , \wRegOut_7_52[15] , \wRegInTop_7_110[0] , 
        \wRegEnTop_7_42[0] , \wRegOut_7_27[25] , \wRegOut_7_71[24] , 
        \wRegInBot_6_4[5] , \wRegInTop_6_5[3] , \wRegInTop_6_6[10] , 
        \ScanLink193[9] , \wRegInTop_7_113[3] , \ScanLink62[2] , 
        \wRegOut_5_31[10] , \wRegInTop_6_33[8] , \ScanLink217[15] , 
        \ScanLink69[21] , \ScanLink191[23] , \ScanLink234[24] , 
        \ScanLink241[14] , \wRegOut_4_2[3] , \wRegInTop_4_12[26] , 
        \wRegOut_6_21[0] , \wRegInBot_6_63[2] , \ScanLink184[17] , 
        \ScanLink221[10] , \ScanLink254[20] , \wRegInBot_6_59[19] , 
        \ScanLink202[21] , \wRegInTop_7_84[12] , \wRegInBot_5_5[9] , 
        \wRegInBot_4_12[21] , \wRegOut_5_9[15] , \wRegInTop_7_91[26] , 
        \wRegInBot_5_0[11] , \wRegOut_6_22[19] , \wRegInTop_6_52[1] , 
        \ScanLink120[6] , \wRegInTop_7_73[7] , \wRegOut_6_57[29] , 
        \wRegOut_7_59[19] , \wRegInTop_3_2[11] , \wRegOut_6_40[9] , 
        \wRegOut_6_57[30] , \ScanLink240[3] , \wRegInTop_3_7[8] , 
        \wRegOut_4_6[16] , \wRegInTop_6_51[2] , \ScanLink123[5] , 
        \wRegInTop_7_70[4] , \wRegInBot_6_8[16] , \wRegOut_7_81[29] , 
        \wRegInTop_7_101[29] , \ScanLink243[0] , \wRegInBot_6_11[20] , 
        \wRegInTop_6_27[22] , \wRegInBot_6_32[11] , \wRegInTop_6_52[12] , 
        \wRegOut_7_81[30] , \wRegInTop_7_101[30] , \wRegInTop_7_122[18] , 
        \wRegInTop_7_29[12] , \wRegInBot_6_47[21] , \wRegOut_7_117[25] , 
        \wRegOut_4_1[0] , \wRegEnBot_5_3[0] , \ScanLink54[31] , 
        \ScanLink77[19] , \ScanLink5[20] , \ScanLink21[18] , \ScanLink54[28] , 
        \wRegInTop_6_11[27] , \wRegOut_7_121[20] , \wRegInBot_6_27[25] , 
        \wRegInTop_6_47[26] , \wRegOut_7_102[11] , \wRegOut_5_12[8] , 
        \wRegOut_6_1[12] , \wRegInBot_6_52[15] , \wRegInTop_7_49[16] , 
        \wRegInTop_6_32[16] , \wRegInTop_6_36[5] , \wRegInTop_7_17[3] , 
        \ScanLink144[2] , \wRegInTop_3_2[22] , \wRegInBot_3_7[31] , 
        \wRegInBot_3_7[28] , \wRegInTop_4_12[15] , \wRegInBot_4_12[12] , 
        \wRegInBot_5_0[22] , \wRegInTop_5_5[31] , \wRegInTop_5_5[28] , 
        \ScanLink224[7] , \wRegOut_7_121[1] , \wRegOut_5_9[26] , 
        \wRegInBot_6_1[8] , \ScanLink122[28] , \ScanLink157[18] , 
        \ScanLink174[30] , \ScanLink196[4] , \ScanLink101[19] , 
        \ScanLink122[31] , \ScanLink174[29] , \wRegInTop_7_91[15] , 
        \wRegOut_6_39[2] , \wRegOut_7_18[4] , \ScanLink239[8] , 
        \wRegInBot_4_15[8] , \wRegOut_6_1[21] , \wRegInTop_6_11[14] , 
        \wRegOut_7_6[2] , \wRegInTop_7_84[21] , \wRegOut_7_121[13] , 
        \wRegInBot_6_52[26] , \wRegInTop_6_27[11] , \wRegInBot_6_27[16] , 
        \wRegInTop_6_32[25] , \wRegInTop_7_49[25] , \wRegOut_7_102[22] , 
        \wRegInTop_6_28[9] , \wRegInTop_6_47[15] , \ScanLink195[7] , 
        \wRegInBot_6_11[13] , \wRegInBot_6_32[22] , \wRegInBot_6_47[12] , 
        \wRegOut_7_117[16] , \wRegInTop_6_52[21] , \wRegOut_7_5[1] , 
        \wRegInTop_7_29[21] , \wRegOut_4_6[25] , \wRegInBot_5_29[1] , 
        \wRegInBot_6_8[25] , \wRegInTop_6_35[6] , \wRegInTop_7_14[0] , 
        \ScanLink147[1] , \ScanLink188[8] , \wRegInTop_7_108[2] , 
        \wRegOut_7_122[2] , \ScanLink79[3] , \wRegInTop_6_60[15] , 
        \ScanLink227[4] , \wRegInTop_1_1[17] , \wRegInBot_5_10[8] , 
        \wRegInTop_6_15[25] , \wRegOut_7_125[22] , \wRegInBot_6_23[27] , 
        \wRegInTop_7_38[24] , \wRegOut_6_5[10] , \wRegInTop_6_43[24] , 
        \wRegOut_7_106[13] , \wRegInBot_6_15[22] , \wRegInTop_6_23[20] , 
        \wRegInTop_6_36[14] , \wRegInBot_6_56[17] , \wRegInBot_6_36[13] , 
        \wRegInTop_6_56[10] , \wRegInBot_6_43[23] , \wRegInTop_7_58[20] , 
        \wRegOut_7_113[27] , \wRegInBot_3_3[19] , \wRegOut_4_2[14] , 
        \wRegInBot_6_60[12] , \ScanLink203[2] , \wRegInTop_3_6[13] , 
        \wRegOut_7_106[4] , \wRegInBot_5_4[13] , \wRegInTop_6_11[0] , 
        \wRegInTop_7_30[6] , \ScanLink163[7] , \wRegOut_7_105[7] , 
        \wRegInBot_6_42[9] , \ScanLink2[5] , \wRegInTop_5_1[19] , 
        \wRegInTop_6_12[3] , \ScanLink160[4] , \ScanLink200[1] , 
        \wRegEnTop_7_125[0] , \ScanLink43[9] , \ScanLink105[31] , 
        \wRegInTop_7_33[5] , \wRegOut_7_118[8] , \ScanLink126[19] , 
        \ScanLink153[29] , \wRegInTop_7_95[24] , \wRegInTop_1_1[24] , 
        \wRegInTop_3_6[20] , \ScanLink39[1] , \wRegInTop_5_18[14] , 
        \wRegInBot_5_18[13] , \ScanLink105[28] , \ScanLink153[30] , 
        \ScanLink170[18] , \wRegInTop_7_80[10] , \wRegOut_4_2[27] , 
        \wRegOut_7_89[3] , \wRegInTop_7_105[18] , \wRegInTop_7_126[30] , 
        \wRegInTop_6_23[13] , \ScanLink107[3] , \wRegOut_7_85[18] , 
        \wRegInTop_7_126[29] , \wRegInTop_7_54[2] , \wRegInBot_6_36[20] , 
        \wRegInBot_6_43[10] , \wRegInTop_7_58[13] , \wRegOut_7_113[14] , 
        \wRegInTop_6_56[23] , \ScanLink218[28] , \wRegInBot_6_38[1] , 
        \wRegInBot_6_60[21] , \ScanLink218[31] , \wRegInBot_4_8[3] , 
        \wRegInTop_4_9[5] , \ScanLink25[30] , \wRegInBot_6_15[11] , 
        \wRegOut_7_125[11] , \ScanLink25[29] , \wRegInTop_5_24[6] , 
        \ScanLink73[28] , \wRegInTop_6_15[16] , \wRegInTop_6_60[26] , 
        \wRegOut_6_5[23] , \wRegInBot_6_56[24] , \wRegInTop_5_18[27] , 
        \ScanLink50[19] , \wRegInTop_6_36[27] , \wRegOut_7_106[20] , 
        \wRegInTop_7_86[4] , \ScanLink73[31] , \wRegInBot_6_23[14] , 
        \wRegInTop_7_38[17] , \wRegInTop_6_43[17] , \wRegInBot_5_18[20] , 
        \wRegInTop_5_27[5] , \ScanLink88[30] , \wRegOut_7_58[6] , 
        \wRegInTop_7_80[23] , \ScanLink88[29] , \wRegInTop_7_85[7] , 
        \wRegInTop_7_95[17] , \wRegOut_7_45[9] , \wRegOut_5_28[2] , 
        \wRegOut_6_26[28] , \wRegOut_6_53[18] , \wRegOut_7_28[18] , 
        \wRegInTop_7_57[1] , \ScanLink104[0] , \wRegInTop_7_98[8] , 
        \ScanLink7[8] , \wRegInBot_5_4[20] , \ScanLink46[4] , 
        \wRegInBot_5_16[6] , \wRegOut_6_26[31] , \wRegOut_5_20[15] , 
        \wRegOut_3_1[22] , \ScanLink18[20] , \wRegInTop_4_5[25] , 
        \wRegOut_5_16[10] , \wRegInTop_6_2[21] , \wRegOut_6_18[9] , 
        \ScanLink218[3] , \ScanLink178[6] , \ScanLink94[2] , \ScanLink213[24] , 
        \wRegOut_7_118[18] , \wRegInBot_6_47[4] , \ScanLink245[25] , 
        \ScanLink78[24] , \wRegOut_7_24[0] , \ScanLink195[12] , 
        \ScanLink230[15] , \ScanLink250[11] , \wRegOut_5_6[31] , 
        \wRegInBot_5_25[30] , \wRegInBot_6_28[18] , \wRegInTop_7_8[9] , 
        \ScanLink180[26] , \ScanLink225[21] , \wRegInTop_7_36[8] , 
        \ScanLink96[11] , \wRegInBot_6_44[7] , \ScanLink165[9] , 
        \ScanLink206[10] , \wRegInBot_5_25[29] , \ScanLink58[8] , 
        \wRegOut_7_27[3] , \wRegOut_7_103[9] , \ScanLink97[1] , 
        \ScanLink138[12] , \wRegOut_5_6[28] , \ScanLink158[16] , 
        \ScanLink45[7] , \wRegInBot_5_15[5] , \ScanLink83[25] , 
        \wRegInBot_6_59[8] , \wRegOut_7_15[11] , \wRegOut_7_60[21] , 
        \wRegEnTop_6_47[0] , \wRegOut_7_36[20] , \wRegOut_7_43[10] , 
        \wRegOut_6_38[10] , \wRegOut_6_58[14] , \wRegInBot_0_0[12] , 
        \wRegOut_3_1[11] , \ScanLink78[17] , \wRegOut_7_23[14] , 
        \wRegInTop_7_28[4] , \wRegOut_7_56[24] , \wRegOut_7_75[15] , 
        \wRegInTop_7_10[19] , \ScanLink18[13] , \wRegInTop_4_5[16] , 
        \wRegInBot_6_23[0] , \wRegInTop_7_33[31] , \wRegInTop_6_48[31] , 
        \ScanLink180[15] , \ScanLink225[12] , \wRegInTop_6_48[28] , 
        \wRegOut_6_61[2] , \wRegOut_7_40[4] , \wRegInTop_7_65[29] , 
        \ScanLink250[22] , \wRegInTop_7_33[28] , \ScanLink206[23] , 
        \wRegInTop_7_46[18] , \wRegInTop_7_65[30] , \ScanLink213[17] , 
        \ScanLink195[21] , \ScanLink230[26] , \ScanLink245[16] , 
        \ScanLink22[0] , \wRegOut_4_9[18] , \wRegOut_5_16[23] , 
        \wRegOut_7_92[2] , \wRegInBot_6_7[18] , \wRegOut_4_11[6] , 
        \wRegOut_4_12[5] , \wRegOut_5_20[26] , \wRegOut_5_30[0] , 
        \wRegInTop_5_22[8] , \wRegInTop_6_2[12] , \wRegOut_7_56[17] , 
        \ScanLink0[31] , \ScanLink0[28] , \ScanLink21[3] , \wRegOut_6_58[27] , 
        \wRegInTop_5_0[20] , \wRegOut_5_9[7] , \ScanLink83[16] , 
        \wRegInBot_6_20[3] , \wRegOut_6_38[23] , \wRegOut_7_15[22] , 
        \wRegOut_7_23[27] , \wRegOut_7_60[12] , \wRegOut_7_75[26] , 
        \wRegOut_7_91[1] , \wRegOut_7_43[23] , \ScanLink158[25] , 
        \wRegOut_7_36[13] , \wRegInTop_7_83[9] , \wRegOut_7_43[7] , 
        \wRegOut_6_62[1] , \wRegInTop_5_13[18] , \wRegInTop_5_30[30] , 
        \wRegInTop_5_30[29] , \ScanLink96[22] , \ScanLink138[21] , 
        \wRegOut_6_47[26] , \wRegOut_6_11[27] , \wRegOut_6_32[16] , 
        \wRegOut_7_49[16] , \wRegInBot_6_36[7] , \wRegOut_7_55[3] , 
        \wRegInTop_1_0[5] , \wRegInBot_1_1[3] , \wRegOut_3_2[8] , 
        \wRegInTop_4_4[0] , \ScanLink37[7] , \wRegOut_5_25[7] , 
        \wRegOut_6_27[22] , \wRegOut_6_52[12] , \wRegOut_7_29[12] , 
        \ScanLink132[14] , \ScanLink147[24] , \wRegInTop_7_88[2] , 
        \wRegEnTop_6_35[0] , \wRegInTop_7_81[30] , \ScanLink164[15] , 
        \wRegInBot_4_5[6] , \ScanLink111[25] , \wRegInTop_7_7[24] , 
        \wRegInTop_7_81[29] , \wRegOut_7_87[5] , \wRegInBot_3_2[20] , 
        \ScanLink12[26] , \ScanLink89[23] , \ScanLink104[11] , 
        \ScanLink171[21] , \ScanLink109[5] , \ScanLink152[10] , 
        \ScanLink127[20] , \wRegInBot_4_6[5] , \wRegInTop_4_7[3] , 
        \wRegInTop_6_57[30] , \wRegOut_7_84[6] , \ScanLink24[23] , 
        \ScanLink31[17] , \ScanLink67[16] , \wRegInTop_6_22[19] , 
        \ScanLink34[4] , \wRegInTop_6_57[29] , \wRegInTop_7_59[19] , 
        \ScanLink44[27] , \ScanLink219[22] , \wRegOut_5_26[4] , 
        \ScanLink51[13] , \wRegOut_6_4[29] , \wRegOut_6_4[30] , 
        \wRegInTop_7_59[7] , \wRegInTop_6_8[27] , \ScanLink72[22] , 
        \wRegInBot_6_35[4] , \wRegOut_7_91[26] , \wRegInTop_7_111[26] , 
        \ScanLink117[9] , \wRegOut_7_56[0] , \wRegOut_7_99[9] , 
        \wRegInTop_7_127[23] , \wRegInTop_7_44[8] , \wRegOut_4_12[26] , 
        \wRegInTop_7_104[12] , \wRegInBot_5_19[19] , \wRegInTop_5_29[3] , 
        \wRegOut_7_84[12] , \ScanLink89[10] , \ScanLink104[22] , 
        \ScanLink171[12] , \ScanLink53[3] , \ScanLink127[13] , 
        \wRegOut_7_108[2] , \wRegInTop_7_122[2] , \wRegInTop_2_1[9] , 
        \wRegInTop_2_3[16] , \wRegInBot_3_2[13] , \wRegOut_4_12[15] , 
        \wRegInTop_5_0[13] , \wRegInBot_5_5[19] , \ScanLink111[16] , 
        \wRegInTop_7_0[1] , \ScanLink152[23] , \ScanLink132[27] , 
        \ScanLink147[17] , \wRegInBot_6_52[3] , \wRegInTop_7_7[17] , 
        \ScanLink164[26] , \wRegOut_6_10[1] , \ScanLink81[5] , 
        \wRegOut_6_27[11] , \wRegOut_7_31[7] , \wRegOut_6_52[21] , 
        \wRegOut_7_29[21] , \wRegOut_6_32[25] , \wRegOut_7_49[25] , 
        \wRegOut_6_11[14] , \wRegOut_6_47[15] , \wRegOut_6_13[2] , 
        \ScanLink82[6] , \wRegInTop_7_127[10] , \wRegInBot_6_51[0] , 
        \wRegInTop_7_104[21] , \wRegOut_7_32[4] , \ScanLink12[15] , 
        \wRegInTop_3_7[19] , \wRegInTop_6_8[14] , \wRegOut_7_84[21] , 
        \ScanLink213[8] , \wRegOut_7_91[15] , \wRegInTop_7_111[15] , 
        \ScanLink24[10] , \ScanLink51[20] , \wRegInTop_7_121[1] , 
        \wRegOut_7_124[31] , \ScanLink50[0] , \wRegOut_7_107[19] , 
        \ScanLink67[25] , \ScanLink72[11] , \wRegOut_7_124[28] , 
        \wRegInBot_6_14[28] , \wRegInBot_6_42[30] , \wRegInBot_6_61[18] , 
        \wRegEnBot_4_13[0] , \ScanLink31[24] , \ScanLink44[14] , 
        \wRegInBot_6_14[31] , \wRegInBot_6_37[19] , \wRegInTop_7_3[2] , 
        \ScanLink219[11] , \wRegOut_5_7[11] , \wRegInBot_5_12[15] , 
        \wRegInBot_6_30[9] , \wRegInBot_6_42[29] , \wRegInTop_5_24[17] , 
        \wRegInBot_5_31[24] , \wRegInBot_5_24[10] , \wRegOut_3_4[6] , 
        \wRegInTop_5_12[12] , \wRegInTop_5_31[23] , \ScanLink97[31] , 
        \wRegInTop_6_60[3] , \wRegInTop_7_41[5] , \ScanLink97[28] , 
        \ScanLink112[4] , \wRegOut_3_7[5] , \wRegInBot_4_3[8] , 
        \wRegInTop_4_10[7] , \ScanLink31[9] , \wRegOut_5_23[9] , 
        \wRegOut_7_0[15] , \wRegOut_5_4[2] , \wRegOut_6_39[29] , 
        \wRegOut_7_42[29] , \wRegOut_7_14[31] , \wRegOut_7_37[19] , 
        \wRegOut_7_42[30] , \wRegInTop_7_93[3] , \wRegOut_6_39[30] , 
        \wRegOut_7_61[18] , \wRegOut_7_14[28] , \wRegOut_5_17[30] , 
        \wRegInTop_5_31[1] , \wRegInBot_6_6[12] , \wRegOut_5_17[29] , 
        \wRegOut_4_8[12] , \wRegOut_5_7[1] , \wRegOut_7_82[8] , 
        \wRegInBot_4_1[16] , \wRegInTop_4_13[4] , \wRegInTop_6_3[18] , 
        \wRegInBot_6_29[21] , \wRegInTop_7_32[22] , \wRegInTop_7_90[0] , 
        \wRegInTop_6_49[22] , \wRegInTop_7_47[12] , \ScanLink207[29] , 
        \ScanLink251[31] , \ScanLink19[19] , \wRegInTop_7_11[13] , 
        \wRegInTop_7_64[23] , \ScanLink207[30] , \ScanLink224[18] , 
        \ScanLink251[28] , \wRegOut_6_0[3] , \wRegInTop_6_29[26] , 
        \wRegInTop_7_27[16] , \wRegInTop_7_71[17] , \ScanLink111[7] , 
        \wRegInBot_6_49[25] , \wRegInTop_7_42[6] , \wRegInTop_7_52[26] , 
        \wRegOut_7_119[21] , \wRegInTop_6_63[0] , \wRegInBot_6_49[2] , 
        \wRegOut_7_0[26] , \wRegInBot_1_1[26] , \wRegInTop_2_3[25] , 
        \ScanLink48[2] , \wRegInBot_5_18[0] , \wRegInTop_6_19[8] , 
        \wRegInBot_5_24[23] , \wRegInTop_5_31[10] , \wRegOut_7_113[3] , 
        \ScanLink139[18] , \wRegOut_3_0[31] , \wRegOut_5_7[22] , 
        \wRegInTop_5_12[21] , \wRegOut_7_37[9] , \ScanLink216[5] , 
        \wRegInBot_5_12[26] , \wRegInTop_5_24[24] , \wRegInBot_5_31[17] , 
        \ScanLink176[0] , \ScanLink84[8] , \wRegInTop_6_29[15] , 
        \wRegInTop_7_25[1] , \ScanLink194[18] , \wRegInTop_7_71[24] , 
        \ScanLink215[6] , \wRegInBot_6_49[16] , \wRegInTop_7_52[15] , 
        \wRegOut_7_110[0] , \wRegOut_7_119[12] , \wRegInBot_6_29[12] , 
        \wRegInTop_7_27[25] , \wRegInTop_7_47[21] , \wRegEnTop_7_68[0] , 
        \wRegOut_3_0[28] , \wRegInBot_4_1[25] , \wRegInTop_6_49[11] , 
        \wRegInTop_7_26[2] , \wRegInTop_7_32[11] , \ScanLink175[3] , 
        \wRegInTop_7_11[20] , \wRegInTop_7_64[10] , \wRegInTop_3_3[31] , 
        \wRegOut_3_4[19] , \wRegOut_4_8[21] , \wRegOut_6_3[0] , 
        \wRegOut_7_29[5] , \ScanLink208[9] , \wRegInBot_6_6[21] , 
        \ScanLink99[7] , \wRegInTop_6_8[6] , \wRegInBot_6_9[0] , 
        \wRegInBot_6_38[17] , \wRegInTop_6_58[14] , \ScanLink190[29] , 
        \wRegInTop_7_75[15] , \ScanLink190[30] , \wRegInTop_7_23[14] , 
        \wRegInTop_6_23[2] , \ScanLink151[5] , \wRegInTop_7_56[24] , 
        \wRegInTop_6_38[10] , \wRegInBot_6_58[13] , \wRegInTop_7_36[20] , 
        \wRegInTop_7_43[10] , \wRegOut_7_108[17] , \wRegInBot_3_6[22] , 
        \wRegInBot_4_5[27] , \wRegInBot_4_5[14] , \wRegOut_5_3[13] , 
        \wRegInTop_5_16[10] , \wRegInBot_5_20[12] , \wRegInBot_5_21[9] , 
        \wRegInBot_6_2[10] , \wRegInTop_7_15[11] , \ScanLink183[3] , 
        \wRegInTop_7_60[21] , \ScanLink231[0] , \ScanLink72[8] , 
        \wRegInTop_7_103[9] , \ScanLink180[0] , \wRegOut_7_4[17] , 
        \wRegInTop_6_20[1] , \ScanLink148[19] , \ScanLink152[6] , 
        \wRegInBot_5_16[17] , \wRegInTop_7_8[19] , \wRegOut_5_13[18] , 
        \wRegInTop_5_16[4] , \wRegInTop_5_20[15] , \wRegOut_6_32[9] , 
        \ScanLink232[3] , \wRegOut_5_30[29] , \wRegInBot_6_2[23] , 
        \wRegOut_5_30[30] , \wRegInTop_6_7[30] , \wRegInTop_6_7[29] , 
        \wRegOut_6_48[1] , \wRegOut_7_69[7] , \wRegInTop_6_38[23] , 
        \wRegInBot_6_58[20] , \wRegInTop_7_43[23] , \wRegOut_7_108[24] , 
        \wRegInTop_6_47[6] , \ScanLink135[1] , \wRegInTop_7_36[13] , 
        \wRegInTop_7_66[0] , \wRegInTop_7_15[22] , \wRegInTop_7_60[12] , 
        \ScanLink203[18] , \ScanLink220[30] , \ScanLink255[19] , 
        \wRegOut_4_9[8] , \wRegOut_5_3[20] , \wRegOut_5_19[3] , 
        \ScanLink68[18] , \wRegOut_7_74[8] , \wRegInTop_7_75[26] , 
        \ScanLink220[29] , \ScanLink255[4] , \wRegInTop_6_58[27] , 
        \wRegInTop_7_56[17] , \wRegInBot_6_38[24] , \wRegInTop_7_23[27] , 
        \wRegInBot_5_16[24] , \wRegInTop_5_15[7] , \wRegInTop_5_16[23] , 
        \wRegEnBot_5_16[0] , \wRegInTop_5_20[26] , \wRegInBot_5_20[21] , 
        \wRegInTop_6_44[5] , \ScanLink136[2] , \wRegInTop_7_65[3] , 
        \ScanLink93[19] , \wRegOut_6_48[31] , \wRegOut_6_48[28] , 
        \wRegOut_7_4[24] , \wRegOut_7_33[28] , \wRegOut_7_10[19] , 
        \wRegOut_7_33[31] , \wRegOut_7_46[18] , \wRegOut_7_65[30] , 
        \wRegOut_7_65[29] , \ScanLink198[2] , \wRegInTop_7_123[21] , 
        \wRegOut_5_18[14] , \wRegOut_7_80[10] , \wRegInTop_7_100[10] , 
        \wRegOut_6_37[4] , \wRegOut_7_16[2] , \wRegOut_7_95[24] , 
        \wRegInTop_7_115[24] , \wRegInTop_3_3[28] , \ScanLink69[9] , 
        \wRegOut_7_8[4] , \wRegInTop_7_118[8] , \ScanLink20[21] , 
        \wRegOut_7_103[28] , \wRegInBot_1_1[15] , \wRegOut_2_0[25] , 
        \ScanLink16[24] , \ScanLink55[11] , \ScanLink76[20] , 
        \wRegInTop_6_38[3] , \wRegInTop_7_19[5] , \ScanLink208[14] , 
        \wRegOut_7_103[31] , \wRegOut_7_120[19] , \wRegInBot_4_13[18] , 
        \ScanLink35[15] , \wRegInBot_5_24[4] , \ScanLink63[14] , 
        \wRegInBot_6_10[19] , \wRegInBot_6_33[31] , \wRegInTop_7_105[7] , 
        \wRegInBot_6_46[18] , \ScanLink40[25] , \ScanLink74[6] , 
        \wRegInBot_6_33[28] , \wRegInBot_5_1[28] , \wRegInBot_5_27[7] , 
        \ScanLink100[13] , \ScanLink175[23] , \ScanLink123[22] , 
        \ScanLink156[12] , \ScanLink143[26] , \ScanLink149[7] , 
        \wRegInTop_7_106[4] , \ScanLink77[5] , \ScanLink136[16] , 
        \wRegOut_6_29[8] , \ScanLink98[15] , \ScanLink160[17] , 
        \wRegInTop_7_3[26] , \ScanLink115[27] , \ScanLink229[2] , 
        \ScanLink16[17] , \wRegInBot_5_1[31] , \wRegOut_6_23[20] , 
        \wRegOut_6_56[10] , \wRegInTop_5_4[22] , \wRegOut_6_43[24] , 
        \ScanLink154[8] , \wRegOut_7_58[20] , \wRegOut_7_38[24] , 
        \wRegEnTop_5_24[0] , \wRegOut_6_15[25] , \wRegOut_6_34[7] , 
        \wRegOut_6_36[14] , \wRegOut_6_60[15] , \wRegOut_7_15[1] , 
        \ScanLink63[27] , \wRegInTop_6_26[31] , \ScanLink35[26] , 
        \ScanLink40[16] , \wRegInTop_6_53[18] , \wRegInTop_6_26[28] , 
        \wRegInTop_7_28[18] , \ScanLink55[22] , \wRegOut_6_0[18] , 
        \ScanLink208[27] , \wRegOut_2_0[16] , \ScanLink10[2] , 
        \ScanLink20[12] , \wRegInBot_3_6[11] , \wRegOut_5_18[27] , 
        \wRegInBot_6_11[2] , \ScanLink76[13] , \wRegInTop_6_41[8] , 
        \wRegOut_7_95[17] , \wCtrlOut_7[0] , \wRegInTop_7_115[17] , 
        \wRegInTop_7_123[12] , \wRegOut_6_53[0] , \wRegInTop_7_100[23] , 
        \wRegOut_7_72[6] , \wRegInTop_5_4[11] , \wRegOut_6_36[27] , 
        \wRegOut_7_80[23] , \wRegOut_7_38[17] , \wRegInBot_6_12[1] , 
        \wRegOut_6_15[16] , \wRegOut_6_43[17] , \wRegOut_6_60[26] , 
        \ScanLink4[19] , \wRegInTop_5_13[9] , \wRegOut_6_23[13] , 
        \wRegOut_6_50[3] , \wRegOut_7_71[5] , \ScanLink250[9] , 
        \ScanLink98[26] , \ScanLink115[14] , \wRegOut_6_56[23] , 
        \wRegOut_7_58[13] , \ScanLink136[25] , \ScanLink143[15] , 
        \ScanLink160[24] , \wRegInTop_7_85[18] , \wRegInTop_7_3[15] , 
        \ScanLink100[20] , \ScanLink123[11] , \ScanLink175[10] , 
        \ScanLink13[1] , \ScanLink156[21] , \wRegEnTop_7_30[0] ;
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink13[31] , \ScanLink13[30] , \ScanLink13[29] , 
        \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , \ScanLink13[25] , 
        \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , \ScanLink13[21] , 
        \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , \ScanLink13[17] , 
        \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , \ScanLink13[13] , 
        \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , \ScanLink13[9] , 
        \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , \ScanLink13[5] , 
        \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , \ScanLink13[1] , 
        \ScanLink13[0] }), .ScanOut({\ScanLink12[31] , \ScanLink12[30] , 
        \ScanLink12[29] , \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , 
        \ScanLink12[25] , \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , 
        \ScanLink12[21] , \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , 
        \ScanLink12[17] , \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , 
        \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , 
        \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , 
        \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , 
        \ScanLink12[1] , \ScanLink12[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_5[31] , \wRegOut_3_5[30] , \wRegOut_3_5[29] , 
        \wRegOut_3_5[28] , \wRegOut_3_5[27] , \wRegOut_3_5[26] , 
        \wRegOut_3_5[25] , \wRegOut_3_5[24] , \wRegOut_3_5[23] , 
        \wRegOut_3_5[22] , \wRegOut_3_5[21] , \wRegOut_3_5[20] , 
        \wRegOut_3_5[19] , \wRegOut_3_5[18] , \wRegOut_3_5[17] , 
        \wRegOut_3_5[16] , \wRegOut_3_5[15] , \wRegOut_3_5[14] , 
        \wRegOut_3_5[13] , \wRegOut_3_5[12] , \wRegOut_3_5[11] , 
        \wRegOut_3_5[10] , \wRegOut_3_5[9] , \wRegOut_3_5[8] , 
        \wRegOut_3_5[7] , \wRegOut_3_5[6] , \wRegOut_3_5[5] , \wRegOut_3_5[4] , 
        \wRegOut_3_5[3] , \wRegOut_3_5[2] , \wRegOut_3_5[1] , \wRegOut_3_5[0] 
        }), .Enable1(\wRegEnTop_3_5[0] ), .Enable2(\wRegEnBot_3_5[0] ), .In1({
        \wRegInTop_3_5[31] , \wRegInTop_3_5[30] , \wRegInTop_3_5[29] , 
        \wRegInTop_3_5[28] , \wRegInTop_3_5[27] , \wRegInTop_3_5[26] , 
        \wRegInTop_3_5[25] , \wRegInTop_3_5[24] , \wRegInTop_3_5[23] , 
        \wRegInTop_3_5[22] , \wRegInTop_3_5[21] , \wRegInTop_3_5[20] , 
        \wRegInTop_3_5[19] , \wRegInTop_3_5[18] , \wRegInTop_3_5[17] , 
        \wRegInTop_3_5[16] , \wRegInTop_3_5[15] , \wRegInTop_3_5[14] , 
        \wRegInTop_3_5[13] , \wRegInTop_3_5[12] , \wRegInTop_3_5[11] , 
        \wRegInTop_3_5[10] , \wRegInTop_3_5[9] , \wRegInTop_3_5[8] , 
        \wRegInTop_3_5[7] , \wRegInTop_3_5[6] , \wRegInTop_3_5[5] , 
        \wRegInTop_3_5[4] , \wRegInTop_3_5[3] , \wRegInTop_3_5[2] , 
        \wRegInTop_3_5[1] , \wRegInTop_3_5[0] }), .In2({\wRegInBot_3_5[31] , 
        \wRegInBot_3_5[30] , \wRegInBot_3_5[29] , \wRegInBot_3_5[28] , 
        \wRegInBot_3_5[27] , \wRegInBot_3_5[26] , \wRegInBot_3_5[25] , 
        \wRegInBot_3_5[24] , \wRegInBot_3_5[23] , \wRegInBot_3_5[22] , 
        \wRegInBot_3_5[21] , \wRegInBot_3_5[20] , \wRegInBot_3_5[19] , 
        \wRegInBot_3_5[18] , \wRegInBot_3_5[17] , \wRegInBot_3_5[16] , 
        \wRegInBot_3_5[15] , \wRegInBot_3_5[14] , \wRegInBot_3_5[13] , 
        \wRegInBot_3_5[12] , \wRegInBot_3_5[11] , \wRegInBot_3_5[10] , 
        \wRegInBot_3_5[9] , \wRegInBot_3_5[8] , \wRegInBot_3_5[7] , 
        \wRegInBot_3_5[6] , \wRegInBot_3_5[5] , \wRegInBot_3_5[4] , 
        \wRegInBot_3_5[3] , \wRegInBot_3_5[2] , \wRegInBot_3_5[1] , 
        \wRegInBot_3_5[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_26 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink58[31] , \ScanLink58[30] , \ScanLink58[29] , 
        \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , \ScanLink58[25] , 
        \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , \ScanLink58[21] , 
        \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , \ScanLink58[17] , 
        \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , \ScanLink58[13] , 
        \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , \ScanLink58[9] , 
        \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , \ScanLink58[5] , 
        \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , \ScanLink58[1] , 
        \ScanLink58[0] }), .ScanOut({\ScanLink57[31] , \ScanLink57[30] , 
        \ScanLink57[29] , \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , 
        \ScanLink57[25] , \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , 
        \ScanLink57[21] , \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , 
        \ScanLink57[17] , \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , 
        \ScanLink57[13] , \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , 
        \ScanLink57[9] , \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , 
        \ScanLink57[5] , \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , 
        \ScanLink57[1] , \ScanLink57[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_26[31] , \wRegOut_5_26[30] , 
        \wRegOut_5_26[29] , \wRegOut_5_26[28] , \wRegOut_5_26[27] , 
        \wRegOut_5_26[26] , \wRegOut_5_26[25] , \wRegOut_5_26[24] , 
        \wRegOut_5_26[23] , \wRegOut_5_26[22] , \wRegOut_5_26[21] , 
        \wRegOut_5_26[20] , \wRegOut_5_26[19] , \wRegOut_5_26[18] , 
        \wRegOut_5_26[17] , \wRegOut_5_26[16] , \wRegOut_5_26[15] , 
        \wRegOut_5_26[14] , \wRegOut_5_26[13] , \wRegOut_5_26[12] , 
        \wRegOut_5_26[11] , \wRegOut_5_26[10] , \wRegOut_5_26[9] , 
        \wRegOut_5_26[8] , \wRegOut_5_26[7] , \wRegOut_5_26[6] , 
        \wRegOut_5_26[5] , \wRegOut_5_26[4] , \wRegOut_5_26[3] , 
        \wRegOut_5_26[2] , \wRegOut_5_26[1] , \wRegOut_5_26[0] }), .Enable1(
        \wRegEnTop_5_26[0] ), .Enable2(\wRegEnBot_5_26[0] ), .In1({
        \wRegInTop_5_26[31] , \wRegInTop_5_26[30] , \wRegInTop_5_26[29] , 
        \wRegInTop_5_26[28] , \wRegInTop_5_26[27] , \wRegInTop_5_26[26] , 
        \wRegInTop_5_26[25] , \wRegInTop_5_26[24] , \wRegInTop_5_26[23] , 
        \wRegInTop_5_26[22] , \wRegInTop_5_26[21] , \wRegInTop_5_26[20] , 
        \wRegInTop_5_26[19] , \wRegInTop_5_26[18] , \wRegInTop_5_26[17] , 
        \wRegInTop_5_26[16] , \wRegInTop_5_26[15] , \wRegInTop_5_26[14] , 
        \wRegInTop_5_26[13] , \wRegInTop_5_26[12] , \wRegInTop_5_26[11] , 
        \wRegInTop_5_26[10] , \wRegInTop_5_26[9] , \wRegInTop_5_26[8] , 
        \wRegInTop_5_26[7] , \wRegInTop_5_26[6] , \wRegInTop_5_26[5] , 
        \wRegInTop_5_26[4] , \wRegInTop_5_26[3] , \wRegInTop_5_26[2] , 
        \wRegInTop_5_26[1] , \wRegInTop_5_26[0] }), .In2({\wRegInBot_5_26[31] , 
        \wRegInBot_5_26[30] , \wRegInBot_5_26[29] , \wRegInBot_5_26[28] , 
        \wRegInBot_5_26[27] , \wRegInBot_5_26[26] , \wRegInBot_5_26[25] , 
        \wRegInBot_5_26[24] , \wRegInBot_5_26[23] , \wRegInBot_5_26[22] , 
        \wRegInBot_5_26[21] , \wRegInBot_5_26[20] , \wRegInBot_5_26[19] , 
        \wRegInBot_5_26[18] , \wRegInBot_5_26[17] , \wRegInBot_5_26[16] , 
        \wRegInBot_5_26[15] , \wRegInBot_5_26[14] , \wRegInBot_5_26[13] , 
        \wRegInBot_5_26[12] , \wRegInBot_5_26[11] , \wRegInBot_5_26[10] , 
        \wRegInBot_5_26[9] , \wRegInBot_5_26[8] , \wRegInBot_5_26[7] , 
        \wRegInBot_5_26[6] , \wRegInBot_5_26[5] , \wRegInBot_5_26[4] , 
        \wRegInBot_5_26[3] , \wRegInBot_5_26[2] , \wRegInBot_5_26[1] , 
        \wRegInBot_5_26[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_16 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink80[31] , \ScanLink80[30] , \ScanLink80[29] , 
        \ScanLink80[28] , \ScanLink80[27] , \ScanLink80[26] , \ScanLink80[25] , 
        \ScanLink80[24] , \ScanLink80[23] , \ScanLink80[22] , \ScanLink80[21] , 
        \ScanLink80[20] , \ScanLink80[19] , \ScanLink80[18] , \ScanLink80[17] , 
        \ScanLink80[16] , \ScanLink80[15] , \ScanLink80[14] , \ScanLink80[13] , 
        \ScanLink80[12] , \ScanLink80[11] , \ScanLink80[10] , \ScanLink80[9] , 
        \ScanLink80[8] , \ScanLink80[7] , \ScanLink80[6] , \ScanLink80[5] , 
        \ScanLink80[4] , \ScanLink80[3] , \ScanLink80[2] , \ScanLink80[1] , 
        \ScanLink80[0] }), .ScanOut({\ScanLink79[31] , \ScanLink79[30] , 
        \ScanLink79[29] , \ScanLink79[28] , \ScanLink79[27] , \ScanLink79[26] , 
        \ScanLink79[25] , \ScanLink79[24] , \ScanLink79[23] , \ScanLink79[22] , 
        \ScanLink79[21] , \ScanLink79[20] , \ScanLink79[19] , \ScanLink79[18] , 
        \ScanLink79[17] , \ScanLink79[16] , \ScanLink79[15] , \ScanLink79[14] , 
        \ScanLink79[13] , \ScanLink79[12] , \ScanLink79[11] , \ScanLink79[10] , 
        \ScanLink79[9] , \ScanLink79[8] , \ScanLink79[7] , \ScanLink79[6] , 
        \ScanLink79[5] , \ScanLink79[4] , \ScanLink79[3] , \ScanLink79[2] , 
        \ScanLink79[1] , \ScanLink79[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_16[31] , \wRegOut_6_16[30] , 
        \wRegOut_6_16[29] , \wRegOut_6_16[28] , \wRegOut_6_16[27] , 
        \wRegOut_6_16[26] , \wRegOut_6_16[25] , \wRegOut_6_16[24] , 
        \wRegOut_6_16[23] , \wRegOut_6_16[22] , \wRegOut_6_16[21] , 
        \wRegOut_6_16[20] , \wRegOut_6_16[19] , \wRegOut_6_16[18] , 
        \wRegOut_6_16[17] , \wRegOut_6_16[16] , \wRegOut_6_16[15] , 
        \wRegOut_6_16[14] , \wRegOut_6_16[13] , \wRegOut_6_16[12] , 
        \wRegOut_6_16[11] , \wRegOut_6_16[10] , \wRegOut_6_16[9] , 
        \wRegOut_6_16[8] , \wRegOut_6_16[7] , \wRegOut_6_16[6] , 
        \wRegOut_6_16[5] , \wRegOut_6_16[4] , \wRegOut_6_16[3] , 
        \wRegOut_6_16[2] , \wRegOut_6_16[1] , \wRegOut_6_16[0] }), .Enable1(
        \wRegEnTop_6_16[0] ), .Enable2(\wRegEnBot_6_16[0] ), .In1({
        \wRegInTop_6_16[31] , \wRegInTop_6_16[30] , \wRegInTop_6_16[29] , 
        \wRegInTop_6_16[28] , \wRegInTop_6_16[27] , \wRegInTop_6_16[26] , 
        \wRegInTop_6_16[25] , \wRegInTop_6_16[24] , \wRegInTop_6_16[23] , 
        \wRegInTop_6_16[22] , \wRegInTop_6_16[21] , \wRegInTop_6_16[20] , 
        \wRegInTop_6_16[19] , \wRegInTop_6_16[18] , \wRegInTop_6_16[17] , 
        \wRegInTop_6_16[16] , \wRegInTop_6_16[15] , \wRegInTop_6_16[14] , 
        \wRegInTop_6_16[13] , \wRegInTop_6_16[12] , \wRegInTop_6_16[11] , 
        \wRegInTop_6_16[10] , \wRegInTop_6_16[9] , \wRegInTop_6_16[8] , 
        \wRegInTop_6_16[7] , \wRegInTop_6_16[6] , \wRegInTop_6_16[5] , 
        \wRegInTop_6_16[4] , \wRegInTop_6_16[3] , \wRegInTop_6_16[2] , 
        \wRegInTop_6_16[1] , \wRegInTop_6_16[0] }), .In2({\wRegInBot_6_16[31] , 
        \wRegInBot_6_16[30] , \wRegInBot_6_16[29] , \wRegInBot_6_16[28] , 
        \wRegInBot_6_16[27] , \wRegInBot_6_16[26] , \wRegInBot_6_16[25] , 
        \wRegInBot_6_16[24] , \wRegInBot_6_16[23] , \wRegInBot_6_16[22] , 
        \wRegInBot_6_16[21] , \wRegInBot_6_16[20] , \wRegInBot_6_16[19] , 
        \wRegInBot_6_16[18] , \wRegInBot_6_16[17] , \wRegInBot_6_16[16] , 
        \wRegInBot_6_16[15] , \wRegInBot_6_16[14] , \wRegInBot_6_16[13] , 
        \wRegInBot_6_16[12] , \wRegInBot_6_16[11] , \wRegInBot_6_16[10] , 
        \wRegInBot_6_16[9] , \wRegInBot_6_16[8] , \wRegInBot_6_16[7] , 
        \wRegInBot_6_16[6] , \wRegInBot_6_16[5] , \wRegInBot_6_16[4] , 
        \wRegInBot_6_16[3] , \wRegInBot_6_16[2] , \wRegInBot_6_16[1] , 
        \wRegInBot_6_16[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_62 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink190[31] , \ScanLink190[30] , \ScanLink190[29] , 
        \ScanLink190[28] , \ScanLink190[27] , \ScanLink190[26] , 
        \ScanLink190[25] , \ScanLink190[24] , \ScanLink190[23] , 
        \ScanLink190[22] , \ScanLink190[21] , \ScanLink190[20] , 
        \ScanLink190[19] , \ScanLink190[18] , \ScanLink190[17] , 
        \ScanLink190[16] , \ScanLink190[15] , \ScanLink190[14] , 
        \ScanLink190[13] , \ScanLink190[12] , \ScanLink190[11] , 
        \ScanLink190[10] , \ScanLink190[9] , \ScanLink190[8] , 
        \ScanLink190[7] , \ScanLink190[6] , \ScanLink190[5] , \ScanLink190[4] , 
        \ScanLink190[3] , \ScanLink190[2] , \ScanLink190[1] , \ScanLink190[0] 
        }), .ScanOut({\ScanLink189[31] , \ScanLink189[30] , \ScanLink189[29] , 
        \ScanLink189[28] , \ScanLink189[27] , \ScanLink189[26] , 
        \ScanLink189[25] , \ScanLink189[24] , \ScanLink189[23] , 
        \ScanLink189[22] , \ScanLink189[21] , \ScanLink189[20] , 
        \ScanLink189[19] , \ScanLink189[18] , \ScanLink189[17] , 
        \ScanLink189[16] , \ScanLink189[15] , \ScanLink189[14] , 
        \ScanLink189[13] , \ScanLink189[12] , \ScanLink189[11] , 
        \ScanLink189[10] , \ScanLink189[9] , \ScanLink189[8] , 
        \ScanLink189[7] , \ScanLink189[6] , \ScanLink189[5] , \ScanLink189[4] , 
        \ScanLink189[3] , \ScanLink189[2] , \ScanLink189[1] , \ScanLink189[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_62[31] , 
        \wRegOut_7_62[30] , \wRegOut_7_62[29] , \wRegOut_7_62[28] , 
        \wRegOut_7_62[27] , \wRegOut_7_62[26] , \wRegOut_7_62[25] , 
        \wRegOut_7_62[24] , \wRegOut_7_62[23] , \wRegOut_7_62[22] , 
        \wRegOut_7_62[21] , \wRegOut_7_62[20] , \wRegOut_7_62[19] , 
        \wRegOut_7_62[18] , \wRegOut_7_62[17] , \wRegOut_7_62[16] , 
        \wRegOut_7_62[15] , \wRegOut_7_62[14] , \wRegOut_7_62[13] , 
        \wRegOut_7_62[12] , \wRegOut_7_62[11] , \wRegOut_7_62[10] , 
        \wRegOut_7_62[9] , \wRegOut_7_62[8] , \wRegOut_7_62[7] , 
        \wRegOut_7_62[6] , \wRegOut_7_62[5] , \wRegOut_7_62[4] , 
        \wRegOut_7_62[3] , \wRegOut_7_62[2] , \wRegOut_7_62[1] , 
        \wRegOut_7_62[0] }), .Enable1(\wRegEnTop_7_62[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_62[31] , \wRegInTop_7_62[30] , \wRegInTop_7_62[29] , 
        \wRegInTop_7_62[28] , \wRegInTop_7_62[27] , \wRegInTop_7_62[26] , 
        \wRegInTop_7_62[25] , \wRegInTop_7_62[24] , \wRegInTop_7_62[23] , 
        \wRegInTop_7_62[22] , \wRegInTop_7_62[21] , \wRegInTop_7_62[20] , 
        \wRegInTop_7_62[19] , \wRegInTop_7_62[18] , \wRegInTop_7_62[17] , 
        \wRegInTop_7_62[16] , \wRegInTop_7_62[15] , \wRegInTop_7_62[14] , 
        \wRegInTop_7_62[13] , \wRegInTop_7_62[12] , \wRegInTop_7_62[11] , 
        \wRegInTop_7_62[10] , \wRegInTop_7_62[9] , \wRegInTop_7_62[8] , 
        \wRegInTop_7_62[7] , \wRegInTop_7_62[6] , \wRegInTop_7_62[5] , 
        \wRegInTop_7_62[4] , \wRegInTop_7_62[3] , \wRegInTop_7_62[2] , 
        \wRegInTop_7_62[1] , \wRegInTop_7_62[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink67[31] , \ScanLink67[30] , \ScanLink67[29] , 
        \ScanLink67[28] , \ScanLink67[27] , \ScanLink67[26] , \ScanLink67[25] , 
        \ScanLink67[24] , \ScanLink67[23] , \ScanLink67[22] , \ScanLink67[21] , 
        \ScanLink67[20] , \ScanLink67[19] , \ScanLink67[18] , \ScanLink67[17] , 
        \ScanLink67[16] , \ScanLink67[15] , \ScanLink67[14] , \ScanLink67[13] , 
        \ScanLink67[12] , \ScanLink67[11] , \ScanLink67[10] , \ScanLink67[9] , 
        \ScanLink67[8] , \ScanLink67[7] , \ScanLink67[6] , \ScanLink67[5] , 
        \ScanLink67[4] , \ScanLink67[3] , \ScanLink67[2] , \ScanLink67[1] , 
        \ScanLink67[0] }), .ScanOut({\ScanLink66[31] , \ScanLink66[30] , 
        \ScanLink66[29] , \ScanLink66[28] , \ScanLink66[27] , \ScanLink66[26] , 
        \ScanLink66[25] , \ScanLink66[24] , \ScanLink66[23] , \ScanLink66[22] , 
        \ScanLink66[21] , \ScanLink66[20] , \ScanLink66[19] , \ScanLink66[18] , 
        \ScanLink66[17] , \ScanLink66[16] , \ScanLink66[15] , \ScanLink66[14] , 
        \ScanLink66[13] , \ScanLink66[12] , \ScanLink66[11] , \ScanLink66[10] , 
        \ScanLink66[9] , \ScanLink66[8] , \ScanLink66[7] , \ScanLink66[6] , 
        \ScanLink66[5] , \ScanLink66[4] , \ScanLink66[3] , \ScanLink66[2] , 
        \ScanLink66[1] , \ScanLink66[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_3[31] , \wRegOut_6_3[30] , \wRegOut_6_3[29] , 
        \wRegOut_6_3[28] , \wRegOut_6_3[27] , \wRegOut_6_3[26] , 
        \wRegOut_6_3[25] , \wRegOut_6_3[24] , \wRegOut_6_3[23] , 
        \wRegOut_6_3[22] , \wRegOut_6_3[21] , \wRegOut_6_3[20] , 
        \wRegOut_6_3[19] , \wRegOut_6_3[18] , \wRegOut_6_3[17] , 
        \wRegOut_6_3[16] , \wRegOut_6_3[15] , \wRegOut_6_3[14] , 
        \wRegOut_6_3[13] , \wRegOut_6_3[12] , \wRegOut_6_3[11] , 
        \wRegOut_6_3[10] , \wRegOut_6_3[9] , \wRegOut_6_3[8] , 
        \wRegOut_6_3[7] , \wRegOut_6_3[6] , \wRegOut_6_3[5] , \wRegOut_6_3[4] , 
        \wRegOut_6_3[3] , \wRegOut_6_3[2] , \wRegOut_6_3[1] , \wRegOut_6_3[0] 
        }), .Enable1(\wRegEnTop_6_3[0] ), .Enable2(\wRegEnBot_6_3[0] ), .In1({
        \wRegInTop_6_3[31] , \wRegInTop_6_3[30] , \wRegInTop_6_3[29] , 
        \wRegInTop_6_3[28] , \wRegInTop_6_3[27] , \wRegInTop_6_3[26] , 
        \wRegInTop_6_3[25] , \wRegInTop_6_3[24] , \wRegInTop_6_3[23] , 
        \wRegInTop_6_3[22] , \wRegInTop_6_3[21] , \wRegInTop_6_3[20] , 
        \wRegInTop_6_3[19] , \wRegInTop_6_3[18] , \wRegInTop_6_3[17] , 
        \wRegInTop_6_3[16] , \wRegInTop_6_3[15] , \wRegInTop_6_3[14] , 
        \wRegInTop_6_3[13] , \wRegInTop_6_3[12] , \wRegInTop_6_3[11] , 
        \wRegInTop_6_3[10] , \wRegInTop_6_3[9] , \wRegInTop_6_3[8] , 
        \wRegInTop_6_3[7] , \wRegInTop_6_3[6] , \wRegInTop_6_3[5] , 
        \wRegInTop_6_3[4] , \wRegInTop_6_3[3] , \wRegInTop_6_3[2] , 
        \wRegInTop_6_3[1] , \wRegInTop_6_3[0] }), .In2({\wRegInBot_6_3[31] , 
        \wRegInBot_6_3[30] , \wRegInBot_6_3[29] , \wRegInBot_6_3[28] , 
        \wRegInBot_6_3[27] , \wRegInBot_6_3[26] , \wRegInBot_6_3[25] , 
        \wRegInBot_6_3[24] , \wRegInBot_6_3[23] , \wRegInBot_6_3[22] , 
        \wRegInBot_6_3[21] , \wRegInBot_6_3[20] , \wRegInBot_6_3[19] , 
        \wRegInBot_6_3[18] , \wRegInBot_6_3[17] , \wRegInBot_6_3[16] , 
        \wRegInBot_6_3[15] , \wRegInBot_6_3[14] , \wRegInBot_6_3[13] , 
        \wRegInBot_6_3[12] , \wRegInBot_6_3[11] , \wRegInBot_6_3[10] , 
        \wRegInBot_6_3[9] , \wRegInBot_6_3[8] , \wRegInBot_6_3[7] , 
        \wRegInBot_6_3[6] , \wRegInBot_6_3[5] , \wRegInBot_6_3[4] , 
        \wRegInBot_6_3[3] , \wRegInBot_6_3[2] , \wRegInBot_6_3[1] , 
        \wRegInBot_6_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_31 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink95[31] , \ScanLink95[30] , \ScanLink95[29] , 
        \ScanLink95[28] , \ScanLink95[27] , \ScanLink95[26] , \ScanLink95[25] , 
        \ScanLink95[24] , \ScanLink95[23] , \ScanLink95[22] , \ScanLink95[21] , 
        \ScanLink95[20] , \ScanLink95[19] , \ScanLink95[18] , \ScanLink95[17] , 
        \ScanLink95[16] , \ScanLink95[15] , \ScanLink95[14] , \ScanLink95[13] , 
        \ScanLink95[12] , \ScanLink95[11] , \ScanLink95[10] , \ScanLink95[9] , 
        \ScanLink95[8] , \ScanLink95[7] , \ScanLink95[6] , \ScanLink95[5] , 
        \ScanLink95[4] , \ScanLink95[3] , \ScanLink95[2] , \ScanLink95[1] , 
        \ScanLink95[0] }), .ScanOut({\ScanLink94[31] , \ScanLink94[30] , 
        \ScanLink94[29] , \ScanLink94[28] , \ScanLink94[27] , \ScanLink94[26] , 
        \ScanLink94[25] , \ScanLink94[24] , \ScanLink94[23] , \ScanLink94[22] , 
        \ScanLink94[21] , \ScanLink94[20] , \ScanLink94[19] , \ScanLink94[18] , 
        \ScanLink94[17] , \ScanLink94[16] , \ScanLink94[15] , \ScanLink94[14] , 
        \ScanLink94[13] , \ScanLink94[12] , \ScanLink94[11] , \ScanLink94[10] , 
        \ScanLink94[9] , \ScanLink94[8] , \ScanLink94[7] , \ScanLink94[6] , 
        \ScanLink94[5] , \ScanLink94[4] , \ScanLink94[3] , \ScanLink94[2] , 
        \ScanLink94[1] , \ScanLink94[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_31[31] , \wRegOut_6_31[30] , 
        \wRegOut_6_31[29] , \wRegOut_6_31[28] , \wRegOut_6_31[27] , 
        \wRegOut_6_31[26] , \wRegOut_6_31[25] , \wRegOut_6_31[24] , 
        \wRegOut_6_31[23] , \wRegOut_6_31[22] , \wRegOut_6_31[21] , 
        \wRegOut_6_31[20] , \wRegOut_6_31[19] , \wRegOut_6_31[18] , 
        \wRegOut_6_31[17] , \wRegOut_6_31[16] , \wRegOut_6_31[15] , 
        \wRegOut_6_31[14] , \wRegOut_6_31[13] , \wRegOut_6_31[12] , 
        \wRegOut_6_31[11] , \wRegOut_6_31[10] , \wRegOut_6_31[9] , 
        \wRegOut_6_31[8] , \wRegOut_6_31[7] , \wRegOut_6_31[6] , 
        \wRegOut_6_31[5] , \wRegOut_6_31[4] , \wRegOut_6_31[3] , 
        \wRegOut_6_31[2] , \wRegOut_6_31[1] , \wRegOut_6_31[0] }), .Enable1(
        \wRegEnTop_6_31[0] ), .Enable2(\wRegEnBot_6_31[0] ), .In1({
        \wRegInTop_6_31[31] , \wRegInTop_6_31[30] , \wRegInTop_6_31[29] , 
        \wRegInTop_6_31[28] , \wRegInTop_6_31[27] , \wRegInTop_6_31[26] , 
        \wRegInTop_6_31[25] , \wRegInTop_6_31[24] , \wRegInTop_6_31[23] , 
        \wRegInTop_6_31[22] , \wRegInTop_6_31[21] , \wRegInTop_6_31[20] , 
        \wRegInTop_6_31[19] , \wRegInTop_6_31[18] , \wRegInTop_6_31[17] , 
        \wRegInTop_6_31[16] , \wRegInTop_6_31[15] , \wRegInTop_6_31[14] , 
        \wRegInTop_6_31[13] , \wRegInTop_6_31[12] , \wRegInTop_6_31[11] , 
        \wRegInTop_6_31[10] , \wRegInTop_6_31[9] , \wRegInTop_6_31[8] , 
        \wRegInTop_6_31[7] , \wRegInTop_6_31[6] , \wRegInTop_6_31[5] , 
        \wRegInTop_6_31[4] , \wRegInTop_6_31[3] , \wRegInTop_6_31[2] , 
        \wRegInTop_6_31[1] , \wRegInTop_6_31[0] }), .In2({\wRegInBot_6_31[31] , 
        \wRegInBot_6_31[30] , \wRegInBot_6_31[29] , \wRegInBot_6_31[28] , 
        \wRegInBot_6_31[27] , \wRegInBot_6_31[26] , \wRegInBot_6_31[25] , 
        \wRegInBot_6_31[24] , \wRegInBot_6_31[23] , \wRegInBot_6_31[22] , 
        \wRegInBot_6_31[21] , \wRegInBot_6_31[20] , \wRegInBot_6_31[19] , 
        \wRegInBot_6_31[18] , \wRegInBot_6_31[17] , \wRegInBot_6_31[16] , 
        \wRegInBot_6_31[15] , \wRegInBot_6_31[14] , \wRegInBot_6_31[13] , 
        \wRegInBot_6_31[12] , \wRegInBot_6_31[11] , \wRegInBot_6_31[10] , 
        \wRegInBot_6_31[9] , \wRegInBot_6_31[8] , \wRegInBot_6_31[7] , 
        \wRegInBot_6_31[6] , \wRegInBot_6_31[5] , \wRegInBot_6_31[4] , 
        \wRegInBot_6_31[3] , \wRegInBot_6_31[2] , \wRegInBot_6_31[1] , 
        \wRegInBot_6_31[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_44 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink108[31] , \ScanLink108[30] , \ScanLink108[29] , 
        \ScanLink108[28] , \ScanLink108[27] , \ScanLink108[26] , 
        \ScanLink108[25] , \ScanLink108[24] , \ScanLink108[23] , 
        \ScanLink108[22] , \ScanLink108[21] , \ScanLink108[20] , 
        \ScanLink108[19] , \ScanLink108[18] , \ScanLink108[17] , 
        \ScanLink108[16] , \ScanLink108[15] , \ScanLink108[14] , 
        \ScanLink108[13] , \ScanLink108[12] , \ScanLink108[11] , 
        \ScanLink108[10] , \ScanLink108[9] , \ScanLink108[8] , 
        \ScanLink108[7] , \ScanLink108[6] , \ScanLink108[5] , \ScanLink108[4] , 
        \ScanLink108[3] , \ScanLink108[2] , \ScanLink108[1] , \ScanLink108[0] 
        }), .ScanOut({\ScanLink107[31] , \ScanLink107[30] , \ScanLink107[29] , 
        \ScanLink107[28] , \ScanLink107[27] , \ScanLink107[26] , 
        \ScanLink107[25] , \ScanLink107[24] , \ScanLink107[23] , 
        \ScanLink107[22] , \ScanLink107[21] , \ScanLink107[20] , 
        \ScanLink107[19] , \ScanLink107[18] , \ScanLink107[17] , 
        \ScanLink107[16] , \ScanLink107[15] , \ScanLink107[14] , 
        \ScanLink107[13] , \ScanLink107[12] , \ScanLink107[11] , 
        \ScanLink107[10] , \ScanLink107[9] , \ScanLink107[8] , 
        \ScanLink107[7] , \ScanLink107[6] , \ScanLink107[5] , \ScanLink107[4] , 
        \ScanLink107[3] , \ScanLink107[2] , \ScanLink107[1] , \ScanLink107[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_44[31] , 
        \wRegOut_6_44[30] , \wRegOut_6_44[29] , \wRegOut_6_44[28] , 
        \wRegOut_6_44[27] , \wRegOut_6_44[26] , \wRegOut_6_44[25] , 
        \wRegOut_6_44[24] , \wRegOut_6_44[23] , \wRegOut_6_44[22] , 
        \wRegOut_6_44[21] , \wRegOut_6_44[20] , \wRegOut_6_44[19] , 
        \wRegOut_6_44[18] , \wRegOut_6_44[17] , \wRegOut_6_44[16] , 
        \wRegOut_6_44[15] , \wRegOut_6_44[14] , \wRegOut_6_44[13] , 
        \wRegOut_6_44[12] , \wRegOut_6_44[11] , \wRegOut_6_44[10] , 
        \wRegOut_6_44[9] , \wRegOut_6_44[8] , \wRegOut_6_44[7] , 
        \wRegOut_6_44[6] , \wRegOut_6_44[5] , \wRegOut_6_44[4] , 
        \wRegOut_6_44[3] , \wRegOut_6_44[2] , \wRegOut_6_44[1] , 
        \wRegOut_6_44[0] }), .Enable1(\wRegEnTop_6_44[0] ), .Enable2(
        \wRegEnBot_6_44[0] ), .In1({\wRegInTop_6_44[31] , \wRegInTop_6_44[30] , 
        \wRegInTop_6_44[29] , \wRegInTop_6_44[28] , \wRegInTop_6_44[27] , 
        \wRegInTop_6_44[26] , \wRegInTop_6_44[25] , \wRegInTop_6_44[24] , 
        \wRegInTop_6_44[23] , \wRegInTop_6_44[22] , \wRegInTop_6_44[21] , 
        \wRegInTop_6_44[20] , \wRegInTop_6_44[19] , \wRegInTop_6_44[18] , 
        \wRegInTop_6_44[17] , \wRegInTop_6_44[16] , \wRegInTop_6_44[15] , 
        \wRegInTop_6_44[14] , \wRegInTop_6_44[13] , \wRegInTop_6_44[12] , 
        \wRegInTop_6_44[11] , \wRegInTop_6_44[10] , \wRegInTop_6_44[9] , 
        \wRegInTop_6_44[8] , \wRegInTop_6_44[7] , \wRegInTop_6_44[6] , 
        \wRegInTop_6_44[5] , \wRegInTop_6_44[4] , \wRegInTop_6_44[3] , 
        \wRegInTop_6_44[2] , \wRegInTop_6_44[1] , \wRegInTop_6_44[0] }), .In2(
        {\wRegInBot_6_44[31] , \wRegInBot_6_44[30] , \wRegInBot_6_44[29] , 
        \wRegInBot_6_44[28] , \wRegInBot_6_44[27] , \wRegInBot_6_44[26] , 
        \wRegInBot_6_44[25] , \wRegInBot_6_44[24] , \wRegInBot_6_44[23] , 
        \wRegInBot_6_44[22] , \wRegInBot_6_44[21] , \wRegInBot_6_44[20] , 
        \wRegInBot_6_44[19] , \wRegInBot_6_44[18] , \wRegInBot_6_44[17] , 
        \wRegInBot_6_44[16] , \wRegInBot_6_44[15] , \wRegInBot_6_44[14] , 
        \wRegInBot_6_44[13] , \wRegInBot_6_44[12] , \wRegInBot_6_44[11] , 
        \wRegInBot_6_44[10] , \wRegInBot_6_44[9] , \wRegInBot_6_44[8] , 
        \wRegInBot_6_44[7] , \wRegInBot_6_44[6] , \wRegInBot_6_44[5] , 
        \wRegInBot_6_44[4] , \wRegInBot_6_44[3] , \wRegInBot_6_44[2] , 
        \wRegInBot_6_44[1] , \wRegInBot_6_44[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_63 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink127[31] , \ScanLink127[30] , \ScanLink127[29] , 
        \ScanLink127[28] , \ScanLink127[27] , \ScanLink127[26] , 
        \ScanLink127[25] , \ScanLink127[24] , \ScanLink127[23] , 
        \ScanLink127[22] , \ScanLink127[21] , \ScanLink127[20] , 
        \ScanLink127[19] , \ScanLink127[18] , \ScanLink127[17] , 
        \ScanLink127[16] , \ScanLink127[15] , \ScanLink127[14] , 
        \ScanLink127[13] , \ScanLink127[12] , \ScanLink127[11] , 
        \ScanLink127[10] , \ScanLink127[9] , \ScanLink127[8] , 
        \ScanLink127[7] , \ScanLink127[6] , \ScanLink127[5] , \ScanLink127[4] , 
        \ScanLink127[3] , \ScanLink127[2] , \ScanLink127[1] , \ScanLink127[0] 
        }), .ScanOut({\ScanLink126[31] , \ScanLink126[30] , \ScanLink126[29] , 
        \ScanLink126[28] , \ScanLink126[27] , \ScanLink126[26] , 
        \ScanLink126[25] , \ScanLink126[24] , \ScanLink126[23] , 
        \ScanLink126[22] , \ScanLink126[21] , \ScanLink126[20] , 
        \ScanLink126[19] , \ScanLink126[18] , \ScanLink126[17] , 
        \ScanLink126[16] , \ScanLink126[15] , \ScanLink126[14] , 
        \ScanLink126[13] , \ScanLink126[12] , \ScanLink126[11] , 
        \ScanLink126[10] , \ScanLink126[9] , \ScanLink126[8] , 
        \ScanLink126[7] , \ScanLink126[6] , \ScanLink126[5] , \ScanLink126[4] , 
        \ScanLink126[3] , \ScanLink126[2] , \ScanLink126[1] , \ScanLink126[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_63[31] , 
        \wRegOut_6_63[30] , \wRegOut_6_63[29] , \wRegOut_6_63[28] , 
        \wRegOut_6_63[27] , \wRegOut_6_63[26] , \wRegOut_6_63[25] , 
        \wRegOut_6_63[24] , \wRegOut_6_63[23] , \wRegOut_6_63[22] , 
        \wRegOut_6_63[21] , \wRegOut_6_63[20] , \wRegOut_6_63[19] , 
        \wRegOut_6_63[18] , \wRegOut_6_63[17] , \wRegOut_6_63[16] , 
        \wRegOut_6_63[15] , \wRegOut_6_63[14] , \wRegOut_6_63[13] , 
        \wRegOut_6_63[12] , \wRegOut_6_63[11] , \wRegOut_6_63[10] , 
        \wRegOut_6_63[9] , \wRegOut_6_63[8] , \wRegOut_6_63[7] , 
        \wRegOut_6_63[6] , \wRegOut_6_63[5] , \wRegOut_6_63[4] , 
        \wRegOut_6_63[3] , \wRegOut_6_63[2] , \wRegOut_6_63[1] , 
        \wRegOut_6_63[0] }), .Enable1(\wRegEnTop_6_63[0] ), .Enable2(
        \wRegEnBot_6_63[0] ), .In1({\wRegInTop_6_63[31] , \wRegInTop_6_63[30] , 
        \wRegInTop_6_63[29] , \wRegInTop_6_63[28] , \wRegInTop_6_63[27] , 
        \wRegInTop_6_63[26] , \wRegInTop_6_63[25] , \wRegInTop_6_63[24] , 
        \wRegInTop_6_63[23] , \wRegInTop_6_63[22] , \wRegInTop_6_63[21] , 
        \wRegInTop_6_63[20] , \wRegInTop_6_63[19] , \wRegInTop_6_63[18] , 
        \wRegInTop_6_63[17] , \wRegInTop_6_63[16] , \wRegInTop_6_63[15] , 
        \wRegInTop_6_63[14] , \wRegInTop_6_63[13] , \wRegInTop_6_63[12] , 
        \wRegInTop_6_63[11] , \wRegInTop_6_63[10] , \wRegInTop_6_63[9] , 
        \wRegInTop_6_63[8] , \wRegInTop_6_63[7] , \wRegInTop_6_63[6] , 
        \wRegInTop_6_63[5] , \wRegInTop_6_63[4] , \wRegInTop_6_63[3] , 
        \wRegInTop_6_63[2] , \wRegInTop_6_63[1] , \wRegInTop_6_63[0] }), .In2(
        {\wRegInBot_6_63[31] , \wRegInBot_6_63[30] , \wRegInBot_6_63[29] , 
        \wRegInBot_6_63[28] , \wRegInBot_6_63[27] , \wRegInBot_6_63[26] , 
        \wRegInBot_6_63[25] , \wRegInBot_6_63[24] , \wRegInBot_6_63[23] , 
        \wRegInBot_6_63[22] , \wRegInBot_6_63[21] , \wRegInBot_6_63[20] , 
        \wRegInBot_6_63[19] , \wRegInBot_6_63[18] , \wRegInBot_6_63[17] , 
        \wRegInBot_6_63[16] , \wRegInBot_6_63[15] , \wRegInBot_6_63[14] , 
        \wRegInBot_6_63[13] , \wRegInBot_6_63[12] , \wRegInBot_6_63[11] , 
        \wRegInBot_6_63[10] , \wRegInBot_6_63[9] , \wRegInBot_6_63[8] , 
        \wRegInBot_6_63[7] , \wRegInBot_6_63[6] , \wRegInBot_6_63[5] , 
        \wRegInBot_6_63[4] , \wRegInBot_6_63[3] , \wRegInBot_6_63[2] , 
        \wRegInBot_6_63[1] , \wRegInBot_6_63[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink131[31] , \ScanLink131[30] , \ScanLink131[29] , 
        \ScanLink131[28] , \ScanLink131[27] , \ScanLink131[26] , 
        \ScanLink131[25] , \ScanLink131[24] , \ScanLink131[23] , 
        \ScanLink131[22] , \ScanLink131[21] , \ScanLink131[20] , 
        \ScanLink131[19] , \ScanLink131[18] , \ScanLink131[17] , 
        \ScanLink131[16] , \ScanLink131[15] , \ScanLink131[14] , 
        \ScanLink131[13] , \ScanLink131[12] , \ScanLink131[11] , 
        \ScanLink131[10] , \ScanLink131[9] , \ScanLink131[8] , 
        \ScanLink131[7] , \ScanLink131[6] , \ScanLink131[5] , \ScanLink131[4] , 
        \ScanLink131[3] , \ScanLink131[2] , \ScanLink131[1] , \ScanLink131[0] 
        }), .ScanOut({\ScanLink130[31] , \ScanLink130[30] , \ScanLink130[29] , 
        \ScanLink130[28] , \ScanLink130[27] , \ScanLink130[26] , 
        \ScanLink130[25] , \ScanLink130[24] , \ScanLink130[23] , 
        \ScanLink130[22] , \ScanLink130[21] , \ScanLink130[20] , 
        \ScanLink130[19] , \ScanLink130[18] , \ScanLink130[17] , 
        \ScanLink130[16] , \ScanLink130[15] , \ScanLink130[14] , 
        \ScanLink130[13] , \ScanLink130[12] , \ScanLink130[11] , 
        \ScanLink130[10] , \ScanLink130[9] , \ScanLink130[8] , 
        \ScanLink130[7] , \ScanLink130[6] , \ScanLink130[5] , \ScanLink130[4] , 
        \ScanLink130[3] , \ScanLink130[2] , \ScanLink130[1] , \ScanLink130[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_3[31] , 
        \wRegOut_7_3[30] , \wRegOut_7_3[29] , \wRegOut_7_3[28] , 
        \wRegOut_7_3[27] , \wRegOut_7_3[26] , \wRegOut_7_3[25] , 
        \wRegOut_7_3[24] , \wRegOut_7_3[23] , \wRegOut_7_3[22] , 
        \wRegOut_7_3[21] , \wRegOut_7_3[20] , \wRegOut_7_3[19] , 
        \wRegOut_7_3[18] , \wRegOut_7_3[17] , \wRegOut_7_3[16] , 
        \wRegOut_7_3[15] , \wRegOut_7_3[14] , \wRegOut_7_3[13] , 
        \wRegOut_7_3[12] , \wRegOut_7_3[11] , \wRegOut_7_3[10] , 
        \wRegOut_7_3[9] , \wRegOut_7_3[8] , \wRegOut_7_3[7] , \wRegOut_7_3[6] , 
        \wRegOut_7_3[5] , \wRegOut_7_3[4] , \wRegOut_7_3[3] , \wRegOut_7_3[2] , 
        \wRegOut_7_3[1] , \wRegOut_7_3[0] }), .Enable1(\wRegEnTop_7_3[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_3[31] , \wRegInTop_7_3[30] , 
        \wRegInTop_7_3[29] , \wRegInTop_7_3[28] , \wRegInTop_7_3[27] , 
        \wRegInTop_7_3[26] , \wRegInTop_7_3[25] , \wRegInTop_7_3[24] , 
        \wRegInTop_7_3[23] , \wRegInTop_7_3[22] , \wRegInTop_7_3[21] , 
        \wRegInTop_7_3[20] , \wRegInTop_7_3[19] , \wRegInTop_7_3[18] , 
        \wRegInTop_7_3[17] , \wRegInTop_7_3[16] , \wRegInTop_7_3[15] , 
        \wRegInTop_7_3[14] , \wRegInTop_7_3[13] , \wRegInTop_7_3[12] , 
        \wRegInTop_7_3[11] , \wRegInTop_7_3[10] , \wRegInTop_7_3[9] , 
        \wRegInTop_7_3[8] , \wRegInTop_7_3[7] , \wRegInTop_7_3[6] , 
        \wRegInTop_7_3[5] , \wRegInTop_7_3[4] , \wRegInTop_7_3[3] , 
        \wRegInTop_7_3[2] , \wRegInTop_7_3[1] , \wRegInTop_7_3[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_45 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink173[31] , \ScanLink173[30] , \ScanLink173[29] , 
        \ScanLink173[28] , \ScanLink173[27] , \ScanLink173[26] , 
        \ScanLink173[25] , \ScanLink173[24] , \ScanLink173[23] , 
        \ScanLink173[22] , \ScanLink173[21] , \ScanLink173[20] , 
        \ScanLink173[19] , \ScanLink173[18] , \ScanLink173[17] , 
        \ScanLink173[16] , \ScanLink173[15] , \ScanLink173[14] , 
        \ScanLink173[13] , \ScanLink173[12] , \ScanLink173[11] , 
        \ScanLink173[10] , \ScanLink173[9] , \ScanLink173[8] , 
        \ScanLink173[7] , \ScanLink173[6] , \ScanLink173[5] , \ScanLink173[4] , 
        \ScanLink173[3] , \ScanLink173[2] , \ScanLink173[1] , \ScanLink173[0] 
        }), .ScanOut({\ScanLink172[31] , \ScanLink172[30] , \ScanLink172[29] , 
        \ScanLink172[28] , \ScanLink172[27] , \ScanLink172[26] , 
        \ScanLink172[25] , \ScanLink172[24] , \ScanLink172[23] , 
        \ScanLink172[22] , \ScanLink172[21] , \ScanLink172[20] , 
        \ScanLink172[19] , \ScanLink172[18] , \ScanLink172[17] , 
        \ScanLink172[16] , \ScanLink172[15] , \ScanLink172[14] , 
        \ScanLink172[13] , \ScanLink172[12] , \ScanLink172[11] , 
        \ScanLink172[10] , \ScanLink172[9] , \ScanLink172[8] , 
        \ScanLink172[7] , \ScanLink172[6] , \ScanLink172[5] , \ScanLink172[4] , 
        \ScanLink172[3] , \ScanLink172[2] , \ScanLink172[1] , \ScanLink172[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_45[31] , 
        \wRegOut_7_45[30] , \wRegOut_7_45[29] , \wRegOut_7_45[28] , 
        \wRegOut_7_45[27] , \wRegOut_7_45[26] , \wRegOut_7_45[25] , 
        \wRegOut_7_45[24] , \wRegOut_7_45[23] , \wRegOut_7_45[22] , 
        \wRegOut_7_45[21] , \wRegOut_7_45[20] , \wRegOut_7_45[19] , 
        \wRegOut_7_45[18] , \wRegOut_7_45[17] , \wRegOut_7_45[16] , 
        \wRegOut_7_45[15] , \wRegOut_7_45[14] , \wRegOut_7_45[13] , 
        \wRegOut_7_45[12] , \wRegOut_7_45[11] , \wRegOut_7_45[10] , 
        \wRegOut_7_45[9] , \wRegOut_7_45[8] , \wRegOut_7_45[7] , 
        \wRegOut_7_45[6] , \wRegOut_7_45[5] , \wRegOut_7_45[4] , 
        \wRegOut_7_45[3] , \wRegOut_7_45[2] , \wRegOut_7_45[1] , 
        \wRegOut_7_45[0] }), .Enable1(\wRegEnTop_7_45[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_45[31] , \wRegInTop_7_45[30] , \wRegInTop_7_45[29] , 
        \wRegInTop_7_45[28] , \wRegInTop_7_45[27] , \wRegInTop_7_45[26] , 
        \wRegInTop_7_45[25] , \wRegInTop_7_45[24] , \wRegInTop_7_45[23] , 
        \wRegInTop_7_45[22] , \wRegInTop_7_45[21] , \wRegInTop_7_45[20] , 
        \wRegInTop_7_45[19] , \wRegInTop_7_45[18] , \wRegInTop_7_45[17] , 
        \wRegInTop_7_45[16] , \wRegInTop_7_45[15] , \wRegInTop_7_45[14] , 
        \wRegInTop_7_45[13] , \wRegInTop_7_45[12] , \wRegInTop_7_45[11] , 
        \wRegInTop_7_45[10] , \wRegInTop_7_45[9] , \wRegInTop_7_45[8] , 
        \wRegInTop_7_45[7] , \wRegInTop_7_45[6] , \wRegInTop_7_45[5] , 
        \wRegInTop_7_45[4] , \wRegInTop_7_45[3] , \wRegInTop_7_45[2] , 
        \wRegInTop_7_45[1] , \wRegInTop_7_45[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_29[0] ), .P_In({\wRegOut_5_29[31] , 
        \wRegOut_5_29[30] , \wRegOut_5_29[29] , \wRegOut_5_29[28] , 
        \wRegOut_5_29[27] , \wRegOut_5_29[26] , \wRegOut_5_29[25] , 
        \wRegOut_5_29[24] , \wRegOut_5_29[23] , \wRegOut_5_29[22] , 
        \wRegOut_5_29[21] , \wRegOut_5_29[20] , \wRegOut_5_29[19] , 
        \wRegOut_5_29[18] , \wRegOut_5_29[17] , \wRegOut_5_29[16] , 
        \wRegOut_5_29[15] , \wRegOut_5_29[14] , \wRegOut_5_29[13] , 
        \wRegOut_5_29[12] , \wRegOut_5_29[11] , \wRegOut_5_29[10] , 
        \wRegOut_5_29[9] , \wRegOut_5_29[8] , \wRegOut_5_29[7] , 
        \wRegOut_5_29[6] , \wRegOut_5_29[5] , \wRegOut_5_29[4] , 
        \wRegOut_5_29[3] , \wRegOut_5_29[2] , \wRegOut_5_29[1] , 
        \wRegOut_5_29[0] }), .P_Out({\wRegInBot_5_29[31] , 
        \wRegInBot_5_29[30] , \wRegInBot_5_29[29] , \wRegInBot_5_29[28] , 
        \wRegInBot_5_29[27] , \wRegInBot_5_29[26] , \wRegInBot_5_29[25] , 
        \wRegInBot_5_29[24] , \wRegInBot_5_29[23] , \wRegInBot_5_29[22] , 
        \wRegInBot_5_29[21] , \wRegInBot_5_29[20] , \wRegInBot_5_29[19] , 
        \wRegInBot_5_29[18] , \wRegInBot_5_29[17] , \wRegInBot_5_29[16] , 
        \wRegInBot_5_29[15] , \wRegInBot_5_29[14] , \wRegInBot_5_29[13] , 
        \wRegInBot_5_29[12] , \wRegInBot_5_29[11] , \wRegInBot_5_29[10] , 
        \wRegInBot_5_29[9] , \wRegInBot_5_29[8] , \wRegInBot_5_29[7] , 
        \wRegInBot_5_29[6] , \wRegInBot_5_29[5] , \wRegInBot_5_29[4] , 
        \wRegInBot_5_29[3] , \wRegInBot_5_29[2] , \wRegInBot_5_29[1] , 
        \wRegInBot_5_29[0] }), .L_WR(\wRegEnTop_6_58[0] ), .L_In({
        \wRegOut_6_58[31] , \wRegOut_6_58[30] , \wRegOut_6_58[29] , 
        \wRegOut_6_58[28] , \wRegOut_6_58[27] , \wRegOut_6_58[26] , 
        \wRegOut_6_58[25] , \wRegOut_6_58[24] , \wRegOut_6_58[23] , 
        \wRegOut_6_58[22] , \wRegOut_6_58[21] , \wRegOut_6_58[20] , 
        \wRegOut_6_58[19] , \wRegOut_6_58[18] , \wRegOut_6_58[17] , 
        \wRegOut_6_58[16] , \wRegOut_6_58[15] , \wRegOut_6_58[14] , 
        \wRegOut_6_58[13] , \wRegOut_6_58[12] , \wRegOut_6_58[11] , 
        \wRegOut_6_58[10] , \wRegOut_6_58[9] , \wRegOut_6_58[8] , 
        \wRegOut_6_58[7] , \wRegOut_6_58[6] , \wRegOut_6_58[5] , 
        \wRegOut_6_58[4] , \wRegOut_6_58[3] , \wRegOut_6_58[2] , 
        \wRegOut_6_58[1] , \wRegOut_6_58[0] }), .L_Out({\wRegInTop_6_58[31] , 
        \wRegInTop_6_58[30] , \wRegInTop_6_58[29] , \wRegInTop_6_58[28] , 
        \wRegInTop_6_58[27] , \wRegInTop_6_58[26] , \wRegInTop_6_58[25] , 
        \wRegInTop_6_58[24] , \wRegInTop_6_58[23] , \wRegInTop_6_58[22] , 
        \wRegInTop_6_58[21] , \wRegInTop_6_58[20] , \wRegInTop_6_58[19] , 
        \wRegInTop_6_58[18] , \wRegInTop_6_58[17] , \wRegInTop_6_58[16] , 
        \wRegInTop_6_58[15] , \wRegInTop_6_58[14] , \wRegInTop_6_58[13] , 
        \wRegInTop_6_58[12] , \wRegInTop_6_58[11] , \wRegInTop_6_58[10] , 
        \wRegInTop_6_58[9] , \wRegInTop_6_58[8] , \wRegInTop_6_58[7] , 
        \wRegInTop_6_58[6] , \wRegInTop_6_58[5] , \wRegInTop_6_58[4] , 
        \wRegInTop_6_58[3] , \wRegInTop_6_58[2] , \wRegInTop_6_58[1] , 
        \wRegInTop_6_58[0] }), .R_WR(\wRegEnTop_6_59[0] ), .R_In({
        \wRegOut_6_59[31] , \wRegOut_6_59[30] , \wRegOut_6_59[29] , 
        \wRegOut_6_59[28] , \wRegOut_6_59[27] , \wRegOut_6_59[26] , 
        \wRegOut_6_59[25] , \wRegOut_6_59[24] , \wRegOut_6_59[23] , 
        \wRegOut_6_59[22] , \wRegOut_6_59[21] , \wRegOut_6_59[20] , 
        \wRegOut_6_59[19] , \wRegOut_6_59[18] , \wRegOut_6_59[17] , 
        \wRegOut_6_59[16] , \wRegOut_6_59[15] , \wRegOut_6_59[14] , 
        \wRegOut_6_59[13] , \wRegOut_6_59[12] , \wRegOut_6_59[11] , 
        \wRegOut_6_59[10] , \wRegOut_6_59[9] , \wRegOut_6_59[8] , 
        \wRegOut_6_59[7] , \wRegOut_6_59[6] , \wRegOut_6_59[5] , 
        \wRegOut_6_59[4] , \wRegOut_6_59[3] , \wRegOut_6_59[2] , 
        \wRegOut_6_59[1] , \wRegOut_6_59[0] }), .R_Out({\wRegInTop_6_59[31] , 
        \wRegInTop_6_59[30] , \wRegInTop_6_59[29] , \wRegInTop_6_59[28] , 
        \wRegInTop_6_59[27] , \wRegInTop_6_59[26] , \wRegInTop_6_59[25] , 
        \wRegInTop_6_59[24] , \wRegInTop_6_59[23] , \wRegInTop_6_59[22] , 
        \wRegInTop_6_59[21] , \wRegInTop_6_59[20] , \wRegInTop_6_59[19] , 
        \wRegInTop_6_59[18] , \wRegInTop_6_59[17] , \wRegInTop_6_59[16] , 
        \wRegInTop_6_59[15] , \wRegInTop_6_59[14] , \wRegInTop_6_59[13] , 
        \wRegInTop_6_59[12] , \wRegInTop_6_59[11] , \wRegInTop_6_59[10] , 
        \wRegInTop_6_59[9] , \wRegInTop_6_59[8] , \wRegInTop_6_59[7] , 
        \wRegInTop_6_59[6] , \wRegInTop_6_59[5] , \wRegInTop_6_59[4] , 
        \wRegInTop_6_59[3] , \wRegInTop_6_59[2] , \wRegInTop_6_59[1] , 
        \wRegInTop_6_59[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_17 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink145[31] , \ScanLink145[30] , \ScanLink145[29] , 
        \ScanLink145[28] , \ScanLink145[27] , \ScanLink145[26] , 
        \ScanLink145[25] , \ScanLink145[24] , \ScanLink145[23] , 
        \ScanLink145[22] , \ScanLink145[21] , \ScanLink145[20] , 
        \ScanLink145[19] , \ScanLink145[18] , \ScanLink145[17] , 
        \ScanLink145[16] , \ScanLink145[15] , \ScanLink145[14] , 
        \ScanLink145[13] , \ScanLink145[12] , \ScanLink145[11] , 
        \ScanLink145[10] , \ScanLink145[9] , \ScanLink145[8] , 
        \ScanLink145[7] , \ScanLink145[6] , \ScanLink145[5] , \ScanLink145[4] , 
        \ScanLink145[3] , \ScanLink145[2] , \ScanLink145[1] , \ScanLink145[0] 
        }), .ScanOut({\ScanLink144[31] , \ScanLink144[30] , \ScanLink144[29] , 
        \ScanLink144[28] , \ScanLink144[27] , \ScanLink144[26] , 
        \ScanLink144[25] , \ScanLink144[24] , \ScanLink144[23] , 
        \ScanLink144[22] , \ScanLink144[21] , \ScanLink144[20] , 
        \ScanLink144[19] , \ScanLink144[18] , \ScanLink144[17] , 
        \ScanLink144[16] , \ScanLink144[15] , \ScanLink144[14] , 
        \ScanLink144[13] , \ScanLink144[12] , \ScanLink144[11] , 
        \ScanLink144[10] , \ScanLink144[9] , \ScanLink144[8] , 
        \ScanLink144[7] , \ScanLink144[6] , \ScanLink144[5] , \ScanLink144[4] , 
        \ScanLink144[3] , \ScanLink144[2] , \ScanLink144[1] , \ScanLink144[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_17[31] , 
        \wRegOut_7_17[30] , \wRegOut_7_17[29] , \wRegOut_7_17[28] , 
        \wRegOut_7_17[27] , \wRegOut_7_17[26] , \wRegOut_7_17[25] , 
        \wRegOut_7_17[24] , \wRegOut_7_17[23] , \wRegOut_7_17[22] , 
        \wRegOut_7_17[21] , \wRegOut_7_17[20] , \wRegOut_7_17[19] , 
        \wRegOut_7_17[18] , \wRegOut_7_17[17] , \wRegOut_7_17[16] , 
        \wRegOut_7_17[15] , \wRegOut_7_17[14] , \wRegOut_7_17[13] , 
        \wRegOut_7_17[12] , \wRegOut_7_17[11] , \wRegOut_7_17[10] , 
        \wRegOut_7_17[9] , \wRegOut_7_17[8] , \wRegOut_7_17[7] , 
        \wRegOut_7_17[6] , \wRegOut_7_17[5] , \wRegOut_7_17[4] , 
        \wRegOut_7_17[3] , \wRegOut_7_17[2] , \wRegOut_7_17[1] , 
        \wRegOut_7_17[0] }), .Enable1(\wRegEnTop_7_17[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_17[31] , \wRegInTop_7_17[30] , \wRegInTop_7_17[29] , 
        \wRegInTop_7_17[28] , \wRegInTop_7_17[27] , \wRegInTop_7_17[26] , 
        \wRegInTop_7_17[25] , \wRegInTop_7_17[24] , \wRegInTop_7_17[23] , 
        \wRegInTop_7_17[22] , \wRegInTop_7_17[21] , \wRegInTop_7_17[20] , 
        \wRegInTop_7_17[19] , \wRegInTop_7_17[18] , \wRegInTop_7_17[17] , 
        \wRegInTop_7_17[16] , \wRegInTop_7_17[15] , \wRegInTop_7_17[14] , 
        \wRegInTop_7_17[13] , \wRegInTop_7_17[12] , \wRegInTop_7_17[11] , 
        \wRegInTop_7_17[10] , \wRegInTop_7_17[9] , \wRegInTop_7_17[8] , 
        \wRegInTop_7_17[7] , \wRegInTop_7_17[6] , \wRegInTop_7_17[5] , 
        \wRegInTop_7_17[4] , \wRegInTop_7_17[3] , \wRegInTop_7_17[2] , 
        \wRegInTop_7_17[1] , \wRegInTop_7_17[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_87 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink215[31] , \ScanLink215[30] , \ScanLink215[29] , 
        \ScanLink215[28] , \ScanLink215[27] , \ScanLink215[26] , 
        \ScanLink215[25] , \ScanLink215[24] , \ScanLink215[23] , 
        \ScanLink215[22] , \ScanLink215[21] , \ScanLink215[20] , 
        \ScanLink215[19] , \ScanLink215[18] , \ScanLink215[17] , 
        \ScanLink215[16] , \ScanLink215[15] , \ScanLink215[14] , 
        \ScanLink215[13] , \ScanLink215[12] , \ScanLink215[11] , 
        \ScanLink215[10] , \ScanLink215[9] , \ScanLink215[8] , 
        \ScanLink215[7] , \ScanLink215[6] , \ScanLink215[5] , \ScanLink215[4] , 
        \ScanLink215[3] , \ScanLink215[2] , \ScanLink215[1] , \ScanLink215[0] 
        }), .ScanOut({\ScanLink214[31] , \ScanLink214[30] , \ScanLink214[29] , 
        \ScanLink214[28] , \ScanLink214[27] , \ScanLink214[26] , 
        \ScanLink214[25] , \ScanLink214[24] , \ScanLink214[23] , 
        \ScanLink214[22] , \ScanLink214[21] , \ScanLink214[20] , 
        \ScanLink214[19] , \ScanLink214[18] , \ScanLink214[17] , 
        \ScanLink214[16] , \ScanLink214[15] , \ScanLink214[14] , 
        \ScanLink214[13] , \ScanLink214[12] , \ScanLink214[11] , 
        \ScanLink214[10] , \ScanLink214[9] , \ScanLink214[8] , 
        \ScanLink214[7] , \ScanLink214[6] , \ScanLink214[5] , \ScanLink214[4] , 
        \ScanLink214[3] , \ScanLink214[2] , \ScanLink214[1] , \ScanLink214[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_87[31] , 
        \wRegOut_7_87[30] , \wRegOut_7_87[29] , \wRegOut_7_87[28] , 
        \wRegOut_7_87[27] , \wRegOut_7_87[26] , \wRegOut_7_87[25] , 
        \wRegOut_7_87[24] , \wRegOut_7_87[23] , \wRegOut_7_87[22] , 
        \wRegOut_7_87[21] , \wRegOut_7_87[20] , \wRegOut_7_87[19] , 
        \wRegOut_7_87[18] , \wRegOut_7_87[17] , \wRegOut_7_87[16] , 
        \wRegOut_7_87[15] , \wRegOut_7_87[14] , \wRegOut_7_87[13] , 
        \wRegOut_7_87[12] , \wRegOut_7_87[11] , \wRegOut_7_87[10] , 
        \wRegOut_7_87[9] , \wRegOut_7_87[8] , \wRegOut_7_87[7] , 
        \wRegOut_7_87[6] , \wRegOut_7_87[5] , \wRegOut_7_87[4] , 
        \wRegOut_7_87[3] , \wRegOut_7_87[2] , \wRegOut_7_87[1] , 
        \wRegOut_7_87[0] }), .Enable1(\wRegEnTop_7_87[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_87[31] , \wRegInTop_7_87[30] , \wRegInTop_7_87[29] , 
        \wRegInTop_7_87[28] , \wRegInTop_7_87[27] , \wRegInTop_7_87[26] , 
        \wRegInTop_7_87[25] , \wRegInTop_7_87[24] , \wRegInTop_7_87[23] , 
        \wRegInTop_7_87[22] , \wRegInTop_7_87[21] , \wRegInTop_7_87[20] , 
        \wRegInTop_7_87[19] , \wRegInTop_7_87[18] , \wRegInTop_7_87[17] , 
        \wRegInTop_7_87[16] , \wRegInTop_7_87[15] , \wRegInTop_7_87[14] , 
        \wRegInTop_7_87[13] , \wRegInTop_7_87[12] , \wRegInTop_7_87[11] , 
        \wRegInTop_7_87[10] , \wRegInTop_7_87[9] , \wRegInTop_7_87[8] , 
        \wRegInTop_7_87[7] , \wRegInTop_7_87[6] , \wRegInTop_7_87[5] , 
        \wRegInTop_7_87[4] , \wRegInTop_7_87[3] , \wRegInTop_7_87[2] , 
        \wRegInTop_7_87[1] , \wRegInTop_7_87[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_1[0] ), .P_In({\wRegOut_6_1[31] , 
        \wRegOut_6_1[30] , \wRegOut_6_1[29] , \wRegOut_6_1[28] , 
        \wRegOut_6_1[27] , \wRegOut_6_1[26] , \wRegOut_6_1[25] , 
        \wRegOut_6_1[24] , \wRegOut_6_1[23] , \wRegOut_6_1[22] , 
        \wRegOut_6_1[21] , \wRegOut_6_1[20] , \wRegOut_6_1[19] , 
        \wRegOut_6_1[18] , \wRegOut_6_1[17] , \wRegOut_6_1[16] , 
        \wRegOut_6_1[15] , \wRegOut_6_1[14] , \wRegOut_6_1[13] , 
        \wRegOut_6_1[12] , \wRegOut_6_1[11] , \wRegOut_6_1[10] , 
        \wRegOut_6_1[9] , \wRegOut_6_1[8] , \wRegOut_6_1[7] , \wRegOut_6_1[6] , 
        \wRegOut_6_1[5] , \wRegOut_6_1[4] , \wRegOut_6_1[3] , \wRegOut_6_1[2] , 
        \wRegOut_6_1[1] , \wRegOut_6_1[0] }), .P_Out({\wRegInBot_6_1[31] , 
        \wRegInBot_6_1[30] , \wRegInBot_6_1[29] , \wRegInBot_6_1[28] , 
        \wRegInBot_6_1[27] , \wRegInBot_6_1[26] , \wRegInBot_6_1[25] , 
        \wRegInBot_6_1[24] , \wRegInBot_6_1[23] , \wRegInBot_6_1[22] , 
        \wRegInBot_6_1[21] , \wRegInBot_6_1[20] , \wRegInBot_6_1[19] , 
        \wRegInBot_6_1[18] , \wRegInBot_6_1[17] , \wRegInBot_6_1[16] , 
        \wRegInBot_6_1[15] , \wRegInBot_6_1[14] , \wRegInBot_6_1[13] , 
        \wRegInBot_6_1[12] , \wRegInBot_6_1[11] , \wRegInBot_6_1[10] , 
        \wRegInBot_6_1[9] , \wRegInBot_6_1[8] , \wRegInBot_6_1[7] , 
        \wRegInBot_6_1[6] , \wRegInBot_6_1[5] , \wRegInBot_6_1[4] , 
        \wRegInBot_6_1[3] , \wRegInBot_6_1[2] , \wRegInBot_6_1[1] , 
        \wRegInBot_6_1[0] }), .L_WR(\wRegEnTop_7_2[0] ), .L_In({
        \wRegOut_7_2[31] , \wRegOut_7_2[30] , \wRegOut_7_2[29] , 
        \wRegOut_7_2[28] , \wRegOut_7_2[27] , \wRegOut_7_2[26] , 
        \wRegOut_7_2[25] , \wRegOut_7_2[24] , \wRegOut_7_2[23] , 
        \wRegOut_7_2[22] , \wRegOut_7_2[21] , \wRegOut_7_2[20] , 
        \wRegOut_7_2[19] , \wRegOut_7_2[18] , \wRegOut_7_2[17] , 
        \wRegOut_7_2[16] , \wRegOut_7_2[15] , \wRegOut_7_2[14] , 
        \wRegOut_7_2[13] , \wRegOut_7_2[12] , \wRegOut_7_2[11] , 
        \wRegOut_7_2[10] , \wRegOut_7_2[9] , \wRegOut_7_2[8] , 
        \wRegOut_7_2[7] , \wRegOut_7_2[6] , \wRegOut_7_2[5] , \wRegOut_7_2[4] , 
        \wRegOut_7_2[3] , \wRegOut_7_2[2] , \wRegOut_7_2[1] , \wRegOut_7_2[0] 
        }), .L_Out({\wRegInTop_7_2[31] , \wRegInTop_7_2[30] , 
        \wRegInTop_7_2[29] , \wRegInTop_7_2[28] , \wRegInTop_7_2[27] , 
        \wRegInTop_7_2[26] , \wRegInTop_7_2[25] , \wRegInTop_7_2[24] , 
        \wRegInTop_7_2[23] , \wRegInTop_7_2[22] , \wRegInTop_7_2[21] , 
        \wRegInTop_7_2[20] , \wRegInTop_7_2[19] , \wRegInTop_7_2[18] , 
        \wRegInTop_7_2[17] , \wRegInTop_7_2[16] , \wRegInTop_7_2[15] , 
        \wRegInTop_7_2[14] , \wRegInTop_7_2[13] , \wRegInTop_7_2[12] , 
        \wRegInTop_7_2[11] , \wRegInTop_7_2[10] , \wRegInTop_7_2[9] , 
        \wRegInTop_7_2[8] , \wRegInTop_7_2[7] , \wRegInTop_7_2[6] , 
        \wRegInTop_7_2[5] , \wRegInTop_7_2[4] , \wRegInTop_7_2[3] , 
        \wRegInTop_7_2[2] , \wRegInTop_7_2[1] , \wRegInTop_7_2[0] }), .R_WR(
        \wRegEnTop_7_3[0] ), .R_In({\wRegOut_7_3[31] , \wRegOut_7_3[30] , 
        \wRegOut_7_3[29] , \wRegOut_7_3[28] , \wRegOut_7_3[27] , 
        \wRegOut_7_3[26] , \wRegOut_7_3[25] , \wRegOut_7_3[24] , 
        \wRegOut_7_3[23] , \wRegOut_7_3[22] , \wRegOut_7_3[21] , 
        \wRegOut_7_3[20] , \wRegOut_7_3[19] , \wRegOut_7_3[18] , 
        \wRegOut_7_3[17] , \wRegOut_7_3[16] , \wRegOut_7_3[15] , 
        \wRegOut_7_3[14] , \wRegOut_7_3[13] , \wRegOut_7_3[12] , 
        \wRegOut_7_3[11] , \wRegOut_7_3[10] , \wRegOut_7_3[9] , 
        \wRegOut_7_3[8] , \wRegOut_7_3[7] , \wRegOut_7_3[6] , \wRegOut_7_3[5] , 
        \wRegOut_7_3[4] , \wRegOut_7_3[3] , \wRegOut_7_3[2] , \wRegOut_7_3[1] , 
        \wRegOut_7_3[0] }), .R_Out({\wRegInTop_7_3[31] , \wRegInTop_7_3[30] , 
        \wRegInTop_7_3[29] , \wRegInTop_7_3[28] , \wRegInTop_7_3[27] , 
        \wRegInTop_7_3[26] , \wRegInTop_7_3[25] , \wRegInTop_7_3[24] , 
        \wRegInTop_7_3[23] , \wRegInTop_7_3[22] , \wRegInTop_7_3[21] , 
        \wRegInTop_7_3[20] , \wRegInTop_7_3[19] , \wRegInTop_7_3[18] , 
        \wRegInTop_7_3[17] , \wRegInTop_7_3[16] , \wRegInTop_7_3[15] , 
        \wRegInTop_7_3[14] , \wRegInTop_7_3[13] , \wRegInTop_7_3[12] , 
        \wRegInTop_7_3[11] , \wRegInTop_7_3[10] , \wRegInTop_7_3[9] , 
        \wRegInTop_7_3[8] , \wRegInTop_7_3[7] , \wRegInTop_7_3[6] , 
        \wRegInTop_7_3[5] , \wRegInTop_7_3[4] , \wRegInTop_7_3[3] , 
        \wRegInTop_7_3[2] , \wRegInTop_7_3[1] , \wRegInTop_7_3[0] }) );
    BHeap_Node_WIDTH32 BHN_6_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_19[0] ), .P_In({\wRegOut_6_19[31] , 
        \wRegOut_6_19[30] , \wRegOut_6_19[29] , \wRegOut_6_19[28] , 
        \wRegOut_6_19[27] , \wRegOut_6_19[26] , \wRegOut_6_19[25] , 
        \wRegOut_6_19[24] , \wRegOut_6_19[23] , \wRegOut_6_19[22] , 
        \wRegOut_6_19[21] , \wRegOut_6_19[20] , \wRegOut_6_19[19] , 
        \wRegOut_6_19[18] , \wRegOut_6_19[17] , \wRegOut_6_19[16] , 
        \wRegOut_6_19[15] , \wRegOut_6_19[14] , \wRegOut_6_19[13] , 
        \wRegOut_6_19[12] , \wRegOut_6_19[11] , \wRegOut_6_19[10] , 
        \wRegOut_6_19[9] , \wRegOut_6_19[8] , \wRegOut_6_19[7] , 
        \wRegOut_6_19[6] , \wRegOut_6_19[5] , \wRegOut_6_19[4] , 
        \wRegOut_6_19[3] , \wRegOut_6_19[2] , \wRegOut_6_19[1] , 
        \wRegOut_6_19[0] }), .P_Out({\wRegInBot_6_19[31] , 
        \wRegInBot_6_19[30] , \wRegInBot_6_19[29] , \wRegInBot_6_19[28] , 
        \wRegInBot_6_19[27] , \wRegInBot_6_19[26] , \wRegInBot_6_19[25] , 
        \wRegInBot_6_19[24] , \wRegInBot_6_19[23] , \wRegInBot_6_19[22] , 
        \wRegInBot_6_19[21] , \wRegInBot_6_19[20] , \wRegInBot_6_19[19] , 
        \wRegInBot_6_19[18] , \wRegInBot_6_19[17] , \wRegInBot_6_19[16] , 
        \wRegInBot_6_19[15] , \wRegInBot_6_19[14] , \wRegInBot_6_19[13] , 
        \wRegInBot_6_19[12] , \wRegInBot_6_19[11] , \wRegInBot_6_19[10] , 
        \wRegInBot_6_19[9] , \wRegInBot_6_19[8] , \wRegInBot_6_19[7] , 
        \wRegInBot_6_19[6] , \wRegInBot_6_19[5] , \wRegInBot_6_19[4] , 
        \wRegInBot_6_19[3] , \wRegInBot_6_19[2] , \wRegInBot_6_19[1] , 
        \wRegInBot_6_19[0] }), .L_WR(\wRegEnTop_7_38[0] ), .L_In({
        \wRegOut_7_38[31] , \wRegOut_7_38[30] , \wRegOut_7_38[29] , 
        \wRegOut_7_38[28] , \wRegOut_7_38[27] , \wRegOut_7_38[26] , 
        \wRegOut_7_38[25] , \wRegOut_7_38[24] , \wRegOut_7_38[23] , 
        \wRegOut_7_38[22] , \wRegOut_7_38[21] , \wRegOut_7_38[20] , 
        \wRegOut_7_38[19] , \wRegOut_7_38[18] , \wRegOut_7_38[17] , 
        \wRegOut_7_38[16] , \wRegOut_7_38[15] , \wRegOut_7_38[14] , 
        \wRegOut_7_38[13] , \wRegOut_7_38[12] , \wRegOut_7_38[11] , 
        \wRegOut_7_38[10] , \wRegOut_7_38[9] , \wRegOut_7_38[8] , 
        \wRegOut_7_38[7] , \wRegOut_7_38[6] , \wRegOut_7_38[5] , 
        \wRegOut_7_38[4] , \wRegOut_7_38[3] , \wRegOut_7_38[2] , 
        \wRegOut_7_38[1] , \wRegOut_7_38[0] }), .L_Out({\wRegInTop_7_38[31] , 
        \wRegInTop_7_38[30] , \wRegInTop_7_38[29] , \wRegInTop_7_38[28] , 
        \wRegInTop_7_38[27] , \wRegInTop_7_38[26] , \wRegInTop_7_38[25] , 
        \wRegInTop_7_38[24] , \wRegInTop_7_38[23] , \wRegInTop_7_38[22] , 
        \wRegInTop_7_38[21] , \wRegInTop_7_38[20] , \wRegInTop_7_38[19] , 
        \wRegInTop_7_38[18] , \wRegInTop_7_38[17] , \wRegInTop_7_38[16] , 
        \wRegInTop_7_38[15] , \wRegInTop_7_38[14] , \wRegInTop_7_38[13] , 
        \wRegInTop_7_38[12] , \wRegInTop_7_38[11] , \wRegInTop_7_38[10] , 
        \wRegInTop_7_38[9] , \wRegInTop_7_38[8] , \wRegInTop_7_38[7] , 
        \wRegInTop_7_38[6] , \wRegInTop_7_38[5] , \wRegInTop_7_38[4] , 
        \wRegInTop_7_38[3] , \wRegInTop_7_38[2] , \wRegInTop_7_38[1] , 
        \wRegInTop_7_38[0] }), .R_WR(\wRegEnTop_7_39[0] ), .R_In({
        \wRegOut_7_39[31] , \wRegOut_7_39[30] , \wRegOut_7_39[29] , 
        \wRegOut_7_39[28] , \wRegOut_7_39[27] , \wRegOut_7_39[26] , 
        \wRegOut_7_39[25] , \wRegOut_7_39[24] , \wRegOut_7_39[23] , 
        \wRegOut_7_39[22] , \wRegOut_7_39[21] , \wRegOut_7_39[20] , 
        \wRegOut_7_39[19] , \wRegOut_7_39[18] , \wRegOut_7_39[17] , 
        \wRegOut_7_39[16] , \wRegOut_7_39[15] , \wRegOut_7_39[14] , 
        \wRegOut_7_39[13] , \wRegOut_7_39[12] , \wRegOut_7_39[11] , 
        \wRegOut_7_39[10] , \wRegOut_7_39[9] , \wRegOut_7_39[8] , 
        \wRegOut_7_39[7] , \wRegOut_7_39[6] , \wRegOut_7_39[5] , 
        \wRegOut_7_39[4] , \wRegOut_7_39[3] , \wRegOut_7_39[2] , 
        \wRegOut_7_39[1] , \wRegOut_7_39[0] }), .R_Out({\wRegInTop_7_39[31] , 
        \wRegInTop_7_39[30] , \wRegInTop_7_39[29] , \wRegInTop_7_39[28] , 
        \wRegInTop_7_39[27] , \wRegInTop_7_39[26] , \wRegInTop_7_39[25] , 
        \wRegInTop_7_39[24] , \wRegInTop_7_39[23] , \wRegInTop_7_39[22] , 
        \wRegInTop_7_39[21] , \wRegInTop_7_39[20] , \wRegInTop_7_39[19] , 
        \wRegInTop_7_39[18] , \wRegInTop_7_39[17] , \wRegInTop_7_39[16] , 
        \wRegInTop_7_39[15] , \wRegInTop_7_39[14] , \wRegInTop_7_39[13] , 
        \wRegInTop_7_39[12] , \wRegInTop_7_39[11] , \wRegInTop_7_39[10] , 
        \wRegInTop_7_39[9] , \wRegInTop_7_39[8] , \wRegInTop_7_39[7] , 
        \wRegInTop_7_39[6] , \wRegInTop_7_39[5] , \wRegInTop_7_39[4] , 
        \wRegInTop_7_39[3] , \wRegInTop_7_39[2] , \wRegInTop_7_39[1] , 
        \wRegInTop_7_39[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_118 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink246[31] , \ScanLink246[30] , \ScanLink246[29] , 
        \ScanLink246[28] , \ScanLink246[27] , \ScanLink246[26] , 
        \ScanLink246[25] , \ScanLink246[24] , \ScanLink246[23] , 
        \ScanLink246[22] , \ScanLink246[21] , \ScanLink246[20] , 
        \ScanLink246[19] , \ScanLink246[18] , \ScanLink246[17] , 
        \ScanLink246[16] , \ScanLink246[15] , \ScanLink246[14] , 
        \ScanLink246[13] , \ScanLink246[12] , \ScanLink246[11] , 
        \ScanLink246[10] , \ScanLink246[9] , \ScanLink246[8] , 
        \ScanLink246[7] , \ScanLink246[6] , \ScanLink246[5] , \ScanLink246[4] , 
        \ScanLink246[3] , \ScanLink246[2] , \ScanLink246[1] , \ScanLink246[0] 
        }), .ScanOut({\ScanLink245[31] , \ScanLink245[30] , \ScanLink245[29] , 
        \ScanLink245[28] , \ScanLink245[27] , \ScanLink245[26] , 
        \ScanLink245[25] , \ScanLink245[24] , \ScanLink245[23] , 
        \ScanLink245[22] , \ScanLink245[21] , \ScanLink245[20] , 
        \ScanLink245[19] , \ScanLink245[18] , \ScanLink245[17] , 
        \ScanLink245[16] , \ScanLink245[15] , \ScanLink245[14] , 
        \ScanLink245[13] , \ScanLink245[12] , \ScanLink245[11] , 
        \ScanLink245[10] , \ScanLink245[9] , \ScanLink245[8] , 
        \ScanLink245[7] , \ScanLink245[6] , \ScanLink245[5] , \ScanLink245[4] , 
        \ScanLink245[3] , \ScanLink245[2] , \ScanLink245[1] , \ScanLink245[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_118[31] , 
        \wRegOut_7_118[30] , \wRegOut_7_118[29] , \wRegOut_7_118[28] , 
        \wRegOut_7_118[27] , \wRegOut_7_118[26] , \wRegOut_7_118[25] , 
        \wRegOut_7_118[24] , \wRegOut_7_118[23] , \wRegOut_7_118[22] , 
        \wRegOut_7_118[21] , \wRegOut_7_118[20] , \wRegOut_7_118[19] , 
        \wRegOut_7_118[18] , \wRegOut_7_118[17] , \wRegOut_7_118[16] , 
        \wRegOut_7_118[15] , \wRegOut_7_118[14] , \wRegOut_7_118[13] , 
        \wRegOut_7_118[12] , \wRegOut_7_118[11] , \wRegOut_7_118[10] , 
        \wRegOut_7_118[9] , \wRegOut_7_118[8] , \wRegOut_7_118[7] , 
        \wRegOut_7_118[6] , \wRegOut_7_118[5] , \wRegOut_7_118[4] , 
        \wRegOut_7_118[3] , \wRegOut_7_118[2] , \wRegOut_7_118[1] , 
        \wRegOut_7_118[0] }), .Enable1(\wRegEnTop_7_118[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_118[31] , \wRegInTop_7_118[30] , 
        \wRegInTop_7_118[29] , \wRegInTop_7_118[28] , \wRegInTop_7_118[27] , 
        \wRegInTop_7_118[26] , \wRegInTop_7_118[25] , \wRegInTop_7_118[24] , 
        \wRegInTop_7_118[23] , \wRegInTop_7_118[22] , \wRegInTop_7_118[21] , 
        \wRegInTop_7_118[20] , \wRegInTop_7_118[19] , \wRegInTop_7_118[18] , 
        \wRegInTop_7_118[17] , \wRegInTop_7_118[16] , \wRegInTop_7_118[15] , 
        \wRegInTop_7_118[14] , \wRegInTop_7_118[13] , \wRegInTop_7_118[12] , 
        \wRegInTop_7_118[11] , \wRegInTop_7_118[10] , \wRegInTop_7_118[9] , 
        \wRegInTop_7_118[8] , \wRegInTop_7_118[7] , \wRegInTop_7_118[6] , 
        \wRegInTop_7_118[5] , \wRegInTop_7_118[4] , \wRegInTop_7_118[3] , 
        \wRegInTop_7_118[2] , \wRegInTop_7_118[1] , \wRegInTop_7_118[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_7[0] ), .P_In({\wRegOut_3_7[31] , 
        \wRegOut_3_7[30] , \wRegOut_3_7[29] , \wRegOut_3_7[28] , 
        \wRegOut_3_7[27] , \wRegOut_3_7[26] , \wRegOut_3_7[25] , 
        \wRegOut_3_7[24] , \wRegOut_3_7[23] , \wRegOut_3_7[22] , 
        \wRegOut_3_7[21] , \wRegOut_3_7[20] , \wRegOut_3_7[19] , 
        \wRegOut_3_7[18] , \wRegOut_3_7[17] , \wRegOut_3_7[16] , 
        \wRegOut_3_7[15] , \wRegOut_3_7[14] , \wRegOut_3_7[13] , 
        \wRegOut_3_7[12] , \wRegOut_3_7[11] , \wRegOut_3_7[10] , 
        \wRegOut_3_7[9] , \wRegOut_3_7[8] , \wRegOut_3_7[7] , \wRegOut_3_7[6] , 
        \wRegOut_3_7[5] , \wRegOut_3_7[4] , \wRegOut_3_7[3] , \wRegOut_3_7[2] , 
        \wRegOut_3_7[1] , \wRegOut_3_7[0] }), .P_Out({\wRegInBot_3_7[31] , 
        \wRegInBot_3_7[30] , \wRegInBot_3_7[29] , \wRegInBot_3_7[28] , 
        \wRegInBot_3_7[27] , \wRegInBot_3_7[26] , \wRegInBot_3_7[25] , 
        \wRegInBot_3_7[24] , \wRegInBot_3_7[23] , \wRegInBot_3_7[22] , 
        \wRegInBot_3_7[21] , \wRegInBot_3_7[20] , \wRegInBot_3_7[19] , 
        \wRegInBot_3_7[18] , \wRegInBot_3_7[17] , \wRegInBot_3_7[16] , 
        \wRegInBot_3_7[15] , \wRegInBot_3_7[14] , \wRegInBot_3_7[13] , 
        \wRegInBot_3_7[12] , \wRegInBot_3_7[11] , \wRegInBot_3_7[10] , 
        \wRegInBot_3_7[9] , \wRegInBot_3_7[8] , \wRegInBot_3_7[7] , 
        \wRegInBot_3_7[6] , \wRegInBot_3_7[5] , \wRegInBot_3_7[4] , 
        \wRegInBot_3_7[3] , \wRegInBot_3_7[2] , \wRegInBot_3_7[1] , 
        \wRegInBot_3_7[0] }), .L_WR(\wRegEnTop_4_14[0] ), .L_In({
        \wRegOut_4_14[31] , \wRegOut_4_14[30] , \wRegOut_4_14[29] , 
        \wRegOut_4_14[28] , \wRegOut_4_14[27] , \wRegOut_4_14[26] , 
        \wRegOut_4_14[25] , \wRegOut_4_14[24] , \wRegOut_4_14[23] , 
        \wRegOut_4_14[22] , \wRegOut_4_14[21] , \wRegOut_4_14[20] , 
        \wRegOut_4_14[19] , \wRegOut_4_14[18] , \wRegOut_4_14[17] , 
        \wRegOut_4_14[16] , \wRegOut_4_14[15] , \wRegOut_4_14[14] , 
        \wRegOut_4_14[13] , \wRegOut_4_14[12] , \wRegOut_4_14[11] , 
        \wRegOut_4_14[10] , \wRegOut_4_14[9] , \wRegOut_4_14[8] , 
        \wRegOut_4_14[7] , \wRegOut_4_14[6] , \wRegOut_4_14[5] , 
        \wRegOut_4_14[4] , \wRegOut_4_14[3] , \wRegOut_4_14[2] , 
        \wRegOut_4_14[1] , \wRegOut_4_14[0] }), .L_Out({\wRegInTop_4_14[31] , 
        \wRegInTop_4_14[30] , \wRegInTop_4_14[29] , \wRegInTop_4_14[28] , 
        \wRegInTop_4_14[27] , \wRegInTop_4_14[26] , \wRegInTop_4_14[25] , 
        \wRegInTop_4_14[24] , \wRegInTop_4_14[23] , \wRegInTop_4_14[22] , 
        \wRegInTop_4_14[21] , \wRegInTop_4_14[20] , \wRegInTop_4_14[19] , 
        \wRegInTop_4_14[18] , \wRegInTop_4_14[17] , \wRegInTop_4_14[16] , 
        \wRegInTop_4_14[15] , \wRegInTop_4_14[14] , \wRegInTop_4_14[13] , 
        \wRegInTop_4_14[12] , \wRegInTop_4_14[11] , \wRegInTop_4_14[10] , 
        \wRegInTop_4_14[9] , \wRegInTop_4_14[8] , \wRegInTop_4_14[7] , 
        \wRegInTop_4_14[6] , \wRegInTop_4_14[5] , \wRegInTop_4_14[4] , 
        \wRegInTop_4_14[3] , \wRegInTop_4_14[2] , \wRegInTop_4_14[1] , 
        \wRegInTop_4_14[0] }), .R_WR(\wRegEnTop_4_15[0] ), .R_In({
        \wRegOut_4_15[31] , \wRegOut_4_15[30] , \wRegOut_4_15[29] , 
        \wRegOut_4_15[28] , \wRegOut_4_15[27] , \wRegOut_4_15[26] , 
        \wRegOut_4_15[25] , \wRegOut_4_15[24] , \wRegOut_4_15[23] , 
        \wRegOut_4_15[22] , \wRegOut_4_15[21] , \wRegOut_4_15[20] , 
        \wRegOut_4_15[19] , \wRegOut_4_15[18] , \wRegOut_4_15[17] , 
        \wRegOut_4_15[16] , \wRegOut_4_15[15] , \wRegOut_4_15[14] , 
        \wRegOut_4_15[13] , \wRegOut_4_15[12] , \wRegOut_4_15[11] , 
        \wRegOut_4_15[10] , \wRegOut_4_15[9] , \wRegOut_4_15[8] , 
        \wRegOut_4_15[7] , \wRegOut_4_15[6] , \wRegOut_4_15[5] , 
        \wRegOut_4_15[4] , \wRegOut_4_15[3] , \wRegOut_4_15[2] , 
        \wRegOut_4_15[1] , \wRegOut_4_15[0] }), .R_Out({\wRegInTop_4_15[31] , 
        \wRegInTop_4_15[30] , \wRegInTop_4_15[29] , \wRegInTop_4_15[28] , 
        \wRegInTop_4_15[27] , \wRegInTop_4_15[26] , \wRegInTop_4_15[25] , 
        \wRegInTop_4_15[24] , \wRegInTop_4_15[23] , \wRegInTop_4_15[22] , 
        \wRegInTop_4_15[21] , \wRegInTop_4_15[20] , \wRegInTop_4_15[19] , 
        \wRegInTop_4_15[18] , \wRegInTop_4_15[17] , \wRegInTop_4_15[16] , 
        \wRegInTop_4_15[15] , \wRegInTop_4_15[14] , \wRegInTop_4_15[13] , 
        \wRegInTop_4_15[12] , \wRegInTop_4_15[11] , \wRegInTop_4_15[10] , 
        \wRegInTop_4_15[9] , \wRegInTop_4_15[8] , \wRegInTop_4_15[7] , 
        \wRegInTop_4_15[6] , \wRegInTop_4_15[5] , \wRegInTop_4_15[4] , 
        \wRegInTop_4_15[3] , \wRegInTop_4_15[2] , \wRegInTop_4_15[1] , 
        \wRegInTop_4_15[0] }) );
    BHeap_Node_WIDTH32 BHN_4_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_14[0] ), .P_In({\wRegOut_4_14[31] , 
        \wRegOut_4_14[30] , \wRegOut_4_14[29] , \wRegOut_4_14[28] , 
        \wRegOut_4_14[27] , \wRegOut_4_14[26] , \wRegOut_4_14[25] , 
        \wRegOut_4_14[24] , \wRegOut_4_14[23] , \wRegOut_4_14[22] , 
        \wRegOut_4_14[21] , \wRegOut_4_14[20] , \wRegOut_4_14[19] , 
        \wRegOut_4_14[18] , \wRegOut_4_14[17] , \wRegOut_4_14[16] , 
        \wRegOut_4_14[15] , \wRegOut_4_14[14] , \wRegOut_4_14[13] , 
        \wRegOut_4_14[12] , \wRegOut_4_14[11] , \wRegOut_4_14[10] , 
        \wRegOut_4_14[9] , \wRegOut_4_14[8] , \wRegOut_4_14[7] , 
        \wRegOut_4_14[6] , \wRegOut_4_14[5] , \wRegOut_4_14[4] , 
        \wRegOut_4_14[3] , \wRegOut_4_14[2] , \wRegOut_4_14[1] , 
        \wRegOut_4_14[0] }), .P_Out({\wRegInBot_4_14[31] , 
        \wRegInBot_4_14[30] , \wRegInBot_4_14[29] , \wRegInBot_4_14[28] , 
        \wRegInBot_4_14[27] , \wRegInBot_4_14[26] , \wRegInBot_4_14[25] , 
        \wRegInBot_4_14[24] , \wRegInBot_4_14[23] , \wRegInBot_4_14[22] , 
        \wRegInBot_4_14[21] , \wRegInBot_4_14[20] , \wRegInBot_4_14[19] , 
        \wRegInBot_4_14[18] , \wRegInBot_4_14[17] , \wRegInBot_4_14[16] , 
        \wRegInBot_4_14[15] , \wRegInBot_4_14[14] , \wRegInBot_4_14[13] , 
        \wRegInBot_4_14[12] , \wRegInBot_4_14[11] , \wRegInBot_4_14[10] , 
        \wRegInBot_4_14[9] , \wRegInBot_4_14[8] , \wRegInBot_4_14[7] , 
        \wRegInBot_4_14[6] , \wRegInBot_4_14[5] , \wRegInBot_4_14[4] , 
        \wRegInBot_4_14[3] , \wRegInBot_4_14[2] , \wRegInBot_4_14[1] , 
        \wRegInBot_4_14[0] }), .L_WR(\wRegEnTop_5_28[0] ), .L_In({
        \wRegOut_5_28[31] , \wRegOut_5_28[30] , \wRegOut_5_28[29] , 
        \wRegOut_5_28[28] , \wRegOut_5_28[27] , \wRegOut_5_28[26] , 
        \wRegOut_5_28[25] , \wRegOut_5_28[24] , \wRegOut_5_28[23] , 
        \wRegOut_5_28[22] , \wRegOut_5_28[21] , \wRegOut_5_28[20] , 
        \wRegOut_5_28[19] , \wRegOut_5_28[18] , \wRegOut_5_28[17] , 
        \wRegOut_5_28[16] , \wRegOut_5_28[15] , \wRegOut_5_28[14] , 
        \wRegOut_5_28[13] , \wRegOut_5_28[12] , \wRegOut_5_28[11] , 
        \wRegOut_5_28[10] , \wRegOut_5_28[9] , \wRegOut_5_28[8] , 
        \wRegOut_5_28[7] , \wRegOut_5_28[6] , \wRegOut_5_28[5] , 
        \wRegOut_5_28[4] , \wRegOut_5_28[3] , \wRegOut_5_28[2] , 
        \wRegOut_5_28[1] , \wRegOut_5_28[0] }), .L_Out({\wRegInTop_5_28[31] , 
        \wRegInTop_5_28[30] , \wRegInTop_5_28[29] , \wRegInTop_5_28[28] , 
        \wRegInTop_5_28[27] , \wRegInTop_5_28[26] , \wRegInTop_5_28[25] , 
        \wRegInTop_5_28[24] , \wRegInTop_5_28[23] , \wRegInTop_5_28[22] , 
        \wRegInTop_5_28[21] , \wRegInTop_5_28[20] , \wRegInTop_5_28[19] , 
        \wRegInTop_5_28[18] , \wRegInTop_5_28[17] , \wRegInTop_5_28[16] , 
        \wRegInTop_5_28[15] , \wRegInTop_5_28[14] , \wRegInTop_5_28[13] , 
        \wRegInTop_5_28[12] , \wRegInTop_5_28[11] , \wRegInTop_5_28[10] , 
        \wRegInTop_5_28[9] , \wRegInTop_5_28[8] , \wRegInTop_5_28[7] , 
        \wRegInTop_5_28[6] , \wRegInTop_5_28[5] , \wRegInTop_5_28[4] , 
        \wRegInTop_5_28[3] , \wRegInTop_5_28[2] , \wRegInTop_5_28[1] , 
        \wRegInTop_5_28[0] }), .R_WR(\wRegEnTop_5_29[0] ), .R_In({
        \wRegOut_5_29[31] , \wRegOut_5_29[30] , \wRegOut_5_29[29] , 
        \wRegOut_5_29[28] , \wRegOut_5_29[27] , \wRegOut_5_29[26] , 
        \wRegOut_5_29[25] , \wRegOut_5_29[24] , \wRegOut_5_29[23] , 
        \wRegOut_5_29[22] , \wRegOut_5_29[21] , \wRegOut_5_29[20] , 
        \wRegOut_5_29[19] , \wRegOut_5_29[18] , \wRegOut_5_29[17] , 
        \wRegOut_5_29[16] , \wRegOut_5_29[15] , \wRegOut_5_29[14] , 
        \wRegOut_5_29[13] , \wRegOut_5_29[12] , \wRegOut_5_29[11] , 
        \wRegOut_5_29[10] , \wRegOut_5_29[9] , \wRegOut_5_29[8] , 
        \wRegOut_5_29[7] , \wRegOut_5_29[6] , \wRegOut_5_29[5] , 
        \wRegOut_5_29[4] , \wRegOut_5_29[3] , \wRegOut_5_29[2] , 
        \wRegOut_5_29[1] , \wRegOut_5_29[0] }), .R_Out({\wRegInTop_5_29[31] , 
        \wRegInTop_5_29[30] , \wRegInTop_5_29[29] , \wRegInTop_5_29[28] , 
        \wRegInTop_5_29[27] , \wRegInTop_5_29[26] , \wRegInTop_5_29[25] , 
        \wRegInTop_5_29[24] , \wRegInTop_5_29[23] , \wRegInTop_5_29[22] , 
        \wRegInTop_5_29[21] , \wRegInTop_5_29[20] , \wRegInTop_5_29[19] , 
        \wRegInTop_5_29[18] , \wRegInTop_5_29[17] , \wRegInTop_5_29[16] , 
        \wRegInTop_5_29[15] , \wRegInTop_5_29[14] , \wRegInTop_5_29[13] , 
        \wRegInTop_5_29[12] , \wRegInTop_5_29[11] , \wRegInTop_5_29[10] , 
        \wRegInTop_5_29[9] , \wRegInTop_5_29[8] , \wRegInTop_5_29[7] , 
        \wRegInTop_5_29[6] , \wRegInTop_5_29[5] , \wRegInTop_5_29[4] , 
        \wRegInTop_5_29[3] , \wRegInTop_5_29[2] , \wRegInTop_5_29[1] , 
        \wRegInTop_5_29[0] }) );
    BHeap_Node_WIDTH32 BHN_6_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_50[0] ), .P_In({\wRegOut_6_50[31] , 
        \wRegOut_6_50[30] , \wRegOut_6_50[29] , \wRegOut_6_50[28] , 
        \wRegOut_6_50[27] , \wRegOut_6_50[26] , \wRegOut_6_50[25] , 
        \wRegOut_6_50[24] , \wRegOut_6_50[23] , \wRegOut_6_50[22] , 
        \wRegOut_6_50[21] , \wRegOut_6_50[20] , \wRegOut_6_50[19] , 
        \wRegOut_6_50[18] , \wRegOut_6_50[17] , \wRegOut_6_50[16] , 
        \wRegOut_6_50[15] , \wRegOut_6_50[14] , \wRegOut_6_50[13] , 
        \wRegOut_6_50[12] , \wRegOut_6_50[11] , \wRegOut_6_50[10] , 
        \wRegOut_6_50[9] , \wRegOut_6_50[8] , \wRegOut_6_50[7] , 
        \wRegOut_6_50[6] , \wRegOut_6_50[5] , \wRegOut_6_50[4] , 
        \wRegOut_6_50[3] , \wRegOut_6_50[2] , \wRegOut_6_50[1] , 
        \wRegOut_6_50[0] }), .P_Out({\wRegInBot_6_50[31] , 
        \wRegInBot_6_50[30] , \wRegInBot_6_50[29] , \wRegInBot_6_50[28] , 
        \wRegInBot_6_50[27] , \wRegInBot_6_50[26] , \wRegInBot_6_50[25] , 
        \wRegInBot_6_50[24] , \wRegInBot_6_50[23] , \wRegInBot_6_50[22] , 
        \wRegInBot_6_50[21] , \wRegInBot_6_50[20] , \wRegInBot_6_50[19] , 
        \wRegInBot_6_50[18] , \wRegInBot_6_50[17] , \wRegInBot_6_50[16] , 
        \wRegInBot_6_50[15] , \wRegInBot_6_50[14] , \wRegInBot_6_50[13] , 
        \wRegInBot_6_50[12] , \wRegInBot_6_50[11] , \wRegInBot_6_50[10] , 
        \wRegInBot_6_50[9] , \wRegInBot_6_50[8] , \wRegInBot_6_50[7] , 
        \wRegInBot_6_50[6] , \wRegInBot_6_50[5] , \wRegInBot_6_50[4] , 
        \wRegInBot_6_50[3] , \wRegInBot_6_50[2] , \wRegInBot_6_50[1] , 
        \wRegInBot_6_50[0] }), .L_WR(\wRegEnTop_7_100[0] ), .L_In({
        \wRegOut_7_100[31] , \wRegOut_7_100[30] , \wRegOut_7_100[29] , 
        \wRegOut_7_100[28] , \wRegOut_7_100[27] , \wRegOut_7_100[26] , 
        \wRegOut_7_100[25] , \wRegOut_7_100[24] , \wRegOut_7_100[23] , 
        \wRegOut_7_100[22] , \wRegOut_7_100[21] , \wRegOut_7_100[20] , 
        \wRegOut_7_100[19] , \wRegOut_7_100[18] , \wRegOut_7_100[17] , 
        \wRegOut_7_100[16] , \wRegOut_7_100[15] , \wRegOut_7_100[14] , 
        \wRegOut_7_100[13] , \wRegOut_7_100[12] , \wRegOut_7_100[11] , 
        \wRegOut_7_100[10] , \wRegOut_7_100[9] , \wRegOut_7_100[8] , 
        \wRegOut_7_100[7] , \wRegOut_7_100[6] , \wRegOut_7_100[5] , 
        \wRegOut_7_100[4] , \wRegOut_7_100[3] , \wRegOut_7_100[2] , 
        \wRegOut_7_100[1] , \wRegOut_7_100[0] }), .L_Out({
        \wRegInTop_7_100[31] , \wRegInTop_7_100[30] , \wRegInTop_7_100[29] , 
        \wRegInTop_7_100[28] , \wRegInTop_7_100[27] , \wRegInTop_7_100[26] , 
        \wRegInTop_7_100[25] , \wRegInTop_7_100[24] , \wRegInTop_7_100[23] , 
        \wRegInTop_7_100[22] , \wRegInTop_7_100[21] , \wRegInTop_7_100[20] , 
        \wRegInTop_7_100[19] , \wRegInTop_7_100[18] , \wRegInTop_7_100[17] , 
        \wRegInTop_7_100[16] , \wRegInTop_7_100[15] , \wRegInTop_7_100[14] , 
        \wRegInTop_7_100[13] , \wRegInTop_7_100[12] , \wRegInTop_7_100[11] , 
        \wRegInTop_7_100[10] , \wRegInTop_7_100[9] , \wRegInTop_7_100[8] , 
        \wRegInTop_7_100[7] , \wRegInTop_7_100[6] , \wRegInTop_7_100[5] , 
        \wRegInTop_7_100[4] , \wRegInTop_7_100[3] , \wRegInTop_7_100[2] , 
        \wRegInTop_7_100[1] , \wRegInTop_7_100[0] }), .R_WR(
        \wRegEnTop_7_101[0] ), .R_In({\wRegOut_7_101[31] , \wRegOut_7_101[30] , 
        \wRegOut_7_101[29] , \wRegOut_7_101[28] , \wRegOut_7_101[27] , 
        \wRegOut_7_101[26] , \wRegOut_7_101[25] , \wRegOut_7_101[24] , 
        \wRegOut_7_101[23] , \wRegOut_7_101[22] , \wRegOut_7_101[21] , 
        \wRegOut_7_101[20] , \wRegOut_7_101[19] , \wRegOut_7_101[18] , 
        \wRegOut_7_101[17] , \wRegOut_7_101[16] , \wRegOut_7_101[15] , 
        \wRegOut_7_101[14] , \wRegOut_7_101[13] , \wRegOut_7_101[12] , 
        \wRegOut_7_101[11] , \wRegOut_7_101[10] , \wRegOut_7_101[9] , 
        \wRegOut_7_101[8] , \wRegOut_7_101[7] , \wRegOut_7_101[6] , 
        \wRegOut_7_101[5] , \wRegOut_7_101[4] , \wRegOut_7_101[3] , 
        \wRegOut_7_101[2] , \wRegOut_7_101[1] , \wRegOut_7_101[0] }), .R_Out({
        \wRegInTop_7_101[31] , \wRegInTop_7_101[30] , \wRegInTop_7_101[29] , 
        \wRegInTop_7_101[28] , \wRegInTop_7_101[27] , \wRegInTop_7_101[26] , 
        \wRegInTop_7_101[25] , \wRegInTop_7_101[24] , \wRegInTop_7_101[23] , 
        \wRegInTop_7_101[22] , \wRegInTop_7_101[21] , \wRegInTop_7_101[20] , 
        \wRegInTop_7_101[19] , \wRegInTop_7_101[18] , \wRegInTop_7_101[17] , 
        \wRegInTop_7_101[16] , \wRegInTop_7_101[15] , \wRegInTop_7_101[14] , 
        \wRegInTop_7_101[13] , \wRegInTop_7_101[12] , \wRegInTop_7_101[11] , 
        \wRegInTop_7_101[10] , \wRegInTop_7_101[9] , \wRegInTop_7_101[8] , 
        \wRegInTop_7_101[7] , \wRegInTop_7_101[6] , \wRegInTop_7_101[5] , 
        \wRegInTop_7_101[4] , \wRegInTop_7_101[3] , \wRegInTop_7_101[2] , 
        \wRegInTop_7_101[1] , \wRegInTop_7_101[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_103 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink231[31] , \ScanLink231[30] , \ScanLink231[29] , 
        \ScanLink231[28] , \ScanLink231[27] , \ScanLink231[26] , 
        \ScanLink231[25] , \ScanLink231[24] , \ScanLink231[23] , 
        \ScanLink231[22] , \ScanLink231[21] , \ScanLink231[20] , 
        \ScanLink231[19] , \ScanLink231[18] , \ScanLink231[17] , 
        \ScanLink231[16] , \ScanLink231[15] , \ScanLink231[14] , 
        \ScanLink231[13] , \ScanLink231[12] , \ScanLink231[11] , 
        \ScanLink231[10] , \ScanLink231[9] , \ScanLink231[8] , 
        \ScanLink231[7] , \ScanLink231[6] , \ScanLink231[5] , \ScanLink231[4] , 
        \ScanLink231[3] , \ScanLink231[2] , \ScanLink231[1] , \ScanLink231[0] 
        }), .ScanOut({\ScanLink230[31] , \ScanLink230[30] , \ScanLink230[29] , 
        \ScanLink230[28] , \ScanLink230[27] , \ScanLink230[26] , 
        \ScanLink230[25] , \ScanLink230[24] , \ScanLink230[23] , 
        \ScanLink230[22] , \ScanLink230[21] , \ScanLink230[20] , 
        \ScanLink230[19] , \ScanLink230[18] , \ScanLink230[17] , 
        \ScanLink230[16] , \ScanLink230[15] , \ScanLink230[14] , 
        \ScanLink230[13] , \ScanLink230[12] , \ScanLink230[11] , 
        \ScanLink230[10] , \ScanLink230[9] , \ScanLink230[8] , 
        \ScanLink230[7] , \ScanLink230[6] , \ScanLink230[5] , \ScanLink230[4] , 
        \ScanLink230[3] , \ScanLink230[2] , \ScanLink230[1] , \ScanLink230[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_103[31] , 
        \wRegOut_7_103[30] , \wRegOut_7_103[29] , \wRegOut_7_103[28] , 
        \wRegOut_7_103[27] , \wRegOut_7_103[26] , \wRegOut_7_103[25] , 
        \wRegOut_7_103[24] , \wRegOut_7_103[23] , \wRegOut_7_103[22] , 
        \wRegOut_7_103[21] , \wRegOut_7_103[20] , \wRegOut_7_103[19] , 
        \wRegOut_7_103[18] , \wRegOut_7_103[17] , \wRegOut_7_103[16] , 
        \wRegOut_7_103[15] , \wRegOut_7_103[14] , \wRegOut_7_103[13] , 
        \wRegOut_7_103[12] , \wRegOut_7_103[11] , \wRegOut_7_103[10] , 
        \wRegOut_7_103[9] , \wRegOut_7_103[8] , \wRegOut_7_103[7] , 
        \wRegOut_7_103[6] , \wRegOut_7_103[5] , \wRegOut_7_103[4] , 
        \wRegOut_7_103[3] , \wRegOut_7_103[2] , \wRegOut_7_103[1] , 
        \wRegOut_7_103[0] }), .Enable1(\wRegEnTop_7_103[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_103[31] , \wRegInTop_7_103[30] , 
        \wRegInTop_7_103[29] , \wRegInTop_7_103[28] , \wRegInTop_7_103[27] , 
        \wRegInTop_7_103[26] , \wRegInTop_7_103[25] , \wRegInTop_7_103[24] , 
        \wRegInTop_7_103[23] , \wRegInTop_7_103[22] , \wRegInTop_7_103[21] , 
        \wRegInTop_7_103[20] , \wRegInTop_7_103[19] , \wRegInTop_7_103[18] , 
        \wRegInTop_7_103[17] , \wRegInTop_7_103[16] , \wRegInTop_7_103[15] , 
        \wRegInTop_7_103[14] , \wRegInTop_7_103[13] , \wRegInTop_7_103[12] , 
        \wRegInTop_7_103[11] , \wRegInTop_7_103[10] , \wRegInTop_7_103[9] , 
        \wRegInTop_7_103[8] , \wRegInTop_7_103[7] , \wRegInTop_7_103[6] , 
        \wRegInTop_7_103[5] , \wRegInTop_7_103[4] , \wRegInTop_7_103[3] , 
        \wRegInTop_7_103[2] , \wRegInTop_7_103[1] , \wRegInTop_7_103[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_30 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink158[31] , \ScanLink158[30] , \ScanLink158[29] , 
        \ScanLink158[28] , \ScanLink158[27] , \ScanLink158[26] , 
        \ScanLink158[25] , \ScanLink158[24] , \ScanLink158[23] , 
        \ScanLink158[22] , \ScanLink158[21] , \ScanLink158[20] , 
        \ScanLink158[19] , \ScanLink158[18] , \ScanLink158[17] , 
        \ScanLink158[16] , \ScanLink158[15] , \ScanLink158[14] , 
        \ScanLink158[13] , \ScanLink158[12] , \ScanLink158[11] , 
        \ScanLink158[10] , \ScanLink158[9] , \ScanLink158[8] , 
        \ScanLink158[7] , \ScanLink158[6] , \ScanLink158[5] , \ScanLink158[4] , 
        \ScanLink158[3] , \ScanLink158[2] , \ScanLink158[1] , \ScanLink158[0] 
        }), .ScanOut({\ScanLink157[31] , \ScanLink157[30] , \ScanLink157[29] , 
        \ScanLink157[28] , \ScanLink157[27] , \ScanLink157[26] , 
        \ScanLink157[25] , \ScanLink157[24] , \ScanLink157[23] , 
        \ScanLink157[22] , \ScanLink157[21] , \ScanLink157[20] , 
        \ScanLink157[19] , \ScanLink157[18] , \ScanLink157[17] , 
        \ScanLink157[16] , \ScanLink157[15] , \ScanLink157[14] , 
        \ScanLink157[13] , \ScanLink157[12] , \ScanLink157[11] , 
        \ScanLink157[10] , \ScanLink157[9] , \ScanLink157[8] , 
        \ScanLink157[7] , \ScanLink157[6] , \ScanLink157[5] , \ScanLink157[4] , 
        \ScanLink157[3] , \ScanLink157[2] , \ScanLink157[1] , \ScanLink157[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_30[31] , 
        \wRegOut_7_30[30] , \wRegOut_7_30[29] , \wRegOut_7_30[28] , 
        \wRegOut_7_30[27] , \wRegOut_7_30[26] , \wRegOut_7_30[25] , 
        \wRegOut_7_30[24] , \wRegOut_7_30[23] , \wRegOut_7_30[22] , 
        \wRegOut_7_30[21] , \wRegOut_7_30[20] , \wRegOut_7_30[19] , 
        \wRegOut_7_30[18] , \wRegOut_7_30[17] , \wRegOut_7_30[16] , 
        \wRegOut_7_30[15] , \wRegOut_7_30[14] , \wRegOut_7_30[13] , 
        \wRegOut_7_30[12] , \wRegOut_7_30[11] , \wRegOut_7_30[10] , 
        \wRegOut_7_30[9] , \wRegOut_7_30[8] , \wRegOut_7_30[7] , 
        \wRegOut_7_30[6] , \wRegOut_7_30[5] , \wRegOut_7_30[4] , 
        \wRegOut_7_30[3] , \wRegOut_7_30[2] , \wRegOut_7_30[1] , 
        \wRegOut_7_30[0] }), .Enable1(\wRegEnTop_7_30[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_30[31] , \wRegInTop_7_30[30] , \wRegInTop_7_30[29] , 
        \wRegInTop_7_30[28] , \wRegInTop_7_30[27] , \wRegInTop_7_30[26] , 
        \wRegInTop_7_30[25] , \wRegInTop_7_30[24] , \wRegInTop_7_30[23] , 
        \wRegInTop_7_30[22] , \wRegInTop_7_30[21] , \wRegInTop_7_30[20] , 
        \wRegInTop_7_30[19] , \wRegInTop_7_30[18] , \wRegInTop_7_30[17] , 
        \wRegInTop_7_30[16] , \wRegInTop_7_30[15] , \wRegInTop_7_30[14] , 
        \wRegInTop_7_30[13] , \wRegInTop_7_30[12] , \wRegInTop_7_30[11] , 
        \wRegInTop_7_30[10] , \wRegInTop_7_30[9] , \wRegInTop_7_30[8] , 
        \wRegInTop_7_30[7] , \wRegInTop_7_30[6] , \wRegInTop_7_30[5] , 
        \wRegInTop_7_30[4] , \wRegInTop_7_30[3] , \wRegInTop_7_30[2] , 
        \wRegInTop_7_30[1] , \wRegInTop_7_30[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_CtrlReg_WIDTH32 BHCR_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_4[0] ), 
        .Out(\wCtrlOut_3[0] ), .Enable(\wEnable_3[0] ) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_124 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink252[31] , \ScanLink252[30] , \ScanLink252[29] , 
        \ScanLink252[28] , \ScanLink252[27] , \ScanLink252[26] , 
        \ScanLink252[25] , \ScanLink252[24] , \ScanLink252[23] , 
        \ScanLink252[22] , \ScanLink252[21] , \ScanLink252[20] , 
        \ScanLink252[19] , \ScanLink252[18] , \ScanLink252[17] , 
        \ScanLink252[16] , \ScanLink252[15] , \ScanLink252[14] , 
        \ScanLink252[13] , \ScanLink252[12] , \ScanLink252[11] , 
        \ScanLink252[10] , \ScanLink252[9] , \ScanLink252[8] , 
        \ScanLink252[7] , \ScanLink252[6] , \ScanLink252[5] , \ScanLink252[4] , 
        \ScanLink252[3] , \ScanLink252[2] , \ScanLink252[1] , \ScanLink252[0] 
        }), .ScanOut({\ScanLink251[31] , \ScanLink251[30] , \ScanLink251[29] , 
        \ScanLink251[28] , \ScanLink251[27] , \ScanLink251[26] , 
        \ScanLink251[25] , \ScanLink251[24] , \ScanLink251[23] , 
        \ScanLink251[22] , \ScanLink251[21] , \ScanLink251[20] , 
        \ScanLink251[19] , \ScanLink251[18] , \ScanLink251[17] , 
        \ScanLink251[16] , \ScanLink251[15] , \ScanLink251[14] , 
        \ScanLink251[13] , \ScanLink251[12] , \ScanLink251[11] , 
        \ScanLink251[10] , \ScanLink251[9] , \ScanLink251[8] , 
        \ScanLink251[7] , \ScanLink251[6] , \ScanLink251[5] , \ScanLink251[4] , 
        \ScanLink251[3] , \ScanLink251[2] , \ScanLink251[1] , \ScanLink251[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_124[31] , 
        \wRegOut_7_124[30] , \wRegOut_7_124[29] , \wRegOut_7_124[28] , 
        \wRegOut_7_124[27] , \wRegOut_7_124[26] , \wRegOut_7_124[25] , 
        \wRegOut_7_124[24] , \wRegOut_7_124[23] , \wRegOut_7_124[22] , 
        \wRegOut_7_124[21] , \wRegOut_7_124[20] , \wRegOut_7_124[19] , 
        \wRegOut_7_124[18] , \wRegOut_7_124[17] , \wRegOut_7_124[16] , 
        \wRegOut_7_124[15] , \wRegOut_7_124[14] , \wRegOut_7_124[13] , 
        \wRegOut_7_124[12] , \wRegOut_7_124[11] , \wRegOut_7_124[10] , 
        \wRegOut_7_124[9] , \wRegOut_7_124[8] , \wRegOut_7_124[7] , 
        \wRegOut_7_124[6] , \wRegOut_7_124[5] , \wRegOut_7_124[4] , 
        \wRegOut_7_124[3] , \wRegOut_7_124[2] , \wRegOut_7_124[1] , 
        \wRegOut_7_124[0] }), .Enable1(\wRegEnTop_7_124[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_124[31] , \wRegInTop_7_124[30] , 
        \wRegInTop_7_124[29] , \wRegInTop_7_124[28] , \wRegInTop_7_124[27] , 
        \wRegInTop_7_124[26] , \wRegInTop_7_124[25] , \wRegInTop_7_124[24] , 
        \wRegInTop_7_124[23] , \wRegInTop_7_124[22] , \wRegInTop_7_124[21] , 
        \wRegInTop_7_124[20] , \wRegInTop_7_124[19] , \wRegInTop_7_124[18] , 
        \wRegInTop_7_124[17] , \wRegInTop_7_124[16] , \wRegInTop_7_124[15] , 
        \wRegInTop_7_124[14] , \wRegInTop_7_124[13] , \wRegInTop_7_124[12] , 
        \wRegInTop_7_124[11] , \wRegInTop_7_124[10] , \wRegInTop_7_124[9] , 
        \wRegInTop_7_124[8] , \wRegInTop_7_124[7] , \wRegInTop_7_124[6] , 
        \wRegInTop_7_124[5] , \wRegInTop_7_124[4] , \wRegInTop_7_124[3] , 
        \wRegInTop_7_124[2] , \wRegInTop_7_124[1] , \wRegInTop_7_124[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_38 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink102[31] , \ScanLink102[30] , \ScanLink102[29] , 
        \ScanLink102[28] , \ScanLink102[27] , \ScanLink102[26] , 
        \ScanLink102[25] , \ScanLink102[24] , \ScanLink102[23] , 
        \ScanLink102[22] , \ScanLink102[21] , \ScanLink102[20] , 
        \ScanLink102[19] , \ScanLink102[18] , \ScanLink102[17] , 
        \ScanLink102[16] , \ScanLink102[15] , \ScanLink102[14] , 
        \ScanLink102[13] , \ScanLink102[12] , \ScanLink102[11] , 
        \ScanLink102[10] , \ScanLink102[9] , \ScanLink102[8] , 
        \ScanLink102[7] , \ScanLink102[6] , \ScanLink102[5] , \ScanLink102[4] , 
        \ScanLink102[3] , \ScanLink102[2] , \ScanLink102[1] , \ScanLink102[0] 
        }), .ScanOut({\ScanLink101[31] , \ScanLink101[30] , \ScanLink101[29] , 
        \ScanLink101[28] , \ScanLink101[27] , \ScanLink101[26] , 
        \ScanLink101[25] , \ScanLink101[24] , \ScanLink101[23] , 
        \ScanLink101[22] , \ScanLink101[21] , \ScanLink101[20] , 
        \ScanLink101[19] , \ScanLink101[18] , \ScanLink101[17] , 
        \ScanLink101[16] , \ScanLink101[15] , \ScanLink101[14] , 
        \ScanLink101[13] , \ScanLink101[12] , \ScanLink101[11] , 
        \ScanLink101[10] , \ScanLink101[9] , \ScanLink101[8] , 
        \ScanLink101[7] , \ScanLink101[6] , \ScanLink101[5] , \ScanLink101[4] , 
        \ScanLink101[3] , \ScanLink101[2] , \ScanLink101[1] , \ScanLink101[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_38[31] , 
        \wRegOut_6_38[30] , \wRegOut_6_38[29] , \wRegOut_6_38[28] , 
        \wRegOut_6_38[27] , \wRegOut_6_38[26] , \wRegOut_6_38[25] , 
        \wRegOut_6_38[24] , \wRegOut_6_38[23] , \wRegOut_6_38[22] , 
        \wRegOut_6_38[21] , \wRegOut_6_38[20] , \wRegOut_6_38[19] , 
        \wRegOut_6_38[18] , \wRegOut_6_38[17] , \wRegOut_6_38[16] , 
        \wRegOut_6_38[15] , \wRegOut_6_38[14] , \wRegOut_6_38[13] , 
        \wRegOut_6_38[12] , \wRegOut_6_38[11] , \wRegOut_6_38[10] , 
        \wRegOut_6_38[9] , \wRegOut_6_38[8] , \wRegOut_6_38[7] , 
        \wRegOut_6_38[6] , \wRegOut_6_38[5] , \wRegOut_6_38[4] , 
        \wRegOut_6_38[3] , \wRegOut_6_38[2] , \wRegOut_6_38[1] , 
        \wRegOut_6_38[0] }), .Enable1(\wRegEnTop_6_38[0] ), .Enable2(
        \wRegEnBot_6_38[0] ), .In1({\wRegInTop_6_38[31] , \wRegInTop_6_38[30] , 
        \wRegInTop_6_38[29] , \wRegInTop_6_38[28] , \wRegInTop_6_38[27] , 
        \wRegInTop_6_38[26] , \wRegInTop_6_38[25] , \wRegInTop_6_38[24] , 
        \wRegInTop_6_38[23] , \wRegInTop_6_38[22] , \wRegInTop_6_38[21] , 
        \wRegInTop_6_38[20] , \wRegInTop_6_38[19] , \wRegInTop_6_38[18] , 
        \wRegInTop_6_38[17] , \wRegInTop_6_38[16] , \wRegInTop_6_38[15] , 
        \wRegInTop_6_38[14] , \wRegInTop_6_38[13] , \wRegInTop_6_38[12] , 
        \wRegInTop_6_38[11] , \wRegInTop_6_38[10] , \wRegInTop_6_38[9] , 
        \wRegInTop_6_38[8] , \wRegInTop_6_38[7] , \wRegInTop_6_38[6] , 
        \wRegInTop_6_38[5] , \wRegInTop_6_38[4] , \wRegInTop_6_38[3] , 
        \wRegInTop_6_38[2] , \wRegInTop_6_38[1] , \wRegInTop_6_38[0] }), .In2(
        {\wRegInBot_6_38[31] , \wRegInBot_6_38[30] , \wRegInBot_6_38[29] , 
        \wRegInBot_6_38[28] , \wRegInBot_6_38[27] , \wRegInBot_6_38[26] , 
        \wRegInBot_6_38[25] , \wRegInBot_6_38[24] , \wRegInBot_6_38[23] , 
        \wRegInBot_6_38[22] , \wRegInBot_6_38[21] , \wRegInBot_6_38[20] , 
        \wRegInBot_6_38[19] , \wRegInBot_6_38[18] , \wRegInBot_6_38[17] , 
        \wRegInBot_6_38[16] , \wRegInBot_6_38[15] , \wRegInBot_6_38[14] , 
        \wRegInBot_6_38[13] , \wRegInBot_6_38[12] , \wRegInBot_6_38[11] , 
        \wRegInBot_6_38[10] , \wRegInBot_6_38[9] , \wRegInBot_6_38[8] , 
        \wRegInBot_6_38[7] , \wRegInBot_6_38[6] , \wRegInBot_6_38[5] , 
        \wRegInBot_6_38[4] , \wRegInBot_6_38[3] , \wRegInBot_6_38[2] , 
        \wRegInBot_6_38[1] , \wRegInBot_6_38[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_79 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink207[31] , \ScanLink207[30] , \ScanLink207[29] , 
        \ScanLink207[28] , \ScanLink207[27] , \ScanLink207[26] , 
        \ScanLink207[25] , \ScanLink207[24] , \ScanLink207[23] , 
        \ScanLink207[22] , \ScanLink207[21] , \ScanLink207[20] , 
        \ScanLink207[19] , \ScanLink207[18] , \ScanLink207[17] , 
        \ScanLink207[16] , \ScanLink207[15] , \ScanLink207[14] , 
        \ScanLink207[13] , \ScanLink207[12] , \ScanLink207[11] , 
        \ScanLink207[10] , \ScanLink207[9] , \ScanLink207[8] , 
        \ScanLink207[7] , \ScanLink207[6] , \ScanLink207[5] , \ScanLink207[4] , 
        \ScanLink207[3] , \ScanLink207[2] , \ScanLink207[1] , \ScanLink207[0] 
        }), .ScanOut({\ScanLink206[31] , \ScanLink206[30] , \ScanLink206[29] , 
        \ScanLink206[28] , \ScanLink206[27] , \ScanLink206[26] , 
        \ScanLink206[25] , \ScanLink206[24] , \ScanLink206[23] , 
        \ScanLink206[22] , \ScanLink206[21] , \ScanLink206[20] , 
        \ScanLink206[19] , \ScanLink206[18] , \ScanLink206[17] , 
        \ScanLink206[16] , \ScanLink206[15] , \ScanLink206[14] , 
        \ScanLink206[13] , \ScanLink206[12] , \ScanLink206[11] , 
        \ScanLink206[10] , \ScanLink206[9] , \ScanLink206[8] , 
        \ScanLink206[7] , \ScanLink206[6] , \ScanLink206[5] , \ScanLink206[4] , 
        \ScanLink206[3] , \ScanLink206[2] , \ScanLink206[1] , \ScanLink206[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_79[31] , 
        \wRegOut_7_79[30] , \wRegOut_7_79[29] , \wRegOut_7_79[28] , 
        \wRegOut_7_79[27] , \wRegOut_7_79[26] , \wRegOut_7_79[25] , 
        \wRegOut_7_79[24] , \wRegOut_7_79[23] , \wRegOut_7_79[22] , 
        \wRegOut_7_79[21] , \wRegOut_7_79[20] , \wRegOut_7_79[19] , 
        \wRegOut_7_79[18] , \wRegOut_7_79[17] , \wRegOut_7_79[16] , 
        \wRegOut_7_79[15] , \wRegOut_7_79[14] , \wRegOut_7_79[13] , 
        \wRegOut_7_79[12] , \wRegOut_7_79[11] , \wRegOut_7_79[10] , 
        \wRegOut_7_79[9] , \wRegOut_7_79[8] , \wRegOut_7_79[7] , 
        \wRegOut_7_79[6] , \wRegOut_7_79[5] , \wRegOut_7_79[4] , 
        \wRegOut_7_79[3] , \wRegOut_7_79[2] , \wRegOut_7_79[1] , 
        \wRegOut_7_79[0] }), .Enable1(\wRegEnTop_7_79[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_79[31] , \wRegInTop_7_79[30] , \wRegInTop_7_79[29] , 
        \wRegInTop_7_79[28] , \wRegInTop_7_79[27] , \wRegInTop_7_79[26] , 
        \wRegInTop_7_79[25] , \wRegInTop_7_79[24] , \wRegInTop_7_79[23] , 
        \wRegInTop_7_79[22] , \wRegInTop_7_79[21] , \wRegInTop_7_79[20] , 
        \wRegInTop_7_79[19] , \wRegInTop_7_79[18] , \wRegInTop_7_79[17] , 
        \wRegInTop_7_79[16] , \wRegInTop_7_79[15] , \wRegInTop_7_79[14] , 
        \wRegInTop_7_79[13] , \wRegInTop_7_79[12] , \wRegInTop_7_79[11] , 
        \wRegInTop_7_79[10] , \wRegInTop_7_79[9] , \wRegInTop_7_79[8] , 
        \wRegInTop_7_79[7] , \wRegInTop_7_79[6] , \wRegInTop_7_79[5] , 
        \wRegInTop_7_79[4] , \wRegInTop_7_79[3] , \wRegInTop_7_79[2] , 
        \wRegInTop_7_79[1] , \wRegInTop_7_79[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_25[0] ), .P_In({\wRegOut_6_25[31] , 
        \wRegOut_6_25[30] , \wRegOut_6_25[29] , \wRegOut_6_25[28] , 
        \wRegOut_6_25[27] , \wRegOut_6_25[26] , \wRegOut_6_25[25] , 
        \wRegOut_6_25[24] , \wRegOut_6_25[23] , \wRegOut_6_25[22] , 
        \wRegOut_6_25[21] , \wRegOut_6_25[20] , \wRegOut_6_25[19] , 
        \wRegOut_6_25[18] , \wRegOut_6_25[17] , \wRegOut_6_25[16] , 
        \wRegOut_6_25[15] , \wRegOut_6_25[14] , \wRegOut_6_25[13] , 
        \wRegOut_6_25[12] , \wRegOut_6_25[11] , \wRegOut_6_25[10] , 
        \wRegOut_6_25[9] , \wRegOut_6_25[8] , \wRegOut_6_25[7] , 
        \wRegOut_6_25[6] , \wRegOut_6_25[5] , \wRegOut_6_25[4] , 
        \wRegOut_6_25[3] , \wRegOut_6_25[2] , \wRegOut_6_25[1] , 
        \wRegOut_6_25[0] }), .P_Out({\wRegInBot_6_25[31] , 
        \wRegInBot_6_25[30] , \wRegInBot_6_25[29] , \wRegInBot_6_25[28] , 
        \wRegInBot_6_25[27] , \wRegInBot_6_25[26] , \wRegInBot_6_25[25] , 
        \wRegInBot_6_25[24] , \wRegInBot_6_25[23] , \wRegInBot_6_25[22] , 
        \wRegInBot_6_25[21] , \wRegInBot_6_25[20] , \wRegInBot_6_25[19] , 
        \wRegInBot_6_25[18] , \wRegInBot_6_25[17] , \wRegInBot_6_25[16] , 
        \wRegInBot_6_25[15] , \wRegInBot_6_25[14] , \wRegInBot_6_25[13] , 
        \wRegInBot_6_25[12] , \wRegInBot_6_25[11] , \wRegInBot_6_25[10] , 
        \wRegInBot_6_25[9] , \wRegInBot_6_25[8] , \wRegInBot_6_25[7] , 
        \wRegInBot_6_25[6] , \wRegInBot_6_25[5] , \wRegInBot_6_25[4] , 
        \wRegInBot_6_25[3] , \wRegInBot_6_25[2] , \wRegInBot_6_25[1] , 
        \wRegInBot_6_25[0] }), .L_WR(\wRegEnTop_7_50[0] ), .L_In({
        \wRegOut_7_50[31] , \wRegOut_7_50[30] , \wRegOut_7_50[29] , 
        \wRegOut_7_50[28] , \wRegOut_7_50[27] , \wRegOut_7_50[26] , 
        \wRegOut_7_50[25] , \wRegOut_7_50[24] , \wRegOut_7_50[23] , 
        \wRegOut_7_50[22] , \wRegOut_7_50[21] , \wRegOut_7_50[20] , 
        \wRegOut_7_50[19] , \wRegOut_7_50[18] , \wRegOut_7_50[17] , 
        \wRegOut_7_50[16] , \wRegOut_7_50[15] , \wRegOut_7_50[14] , 
        \wRegOut_7_50[13] , \wRegOut_7_50[12] , \wRegOut_7_50[11] , 
        \wRegOut_7_50[10] , \wRegOut_7_50[9] , \wRegOut_7_50[8] , 
        \wRegOut_7_50[7] , \wRegOut_7_50[6] , \wRegOut_7_50[5] , 
        \wRegOut_7_50[4] , \wRegOut_7_50[3] , \wRegOut_7_50[2] , 
        \wRegOut_7_50[1] , \wRegOut_7_50[0] }), .L_Out({\wRegInTop_7_50[31] , 
        \wRegInTop_7_50[30] , \wRegInTop_7_50[29] , \wRegInTop_7_50[28] , 
        \wRegInTop_7_50[27] , \wRegInTop_7_50[26] , \wRegInTop_7_50[25] , 
        \wRegInTop_7_50[24] , \wRegInTop_7_50[23] , \wRegInTop_7_50[22] , 
        \wRegInTop_7_50[21] , \wRegInTop_7_50[20] , \wRegInTop_7_50[19] , 
        \wRegInTop_7_50[18] , \wRegInTop_7_50[17] , \wRegInTop_7_50[16] , 
        \wRegInTop_7_50[15] , \wRegInTop_7_50[14] , \wRegInTop_7_50[13] , 
        \wRegInTop_7_50[12] , \wRegInTop_7_50[11] , \wRegInTop_7_50[10] , 
        \wRegInTop_7_50[9] , \wRegInTop_7_50[8] , \wRegInTop_7_50[7] , 
        \wRegInTop_7_50[6] , \wRegInTop_7_50[5] , \wRegInTop_7_50[4] , 
        \wRegInTop_7_50[3] , \wRegInTop_7_50[2] , \wRegInTop_7_50[1] , 
        \wRegInTop_7_50[0] }), .R_WR(\wRegEnTop_7_51[0] ), .R_In({
        \wRegOut_7_51[31] , \wRegOut_7_51[30] , \wRegOut_7_51[29] , 
        \wRegOut_7_51[28] , \wRegOut_7_51[27] , \wRegOut_7_51[26] , 
        \wRegOut_7_51[25] , \wRegOut_7_51[24] , \wRegOut_7_51[23] , 
        \wRegOut_7_51[22] , \wRegOut_7_51[21] , \wRegOut_7_51[20] , 
        \wRegOut_7_51[19] , \wRegOut_7_51[18] , \wRegOut_7_51[17] , 
        \wRegOut_7_51[16] , \wRegOut_7_51[15] , \wRegOut_7_51[14] , 
        \wRegOut_7_51[13] , \wRegOut_7_51[12] , \wRegOut_7_51[11] , 
        \wRegOut_7_51[10] , \wRegOut_7_51[9] , \wRegOut_7_51[8] , 
        \wRegOut_7_51[7] , \wRegOut_7_51[6] , \wRegOut_7_51[5] , 
        \wRegOut_7_51[4] , \wRegOut_7_51[3] , \wRegOut_7_51[2] , 
        \wRegOut_7_51[1] , \wRegOut_7_51[0] }), .R_Out({\wRegInTop_7_51[31] , 
        \wRegInTop_7_51[30] , \wRegInTop_7_51[29] , \wRegInTop_7_51[28] , 
        \wRegInTop_7_51[27] , \wRegInTop_7_51[26] , \wRegInTop_7_51[25] , 
        \wRegInTop_7_51[24] , \wRegInTop_7_51[23] , \wRegInTop_7_51[22] , 
        \wRegInTop_7_51[21] , \wRegInTop_7_51[20] , \wRegInTop_7_51[19] , 
        \wRegInTop_7_51[18] , \wRegInTop_7_51[17] , \wRegInTop_7_51[16] , 
        \wRegInTop_7_51[15] , \wRegInTop_7_51[14] , \wRegInTop_7_51[13] , 
        \wRegInTop_7_51[12] , \wRegInTop_7_51[11] , \wRegInTop_7_51[10] , 
        \wRegInTop_7_51[9] , \wRegInTop_7_51[8] , \wRegInTop_7_51[7] , 
        \wRegInTop_7_51[6] , \wRegInTop_7_51[5] , \wRegInTop_7_51[4] , 
        \wRegInTop_7_51[3] , \wRegInTop_7_51[2] , \wRegInTop_7_51[1] , 
        \wRegInTop_7_51[0] }) );
    BHeap_Node_WIDTH32 BHN_5_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_15[0] ), .P_In({\wRegOut_5_15[31] , 
        \wRegOut_5_15[30] , \wRegOut_5_15[29] , \wRegOut_5_15[28] , 
        \wRegOut_5_15[27] , \wRegOut_5_15[26] , \wRegOut_5_15[25] , 
        \wRegOut_5_15[24] , \wRegOut_5_15[23] , \wRegOut_5_15[22] , 
        \wRegOut_5_15[21] , \wRegOut_5_15[20] , \wRegOut_5_15[19] , 
        \wRegOut_5_15[18] , \wRegOut_5_15[17] , \wRegOut_5_15[16] , 
        \wRegOut_5_15[15] , \wRegOut_5_15[14] , \wRegOut_5_15[13] , 
        \wRegOut_5_15[12] , \wRegOut_5_15[11] , \wRegOut_5_15[10] , 
        \wRegOut_5_15[9] , \wRegOut_5_15[8] , \wRegOut_5_15[7] , 
        \wRegOut_5_15[6] , \wRegOut_5_15[5] , \wRegOut_5_15[4] , 
        \wRegOut_5_15[3] , \wRegOut_5_15[2] , \wRegOut_5_15[1] , 
        \wRegOut_5_15[0] }), .P_Out({\wRegInBot_5_15[31] , 
        \wRegInBot_5_15[30] , \wRegInBot_5_15[29] , \wRegInBot_5_15[28] , 
        \wRegInBot_5_15[27] , \wRegInBot_5_15[26] , \wRegInBot_5_15[25] , 
        \wRegInBot_5_15[24] , \wRegInBot_5_15[23] , \wRegInBot_5_15[22] , 
        \wRegInBot_5_15[21] , \wRegInBot_5_15[20] , \wRegInBot_5_15[19] , 
        \wRegInBot_5_15[18] , \wRegInBot_5_15[17] , \wRegInBot_5_15[16] , 
        \wRegInBot_5_15[15] , \wRegInBot_5_15[14] , \wRegInBot_5_15[13] , 
        \wRegInBot_5_15[12] , \wRegInBot_5_15[11] , \wRegInBot_5_15[10] , 
        \wRegInBot_5_15[9] , \wRegInBot_5_15[8] , \wRegInBot_5_15[7] , 
        \wRegInBot_5_15[6] , \wRegInBot_5_15[5] , \wRegInBot_5_15[4] , 
        \wRegInBot_5_15[3] , \wRegInBot_5_15[2] , \wRegInBot_5_15[1] , 
        \wRegInBot_5_15[0] }), .L_WR(\wRegEnTop_6_30[0] ), .L_In({
        \wRegOut_6_30[31] , \wRegOut_6_30[30] , \wRegOut_6_30[29] , 
        \wRegOut_6_30[28] , \wRegOut_6_30[27] , \wRegOut_6_30[26] , 
        \wRegOut_6_30[25] , \wRegOut_6_30[24] , \wRegOut_6_30[23] , 
        \wRegOut_6_30[22] , \wRegOut_6_30[21] , \wRegOut_6_30[20] , 
        \wRegOut_6_30[19] , \wRegOut_6_30[18] , \wRegOut_6_30[17] , 
        \wRegOut_6_30[16] , \wRegOut_6_30[15] , \wRegOut_6_30[14] , 
        \wRegOut_6_30[13] , \wRegOut_6_30[12] , \wRegOut_6_30[11] , 
        \wRegOut_6_30[10] , \wRegOut_6_30[9] , \wRegOut_6_30[8] , 
        \wRegOut_6_30[7] , \wRegOut_6_30[6] , \wRegOut_6_30[5] , 
        \wRegOut_6_30[4] , \wRegOut_6_30[3] , \wRegOut_6_30[2] , 
        \wRegOut_6_30[1] , \wRegOut_6_30[0] }), .L_Out({\wRegInTop_6_30[31] , 
        \wRegInTop_6_30[30] , \wRegInTop_6_30[29] , \wRegInTop_6_30[28] , 
        \wRegInTop_6_30[27] , \wRegInTop_6_30[26] , \wRegInTop_6_30[25] , 
        \wRegInTop_6_30[24] , \wRegInTop_6_30[23] , \wRegInTop_6_30[22] , 
        \wRegInTop_6_30[21] , \wRegInTop_6_30[20] , \wRegInTop_6_30[19] , 
        \wRegInTop_6_30[18] , \wRegInTop_6_30[17] , \wRegInTop_6_30[16] , 
        \wRegInTop_6_30[15] , \wRegInTop_6_30[14] , \wRegInTop_6_30[13] , 
        \wRegInTop_6_30[12] , \wRegInTop_6_30[11] , \wRegInTop_6_30[10] , 
        \wRegInTop_6_30[9] , \wRegInTop_6_30[8] , \wRegInTop_6_30[7] , 
        \wRegInTop_6_30[6] , \wRegInTop_6_30[5] , \wRegInTop_6_30[4] , 
        \wRegInTop_6_30[3] , \wRegInTop_6_30[2] , \wRegInTop_6_30[1] , 
        \wRegInTop_6_30[0] }), .R_WR(\wRegEnTop_6_31[0] ), .R_In({
        \wRegOut_6_31[31] , \wRegOut_6_31[30] , \wRegOut_6_31[29] , 
        \wRegOut_6_31[28] , \wRegOut_6_31[27] , \wRegOut_6_31[26] , 
        \wRegOut_6_31[25] , \wRegOut_6_31[24] , \wRegOut_6_31[23] , 
        \wRegOut_6_31[22] , \wRegOut_6_31[21] , \wRegOut_6_31[20] , 
        \wRegOut_6_31[19] , \wRegOut_6_31[18] , \wRegOut_6_31[17] , 
        \wRegOut_6_31[16] , \wRegOut_6_31[15] , \wRegOut_6_31[14] , 
        \wRegOut_6_31[13] , \wRegOut_6_31[12] , \wRegOut_6_31[11] , 
        \wRegOut_6_31[10] , \wRegOut_6_31[9] , \wRegOut_6_31[8] , 
        \wRegOut_6_31[7] , \wRegOut_6_31[6] , \wRegOut_6_31[5] , 
        \wRegOut_6_31[4] , \wRegOut_6_31[3] , \wRegOut_6_31[2] , 
        \wRegOut_6_31[1] , \wRegOut_6_31[0] }), .R_Out({\wRegInTop_6_31[31] , 
        \wRegInTop_6_31[30] , \wRegInTop_6_31[29] , \wRegInTop_6_31[28] , 
        \wRegInTop_6_31[27] , \wRegInTop_6_31[26] , \wRegInTop_6_31[25] , 
        \wRegInTop_6_31[24] , \wRegInTop_6_31[23] , \wRegInTop_6_31[22] , 
        \wRegInTop_6_31[21] , \wRegInTop_6_31[20] , \wRegInTop_6_31[19] , 
        \wRegInTop_6_31[18] , \wRegInTop_6_31[17] , \wRegInTop_6_31[16] , 
        \wRegInTop_6_31[15] , \wRegInTop_6_31[14] , \wRegInTop_6_31[13] , 
        \wRegInTop_6_31[12] , \wRegInTop_6_31[11] , \wRegInTop_6_31[10] , 
        \wRegInTop_6_31[9] , \wRegInTop_6_31[8] , \wRegInTop_6_31[7] , 
        \wRegInTop_6_31[6] , \wRegInTop_6_31[5] , \wRegInTop_6_31[4] , 
        \wRegInTop_6_31[3] , \wRegInTop_6_31[2] , \wRegInTop_6_31[1] , 
        \wRegInTop_6_31[0] }) );
    BHeap_Node_WIDTH32 BHN_5_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_20[0] ), .P_In({\wRegOut_5_20[31] , 
        \wRegOut_5_20[30] , \wRegOut_5_20[29] , \wRegOut_5_20[28] , 
        \wRegOut_5_20[27] , \wRegOut_5_20[26] , \wRegOut_5_20[25] , 
        \wRegOut_5_20[24] , \wRegOut_5_20[23] , \wRegOut_5_20[22] , 
        \wRegOut_5_20[21] , \wRegOut_5_20[20] , \wRegOut_5_20[19] , 
        \wRegOut_5_20[18] , \wRegOut_5_20[17] , \wRegOut_5_20[16] , 
        \wRegOut_5_20[15] , \wRegOut_5_20[14] , \wRegOut_5_20[13] , 
        \wRegOut_5_20[12] , \wRegOut_5_20[11] , \wRegOut_5_20[10] , 
        \wRegOut_5_20[9] , \wRegOut_5_20[8] , \wRegOut_5_20[7] , 
        \wRegOut_5_20[6] , \wRegOut_5_20[5] , \wRegOut_5_20[4] , 
        \wRegOut_5_20[3] , \wRegOut_5_20[2] , \wRegOut_5_20[1] , 
        \wRegOut_5_20[0] }), .P_Out({\wRegInBot_5_20[31] , 
        \wRegInBot_5_20[30] , \wRegInBot_5_20[29] , \wRegInBot_5_20[28] , 
        \wRegInBot_5_20[27] , \wRegInBot_5_20[26] , \wRegInBot_5_20[25] , 
        \wRegInBot_5_20[24] , \wRegInBot_5_20[23] , \wRegInBot_5_20[22] , 
        \wRegInBot_5_20[21] , \wRegInBot_5_20[20] , \wRegInBot_5_20[19] , 
        \wRegInBot_5_20[18] , \wRegInBot_5_20[17] , \wRegInBot_5_20[16] , 
        \wRegInBot_5_20[15] , \wRegInBot_5_20[14] , \wRegInBot_5_20[13] , 
        \wRegInBot_5_20[12] , \wRegInBot_5_20[11] , \wRegInBot_5_20[10] , 
        \wRegInBot_5_20[9] , \wRegInBot_5_20[8] , \wRegInBot_5_20[7] , 
        \wRegInBot_5_20[6] , \wRegInBot_5_20[5] , \wRegInBot_5_20[4] , 
        \wRegInBot_5_20[3] , \wRegInBot_5_20[2] , \wRegInBot_5_20[1] , 
        \wRegInBot_5_20[0] }), .L_WR(\wRegEnTop_6_40[0] ), .L_In({
        \wRegOut_6_40[31] , \wRegOut_6_40[30] , \wRegOut_6_40[29] , 
        \wRegOut_6_40[28] , \wRegOut_6_40[27] , \wRegOut_6_40[26] , 
        \wRegOut_6_40[25] , \wRegOut_6_40[24] , \wRegOut_6_40[23] , 
        \wRegOut_6_40[22] , \wRegOut_6_40[21] , \wRegOut_6_40[20] , 
        \wRegOut_6_40[19] , \wRegOut_6_40[18] , \wRegOut_6_40[17] , 
        \wRegOut_6_40[16] , \wRegOut_6_40[15] , \wRegOut_6_40[14] , 
        \wRegOut_6_40[13] , \wRegOut_6_40[12] , \wRegOut_6_40[11] , 
        \wRegOut_6_40[10] , \wRegOut_6_40[9] , \wRegOut_6_40[8] , 
        \wRegOut_6_40[7] , \wRegOut_6_40[6] , \wRegOut_6_40[5] , 
        \wRegOut_6_40[4] , \wRegOut_6_40[3] , \wRegOut_6_40[2] , 
        \wRegOut_6_40[1] , \wRegOut_6_40[0] }), .L_Out({\wRegInTop_6_40[31] , 
        \wRegInTop_6_40[30] , \wRegInTop_6_40[29] , \wRegInTop_6_40[28] , 
        \wRegInTop_6_40[27] , \wRegInTop_6_40[26] , \wRegInTop_6_40[25] , 
        \wRegInTop_6_40[24] , \wRegInTop_6_40[23] , \wRegInTop_6_40[22] , 
        \wRegInTop_6_40[21] , \wRegInTop_6_40[20] , \wRegInTop_6_40[19] , 
        \wRegInTop_6_40[18] , \wRegInTop_6_40[17] , \wRegInTop_6_40[16] , 
        \wRegInTop_6_40[15] , \wRegInTop_6_40[14] , \wRegInTop_6_40[13] , 
        \wRegInTop_6_40[12] , \wRegInTop_6_40[11] , \wRegInTop_6_40[10] , 
        \wRegInTop_6_40[9] , \wRegInTop_6_40[8] , \wRegInTop_6_40[7] , 
        \wRegInTop_6_40[6] , \wRegInTop_6_40[5] , \wRegInTop_6_40[4] , 
        \wRegInTop_6_40[3] , \wRegInTop_6_40[2] , \wRegInTop_6_40[1] , 
        \wRegInTop_6_40[0] }), .R_WR(\wRegEnTop_6_41[0] ), .R_In({
        \wRegOut_6_41[31] , \wRegOut_6_41[30] , \wRegOut_6_41[29] , 
        \wRegOut_6_41[28] , \wRegOut_6_41[27] , \wRegOut_6_41[26] , 
        \wRegOut_6_41[25] , \wRegOut_6_41[24] , \wRegOut_6_41[23] , 
        \wRegOut_6_41[22] , \wRegOut_6_41[21] , \wRegOut_6_41[20] , 
        \wRegOut_6_41[19] , \wRegOut_6_41[18] , \wRegOut_6_41[17] , 
        \wRegOut_6_41[16] , \wRegOut_6_41[15] , \wRegOut_6_41[14] , 
        \wRegOut_6_41[13] , \wRegOut_6_41[12] , \wRegOut_6_41[11] , 
        \wRegOut_6_41[10] , \wRegOut_6_41[9] , \wRegOut_6_41[8] , 
        \wRegOut_6_41[7] , \wRegOut_6_41[6] , \wRegOut_6_41[5] , 
        \wRegOut_6_41[4] , \wRegOut_6_41[3] , \wRegOut_6_41[2] , 
        \wRegOut_6_41[1] , \wRegOut_6_41[0] }), .R_Out({\wRegInTop_6_41[31] , 
        \wRegInTop_6_41[30] , \wRegInTop_6_41[29] , \wRegInTop_6_41[28] , 
        \wRegInTop_6_41[27] , \wRegInTop_6_41[26] , \wRegInTop_6_41[25] , 
        \wRegInTop_6_41[24] , \wRegInTop_6_41[23] , \wRegInTop_6_41[22] , 
        \wRegInTop_6_41[21] , \wRegInTop_6_41[20] , \wRegInTop_6_41[19] , 
        \wRegInTop_6_41[18] , \wRegInTop_6_41[17] , \wRegInTop_6_41[16] , 
        \wRegInTop_6_41[15] , \wRegInTop_6_41[14] , \wRegInTop_6_41[13] , 
        \wRegInTop_6_41[12] , \wRegInTop_6_41[11] , \wRegInTop_6_41[10] , 
        \wRegInTop_6_41[9] , \wRegInTop_6_41[8] , \wRegInTop_6_41[7] , 
        \wRegInTop_6_41[6] , \wRegInTop_6_41[5] , \wRegInTop_6_41[4] , 
        \wRegInTop_6_41[3] , \wRegInTop_6_41[2] , \wRegInTop_6_41[1] , 
        \wRegInTop_6_41[0] }) );
    BHeap_Node_WIDTH32 BHN_6_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_10[0] ), .P_In({\wRegOut_6_10[31] , 
        \wRegOut_6_10[30] , \wRegOut_6_10[29] , \wRegOut_6_10[28] , 
        \wRegOut_6_10[27] , \wRegOut_6_10[26] , \wRegOut_6_10[25] , 
        \wRegOut_6_10[24] , \wRegOut_6_10[23] , \wRegOut_6_10[22] , 
        \wRegOut_6_10[21] , \wRegOut_6_10[20] , \wRegOut_6_10[19] , 
        \wRegOut_6_10[18] , \wRegOut_6_10[17] , \wRegOut_6_10[16] , 
        \wRegOut_6_10[15] , \wRegOut_6_10[14] , \wRegOut_6_10[13] , 
        \wRegOut_6_10[12] , \wRegOut_6_10[11] , \wRegOut_6_10[10] , 
        \wRegOut_6_10[9] , \wRegOut_6_10[8] , \wRegOut_6_10[7] , 
        \wRegOut_6_10[6] , \wRegOut_6_10[5] , \wRegOut_6_10[4] , 
        \wRegOut_6_10[3] , \wRegOut_6_10[2] , \wRegOut_6_10[1] , 
        \wRegOut_6_10[0] }), .P_Out({\wRegInBot_6_10[31] , 
        \wRegInBot_6_10[30] , \wRegInBot_6_10[29] , \wRegInBot_6_10[28] , 
        \wRegInBot_6_10[27] , \wRegInBot_6_10[26] , \wRegInBot_6_10[25] , 
        \wRegInBot_6_10[24] , \wRegInBot_6_10[23] , \wRegInBot_6_10[22] , 
        \wRegInBot_6_10[21] , \wRegInBot_6_10[20] , \wRegInBot_6_10[19] , 
        \wRegInBot_6_10[18] , \wRegInBot_6_10[17] , \wRegInBot_6_10[16] , 
        \wRegInBot_6_10[15] , \wRegInBot_6_10[14] , \wRegInBot_6_10[13] , 
        \wRegInBot_6_10[12] , \wRegInBot_6_10[11] , \wRegInBot_6_10[10] , 
        \wRegInBot_6_10[9] , \wRegInBot_6_10[8] , \wRegInBot_6_10[7] , 
        \wRegInBot_6_10[6] , \wRegInBot_6_10[5] , \wRegInBot_6_10[4] , 
        \wRegInBot_6_10[3] , \wRegInBot_6_10[2] , \wRegInBot_6_10[1] , 
        \wRegInBot_6_10[0] }), .L_WR(\wRegEnTop_7_20[0] ), .L_In({
        \wRegOut_7_20[31] , \wRegOut_7_20[30] , \wRegOut_7_20[29] , 
        \wRegOut_7_20[28] , \wRegOut_7_20[27] , \wRegOut_7_20[26] , 
        \wRegOut_7_20[25] , \wRegOut_7_20[24] , \wRegOut_7_20[23] , 
        \wRegOut_7_20[22] , \wRegOut_7_20[21] , \wRegOut_7_20[20] , 
        \wRegOut_7_20[19] , \wRegOut_7_20[18] , \wRegOut_7_20[17] , 
        \wRegOut_7_20[16] , \wRegOut_7_20[15] , \wRegOut_7_20[14] , 
        \wRegOut_7_20[13] , \wRegOut_7_20[12] , \wRegOut_7_20[11] , 
        \wRegOut_7_20[10] , \wRegOut_7_20[9] , \wRegOut_7_20[8] , 
        \wRegOut_7_20[7] , \wRegOut_7_20[6] , \wRegOut_7_20[5] , 
        \wRegOut_7_20[4] , \wRegOut_7_20[3] , \wRegOut_7_20[2] , 
        \wRegOut_7_20[1] , \wRegOut_7_20[0] }), .L_Out({\wRegInTop_7_20[31] , 
        \wRegInTop_7_20[30] , \wRegInTop_7_20[29] , \wRegInTop_7_20[28] , 
        \wRegInTop_7_20[27] , \wRegInTop_7_20[26] , \wRegInTop_7_20[25] , 
        \wRegInTop_7_20[24] , \wRegInTop_7_20[23] , \wRegInTop_7_20[22] , 
        \wRegInTop_7_20[21] , \wRegInTop_7_20[20] , \wRegInTop_7_20[19] , 
        \wRegInTop_7_20[18] , \wRegInTop_7_20[17] , \wRegInTop_7_20[16] , 
        \wRegInTop_7_20[15] , \wRegInTop_7_20[14] , \wRegInTop_7_20[13] , 
        \wRegInTop_7_20[12] , \wRegInTop_7_20[11] , \wRegInTop_7_20[10] , 
        \wRegInTop_7_20[9] , \wRegInTop_7_20[8] , \wRegInTop_7_20[7] , 
        \wRegInTop_7_20[6] , \wRegInTop_7_20[5] , \wRegInTop_7_20[4] , 
        \wRegInTop_7_20[3] , \wRegInTop_7_20[2] , \wRegInTop_7_20[1] , 
        \wRegInTop_7_20[0] }), .R_WR(\wRegEnTop_7_21[0] ), .R_In({
        \wRegOut_7_21[31] , \wRegOut_7_21[30] , \wRegOut_7_21[29] , 
        \wRegOut_7_21[28] , \wRegOut_7_21[27] , \wRegOut_7_21[26] , 
        \wRegOut_7_21[25] , \wRegOut_7_21[24] , \wRegOut_7_21[23] , 
        \wRegOut_7_21[22] , \wRegOut_7_21[21] , \wRegOut_7_21[20] , 
        \wRegOut_7_21[19] , \wRegOut_7_21[18] , \wRegOut_7_21[17] , 
        \wRegOut_7_21[16] , \wRegOut_7_21[15] , \wRegOut_7_21[14] , 
        \wRegOut_7_21[13] , \wRegOut_7_21[12] , \wRegOut_7_21[11] , 
        \wRegOut_7_21[10] , \wRegOut_7_21[9] , \wRegOut_7_21[8] , 
        \wRegOut_7_21[7] , \wRegOut_7_21[6] , \wRegOut_7_21[5] , 
        \wRegOut_7_21[4] , \wRegOut_7_21[3] , \wRegOut_7_21[2] , 
        \wRegOut_7_21[1] , \wRegOut_7_21[0] }), .R_Out({\wRegInTop_7_21[31] , 
        \wRegInTop_7_21[30] , \wRegInTop_7_21[29] , \wRegInTop_7_21[28] , 
        \wRegInTop_7_21[27] , \wRegInTop_7_21[26] , \wRegInTop_7_21[25] , 
        \wRegInTop_7_21[24] , \wRegInTop_7_21[23] , \wRegInTop_7_21[22] , 
        \wRegInTop_7_21[21] , \wRegInTop_7_21[20] , \wRegInTop_7_21[19] , 
        \wRegInTop_7_21[18] , \wRegInTop_7_21[17] , \wRegInTop_7_21[16] , 
        \wRegInTop_7_21[15] , \wRegInTop_7_21[14] , \wRegInTop_7_21[13] , 
        \wRegInTop_7_21[12] , \wRegInTop_7_21[11] , \wRegInTop_7_21[10] , 
        \wRegInTop_7_21[9] , \wRegInTop_7_21[8] , \wRegInTop_7_21[7] , 
        \wRegInTop_7_21[6] , \wRegInTop_7_21[5] , \wRegInTop_7_21[4] , 
        \wRegInTop_7_21[3] , \wRegInTop_7_21[2] , \wRegInTop_7_21[1] , 
        \wRegInTop_7_21[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_0_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink1[31] , \ScanLink1[30] , \ScanLink1[29] , 
        \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , \ScanLink1[25] , 
        \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , \ScanLink1[21] , 
        \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , \ScanLink1[17] , 
        \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , \ScanLink1[13] , 
        \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , \ScanLink1[9] , 
        \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , \ScanLink1[5] , 
        \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , \ScanLink1[1] , 
        \ScanLink1[0] }), .ScanOut({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_0_0[31] , \wRegOut_0_0[30] , \wRegOut_0_0[29] , 
        \wRegOut_0_0[28] , \wRegOut_0_0[27] , \wRegOut_0_0[26] , 
        \wRegOut_0_0[25] , \wRegOut_0_0[24] , \wRegOut_0_0[23] , 
        \wRegOut_0_0[22] , \wRegOut_0_0[21] , \wRegOut_0_0[20] , 
        \wRegOut_0_0[19] , \wRegOut_0_0[18] , \wRegOut_0_0[17] , 
        \wRegOut_0_0[16] , \wRegOut_0_0[15] , \wRegOut_0_0[14] , 
        \wRegOut_0_0[13] , \wRegOut_0_0[12] , \wRegOut_0_0[11] , 
        \wRegOut_0_0[10] , \wRegOut_0_0[9] , \wRegOut_0_0[8] , 
        \wRegOut_0_0[7] , \wRegOut_0_0[6] , \wRegOut_0_0[5] , \wRegOut_0_0[4] , 
        \wRegOut_0_0[3] , \wRegOut_0_0[2] , \wRegOut_0_0[1] , \wRegOut_0_0[0] 
        }), .Enable1(1'b0), .Enable2(\wRegEnBot_0_0[0] ), .In1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .In2({\wRegInBot_0_0[31] , 
        \wRegInBot_0_0[30] , \wRegInBot_0_0[29] , \wRegInBot_0_0[28] , 
        \wRegInBot_0_0[27] , \wRegInBot_0_0[26] , \wRegInBot_0_0[25] , 
        \wRegInBot_0_0[24] , \wRegInBot_0_0[23] , \wRegInBot_0_0[22] , 
        \wRegInBot_0_0[21] , \wRegInBot_0_0[20] , \wRegInBot_0_0[19] , 
        \wRegInBot_0_0[18] , \wRegInBot_0_0[17] , \wRegInBot_0_0[16] , 
        \wRegInBot_0_0[15] , \wRegInBot_0_0[14] , \wRegInBot_0_0[13] , 
        \wRegInBot_0_0[12] , \wRegInBot_0_0[11] , \wRegInBot_0_0[10] , 
        \wRegInBot_0_0[9] , \wRegInBot_0_0[8] , \wRegInBot_0_0[7] , 
        \wRegInBot_0_0[6] , \wRegInBot_0_0[5] , \wRegInBot_0_0[4] , 
        \wRegInBot_0_0[3] , \wRegInBot_0_0[2] , \wRegInBot_0_0[1] , 
        \wRegInBot_0_0[0] }) );
    BHeap_Node_WIDTH32 BHN_6_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_37[0] ), .P_In({\wRegOut_6_37[31] , 
        \wRegOut_6_37[30] , \wRegOut_6_37[29] , \wRegOut_6_37[28] , 
        \wRegOut_6_37[27] , \wRegOut_6_37[26] , \wRegOut_6_37[25] , 
        \wRegOut_6_37[24] , \wRegOut_6_37[23] , \wRegOut_6_37[22] , 
        \wRegOut_6_37[21] , \wRegOut_6_37[20] , \wRegOut_6_37[19] , 
        \wRegOut_6_37[18] , \wRegOut_6_37[17] , \wRegOut_6_37[16] , 
        \wRegOut_6_37[15] , \wRegOut_6_37[14] , \wRegOut_6_37[13] , 
        \wRegOut_6_37[12] , \wRegOut_6_37[11] , \wRegOut_6_37[10] , 
        \wRegOut_6_37[9] , \wRegOut_6_37[8] , \wRegOut_6_37[7] , 
        \wRegOut_6_37[6] , \wRegOut_6_37[5] , \wRegOut_6_37[4] , 
        \wRegOut_6_37[3] , \wRegOut_6_37[2] , \wRegOut_6_37[1] , 
        \wRegOut_6_37[0] }), .P_Out({\wRegInBot_6_37[31] , 
        \wRegInBot_6_37[30] , \wRegInBot_6_37[29] , \wRegInBot_6_37[28] , 
        \wRegInBot_6_37[27] , \wRegInBot_6_37[26] , \wRegInBot_6_37[25] , 
        \wRegInBot_6_37[24] , \wRegInBot_6_37[23] , \wRegInBot_6_37[22] , 
        \wRegInBot_6_37[21] , \wRegInBot_6_37[20] , \wRegInBot_6_37[19] , 
        \wRegInBot_6_37[18] , \wRegInBot_6_37[17] , \wRegInBot_6_37[16] , 
        \wRegInBot_6_37[15] , \wRegInBot_6_37[14] , \wRegInBot_6_37[13] , 
        \wRegInBot_6_37[12] , \wRegInBot_6_37[11] , \wRegInBot_6_37[10] , 
        \wRegInBot_6_37[9] , \wRegInBot_6_37[8] , \wRegInBot_6_37[7] , 
        \wRegInBot_6_37[6] , \wRegInBot_6_37[5] , \wRegInBot_6_37[4] , 
        \wRegInBot_6_37[3] , \wRegInBot_6_37[2] , \wRegInBot_6_37[1] , 
        \wRegInBot_6_37[0] }), .L_WR(\wRegEnTop_7_74[0] ), .L_In({
        \wRegOut_7_74[31] , \wRegOut_7_74[30] , \wRegOut_7_74[29] , 
        \wRegOut_7_74[28] , \wRegOut_7_74[27] , \wRegOut_7_74[26] , 
        \wRegOut_7_74[25] , \wRegOut_7_74[24] , \wRegOut_7_74[23] , 
        \wRegOut_7_74[22] , \wRegOut_7_74[21] , \wRegOut_7_74[20] , 
        \wRegOut_7_74[19] , \wRegOut_7_74[18] , \wRegOut_7_74[17] , 
        \wRegOut_7_74[16] , \wRegOut_7_74[15] , \wRegOut_7_74[14] , 
        \wRegOut_7_74[13] , \wRegOut_7_74[12] , \wRegOut_7_74[11] , 
        \wRegOut_7_74[10] , \wRegOut_7_74[9] , \wRegOut_7_74[8] , 
        \wRegOut_7_74[7] , \wRegOut_7_74[6] , \wRegOut_7_74[5] , 
        \wRegOut_7_74[4] , \wRegOut_7_74[3] , \wRegOut_7_74[2] , 
        \wRegOut_7_74[1] , \wRegOut_7_74[0] }), .L_Out({\wRegInTop_7_74[31] , 
        \wRegInTop_7_74[30] , \wRegInTop_7_74[29] , \wRegInTop_7_74[28] , 
        \wRegInTop_7_74[27] , \wRegInTop_7_74[26] , \wRegInTop_7_74[25] , 
        \wRegInTop_7_74[24] , \wRegInTop_7_74[23] , \wRegInTop_7_74[22] , 
        \wRegInTop_7_74[21] , \wRegInTop_7_74[20] , \wRegInTop_7_74[19] , 
        \wRegInTop_7_74[18] , \wRegInTop_7_74[17] , \wRegInTop_7_74[16] , 
        \wRegInTop_7_74[15] , \wRegInTop_7_74[14] , \wRegInTop_7_74[13] , 
        \wRegInTop_7_74[12] , \wRegInTop_7_74[11] , \wRegInTop_7_74[10] , 
        \wRegInTop_7_74[9] , \wRegInTop_7_74[8] , \wRegInTop_7_74[7] , 
        \wRegInTop_7_74[6] , \wRegInTop_7_74[5] , \wRegInTop_7_74[4] , 
        \wRegInTop_7_74[3] , \wRegInTop_7_74[2] , \wRegInTop_7_74[1] , 
        \wRegInTop_7_74[0] }), .R_WR(\wRegEnTop_7_75[0] ), .R_In({
        \wRegOut_7_75[31] , \wRegOut_7_75[30] , \wRegOut_7_75[29] , 
        \wRegOut_7_75[28] , \wRegOut_7_75[27] , \wRegOut_7_75[26] , 
        \wRegOut_7_75[25] , \wRegOut_7_75[24] , \wRegOut_7_75[23] , 
        \wRegOut_7_75[22] , \wRegOut_7_75[21] , \wRegOut_7_75[20] , 
        \wRegOut_7_75[19] , \wRegOut_7_75[18] , \wRegOut_7_75[17] , 
        \wRegOut_7_75[16] , \wRegOut_7_75[15] , \wRegOut_7_75[14] , 
        \wRegOut_7_75[13] , \wRegOut_7_75[12] , \wRegOut_7_75[11] , 
        \wRegOut_7_75[10] , \wRegOut_7_75[9] , \wRegOut_7_75[8] , 
        \wRegOut_7_75[7] , \wRegOut_7_75[6] , \wRegOut_7_75[5] , 
        \wRegOut_7_75[4] , \wRegOut_7_75[3] , \wRegOut_7_75[2] , 
        \wRegOut_7_75[1] , \wRegOut_7_75[0] }), .R_Out({\wRegInTop_7_75[31] , 
        \wRegInTop_7_75[30] , \wRegInTop_7_75[29] , \wRegInTop_7_75[28] , 
        \wRegInTop_7_75[27] , \wRegInTop_7_75[26] , \wRegInTop_7_75[25] , 
        \wRegInTop_7_75[24] , \wRegInTop_7_75[23] , \wRegInTop_7_75[22] , 
        \wRegInTop_7_75[21] , \wRegInTop_7_75[20] , \wRegInTop_7_75[19] , 
        \wRegInTop_7_75[18] , \wRegInTop_7_75[17] , \wRegInTop_7_75[16] , 
        \wRegInTop_7_75[15] , \wRegInTop_7_75[14] , \wRegInTop_7_75[13] , 
        \wRegInTop_7_75[12] , \wRegInTop_7_75[11] , \wRegInTop_7_75[10] , 
        \wRegInTop_7_75[9] , \wRegInTop_7_75[8] , \wRegInTop_7_75[7] , 
        \wRegInTop_7_75[6] , \wRegInTop_7_75[5] , \wRegInTop_7_75[4] , 
        \wRegInTop_7_75[3] , \wRegInTop_7_75[2] , \wRegInTop_7_75[1] , 
        \wRegInTop_7_75[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_1_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink2[31] , \ScanLink2[30] , \ScanLink2[29] , 
        \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , \ScanLink2[25] , 
        \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , \ScanLink2[21] , 
        \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , \ScanLink2[17] , 
        \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , \ScanLink2[13] , 
        \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , \ScanLink2[9] , 
        \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , \ScanLink2[5] , 
        \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , \ScanLink2[1] , 
        \ScanLink2[0] }), .ScanOut({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_1_0[31] , \wRegOut_1_0[30] , \wRegOut_1_0[29] , 
        \wRegOut_1_0[28] , \wRegOut_1_0[27] , \wRegOut_1_0[26] , 
        \wRegOut_1_0[25] , \wRegOut_1_0[24] , \wRegOut_1_0[23] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[21] , \wRegOut_1_0[20] , 
        \wRegOut_1_0[19] , \wRegOut_1_0[18] , \wRegOut_1_0[17] , 
        \wRegOut_1_0[16] , \wRegOut_1_0[15] , \wRegOut_1_0[14] , 
        \wRegOut_1_0[13] , \wRegOut_1_0[12] , \wRegOut_1_0[11] , 
        \wRegOut_1_0[10] , \wRegOut_1_0[9] , \wRegOut_1_0[8] , 
        \wRegOut_1_0[7] , \wRegOut_1_0[6] , \wRegOut_1_0[5] , \wRegOut_1_0[4] , 
        \wRegOut_1_0[3] , \wRegOut_1_0[2] , \wRegOut_1_0[1] , \wRegOut_1_0[0] 
        }), .Enable1(\wRegEnTop_1_0[0] ), .Enable2(\wRegEnBot_1_0[0] ), .In1({
        \wRegInTop_1_0[31] , \wRegInTop_1_0[30] , \wRegInTop_1_0[29] , 
        \wRegInTop_1_0[28] , \wRegInTop_1_0[27] , \wRegInTop_1_0[26] , 
        \wRegInTop_1_0[25] , \wRegInTop_1_0[24] , \wRegInTop_1_0[23] , 
        \wRegInTop_1_0[22] , \wRegInTop_1_0[21] , \wRegInTop_1_0[20] , 
        \wRegInTop_1_0[19] , \wRegInTop_1_0[18] , \wRegInTop_1_0[17] , 
        \wRegInTop_1_0[16] , \wRegInTop_1_0[15] , \wRegInTop_1_0[14] , 
        \wRegInTop_1_0[13] , \wRegInTop_1_0[12] , \wRegInTop_1_0[11] , 
        \wRegInTop_1_0[10] , \wRegInTop_1_0[9] , \wRegInTop_1_0[8] , 
        \wRegInTop_1_0[7] , \wRegInTop_1_0[6] , \wRegInTop_1_0[5] , 
        \wRegInTop_1_0[4] , \wRegInTop_1_0[3] , \wRegInTop_1_0[2] , 
        \wRegInTop_1_0[1] , \wRegInTop_1_0[0] }), .In2({\wRegInBot_1_0[31] , 
        \wRegInBot_1_0[30] , \wRegInBot_1_0[29] , \wRegInBot_1_0[28] , 
        \wRegInBot_1_0[27] , \wRegInBot_1_0[26] , \wRegInBot_1_0[25] , 
        \wRegInBot_1_0[24] , \wRegInBot_1_0[23] , \wRegInBot_1_0[22] , 
        \wRegInBot_1_0[21] , \wRegInBot_1_0[20] , \wRegInBot_1_0[19] , 
        \wRegInBot_1_0[18] , \wRegInBot_1_0[17] , \wRegInBot_1_0[16] , 
        \wRegInBot_1_0[15] , \wRegInBot_1_0[14] , \wRegInBot_1_0[13] , 
        \wRegInBot_1_0[12] , \wRegInBot_1_0[11] , \wRegInBot_1_0[10] , 
        \wRegInBot_1_0[9] , \wRegInBot_1_0[8] , \wRegInBot_1_0[7] , 
        \wRegInBot_1_0[6] , \wRegInBot_1_0[5] , \wRegInBot_1_0[4] , 
        \wRegInBot_1_0[3] , \wRegInBot_1_0[2] , \wRegInBot_1_0[1] , 
        \wRegInBot_1_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink22[31] , \ScanLink22[30] , \ScanLink22[29] , 
        \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , \ScanLink22[25] , 
        \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , \ScanLink22[21] , 
        \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , \ScanLink22[17] , 
        \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , \ScanLink22[13] , 
        \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , \ScanLink22[9] , 
        \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , \ScanLink22[5] , 
        \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , \ScanLink22[1] , 
        \ScanLink22[0] }), .ScanOut({\ScanLink21[31] , \ScanLink21[30] , 
        \ScanLink21[29] , \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , 
        \ScanLink21[25] , \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , 
        \ScanLink21[21] , \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , 
        \ScanLink21[17] , \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , 
        \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , 
        \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , 
        \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , 
        \ScanLink21[1] , \ScanLink21[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_6[31] , \wRegOut_4_6[30] , \wRegOut_4_6[29] , 
        \wRegOut_4_6[28] , \wRegOut_4_6[27] , \wRegOut_4_6[26] , 
        \wRegOut_4_6[25] , \wRegOut_4_6[24] , \wRegOut_4_6[23] , 
        \wRegOut_4_6[22] , \wRegOut_4_6[21] , \wRegOut_4_6[20] , 
        \wRegOut_4_6[19] , \wRegOut_4_6[18] , \wRegOut_4_6[17] , 
        \wRegOut_4_6[16] , \wRegOut_4_6[15] , \wRegOut_4_6[14] , 
        \wRegOut_4_6[13] , \wRegOut_4_6[12] , \wRegOut_4_6[11] , 
        \wRegOut_4_6[10] , \wRegOut_4_6[9] , \wRegOut_4_6[8] , 
        \wRegOut_4_6[7] , \wRegOut_4_6[6] , \wRegOut_4_6[5] , \wRegOut_4_6[4] , 
        \wRegOut_4_6[3] , \wRegOut_4_6[2] , \wRegOut_4_6[1] , \wRegOut_4_6[0] 
        }), .Enable1(\wRegEnTop_4_6[0] ), .Enable2(\wRegEnBot_4_6[0] ), .In1({
        \wRegInTop_4_6[31] , \wRegInTop_4_6[30] , \wRegInTop_4_6[29] , 
        \wRegInTop_4_6[28] , \wRegInTop_4_6[27] , \wRegInTop_4_6[26] , 
        \wRegInTop_4_6[25] , \wRegInTop_4_6[24] , \wRegInTop_4_6[23] , 
        \wRegInTop_4_6[22] , \wRegInTop_4_6[21] , \wRegInTop_4_6[20] , 
        \wRegInTop_4_6[19] , \wRegInTop_4_6[18] , \wRegInTop_4_6[17] , 
        \wRegInTop_4_6[16] , \wRegInTop_4_6[15] , \wRegInTop_4_6[14] , 
        \wRegInTop_4_6[13] , \wRegInTop_4_6[12] , \wRegInTop_4_6[11] , 
        \wRegInTop_4_6[10] , \wRegInTop_4_6[9] , \wRegInTop_4_6[8] , 
        \wRegInTop_4_6[7] , \wRegInTop_4_6[6] , \wRegInTop_4_6[5] , 
        \wRegInTop_4_6[4] , \wRegInTop_4_6[3] , \wRegInTop_4_6[2] , 
        \wRegInTop_4_6[1] , \wRegInTop_4_6[0] }), .In2({\wRegInBot_4_6[31] , 
        \wRegInBot_4_6[30] , \wRegInBot_4_6[29] , \wRegInBot_4_6[28] , 
        \wRegInBot_4_6[27] , \wRegInBot_4_6[26] , \wRegInBot_4_6[25] , 
        \wRegInBot_4_6[24] , \wRegInBot_4_6[23] , \wRegInBot_4_6[22] , 
        \wRegInBot_4_6[21] , \wRegInBot_4_6[20] , \wRegInBot_4_6[19] , 
        \wRegInBot_4_6[18] , \wRegInBot_4_6[17] , \wRegInBot_4_6[16] , 
        \wRegInBot_4_6[15] , \wRegInBot_4_6[14] , \wRegInBot_4_6[13] , 
        \wRegInBot_4_6[12] , \wRegInBot_4_6[11] , \wRegInBot_4_6[10] , 
        \wRegInBot_4_6[9] , \wRegInBot_4_6[8] , \wRegInBot_4_6[7] , 
        \wRegInBot_4_6[6] , \wRegInBot_4_6[5] , \wRegInBot_4_6[4] , 
        \wRegInBot_4_6[3] , \wRegInBot_4_6[2] , \wRegInBot_4_6[1] , 
        \wRegInBot_4_6[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink28[31] , \ScanLink28[30] , \ScanLink28[29] , 
        \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , \ScanLink28[25] , 
        \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , \ScanLink28[21] , 
        \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , \ScanLink28[17] , 
        \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , \ScanLink28[13] , 
        \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , \ScanLink28[9] , 
        \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , \ScanLink28[5] , 
        \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , \ScanLink28[1] , 
        \ScanLink28[0] }), .ScanOut({\ScanLink27[31] , \ScanLink27[30] , 
        \ScanLink27[29] , \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , 
        \ScanLink27[25] , \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , 
        \ScanLink27[21] , \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , 
        \ScanLink27[17] , \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , 
        \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , 
        \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , 
        \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , 
        \ScanLink27[1] , \ScanLink27[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_12[31] , \wRegOut_4_12[30] , 
        \wRegOut_4_12[29] , \wRegOut_4_12[28] , \wRegOut_4_12[27] , 
        \wRegOut_4_12[26] , \wRegOut_4_12[25] , \wRegOut_4_12[24] , 
        \wRegOut_4_12[23] , \wRegOut_4_12[22] , \wRegOut_4_12[21] , 
        \wRegOut_4_12[20] , \wRegOut_4_12[19] , \wRegOut_4_12[18] , 
        \wRegOut_4_12[17] , \wRegOut_4_12[16] , \wRegOut_4_12[15] , 
        \wRegOut_4_12[14] , \wRegOut_4_12[13] , \wRegOut_4_12[12] , 
        \wRegOut_4_12[11] , \wRegOut_4_12[10] , \wRegOut_4_12[9] , 
        \wRegOut_4_12[8] , \wRegOut_4_12[7] , \wRegOut_4_12[6] , 
        \wRegOut_4_12[5] , \wRegOut_4_12[4] , \wRegOut_4_12[3] , 
        \wRegOut_4_12[2] , \wRegOut_4_12[1] , \wRegOut_4_12[0] }), .Enable1(
        \wRegEnTop_4_12[0] ), .Enable2(\wRegEnBot_4_12[0] ), .In1({
        \wRegInTop_4_12[31] , \wRegInTop_4_12[30] , \wRegInTop_4_12[29] , 
        \wRegInTop_4_12[28] , \wRegInTop_4_12[27] , \wRegInTop_4_12[26] , 
        \wRegInTop_4_12[25] , \wRegInTop_4_12[24] , \wRegInTop_4_12[23] , 
        \wRegInTop_4_12[22] , \wRegInTop_4_12[21] , \wRegInTop_4_12[20] , 
        \wRegInTop_4_12[19] , \wRegInTop_4_12[18] , \wRegInTop_4_12[17] , 
        \wRegInTop_4_12[16] , \wRegInTop_4_12[15] , \wRegInTop_4_12[14] , 
        \wRegInTop_4_12[13] , \wRegInTop_4_12[12] , \wRegInTop_4_12[11] , 
        \wRegInTop_4_12[10] , \wRegInTop_4_12[9] , \wRegInTop_4_12[8] , 
        \wRegInTop_4_12[7] , \wRegInTop_4_12[6] , \wRegInTop_4_12[5] , 
        \wRegInTop_4_12[4] , \wRegInTop_4_12[3] , \wRegInTop_4_12[2] , 
        \wRegInTop_4_12[1] , \wRegInTop_4_12[0] }), .In2({\wRegInBot_4_12[31] , 
        \wRegInBot_4_12[30] , \wRegInBot_4_12[29] , \wRegInBot_4_12[28] , 
        \wRegInBot_4_12[27] , \wRegInBot_4_12[26] , \wRegInBot_4_12[25] , 
        \wRegInBot_4_12[24] , \wRegInBot_4_12[23] , \wRegInBot_4_12[22] , 
        \wRegInBot_4_12[21] , \wRegInBot_4_12[20] , \wRegInBot_4_12[19] , 
        \wRegInBot_4_12[18] , \wRegInBot_4_12[17] , \wRegInBot_4_12[16] , 
        \wRegInBot_4_12[15] , \wRegInBot_4_12[14] , \wRegInBot_4_12[13] , 
        \wRegInBot_4_12[12] , \wRegInBot_4_12[11] , \wRegInBot_4_12[10] , 
        \wRegInBot_4_12[9] , \wRegInBot_4_12[8] , \wRegInBot_4_12[7] , 
        \wRegInBot_4_12[6] , \wRegInBot_4_12[5] , \wRegInBot_4_12[4] , 
        \wRegInBot_4_12[3] , \wRegInBot_4_12[2] , \wRegInBot_4_12[1] , 
        \wRegInBot_4_12[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink38[31] , \ScanLink38[30] , \ScanLink38[29] , 
        \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , \ScanLink38[25] , 
        \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , \ScanLink38[21] , 
        \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , \ScanLink38[17] , 
        \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , \ScanLink38[13] , 
        \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , \ScanLink38[9] , 
        \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , \ScanLink38[5] , 
        \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , \ScanLink38[1] , 
        \ScanLink38[0] }), .ScanOut({\ScanLink37[31] , \ScanLink37[30] , 
        \ScanLink37[29] , \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , 
        \ScanLink37[25] , \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , 
        \ScanLink37[21] , \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , 
        \ScanLink37[17] , \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , 
        \ScanLink37[13] , \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , 
        \ScanLink37[9] , \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , 
        \ScanLink37[5] , \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , 
        \ScanLink37[1] , \ScanLink37[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_6[31] , \wRegOut_5_6[30] , \wRegOut_5_6[29] , 
        \wRegOut_5_6[28] , \wRegOut_5_6[27] , \wRegOut_5_6[26] , 
        \wRegOut_5_6[25] , \wRegOut_5_6[24] , \wRegOut_5_6[23] , 
        \wRegOut_5_6[22] , \wRegOut_5_6[21] , \wRegOut_5_6[20] , 
        \wRegOut_5_6[19] , \wRegOut_5_6[18] , \wRegOut_5_6[17] , 
        \wRegOut_5_6[16] , \wRegOut_5_6[15] , \wRegOut_5_6[14] , 
        \wRegOut_5_6[13] , \wRegOut_5_6[12] , \wRegOut_5_6[11] , 
        \wRegOut_5_6[10] , \wRegOut_5_6[9] , \wRegOut_5_6[8] , 
        \wRegOut_5_6[7] , \wRegOut_5_6[6] , \wRegOut_5_6[5] , \wRegOut_5_6[4] , 
        \wRegOut_5_6[3] , \wRegOut_5_6[2] , \wRegOut_5_6[1] , \wRegOut_5_6[0] 
        }), .Enable1(\wRegEnTop_5_6[0] ), .Enable2(\wRegEnBot_5_6[0] ), .In1({
        \wRegInTop_5_6[31] , \wRegInTop_5_6[30] , \wRegInTop_5_6[29] , 
        \wRegInTop_5_6[28] , \wRegInTop_5_6[27] , \wRegInTop_5_6[26] , 
        \wRegInTop_5_6[25] , \wRegInTop_5_6[24] , \wRegInTop_5_6[23] , 
        \wRegInTop_5_6[22] , \wRegInTop_5_6[21] , \wRegInTop_5_6[20] , 
        \wRegInTop_5_6[19] , \wRegInTop_5_6[18] , \wRegInTop_5_6[17] , 
        \wRegInTop_5_6[16] , \wRegInTop_5_6[15] , \wRegInTop_5_6[14] , 
        \wRegInTop_5_6[13] , \wRegInTop_5_6[12] , \wRegInTop_5_6[11] , 
        \wRegInTop_5_6[10] , \wRegInTop_5_6[9] , \wRegInTop_5_6[8] , 
        \wRegInTop_5_6[7] , \wRegInTop_5_6[6] , \wRegInTop_5_6[5] , 
        \wRegInTop_5_6[4] , \wRegInTop_5_6[3] , \wRegInTop_5_6[2] , 
        \wRegInTop_5_6[1] , \wRegInTop_5_6[0] }), .In2({\wRegInBot_5_6[31] , 
        \wRegInBot_5_6[30] , \wRegInBot_5_6[29] , \wRegInBot_5_6[28] , 
        \wRegInBot_5_6[27] , \wRegInBot_5_6[26] , \wRegInBot_5_6[25] , 
        \wRegInBot_5_6[24] , \wRegInBot_5_6[23] , \wRegInBot_5_6[22] , 
        \wRegInBot_5_6[21] , \wRegInBot_5_6[20] , \wRegInBot_5_6[19] , 
        \wRegInBot_5_6[18] , \wRegInBot_5_6[17] , \wRegInBot_5_6[16] , 
        \wRegInBot_5_6[15] , \wRegInBot_5_6[14] , \wRegInBot_5_6[13] , 
        \wRegInBot_5_6[12] , \wRegInBot_5_6[11] , \wRegInBot_5_6[10] , 
        \wRegInBot_5_6[9] , \wRegInBot_5_6[8] , \wRegInBot_5_6[7] , 
        \wRegInBot_5_6[6] , \wRegInBot_5_6[5] , \wRegInBot_5_6[4] , 
        \wRegInBot_5_6[3] , \wRegInBot_5_6[2] , \wRegInBot_5_6[1] , 
        \wRegInBot_5_6[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_22 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink150[31] , \ScanLink150[30] , \ScanLink150[29] , 
        \ScanLink150[28] , \ScanLink150[27] , \ScanLink150[26] , 
        \ScanLink150[25] , \ScanLink150[24] , \ScanLink150[23] , 
        \ScanLink150[22] , \ScanLink150[21] , \ScanLink150[20] , 
        \ScanLink150[19] , \ScanLink150[18] , \ScanLink150[17] , 
        \ScanLink150[16] , \ScanLink150[15] , \ScanLink150[14] , 
        \ScanLink150[13] , \ScanLink150[12] , \ScanLink150[11] , 
        \ScanLink150[10] , \ScanLink150[9] , \ScanLink150[8] , 
        \ScanLink150[7] , \ScanLink150[6] , \ScanLink150[5] , \ScanLink150[4] , 
        \ScanLink150[3] , \ScanLink150[2] , \ScanLink150[1] , \ScanLink150[0] 
        }), .ScanOut({\ScanLink149[31] , \ScanLink149[30] , \ScanLink149[29] , 
        \ScanLink149[28] , \ScanLink149[27] , \ScanLink149[26] , 
        \ScanLink149[25] , \ScanLink149[24] , \ScanLink149[23] , 
        \ScanLink149[22] , \ScanLink149[21] , \ScanLink149[20] , 
        \ScanLink149[19] , \ScanLink149[18] , \ScanLink149[17] , 
        \ScanLink149[16] , \ScanLink149[15] , \ScanLink149[14] , 
        \ScanLink149[13] , \ScanLink149[12] , \ScanLink149[11] , 
        \ScanLink149[10] , \ScanLink149[9] , \ScanLink149[8] , 
        \ScanLink149[7] , \ScanLink149[6] , \ScanLink149[5] , \ScanLink149[4] , 
        \ScanLink149[3] , \ScanLink149[2] , \ScanLink149[1] , \ScanLink149[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_22[31] , 
        \wRegOut_7_22[30] , \wRegOut_7_22[29] , \wRegOut_7_22[28] , 
        \wRegOut_7_22[27] , \wRegOut_7_22[26] , \wRegOut_7_22[25] , 
        \wRegOut_7_22[24] , \wRegOut_7_22[23] , \wRegOut_7_22[22] , 
        \wRegOut_7_22[21] , \wRegOut_7_22[20] , \wRegOut_7_22[19] , 
        \wRegOut_7_22[18] , \wRegOut_7_22[17] , \wRegOut_7_22[16] , 
        \wRegOut_7_22[15] , \wRegOut_7_22[14] , \wRegOut_7_22[13] , 
        \wRegOut_7_22[12] , \wRegOut_7_22[11] , \wRegOut_7_22[10] , 
        \wRegOut_7_22[9] , \wRegOut_7_22[8] , \wRegOut_7_22[7] , 
        \wRegOut_7_22[6] , \wRegOut_7_22[5] , \wRegOut_7_22[4] , 
        \wRegOut_7_22[3] , \wRegOut_7_22[2] , \wRegOut_7_22[1] , 
        \wRegOut_7_22[0] }), .Enable1(\wRegEnTop_7_22[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_22[31] , \wRegInTop_7_22[30] , \wRegInTop_7_22[29] , 
        \wRegInTop_7_22[28] , \wRegInTop_7_22[27] , \wRegInTop_7_22[26] , 
        \wRegInTop_7_22[25] , \wRegInTop_7_22[24] , \wRegInTop_7_22[23] , 
        \wRegInTop_7_22[22] , \wRegInTop_7_22[21] , \wRegInTop_7_22[20] , 
        \wRegInTop_7_22[19] , \wRegInTop_7_22[18] , \wRegInTop_7_22[17] , 
        \wRegInTop_7_22[16] , \wRegInTop_7_22[15] , \wRegInTop_7_22[14] , 
        \wRegInTop_7_22[13] , \wRegInTop_7_22[12] , \wRegInTop_7_22[11] , 
        \wRegInTop_7_22[10] , \wRegInTop_7_22[9] , \wRegInTop_7_22[8] , 
        \wRegInTop_7_22[7] , \wRegInTop_7_22[6] , \wRegInTop_7_22[5] , 
        \wRegInTop_7_22[4] , \wRegInTop_7_22[3] , \wRegInTop_7_22[2] , 
        \wRegInTop_7_22[1] , \wRegInTop_7_22[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_111 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink239[31] , \ScanLink239[30] , \ScanLink239[29] , 
        \ScanLink239[28] , \ScanLink239[27] , \ScanLink239[26] , 
        \ScanLink239[25] , \ScanLink239[24] , \ScanLink239[23] , 
        \ScanLink239[22] , \ScanLink239[21] , \ScanLink239[20] , 
        \ScanLink239[19] , \ScanLink239[18] , \ScanLink239[17] , 
        \ScanLink239[16] , \ScanLink239[15] , \ScanLink239[14] , 
        \ScanLink239[13] , \ScanLink239[12] , \ScanLink239[11] , 
        \ScanLink239[10] , \ScanLink239[9] , \ScanLink239[8] , 
        \ScanLink239[7] , \ScanLink239[6] , \ScanLink239[5] , \ScanLink239[4] , 
        \ScanLink239[3] , \ScanLink239[2] , \ScanLink239[1] , \ScanLink239[0] 
        }), .ScanOut({\ScanLink238[31] , \ScanLink238[30] , \ScanLink238[29] , 
        \ScanLink238[28] , \ScanLink238[27] , \ScanLink238[26] , 
        \ScanLink238[25] , \ScanLink238[24] , \ScanLink238[23] , 
        \ScanLink238[22] , \ScanLink238[21] , \ScanLink238[20] , 
        \ScanLink238[19] , \ScanLink238[18] , \ScanLink238[17] , 
        \ScanLink238[16] , \ScanLink238[15] , \ScanLink238[14] , 
        \ScanLink238[13] , \ScanLink238[12] , \ScanLink238[11] , 
        \ScanLink238[10] , \ScanLink238[9] , \ScanLink238[8] , 
        \ScanLink238[7] , \ScanLink238[6] , \ScanLink238[5] , \ScanLink238[4] , 
        \ScanLink238[3] , \ScanLink238[2] , \ScanLink238[1] , \ScanLink238[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_111[31] , 
        \wRegOut_7_111[30] , \wRegOut_7_111[29] , \wRegOut_7_111[28] , 
        \wRegOut_7_111[27] , \wRegOut_7_111[26] , \wRegOut_7_111[25] , 
        \wRegOut_7_111[24] , \wRegOut_7_111[23] , \wRegOut_7_111[22] , 
        \wRegOut_7_111[21] , \wRegOut_7_111[20] , \wRegOut_7_111[19] , 
        \wRegOut_7_111[18] , \wRegOut_7_111[17] , \wRegOut_7_111[16] , 
        \wRegOut_7_111[15] , \wRegOut_7_111[14] , \wRegOut_7_111[13] , 
        \wRegOut_7_111[12] , \wRegOut_7_111[11] , \wRegOut_7_111[10] , 
        \wRegOut_7_111[9] , \wRegOut_7_111[8] , \wRegOut_7_111[7] , 
        \wRegOut_7_111[6] , \wRegOut_7_111[5] , \wRegOut_7_111[4] , 
        \wRegOut_7_111[3] , \wRegOut_7_111[2] , \wRegOut_7_111[1] , 
        \wRegOut_7_111[0] }), .Enable1(\wRegEnTop_7_111[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_111[31] , \wRegInTop_7_111[30] , 
        \wRegInTop_7_111[29] , \wRegInTop_7_111[28] , \wRegInTop_7_111[27] , 
        \wRegInTop_7_111[26] , \wRegInTop_7_111[25] , \wRegInTop_7_111[24] , 
        \wRegInTop_7_111[23] , \wRegInTop_7_111[22] , \wRegInTop_7_111[21] , 
        \wRegInTop_7_111[20] , \wRegInTop_7_111[19] , \wRegInTop_7_111[18] , 
        \wRegInTop_7_111[17] , \wRegInTop_7_111[16] , \wRegInTop_7_111[15] , 
        \wRegInTop_7_111[14] , \wRegInTop_7_111[13] , \wRegInTop_7_111[12] , 
        \wRegInTop_7_111[11] , \wRegInTop_7_111[10] , \wRegInTop_7_111[9] , 
        \wRegInTop_7_111[8] , \wRegInTop_7_111[7] , \wRegInTop_7_111[6] , 
        \wRegInTop_7_111[5] , \wRegInTop_7_111[4] , \wRegInTop_7_111[3] , 
        \wRegInTop_7_111[2] , \wRegInTop_7_111[1] , \wRegInTop_7_111[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_4[0] ), .P_In({\wRegOut_4_4[31] , 
        \wRegOut_4_4[30] , \wRegOut_4_4[29] , \wRegOut_4_4[28] , 
        \wRegOut_4_4[27] , \wRegOut_4_4[26] , \wRegOut_4_4[25] , 
        \wRegOut_4_4[24] , \wRegOut_4_4[23] , \wRegOut_4_4[22] , 
        \wRegOut_4_4[21] , \wRegOut_4_4[20] , \wRegOut_4_4[19] , 
        \wRegOut_4_4[18] , \wRegOut_4_4[17] , \wRegOut_4_4[16] , 
        \wRegOut_4_4[15] , \wRegOut_4_4[14] , \wRegOut_4_4[13] , 
        \wRegOut_4_4[12] , \wRegOut_4_4[11] , \wRegOut_4_4[10] , 
        \wRegOut_4_4[9] , \wRegOut_4_4[8] , \wRegOut_4_4[7] , \wRegOut_4_4[6] , 
        \wRegOut_4_4[5] , \wRegOut_4_4[4] , \wRegOut_4_4[3] , \wRegOut_4_4[2] , 
        \wRegOut_4_4[1] , \wRegOut_4_4[0] }), .P_Out({\wRegInBot_4_4[31] , 
        \wRegInBot_4_4[30] , \wRegInBot_4_4[29] , \wRegInBot_4_4[28] , 
        \wRegInBot_4_4[27] , \wRegInBot_4_4[26] , \wRegInBot_4_4[25] , 
        \wRegInBot_4_4[24] , \wRegInBot_4_4[23] , \wRegInBot_4_4[22] , 
        \wRegInBot_4_4[21] , \wRegInBot_4_4[20] , \wRegInBot_4_4[19] , 
        \wRegInBot_4_4[18] , \wRegInBot_4_4[17] , \wRegInBot_4_4[16] , 
        \wRegInBot_4_4[15] , \wRegInBot_4_4[14] , \wRegInBot_4_4[13] , 
        \wRegInBot_4_4[12] , \wRegInBot_4_4[11] , \wRegInBot_4_4[10] , 
        \wRegInBot_4_4[9] , \wRegInBot_4_4[8] , \wRegInBot_4_4[7] , 
        \wRegInBot_4_4[6] , \wRegInBot_4_4[5] , \wRegInBot_4_4[4] , 
        \wRegInBot_4_4[3] , \wRegInBot_4_4[2] , \wRegInBot_4_4[1] , 
        \wRegInBot_4_4[0] }), .L_WR(\wRegEnTop_5_8[0] ), .L_In({
        \wRegOut_5_8[31] , \wRegOut_5_8[30] , \wRegOut_5_8[29] , 
        \wRegOut_5_8[28] , \wRegOut_5_8[27] , \wRegOut_5_8[26] , 
        \wRegOut_5_8[25] , \wRegOut_5_8[24] , \wRegOut_5_8[23] , 
        \wRegOut_5_8[22] , \wRegOut_5_8[21] , \wRegOut_5_8[20] , 
        \wRegOut_5_8[19] , \wRegOut_5_8[18] , \wRegOut_5_8[17] , 
        \wRegOut_5_8[16] , \wRegOut_5_8[15] , \wRegOut_5_8[14] , 
        \wRegOut_5_8[13] , \wRegOut_5_8[12] , \wRegOut_5_8[11] , 
        \wRegOut_5_8[10] , \wRegOut_5_8[9] , \wRegOut_5_8[8] , 
        \wRegOut_5_8[7] , \wRegOut_5_8[6] , \wRegOut_5_8[5] , \wRegOut_5_8[4] , 
        \wRegOut_5_8[3] , \wRegOut_5_8[2] , \wRegOut_5_8[1] , \wRegOut_5_8[0] 
        }), .L_Out({\wRegInTop_5_8[31] , \wRegInTop_5_8[30] , 
        \wRegInTop_5_8[29] , \wRegInTop_5_8[28] , \wRegInTop_5_8[27] , 
        \wRegInTop_5_8[26] , \wRegInTop_5_8[25] , \wRegInTop_5_8[24] , 
        \wRegInTop_5_8[23] , \wRegInTop_5_8[22] , \wRegInTop_5_8[21] , 
        \wRegInTop_5_8[20] , \wRegInTop_5_8[19] , \wRegInTop_5_8[18] , 
        \wRegInTop_5_8[17] , \wRegInTop_5_8[16] , \wRegInTop_5_8[15] , 
        \wRegInTop_5_8[14] , \wRegInTop_5_8[13] , \wRegInTop_5_8[12] , 
        \wRegInTop_5_8[11] , \wRegInTop_5_8[10] , \wRegInTop_5_8[9] , 
        \wRegInTop_5_8[8] , \wRegInTop_5_8[7] , \wRegInTop_5_8[6] , 
        \wRegInTop_5_8[5] , \wRegInTop_5_8[4] , \wRegInTop_5_8[3] , 
        \wRegInTop_5_8[2] , \wRegInTop_5_8[1] , \wRegInTop_5_8[0] }), .R_WR(
        \wRegEnTop_5_9[0] ), .R_In({\wRegOut_5_9[31] , \wRegOut_5_9[30] , 
        \wRegOut_5_9[29] , \wRegOut_5_9[28] , \wRegOut_5_9[27] , 
        \wRegOut_5_9[26] , \wRegOut_5_9[25] , \wRegOut_5_9[24] , 
        \wRegOut_5_9[23] , \wRegOut_5_9[22] , \wRegOut_5_9[21] , 
        \wRegOut_5_9[20] , \wRegOut_5_9[19] , \wRegOut_5_9[18] , 
        \wRegOut_5_9[17] , \wRegOut_5_9[16] , \wRegOut_5_9[15] , 
        \wRegOut_5_9[14] , \wRegOut_5_9[13] , \wRegOut_5_9[12] , 
        \wRegOut_5_9[11] , \wRegOut_5_9[10] , \wRegOut_5_9[9] , 
        \wRegOut_5_9[8] , \wRegOut_5_9[7] , \wRegOut_5_9[6] , \wRegOut_5_9[5] , 
        \wRegOut_5_9[4] , \wRegOut_5_9[3] , \wRegOut_5_9[2] , \wRegOut_5_9[1] , 
        \wRegOut_5_9[0] }), .R_Out({\wRegInTop_5_9[31] , \wRegInTop_5_9[30] , 
        \wRegInTop_5_9[29] , \wRegInTop_5_9[28] , \wRegInTop_5_9[27] , 
        \wRegInTop_5_9[26] , \wRegInTop_5_9[25] , \wRegInTop_5_9[24] , 
        \wRegInTop_5_9[23] , \wRegInTop_5_9[22] , \wRegInTop_5_9[21] , 
        \wRegInTop_5_9[20] , \wRegInTop_5_9[19] , \wRegInTop_5_9[18] , 
        \wRegInTop_5_9[17] , \wRegInTop_5_9[16] , \wRegInTop_5_9[15] , 
        \wRegInTop_5_9[14] , \wRegInTop_5_9[13] , \wRegInTop_5_9[12] , 
        \wRegInTop_5_9[11] , \wRegInTop_5_9[10] , \wRegInTop_5_9[9] , 
        \wRegInTop_5_9[8] , \wRegInTop_5_9[7] , \wRegInTop_5_9[6] , 
        \wRegInTop_5_9[5] , \wRegInTop_5_9[4] , \wRegInTop_5_9[3] , 
        \wRegInTop_5_9[2] , \wRegInTop_5_9[1] , \wRegInTop_5_9[0] }) );
    BHeap_Node_WIDTH32 BHN_6_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_8[0] ), .P_In({\wRegOut_6_8[31] , 
        \wRegOut_6_8[30] , \wRegOut_6_8[29] , \wRegOut_6_8[28] , 
        \wRegOut_6_8[27] , \wRegOut_6_8[26] , \wRegOut_6_8[25] , 
        \wRegOut_6_8[24] , \wRegOut_6_8[23] , \wRegOut_6_8[22] , 
        \wRegOut_6_8[21] , \wRegOut_6_8[20] , \wRegOut_6_8[19] , 
        \wRegOut_6_8[18] , \wRegOut_6_8[17] , \wRegOut_6_8[16] , 
        \wRegOut_6_8[15] , \wRegOut_6_8[14] , \wRegOut_6_8[13] , 
        \wRegOut_6_8[12] , \wRegOut_6_8[11] , \wRegOut_6_8[10] , 
        \wRegOut_6_8[9] , \wRegOut_6_8[8] , \wRegOut_6_8[7] , \wRegOut_6_8[6] , 
        \wRegOut_6_8[5] , \wRegOut_6_8[4] , \wRegOut_6_8[3] , \wRegOut_6_8[2] , 
        \wRegOut_6_8[1] , \wRegOut_6_8[0] }), .P_Out({\wRegInBot_6_8[31] , 
        \wRegInBot_6_8[30] , \wRegInBot_6_8[29] , \wRegInBot_6_8[28] , 
        \wRegInBot_6_8[27] , \wRegInBot_6_8[26] , \wRegInBot_6_8[25] , 
        \wRegInBot_6_8[24] , \wRegInBot_6_8[23] , \wRegInBot_6_8[22] , 
        \wRegInBot_6_8[21] , \wRegInBot_6_8[20] , \wRegInBot_6_8[19] , 
        \wRegInBot_6_8[18] , \wRegInBot_6_8[17] , \wRegInBot_6_8[16] , 
        \wRegInBot_6_8[15] , \wRegInBot_6_8[14] , \wRegInBot_6_8[13] , 
        \wRegInBot_6_8[12] , \wRegInBot_6_8[11] , \wRegInBot_6_8[10] , 
        \wRegInBot_6_8[9] , \wRegInBot_6_8[8] , \wRegInBot_6_8[7] , 
        \wRegInBot_6_8[6] , \wRegInBot_6_8[5] , \wRegInBot_6_8[4] , 
        \wRegInBot_6_8[3] , \wRegInBot_6_8[2] , \wRegInBot_6_8[1] , 
        \wRegInBot_6_8[0] }), .L_WR(\wRegEnTop_7_16[0] ), .L_In({
        \wRegOut_7_16[31] , \wRegOut_7_16[30] , \wRegOut_7_16[29] , 
        \wRegOut_7_16[28] , \wRegOut_7_16[27] , \wRegOut_7_16[26] , 
        \wRegOut_7_16[25] , \wRegOut_7_16[24] , \wRegOut_7_16[23] , 
        \wRegOut_7_16[22] , \wRegOut_7_16[21] , \wRegOut_7_16[20] , 
        \wRegOut_7_16[19] , \wRegOut_7_16[18] , \wRegOut_7_16[17] , 
        \wRegOut_7_16[16] , \wRegOut_7_16[15] , \wRegOut_7_16[14] , 
        \wRegOut_7_16[13] , \wRegOut_7_16[12] , \wRegOut_7_16[11] , 
        \wRegOut_7_16[10] , \wRegOut_7_16[9] , \wRegOut_7_16[8] , 
        \wRegOut_7_16[7] , \wRegOut_7_16[6] , \wRegOut_7_16[5] , 
        \wRegOut_7_16[4] , \wRegOut_7_16[3] , \wRegOut_7_16[2] , 
        \wRegOut_7_16[1] , \wRegOut_7_16[0] }), .L_Out({\wRegInTop_7_16[31] , 
        \wRegInTop_7_16[30] , \wRegInTop_7_16[29] , \wRegInTop_7_16[28] , 
        \wRegInTop_7_16[27] , \wRegInTop_7_16[26] , \wRegInTop_7_16[25] , 
        \wRegInTop_7_16[24] , \wRegInTop_7_16[23] , \wRegInTop_7_16[22] , 
        \wRegInTop_7_16[21] , \wRegInTop_7_16[20] , \wRegInTop_7_16[19] , 
        \wRegInTop_7_16[18] , \wRegInTop_7_16[17] , \wRegInTop_7_16[16] , 
        \wRegInTop_7_16[15] , \wRegInTop_7_16[14] , \wRegInTop_7_16[13] , 
        \wRegInTop_7_16[12] , \wRegInTop_7_16[11] , \wRegInTop_7_16[10] , 
        \wRegInTop_7_16[9] , \wRegInTop_7_16[8] , \wRegInTop_7_16[7] , 
        \wRegInTop_7_16[6] , \wRegInTop_7_16[5] , \wRegInTop_7_16[4] , 
        \wRegInTop_7_16[3] , \wRegInTop_7_16[2] , \wRegInTop_7_16[1] , 
        \wRegInTop_7_16[0] }), .R_WR(\wRegEnTop_7_17[0] ), .R_In({
        \wRegOut_7_17[31] , \wRegOut_7_17[30] , \wRegOut_7_17[29] , 
        \wRegOut_7_17[28] , \wRegOut_7_17[27] , \wRegOut_7_17[26] , 
        \wRegOut_7_17[25] , \wRegOut_7_17[24] , \wRegOut_7_17[23] , 
        \wRegOut_7_17[22] , \wRegOut_7_17[21] , \wRegOut_7_17[20] , 
        \wRegOut_7_17[19] , \wRegOut_7_17[18] , \wRegOut_7_17[17] , 
        \wRegOut_7_17[16] , \wRegOut_7_17[15] , \wRegOut_7_17[14] , 
        \wRegOut_7_17[13] , \wRegOut_7_17[12] , \wRegOut_7_17[11] , 
        \wRegOut_7_17[10] , \wRegOut_7_17[9] , \wRegOut_7_17[8] , 
        \wRegOut_7_17[7] , \wRegOut_7_17[6] , \wRegOut_7_17[5] , 
        \wRegOut_7_17[4] , \wRegOut_7_17[3] , \wRegOut_7_17[2] , 
        \wRegOut_7_17[1] , \wRegOut_7_17[0] }), .R_Out({\wRegInTop_7_17[31] , 
        \wRegInTop_7_17[30] , \wRegInTop_7_17[29] , \wRegInTop_7_17[28] , 
        \wRegInTop_7_17[27] , \wRegInTop_7_17[26] , \wRegInTop_7_17[25] , 
        \wRegInTop_7_17[24] , \wRegInTop_7_17[23] , \wRegInTop_7_17[22] , 
        \wRegInTop_7_17[21] , \wRegInTop_7_17[20] , \wRegInTop_7_17[19] , 
        \wRegInTop_7_17[18] , \wRegInTop_7_17[17] , \wRegInTop_7_17[16] , 
        \wRegInTop_7_17[15] , \wRegInTop_7_17[14] , \wRegInTop_7_17[13] , 
        \wRegInTop_7_17[12] , \wRegInTop_7_17[11] , \wRegInTop_7_17[10] , 
        \wRegInTop_7_17[9] , \wRegInTop_7_17[8] , \wRegInTop_7_17[7] , 
        \wRegInTop_7_17[6] , \wRegInTop_7_17[5] , \wRegInTop_7_17[4] , 
        \wRegInTop_7_17[3] , \wRegInTop_7_17[2] , \wRegInTop_7_17[1] , 
        \wRegInTop_7_17[0] }) );
    BHeap_Node_WIDTH32 BHN_6_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_59[0] ), .P_In({\wRegOut_6_59[31] , 
        \wRegOut_6_59[30] , \wRegOut_6_59[29] , \wRegOut_6_59[28] , 
        \wRegOut_6_59[27] , \wRegOut_6_59[26] , \wRegOut_6_59[25] , 
        \wRegOut_6_59[24] , \wRegOut_6_59[23] , \wRegOut_6_59[22] , 
        \wRegOut_6_59[21] , \wRegOut_6_59[20] , \wRegOut_6_59[19] , 
        \wRegOut_6_59[18] , \wRegOut_6_59[17] , \wRegOut_6_59[16] , 
        \wRegOut_6_59[15] , \wRegOut_6_59[14] , \wRegOut_6_59[13] , 
        \wRegOut_6_59[12] , \wRegOut_6_59[11] , \wRegOut_6_59[10] , 
        \wRegOut_6_59[9] , \wRegOut_6_59[8] , \wRegOut_6_59[7] , 
        \wRegOut_6_59[6] , \wRegOut_6_59[5] , \wRegOut_6_59[4] , 
        \wRegOut_6_59[3] , \wRegOut_6_59[2] , \wRegOut_6_59[1] , 
        \wRegOut_6_59[0] }), .P_Out({\wRegInBot_6_59[31] , 
        \wRegInBot_6_59[30] , \wRegInBot_6_59[29] , \wRegInBot_6_59[28] , 
        \wRegInBot_6_59[27] , \wRegInBot_6_59[26] , \wRegInBot_6_59[25] , 
        \wRegInBot_6_59[24] , \wRegInBot_6_59[23] , \wRegInBot_6_59[22] , 
        \wRegInBot_6_59[21] , \wRegInBot_6_59[20] , \wRegInBot_6_59[19] , 
        \wRegInBot_6_59[18] , \wRegInBot_6_59[17] , \wRegInBot_6_59[16] , 
        \wRegInBot_6_59[15] , \wRegInBot_6_59[14] , \wRegInBot_6_59[13] , 
        \wRegInBot_6_59[12] , \wRegInBot_6_59[11] , \wRegInBot_6_59[10] , 
        \wRegInBot_6_59[9] , \wRegInBot_6_59[8] , \wRegInBot_6_59[7] , 
        \wRegInBot_6_59[6] , \wRegInBot_6_59[5] , \wRegInBot_6_59[4] , 
        \wRegInBot_6_59[3] , \wRegInBot_6_59[2] , \wRegInBot_6_59[1] , 
        \wRegInBot_6_59[0] }), .L_WR(\wRegEnTop_7_118[0] ), .L_In({
        \wRegOut_7_118[31] , \wRegOut_7_118[30] , \wRegOut_7_118[29] , 
        \wRegOut_7_118[28] , \wRegOut_7_118[27] , \wRegOut_7_118[26] , 
        \wRegOut_7_118[25] , \wRegOut_7_118[24] , \wRegOut_7_118[23] , 
        \wRegOut_7_118[22] , \wRegOut_7_118[21] , \wRegOut_7_118[20] , 
        \wRegOut_7_118[19] , \wRegOut_7_118[18] , \wRegOut_7_118[17] , 
        \wRegOut_7_118[16] , \wRegOut_7_118[15] , \wRegOut_7_118[14] , 
        \wRegOut_7_118[13] , \wRegOut_7_118[12] , \wRegOut_7_118[11] , 
        \wRegOut_7_118[10] , \wRegOut_7_118[9] , \wRegOut_7_118[8] , 
        \wRegOut_7_118[7] , \wRegOut_7_118[6] , \wRegOut_7_118[5] , 
        \wRegOut_7_118[4] , \wRegOut_7_118[3] , \wRegOut_7_118[2] , 
        \wRegOut_7_118[1] , \wRegOut_7_118[0] }), .L_Out({
        \wRegInTop_7_118[31] , \wRegInTop_7_118[30] , \wRegInTop_7_118[29] , 
        \wRegInTop_7_118[28] , \wRegInTop_7_118[27] , \wRegInTop_7_118[26] , 
        \wRegInTop_7_118[25] , \wRegInTop_7_118[24] , \wRegInTop_7_118[23] , 
        \wRegInTop_7_118[22] , \wRegInTop_7_118[21] , \wRegInTop_7_118[20] , 
        \wRegInTop_7_118[19] , \wRegInTop_7_118[18] , \wRegInTop_7_118[17] , 
        \wRegInTop_7_118[16] , \wRegInTop_7_118[15] , \wRegInTop_7_118[14] , 
        \wRegInTop_7_118[13] , \wRegInTop_7_118[12] , \wRegInTop_7_118[11] , 
        \wRegInTop_7_118[10] , \wRegInTop_7_118[9] , \wRegInTop_7_118[8] , 
        \wRegInTop_7_118[7] , \wRegInTop_7_118[6] , \wRegInTop_7_118[5] , 
        \wRegInTop_7_118[4] , \wRegInTop_7_118[3] , \wRegInTop_7_118[2] , 
        \wRegInTop_7_118[1] , \wRegInTop_7_118[0] }), .R_WR(
        \wRegEnTop_7_119[0] ), .R_In({\wRegOut_7_119[31] , \wRegOut_7_119[30] , 
        \wRegOut_7_119[29] , \wRegOut_7_119[28] , \wRegOut_7_119[27] , 
        \wRegOut_7_119[26] , \wRegOut_7_119[25] , \wRegOut_7_119[24] , 
        \wRegOut_7_119[23] , \wRegOut_7_119[22] , \wRegOut_7_119[21] , 
        \wRegOut_7_119[20] , \wRegOut_7_119[19] , \wRegOut_7_119[18] , 
        \wRegOut_7_119[17] , \wRegOut_7_119[16] , \wRegOut_7_119[15] , 
        \wRegOut_7_119[14] , \wRegOut_7_119[13] , \wRegOut_7_119[12] , 
        \wRegOut_7_119[11] , \wRegOut_7_119[10] , \wRegOut_7_119[9] , 
        \wRegOut_7_119[8] , \wRegOut_7_119[7] , \wRegOut_7_119[6] , 
        \wRegOut_7_119[5] , \wRegOut_7_119[4] , \wRegOut_7_119[3] , 
        \wRegOut_7_119[2] , \wRegOut_7_119[1] , \wRegOut_7_119[0] }), .R_Out({
        \wRegInTop_7_119[31] , \wRegInTop_7_119[30] , \wRegInTop_7_119[29] , 
        \wRegInTop_7_119[28] , \wRegInTop_7_119[27] , \wRegInTop_7_119[26] , 
        \wRegInTop_7_119[25] , \wRegInTop_7_119[24] , \wRegInTop_7_119[23] , 
        \wRegInTop_7_119[22] , \wRegInTop_7_119[21] , \wRegInTop_7_119[20] , 
        \wRegInTop_7_119[19] , \wRegInTop_7_119[18] , \wRegInTop_7_119[17] , 
        \wRegInTop_7_119[16] , \wRegInTop_7_119[15] , \wRegInTop_7_119[14] , 
        \wRegInTop_7_119[13] , \wRegInTop_7_119[12] , \wRegInTop_7_119[11] , 
        \wRegInTop_7_119[10] , \wRegInTop_7_119[9] , \wRegInTop_7_119[8] , 
        \wRegInTop_7_119[7] , \wRegInTop_7_119[6] , \wRegInTop_7_119[5] , 
        \wRegInTop_7_119[4] , \wRegInTop_7_119[3] , \wRegInTop_7_119[2] , 
        \wRegInTop_7_119[1] , \wRegInTop_7_119[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_56 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink120[31] , \ScanLink120[30] , \ScanLink120[29] , 
        \ScanLink120[28] , \ScanLink120[27] , \ScanLink120[26] , 
        \ScanLink120[25] , \ScanLink120[24] , \ScanLink120[23] , 
        \ScanLink120[22] , \ScanLink120[21] , \ScanLink120[20] , 
        \ScanLink120[19] , \ScanLink120[18] , \ScanLink120[17] , 
        \ScanLink120[16] , \ScanLink120[15] , \ScanLink120[14] , 
        \ScanLink120[13] , \ScanLink120[12] , \ScanLink120[11] , 
        \ScanLink120[10] , \ScanLink120[9] , \ScanLink120[8] , 
        \ScanLink120[7] , \ScanLink120[6] , \ScanLink120[5] , \ScanLink120[4] , 
        \ScanLink120[3] , \ScanLink120[2] , \ScanLink120[1] , \ScanLink120[0] 
        }), .ScanOut({\ScanLink119[31] , \ScanLink119[30] , \ScanLink119[29] , 
        \ScanLink119[28] , \ScanLink119[27] , \ScanLink119[26] , 
        \ScanLink119[25] , \ScanLink119[24] , \ScanLink119[23] , 
        \ScanLink119[22] , \ScanLink119[21] , \ScanLink119[20] , 
        \ScanLink119[19] , \ScanLink119[18] , \ScanLink119[17] , 
        \ScanLink119[16] , \ScanLink119[15] , \ScanLink119[14] , 
        \ScanLink119[13] , \ScanLink119[12] , \ScanLink119[11] , 
        \ScanLink119[10] , \ScanLink119[9] , \ScanLink119[8] , 
        \ScanLink119[7] , \ScanLink119[6] , \ScanLink119[5] , \ScanLink119[4] , 
        \ScanLink119[3] , \ScanLink119[2] , \ScanLink119[1] , \ScanLink119[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_56[31] , 
        \wRegOut_6_56[30] , \wRegOut_6_56[29] , \wRegOut_6_56[28] , 
        \wRegOut_6_56[27] , \wRegOut_6_56[26] , \wRegOut_6_56[25] , 
        \wRegOut_6_56[24] , \wRegOut_6_56[23] , \wRegOut_6_56[22] , 
        \wRegOut_6_56[21] , \wRegOut_6_56[20] , \wRegOut_6_56[19] , 
        \wRegOut_6_56[18] , \wRegOut_6_56[17] , \wRegOut_6_56[16] , 
        \wRegOut_6_56[15] , \wRegOut_6_56[14] , \wRegOut_6_56[13] , 
        \wRegOut_6_56[12] , \wRegOut_6_56[11] , \wRegOut_6_56[10] , 
        \wRegOut_6_56[9] , \wRegOut_6_56[8] , \wRegOut_6_56[7] , 
        \wRegOut_6_56[6] , \wRegOut_6_56[5] , \wRegOut_6_56[4] , 
        \wRegOut_6_56[3] , \wRegOut_6_56[2] , \wRegOut_6_56[1] , 
        \wRegOut_6_56[0] }), .Enable1(\wRegEnTop_6_56[0] ), .Enable2(
        \wRegEnBot_6_56[0] ), .In1({\wRegInTop_6_56[31] , \wRegInTop_6_56[30] , 
        \wRegInTop_6_56[29] , \wRegInTop_6_56[28] , \wRegInTop_6_56[27] , 
        \wRegInTop_6_56[26] , \wRegInTop_6_56[25] , \wRegInTop_6_56[24] , 
        \wRegInTop_6_56[23] , \wRegInTop_6_56[22] , \wRegInTop_6_56[21] , 
        \wRegInTop_6_56[20] , \wRegInTop_6_56[19] , \wRegInTop_6_56[18] , 
        \wRegInTop_6_56[17] , \wRegInTop_6_56[16] , \wRegInTop_6_56[15] , 
        \wRegInTop_6_56[14] , \wRegInTop_6_56[13] , \wRegInTop_6_56[12] , 
        \wRegInTop_6_56[11] , \wRegInTop_6_56[10] , \wRegInTop_6_56[9] , 
        \wRegInTop_6_56[8] , \wRegInTop_6_56[7] , \wRegInTop_6_56[6] , 
        \wRegInTop_6_56[5] , \wRegInTop_6_56[4] , \wRegInTop_6_56[3] , 
        \wRegInTop_6_56[2] , \wRegInTop_6_56[1] , \wRegInTop_6_56[0] }), .In2(
        {\wRegInBot_6_56[31] , \wRegInBot_6_56[30] , \wRegInBot_6_56[29] , 
        \wRegInBot_6_56[28] , \wRegInBot_6_56[27] , \wRegInBot_6_56[26] , 
        \wRegInBot_6_56[25] , \wRegInBot_6_56[24] , \wRegInBot_6_56[23] , 
        \wRegInBot_6_56[22] , \wRegInBot_6_56[21] , \wRegInBot_6_56[20] , 
        \wRegInBot_6_56[19] , \wRegInBot_6_56[18] , \wRegInBot_6_56[17] , 
        \wRegInBot_6_56[16] , \wRegInBot_6_56[15] , \wRegInBot_6_56[14] , 
        \wRegInBot_6_56[13] , \wRegInBot_6_56[12] , \wRegInBot_6_56[11] , 
        \wRegInBot_6_56[10] , \wRegInBot_6_56[9] , \wRegInBot_6_56[8] , 
        \wRegInBot_6_56[7] , \wRegInBot_6_56[6] , \wRegInBot_6_56[5] , 
        \wRegInBot_6_56[4] , \wRegInBot_6_56[3] , \wRegInBot_6_56[2] , 
        \wRegInBot_6_56[1] , \wRegInBot_6_56[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_39 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink167[31] , \ScanLink167[30] , \ScanLink167[29] , 
        \ScanLink167[28] , \ScanLink167[27] , \ScanLink167[26] , 
        \ScanLink167[25] , \ScanLink167[24] , \ScanLink167[23] , 
        \ScanLink167[22] , \ScanLink167[21] , \ScanLink167[20] , 
        \ScanLink167[19] , \ScanLink167[18] , \ScanLink167[17] , 
        \ScanLink167[16] , \ScanLink167[15] , \ScanLink167[14] , 
        \ScanLink167[13] , \ScanLink167[12] , \ScanLink167[11] , 
        \ScanLink167[10] , \ScanLink167[9] , \ScanLink167[8] , 
        \ScanLink167[7] , \ScanLink167[6] , \ScanLink167[5] , \ScanLink167[4] , 
        \ScanLink167[3] , \ScanLink167[2] , \ScanLink167[1] , \ScanLink167[0] 
        }), .ScanOut({\ScanLink166[31] , \ScanLink166[30] , \ScanLink166[29] , 
        \ScanLink166[28] , \ScanLink166[27] , \ScanLink166[26] , 
        \ScanLink166[25] , \ScanLink166[24] , \ScanLink166[23] , 
        \ScanLink166[22] , \ScanLink166[21] , \ScanLink166[20] , 
        \ScanLink166[19] , \ScanLink166[18] , \ScanLink166[17] , 
        \ScanLink166[16] , \ScanLink166[15] , \ScanLink166[14] , 
        \ScanLink166[13] , \ScanLink166[12] , \ScanLink166[11] , 
        \ScanLink166[10] , \ScanLink166[9] , \ScanLink166[8] , 
        \ScanLink166[7] , \ScanLink166[6] , \ScanLink166[5] , \ScanLink166[4] , 
        \ScanLink166[3] , \ScanLink166[2] , \ScanLink166[1] , \ScanLink166[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_39[31] , 
        \wRegOut_7_39[30] , \wRegOut_7_39[29] , \wRegOut_7_39[28] , 
        \wRegOut_7_39[27] , \wRegOut_7_39[26] , \wRegOut_7_39[25] , 
        \wRegOut_7_39[24] , \wRegOut_7_39[23] , \wRegOut_7_39[22] , 
        \wRegOut_7_39[21] , \wRegOut_7_39[20] , \wRegOut_7_39[19] , 
        \wRegOut_7_39[18] , \wRegOut_7_39[17] , \wRegOut_7_39[16] , 
        \wRegOut_7_39[15] , \wRegOut_7_39[14] , \wRegOut_7_39[13] , 
        \wRegOut_7_39[12] , \wRegOut_7_39[11] , \wRegOut_7_39[10] , 
        \wRegOut_7_39[9] , \wRegOut_7_39[8] , \wRegOut_7_39[7] , 
        \wRegOut_7_39[6] , \wRegOut_7_39[5] , \wRegOut_7_39[4] , 
        \wRegOut_7_39[3] , \wRegOut_7_39[2] , \wRegOut_7_39[1] , 
        \wRegOut_7_39[0] }), .Enable1(\wRegEnTop_7_39[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_39[31] , \wRegInTop_7_39[30] , \wRegInTop_7_39[29] , 
        \wRegInTop_7_39[28] , \wRegInTop_7_39[27] , \wRegInTop_7_39[26] , 
        \wRegInTop_7_39[25] , \wRegInTop_7_39[24] , \wRegInTop_7_39[23] , 
        \wRegInTop_7_39[22] , \wRegInTop_7_39[21] , \wRegInTop_7_39[20] , 
        \wRegInTop_7_39[19] , \wRegInTop_7_39[18] , \wRegInTop_7_39[17] , 
        \wRegInTop_7_39[16] , \wRegInTop_7_39[15] , \wRegInTop_7_39[14] , 
        \wRegInTop_7_39[13] , \wRegInTop_7_39[12] , \wRegInTop_7_39[11] , 
        \wRegInTop_7_39[10] , \wRegInTop_7_39[9] , \wRegInTop_7_39[8] , 
        \wRegInTop_7_39[7] , \wRegInTop_7_39[6] , \wRegInTop_7_39[5] , 
        \wRegInTop_7_39[4] , \wRegInTop_7_39[3] , \wRegInTop_7_39[2] , 
        \wRegInTop_7_39[1] , \wRegInTop_7_39[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_70 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink198[31] , \ScanLink198[30] , \ScanLink198[29] , 
        \ScanLink198[28] , \ScanLink198[27] , \ScanLink198[26] , 
        \ScanLink198[25] , \ScanLink198[24] , \ScanLink198[23] , 
        \ScanLink198[22] , \ScanLink198[21] , \ScanLink198[20] , 
        \ScanLink198[19] , \ScanLink198[18] , \ScanLink198[17] , 
        \ScanLink198[16] , \ScanLink198[15] , \ScanLink198[14] , 
        \ScanLink198[13] , \ScanLink198[12] , \ScanLink198[11] , 
        \ScanLink198[10] , \ScanLink198[9] , \ScanLink198[8] , 
        \ScanLink198[7] , \ScanLink198[6] , \ScanLink198[5] , \ScanLink198[4] , 
        \ScanLink198[3] , \ScanLink198[2] , \ScanLink198[1] , \ScanLink198[0] 
        }), .ScanOut({\ScanLink197[31] , \ScanLink197[30] , \ScanLink197[29] , 
        \ScanLink197[28] , \ScanLink197[27] , \ScanLink197[26] , 
        \ScanLink197[25] , \ScanLink197[24] , \ScanLink197[23] , 
        \ScanLink197[22] , \ScanLink197[21] , \ScanLink197[20] , 
        \ScanLink197[19] , \ScanLink197[18] , \ScanLink197[17] , 
        \ScanLink197[16] , \ScanLink197[15] , \ScanLink197[14] , 
        \ScanLink197[13] , \ScanLink197[12] , \ScanLink197[11] , 
        \ScanLink197[10] , \ScanLink197[9] , \ScanLink197[8] , 
        \ScanLink197[7] , \ScanLink197[6] , \ScanLink197[5] , \ScanLink197[4] , 
        \ScanLink197[3] , \ScanLink197[2] , \ScanLink197[1] , \ScanLink197[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_70[31] , 
        \wRegOut_7_70[30] , \wRegOut_7_70[29] , \wRegOut_7_70[28] , 
        \wRegOut_7_70[27] , \wRegOut_7_70[26] , \wRegOut_7_70[25] , 
        \wRegOut_7_70[24] , \wRegOut_7_70[23] , \wRegOut_7_70[22] , 
        \wRegOut_7_70[21] , \wRegOut_7_70[20] , \wRegOut_7_70[19] , 
        \wRegOut_7_70[18] , \wRegOut_7_70[17] , \wRegOut_7_70[16] , 
        \wRegOut_7_70[15] , \wRegOut_7_70[14] , \wRegOut_7_70[13] , 
        \wRegOut_7_70[12] , \wRegOut_7_70[11] , \wRegOut_7_70[10] , 
        \wRegOut_7_70[9] , \wRegOut_7_70[8] , \wRegOut_7_70[7] , 
        \wRegOut_7_70[6] , \wRegOut_7_70[5] , \wRegOut_7_70[4] , 
        \wRegOut_7_70[3] , \wRegOut_7_70[2] , \wRegOut_7_70[1] , 
        \wRegOut_7_70[0] }), .Enable1(\wRegEnTop_7_70[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_70[31] , \wRegInTop_7_70[30] , \wRegInTop_7_70[29] , 
        \wRegInTop_7_70[28] , \wRegInTop_7_70[27] , \wRegInTop_7_70[26] , 
        \wRegInTop_7_70[25] , \wRegInTop_7_70[24] , \wRegInTop_7_70[23] , 
        \wRegInTop_7_70[22] , \wRegInTop_7_70[21] , \wRegInTop_7_70[20] , 
        \wRegInTop_7_70[19] , \wRegInTop_7_70[18] , \wRegInTop_7_70[17] , 
        \wRegInTop_7_70[16] , \wRegInTop_7_70[15] , \wRegInTop_7_70[14] , 
        \wRegInTop_7_70[13] , \wRegInTop_7_70[12] , \wRegInTop_7_70[11] , 
        \wRegInTop_7_70[10] , \wRegInTop_7_70[9] , \wRegInTop_7_70[8] , 
        \wRegInTop_7_70[7] , \wRegInTop_7_70[6] , \wRegInTop_7_70[5] , 
        \wRegInTop_7_70[4] , \wRegInTop_7_70[3] , \wRegInTop_7_70[2] , 
        \wRegInTop_7_70[1] , \wRegInTop_7_70[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_95 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink223[31] , \ScanLink223[30] , \ScanLink223[29] , 
        \ScanLink223[28] , \ScanLink223[27] , \ScanLink223[26] , 
        \ScanLink223[25] , \ScanLink223[24] , \ScanLink223[23] , 
        \ScanLink223[22] , \ScanLink223[21] , \ScanLink223[20] , 
        \ScanLink223[19] , \ScanLink223[18] , \ScanLink223[17] , 
        \ScanLink223[16] , \ScanLink223[15] , \ScanLink223[14] , 
        \ScanLink223[13] , \ScanLink223[12] , \ScanLink223[11] , 
        \ScanLink223[10] , \ScanLink223[9] , \ScanLink223[8] , 
        \ScanLink223[7] , \ScanLink223[6] , \ScanLink223[5] , \ScanLink223[4] , 
        \ScanLink223[3] , \ScanLink223[2] , \ScanLink223[1] , \ScanLink223[0] 
        }), .ScanOut({\ScanLink222[31] , \ScanLink222[30] , \ScanLink222[29] , 
        \ScanLink222[28] , \ScanLink222[27] , \ScanLink222[26] , 
        \ScanLink222[25] , \ScanLink222[24] , \ScanLink222[23] , 
        \ScanLink222[22] , \ScanLink222[21] , \ScanLink222[20] , 
        \ScanLink222[19] , \ScanLink222[18] , \ScanLink222[17] , 
        \ScanLink222[16] , \ScanLink222[15] , \ScanLink222[14] , 
        \ScanLink222[13] , \ScanLink222[12] , \ScanLink222[11] , 
        \ScanLink222[10] , \ScanLink222[9] , \ScanLink222[8] , 
        \ScanLink222[7] , \ScanLink222[6] , \ScanLink222[5] , \ScanLink222[4] , 
        \ScanLink222[3] , \ScanLink222[2] , \ScanLink222[1] , \ScanLink222[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_95[31] , 
        \wRegOut_7_95[30] , \wRegOut_7_95[29] , \wRegOut_7_95[28] , 
        \wRegOut_7_95[27] , \wRegOut_7_95[26] , \wRegOut_7_95[25] , 
        \wRegOut_7_95[24] , \wRegOut_7_95[23] , \wRegOut_7_95[22] , 
        \wRegOut_7_95[21] , \wRegOut_7_95[20] , \wRegOut_7_95[19] , 
        \wRegOut_7_95[18] , \wRegOut_7_95[17] , \wRegOut_7_95[16] , 
        \wRegOut_7_95[15] , \wRegOut_7_95[14] , \wRegOut_7_95[13] , 
        \wRegOut_7_95[12] , \wRegOut_7_95[11] , \wRegOut_7_95[10] , 
        \wRegOut_7_95[9] , \wRegOut_7_95[8] , \wRegOut_7_95[7] , 
        \wRegOut_7_95[6] , \wRegOut_7_95[5] , \wRegOut_7_95[4] , 
        \wRegOut_7_95[3] , \wRegOut_7_95[2] , \wRegOut_7_95[1] , 
        \wRegOut_7_95[0] }), .Enable1(\wRegEnTop_7_95[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_95[31] , \wRegInTop_7_95[30] , \wRegInTop_7_95[29] , 
        \wRegInTop_7_95[28] , \wRegInTop_7_95[27] , \wRegInTop_7_95[26] , 
        \wRegInTop_7_95[25] , \wRegInTop_7_95[24] , \wRegInTop_7_95[23] , 
        \wRegInTop_7_95[22] , \wRegInTop_7_95[21] , \wRegInTop_7_95[20] , 
        \wRegInTop_7_95[19] , \wRegInTop_7_95[18] , \wRegInTop_7_95[17] , 
        \wRegInTop_7_95[16] , \wRegInTop_7_95[15] , \wRegInTop_7_95[14] , 
        \wRegInTop_7_95[13] , \wRegInTop_7_95[12] , \wRegInTop_7_95[11] , 
        \wRegInTop_7_95[10] , \wRegInTop_7_95[9] , \wRegInTop_7_95[8] , 
        \wRegInTop_7_95[7] , \wRegInTop_7_95[6] , \wRegInTop_7_95[5] , 
        \wRegInTop_7_95[4] , \wRegInTop_7_95[3] , \wRegInTop_7_95[2] , 
        \wRegInTop_7_95[1] , \wRegInTop_7_95[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_42[0] ), .P_In({\wRegOut_6_42[31] , 
        \wRegOut_6_42[30] , \wRegOut_6_42[29] , \wRegOut_6_42[28] , 
        \wRegOut_6_42[27] , \wRegOut_6_42[26] , \wRegOut_6_42[25] , 
        \wRegOut_6_42[24] , \wRegOut_6_42[23] , \wRegOut_6_42[22] , 
        \wRegOut_6_42[21] , \wRegOut_6_42[20] , \wRegOut_6_42[19] , 
        \wRegOut_6_42[18] , \wRegOut_6_42[17] , \wRegOut_6_42[16] , 
        \wRegOut_6_42[15] , \wRegOut_6_42[14] , \wRegOut_6_42[13] , 
        \wRegOut_6_42[12] , \wRegOut_6_42[11] , \wRegOut_6_42[10] , 
        \wRegOut_6_42[9] , \wRegOut_6_42[8] , \wRegOut_6_42[7] , 
        \wRegOut_6_42[6] , \wRegOut_6_42[5] , \wRegOut_6_42[4] , 
        \wRegOut_6_42[3] , \wRegOut_6_42[2] , \wRegOut_6_42[1] , 
        \wRegOut_6_42[0] }), .P_Out({\wRegInBot_6_42[31] , 
        \wRegInBot_6_42[30] , \wRegInBot_6_42[29] , \wRegInBot_6_42[28] , 
        \wRegInBot_6_42[27] , \wRegInBot_6_42[26] , \wRegInBot_6_42[25] , 
        \wRegInBot_6_42[24] , \wRegInBot_6_42[23] , \wRegInBot_6_42[22] , 
        \wRegInBot_6_42[21] , \wRegInBot_6_42[20] , \wRegInBot_6_42[19] , 
        \wRegInBot_6_42[18] , \wRegInBot_6_42[17] , \wRegInBot_6_42[16] , 
        \wRegInBot_6_42[15] , \wRegInBot_6_42[14] , \wRegInBot_6_42[13] , 
        \wRegInBot_6_42[12] , \wRegInBot_6_42[11] , \wRegInBot_6_42[10] , 
        \wRegInBot_6_42[9] , \wRegInBot_6_42[8] , \wRegInBot_6_42[7] , 
        \wRegInBot_6_42[6] , \wRegInBot_6_42[5] , \wRegInBot_6_42[4] , 
        \wRegInBot_6_42[3] , \wRegInBot_6_42[2] , \wRegInBot_6_42[1] , 
        \wRegInBot_6_42[0] }), .L_WR(\wRegEnTop_7_84[0] ), .L_In({
        \wRegOut_7_84[31] , \wRegOut_7_84[30] , \wRegOut_7_84[29] , 
        \wRegOut_7_84[28] , \wRegOut_7_84[27] , \wRegOut_7_84[26] , 
        \wRegOut_7_84[25] , \wRegOut_7_84[24] , \wRegOut_7_84[23] , 
        \wRegOut_7_84[22] , \wRegOut_7_84[21] , \wRegOut_7_84[20] , 
        \wRegOut_7_84[19] , \wRegOut_7_84[18] , \wRegOut_7_84[17] , 
        \wRegOut_7_84[16] , \wRegOut_7_84[15] , \wRegOut_7_84[14] , 
        \wRegOut_7_84[13] , \wRegOut_7_84[12] , \wRegOut_7_84[11] , 
        \wRegOut_7_84[10] , \wRegOut_7_84[9] , \wRegOut_7_84[8] , 
        \wRegOut_7_84[7] , \wRegOut_7_84[6] , \wRegOut_7_84[5] , 
        \wRegOut_7_84[4] , \wRegOut_7_84[3] , \wRegOut_7_84[2] , 
        \wRegOut_7_84[1] , \wRegOut_7_84[0] }), .L_Out({\wRegInTop_7_84[31] , 
        \wRegInTop_7_84[30] , \wRegInTop_7_84[29] , \wRegInTop_7_84[28] , 
        \wRegInTop_7_84[27] , \wRegInTop_7_84[26] , \wRegInTop_7_84[25] , 
        \wRegInTop_7_84[24] , \wRegInTop_7_84[23] , \wRegInTop_7_84[22] , 
        \wRegInTop_7_84[21] , \wRegInTop_7_84[20] , \wRegInTop_7_84[19] , 
        \wRegInTop_7_84[18] , \wRegInTop_7_84[17] , \wRegInTop_7_84[16] , 
        \wRegInTop_7_84[15] , \wRegInTop_7_84[14] , \wRegInTop_7_84[13] , 
        \wRegInTop_7_84[12] , \wRegInTop_7_84[11] , \wRegInTop_7_84[10] , 
        \wRegInTop_7_84[9] , \wRegInTop_7_84[8] , \wRegInTop_7_84[7] , 
        \wRegInTop_7_84[6] , \wRegInTop_7_84[5] , \wRegInTop_7_84[4] , 
        \wRegInTop_7_84[3] , \wRegInTop_7_84[2] , \wRegInTop_7_84[1] , 
        \wRegInTop_7_84[0] }), .R_WR(\wRegEnTop_7_85[0] ), .R_In({
        \wRegOut_7_85[31] , \wRegOut_7_85[30] , \wRegOut_7_85[29] , 
        \wRegOut_7_85[28] , \wRegOut_7_85[27] , \wRegOut_7_85[26] , 
        \wRegOut_7_85[25] , \wRegOut_7_85[24] , \wRegOut_7_85[23] , 
        \wRegOut_7_85[22] , \wRegOut_7_85[21] , \wRegOut_7_85[20] , 
        \wRegOut_7_85[19] , \wRegOut_7_85[18] , \wRegOut_7_85[17] , 
        \wRegOut_7_85[16] , \wRegOut_7_85[15] , \wRegOut_7_85[14] , 
        \wRegOut_7_85[13] , \wRegOut_7_85[12] , \wRegOut_7_85[11] , 
        \wRegOut_7_85[10] , \wRegOut_7_85[9] , \wRegOut_7_85[8] , 
        \wRegOut_7_85[7] , \wRegOut_7_85[6] , \wRegOut_7_85[5] , 
        \wRegOut_7_85[4] , \wRegOut_7_85[3] , \wRegOut_7_85[2] , 
        \wRegOut_7_85[1] , \wRegOut_7_85[0] }), .R_Out({\wRegInTop_7_85[31] , 
        \wRegInTop_7_85[30] , \wRegInTop_7_85[29] , \wRegInTop_7_85[28] , 
        \wRegInTop_7_85[27] , \wRegInTop_7_85[26] , \wRegInTop_7_85[25] , 
        \wRegInTop_7_85[24] , \wRegInTop_7_85[23] , \wRegInTop_7_85[22] , 
        \wRegInTop_7_85[21] , \wRegInTop_7_85[20] , \wRegInTop_7_85[19] , 
        \wRegInTop_7_85[18] , \wRegInTop_7_85[17] , \wRegInTop_7_85[16] , 
        \wRegInTop_7_85[15] , \wRegInTop_7_85[14] , \wRegInTop_7_85[13] , 
        \wRegInTop_7_85[12] , \wRegInTop_7_85[11] , \wRegInTop_7_85[10] , 
        \wRegInTop_7_85[9] , \wRegInTop_7_85[8] , \wRegInTop_7_85[7] , 
        \wRegInTop_7_85[6] , \wRegInTop_7_85[5] , \wRegInTop_7_85[4] , 
        \wRegInTop_7_85[3] , \wRegInTop_7_85[2] , \wRegInTop_7_85[1] , 
        \wRegInTop_7_85[0] }) );
    BHeap_Node_WIDTH32 BHN_5_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_4[0] ), .P_In({\wRegOut_5_4[31] , 
        \wRegOut_5_4[30] , \wRegOut_5_4[29] , \wRegOut_5_4[28] , 
        \wRegOut_5_4[27] , \wRegOut_5_4[26] , \wRegOut_5_4[25] , 
        \wRegOut_5_4[24] , \wRegOut_5_4[23] , \wRegOut_5_4[22] , 
        \wRegOut_5_4[21] , \wRegOut_5_4[20] , \wRegOut_5_4[19] , 
        \wRegOut_5_4[18] , \wRegOut_5_4[17] , \wRegOut_5_4[16] , 
        \wRegOut_5_4[15] , \wRegOut_5_4[14] , \wRegOut_5_4[13] , 
        \wRegOut_5_4[12] , \wRegOut_5_4[11] , \wRegOut_5_4[10] , 
        \wRegOut_5_4[9] , \wRegOut_5_4[8] , \wRegOut_5_4[7] , \wRegOut_5_4[6] , 
        \wRegOut_5_4[5] , \wRegOut_5_4[4] , \wRegOut_5_4[3] , \wRegOut_5_4[2] , 
        \wRegOut_5_4[1] , \wRegOut_5_4[0] }), .P_Out({\wRegInBot_5_4[31] , 
        \wRegInBot_5_4[30] , \wRegInBot_5_4[29] , \wRegInBot_5_4[28] , 
        \wRegInBot_5_4[27] , \wRegInBot_5_4[26] , \wRegInBot_5_4[25] , 
        \wRegInBot_5_4[24] , \wRegInBot_5_4[23] , \wRegInBot_5_4[22] , 
        \wRegInBot_5_4[21] , \wRegInBot_5_4[20] , \wRegInBot_5_4[19] , 
        \wRegInBot_5_4[18] , \wRegInBot_5_4[17] , \wRegInBot_5_4[16] , 
        \wRegInBot_5_4[15] , \wRegInBot_5_4[14] , \wRegInBot_5_4[13] , 
        \wRegInBot_5_4[12] , \wRegInBot_5_4[11] , \wRegInBot_5_4[10] , 
        \wRegInBot_5_4[9] , \wRegInBot_5_4[8] , \wRegInBot_5_4[7] , 
        \wRegInBot_5_4[6] , \wRegInBot_5_4[5] , \wRegInBot_5_4[4] , 
        \wRegInBot_5_4[3] , \wRegInBot_5_4[2] , \wRegInBot_5_4[1] , 
        \wRegInBot_5_4[0] }), .L_WR(\wRegEnTop_6_8[0] ), .L_In({
        \wRegOut_6_8[31] , \wRegOut_6_8[30] , \wRegOut_6_8[29] , 
        \wRegOut_6_8[28] , \wRegOut_6_8[27] , \wRegOut_6_8[26] , 
        \wRegOut_6_8[25] , \wRegOut_6_8[24] , \wRegOut_6_8[23] , 
        \wRegOut_6_8[22] , \wRegOut_6_8[21] , \wRegOut_6_8[20] , 
        \wRegOut_6_8[19] , \wRegOut_6_8[18] , \wRegOut_6_8[17] , 
        \wRegOut_6_8[16] , \wRegOut_6_8[15] , \wRegOut_6_8[14] , 
        \wRegOut_6_8[13] , \wRegOut_6_8[12] , \wRegOut_6_8[11] , 
        \wRegOut_6_8[10] , \wRegOut_6_8[9] , \wRegOut_6_8[8] , 
        \wRegOut_6_8[7] , \wRegOut_6_8[6] , \wRegOut_6_8[5] , \wRegOut_6_8[4] , 
        \wRegOut_6_8[3] , \wRegOut_6_8[2] , \wRegOut_6_8[1] , \wRegOut_6_8[0] 
        }), .L_Out({\wRegInTop_6_8[31] , \wRegInTop_6_8[30] , 
        \wRegInTop_6_8[29] , \wRegInTop_6_8[28] , \wRegInTop_6_8[27] , 
        \wRegInTop_6_8[26] , \wRegInTop_6_8[25] , \wRegInTop_6_8[24] , 
        \wRegInTop_6_8[23] , \wRegInTop_6_8[22] , \wRegInTop_6_8[21] , 
        \wRegInTop_6_8[20] , \wRegInTop_6_8[19] , \wRegInTop_6_8[18] , 
        \wRegInTop_6_8[17] , \wRegInTop_6_8[16] , \wRegInTop_6_8[15] , 
        \wRegInTop_6_8[14] , \wRegInTop_6_8[13] , \wRegInTop_6_8[12] , 
        \wRegInTop_6_8[11] , \wRegInTop_6_8[10] , \wRegInTop_6_8[9] , 
        \wRegInTop_6_8[8] , \wRegInTop_6_8[7] , \wRegInTop_6_8[6] , 
        \wRegInTop_6_8[5] , \wRegInTop_6_8[4] , \wRegInTop_6_8[3] , 
        \wRegInTop_6_8[2] , \wRegInTop_6_8[1] , \wRegInTop_6_8[0] }), .R_WR(
        \wRegEnTop_6_9[0] ), .R_In({\wRegOut_6_9[31] , \wRegOut_6_9[30] , 
        \wRegOut_6_9[29] , \wRegOut_6_9[28] , \wRegOut_6_9[27] , 
        \wRegOut_6_9[26] , \wRegOut_6_9[25] , \wRegOut_6_9[24] , 
        \wRegOut_6_9[23] , \wRegOut_6_9[22] , \wRegOut_6_9[21] , 
        \wRegOut_6_9[20] , \wRegOut_6_9[19] , \wRegOut_6_9[18] , 
        \wRegOut_6_9[17] , \wRegOut_6_9[16] , \wRegOut_6_9[15] , 
        \wRegOut_6_9[14] , \wRegOut_6_9[13] , \wRegOut_6_9[12] , 
        \wRegOut_6_9[11] , \wRegOut_6_9[10] , \wRegOut_6_9[9] , 
        \wRegOut_6_9[8] , \wRegOut_6_9[7] , \wRegOut_6_9[6] , \wRegOut_6_9[5] , 
        \wRegOut_6_9[4] , \wRegOut_6_9[3] , \wRegOut_6_9[2] , \wRegOut_6_9[1] , 
        \wRegOut_6_9[0] }), .R_Out({\wRegInTop_6_9[31] , \wRegInTop_6_9[30] , 
        \wRegInTop_6_9[29] , \wRegInTop_6_9[28] , \wRegInTop_6_9[27] , 
        \wRegInTop_6_9[26] , \wRegInTop_6_9[25] , \wRegInTop_6_9[24] , 
        \wRegInTop_6_9[23] , \wRegInTop_6_9[22] , \wRegInTop_6_9[21] , 
        \wRegInTop_6_9[20] , \wRegInTop_6_9[19] , \wRegInTop_6_9[18] , 
        \wRegInTop_6_9[17] , \wRegInTop_6_9[16] , \wRegInTop_6_9[15] , 
        \wRegInTop_6_9[14] , \wRegInTop_6_9[13] , \wRegInTop_6_9[12] , 
        \wRegInTop_6_9[11] , \wRegInTop_6_9[10] , \wRegInTop_6_9[9] , 
        \wRegInTop_6_9[8] , \wRegInTop_6_9[7] , \wRegInTop_6_9[6] , 
        \wRegInTop_6_9[5] , \wRegInTop_6_9[4] , \wRegInTop_6_9[3] , 
        \wRegInTop_6_9[2] , \wRegInTop_6_9[1] , \wRegInTop_6_9[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink45[31] , \ScanLink45[30] , \ScanLink45[29] , 
        \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , \ScanLink45[25] , 
        \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , \ScanLink45[21] , 
        \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , \ScanLink45[17] , 
        \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , \ScanLink45[13] , 
        \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , \ScanLink45[9] , 
        \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , \ScanLink45[5] , 
        \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , \ScanLink45[1] , 
        \ScanLink45[0] }), .ScanOut({\ScanLink44[31] , \ScanLink44[30] , 
        \ScanLink44[29] , \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , 
        \ScanLink44[25] , \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , 
        \ScanLink44[21] , \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , 
        \ScanLink44[17] , \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , 
        \ScanLink44[13] , \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , 
        \ScanLink44[9] , \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , 
        \ScanLink44[5] , \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , 
        \ScanLink44[1] , \ScanLink44[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_13[31] , \wRegOut_5_13[30] , 
        \wRegOut_5_13[29] , \wRegOut_5_13[28] , \wRegOut_5_13[27] , 
        \wRegOut_5_13[26] , \wRegOut_5_13[25] , \wRegOut_5_13[24] , 
        \wRegOut_5_13[23] , \wRegOut_5_13[22] , \wRegOut_5_13[21] , 
        \wRegOut_5_13[20] , \wRegOut_5_13[19] , \wRegOut_5_13[18] , 
        \wRegOut_5_13[17] , \wRegOut_5_13[16] , \wRegOut_5_13[15] , 
        \wRegOut_5_13[14] , \wRegOut_5_13[13] , \wRegOut_5_13[12] , 
        \wRegOut_5_13[11] , \wRegOut_5_13[10] , \wRegOut_5_13[9] , 
        \wRegOut_5_13[8] , \wRegOut_5_13[7] , \wRegOut_5_13[6] , 
        \wRegOut_5_13[5] , \wRegOut_5_13[4] , \wRegOut_5_13[3] , 
        \wRegOut_5_13[2] , \wRegOut_5_13[1] , \wRegOut_5_13[0] }), .Enable1(
        \wRegEnTop_5_13[0] ), .Enable2(\wRegEnBot_5_13[0] ), .In1({
        \wRegInTop_5_13[31] , \wRegInTop_5_13[30] , \wRegInTop_5_13[29] , 
        \wRegInTop_5_13[28] , \wRegInTop_5_13[27] , \wRegInTop_5_13[26] , 
        \wRegInTop_5_13[25] , \wRegInTop_5_13[24] , \wRegInTop_5_13[23] , 
        \wRegInTop_5_13[22] , \wRegInTop_5_13[21] , \wRegInTop_5_13[20] , 
        \wRegInTop_5_13[19] , \wRegInTop_5_13[18] , \wRegInTop_5_13[17] , 
        \wRegInTop_5_13[16] , \wRegInTop_5_13[15] , \wRegInTop_5_13[14] , 
        \wRegInTop_5_13[13] , \wRegInTop_5_13[12] , \wRegInTop_5_13[11] , 
        \wRegInTop_5_13[10] , \wRegInTop_5_13[9] , \wRegInTop_5_13[8] , 
        \wRegInTop_5_13[7] , \wRegInTop_5_13[6] , \wRegInTop_5_13[5] , 
        \wRegInTop_5_13[4] , \wRegInTop_5_13[3] , \wRegInTop_5_13[2] , 
        \wRegInTop_5_13[1] , \wRegInTop_5_13[0] }), .In2({\wRegInBot_5_13[31] , 
        \wRegInBot_5_13[30] , \wRegInBot_5_13[29] , \wRegInBot_5_13[28] , 
        \wRegInBot_5_13[27] , \wRegInBot_5_13[26] , \wRegInBot_5_13[25] , 
        \wRegInBot_5_13[24] , \wRegInBot_5_13[23] , \wRegInBot_5_13[22] , 
        \wRegInBot_5_13[21] , \wRegInBot_5_13[20] , \wRegInBot_5_13[19] , 
        \wRegInBot_5_13[18] , \wRegInBot_5_13[17] , \wRegInBot_5_13[16] , 
        \wRegInBot_5_13[15] , \wRegInBot_5_13[14] , \wRegInBot_5_13[13] , 
        \wRegInBot_5_13[12] , \wRegInBot_5_13[11] , \wRegInBot_5_13[10] , 
        \wRegInBot_5_13[9] , \wRegInBot_5_13[8] , \wRegInBot_5_13[7] , 
        \wRegInBot_5_13[6] , \wRegInBot_5_13[5] , \wRegInBot_5_13[4] , 
        \wRegInBot_5_13[3] , \wRegInBot_5_13[2] , \wRegInBot_5_13[1] , 
        \wRegInBot_5_13[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_23 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink87[31] , \ScanLink87[30] , \ScanLink87[29] , 
        \ScanLink87[28] , \ScanLink87[27] , \ScanLink87[26] , \ScanLink87[25] , 
        \ScanLink87[24] , \ScanLink87[23] , \ScanLink87[22] , \ScanLink87[21] , 
        \ScanLink87[20] , \ScanLink87[19] , \ScanLink87[18] , \ScanLink87[17] , 
        \ScanLink87[16] , \ScanLink87[15] , \ScanLink87[14] , \ScanLink87[13] , 
        \ScanLink87[12] , \ScanLink87[11] , \ScanLink87[10] , \ScanLink87[9] , 
        \ScanLink87[8] , \ScanLink87[7] , \ScanLink87[6] , \ScanLink87[5] , 
        \ScanLink87[4] , \ScanLink87[3] , \ScanLink87[2] , \ScanLink87[1] , 
        \ScanLink87[0] }), .ScanOut({\ScanLink86[31] , \ScanLink86[30] , 
        \ScanLink86[29] , \ScanLink86[28] , \ScanLink86[27] , \ScanLink86[26] , 
        \ScanLink86[25] , \ScanLink86[24] , \ScanLink86[23] , \ScanLink86[22] , 
        \ScanLink86[21] , \ScanLink86[20] , \ScanLink86[19] , \ScanLink86[18] , 
        \ScanLink86[17] , \ScanLink86[16] , \ScanLink86[15] , \ScanLink86[14] , 
        \ScanLink86[13] , \ScanLink86[12] , \ScanLink86[11] , \ScanLink86[10] , 
        \ScanLink86[9] , \ScanLink86[8] , \ScanLink86[7] , \ScanLink86[6] , 
        \ScanLink86[5] , \ScanLink86[4] , \ScanLink86[3] , \ScanLink86[2] , 
        \ScanLink86[1] , \ScanLink86[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_23[31] , \wRegOut_6_23[30] , 
        \wRegOut_6_23[29] , \wRegOut_6_23[28] , \wRegOut_6_23[27] , 
        \wRegOut_6_23[26] , \wRegOut_6_23[25] , \wRegOut_6_23[24] , 
        \wRegOut_6_23[23] , \wRegOut_6_23[22] , \wRegOut_6_23[21] , 
        \wRegOut_6_23[20] , \wRegOut_6_23[19] , \wRegOut_6_23[18] , 
        \wRegOut_6_23[17] , \wRegOut_6_23[16] , \wRegOut_6_23[15] , 
        \wRegOut_6_23[14] , \wRegOut_6_23[13] , \wRegOut_6_23[12] , 
        \wRegOut_6_23[11] , \wRegOut_6_23[10] , \wRegOut_6_23[9] , 
        \wRegOut_6_23[8] , \wRegOut_6_23[7] , \wRegOut_6_23[6] , 
        \wRegOut_6_23[5] , \wRegOut_6_23[4] , \wRegOut_6_23[3] , 
        \wRegOut_6_23[2] , \wRegOut_6_23[1] , \wRegOut_6_23[0] }), .Enable1(
        \wRegEnTop_6_23[0] ), .Enable2(\wRegEnBot_6_23[0] ), .In1({
        \wRegInTop_6_23[31] , \wRegInTop_6_23[30] , \wRegInTop_6_23[29] , 
        \wRegInTop_6_23[28] , \wRegInTop_6_23[27] , \wRegInTop_6_23[26] , 
        \wRegInTop_6_23[25] , \wRegInTop_6_23[24] , \wRegInTop_6_23[23] , 
        \wRegInTop_6_23[22] , \wRegInTop_6_23[21] , \wRegInTop_6_23[20] , 
        \wRegInTop_6_23[19] , \wRegInTop_6_23[18] , \wRegInTop_6_23[17] , 
        \wRegInTop_6_23[16] , \wRegInTop_6_23[15] , \wRegInTop_6_23[14] , 
        \wRegInTop_6_23[13] , \wRegInTop_6_23[12] , \wRegInTop_6_23[11] , 
        \wRegInTop_6_23[10] , \wRegInTop_6_23[9] , \wRegInTop_6_23[8] , 
        \wRegInTop_6_23[7] , \wRegInTop_6_23[6] , \wRegInTop_6_23[5] , 
        \wRegInTop_6_23[4] , \wRegInTop_6_23[3] , \wRegInTop_6_23[2] , 
        \wRegInTop_6_23[1] , \wRegInTop_6_23[0] }), .In2({\wRegInBot_6_23[31] , 
        \wRegInBot_6_23[30] , \wRegInBot_6_23[29] , \wRegInBot_6_23[28] , 
        \wRegInBot_6_23[27] , \wRegInBot_6_23[26] , \wRegInBot_6_23[25] , 
        \wRegInBot_6_23[24] , \wRegInBot_6_23[23] , \wRegInBot_6_23[22] , 
        \wRegInBot_6_23[21] , \wRegInBot_6_23[20] , \wRegInBot_6_23[19] , 
        \wRegInBot_6_23[18] , \wRegInBot_6_23[17] , \wRegInBot_6_23[16] , 
        \wRegInBot_6_23[15] , \wRegInBot_6_23[14] , \wRegInBot_6_23[13] , 
        \wRegInBot_6_23[12] , \wRegInBot_6_23[11] , \wRegInBot_6_23[10] , 
        \wRegInBot_6_23[9] , \wRegInBot_6_23[8] , \wRegInBot_6_23[7] , 
        \wRegInBot_6_23[6] , \wRegInBot_6_23[5] , \wRegInBot_6_23[4] , 
        \wRegInBot_6_23[3] , \wRegInBot_6_23[2] , \wRegInBot_6_23[1] , 
        \wRegInBot_6_23[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_1_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink3[31] , \ScanLink3[30] , \ScanLink3[29] , 
        \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , \ScanLink3[25] , 
        \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , \ScanLink3[21] , 
        \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , \ScanLink3[17] , 
        \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , \ScanLink3[13] , 
        \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , \ScanLink3[9] , 
        \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , \ScanLink3[5] , 
        \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , \ScanLink3[1] , 
        \ScanLink3[0] }), .ScanOut({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_1_1[31] , \wRegOut_1_1[30] , \wRegOut_1_1[29] , 
        \wRegOut_1_1[28] , \wRegOut_1_1[27] , \wRegOut_1_1[26] , 
        \wRegOut_1_1[25] , \wRegOut_1_1[24] , \wRegOut_1_1[23] , 
        \wRegOut_1_1[22] , \wRegOut_1_1[21] , \wRegOut_1_1[20] , 
        \wRegOut_1_1[19] , \wRegOut_1_1[18] , \wRegOut_1_1[17] , 
        \wRegOut_1_1[16] , \wRegOut_1_1[15] , \wRegOut_1_1[14] , 
        \wRegOut_1_1[13] , \wRegOut_1_1[12] , \wRegOut_1_1[11] , 
        \wRegOut_1_1[10] , \wRegOut_1_1[9] , \wRegOut_1_1[8] , 
        \wRegOut_1_1[7] , \wRegOut_1_1[6] , \wRegOut_1_1[5] , \wRegOut_1_1[4] , 
        \wRegOut_1_1[3] , \wRegOut_1_1[2] , \wRegOut_1_1[1] , \wRegOut_1_1[0] 
        }), .Enable1(\wRegEnTop_1_1[0] ), .Enable2(\wRegEnBot_1_1[0] ), .In1({
        \wRegInTop_1_1[31] , \wRegInTop_1_1[30] , \wRegInTop_1_1[29] , 
        \wRegInTop_1_1[28] , \wRegInTop_1_1[27] , \wRegInTop_1_1[26] , 
        \wRegInTop_1_1[25] , \wRegInTop_1_1[24] , \wRegInTop_1_1[23] , 
        \wRegInTop_1_1[22] , \wRegInTop_1_1[21] , \wRegInTop_1_1[20] , 
        \wRegInTop_1_1[19] , \wRegInTop_1_1[18] , \wRegInTop_1_1[17] , 
        \wRegInTop_1_1[16] , \wRegInTop_1_1[15] , \wRegInTop_1_1[14] , 
        \wRegInTop_1_1[13] , \wRegInTop_1_1[12] , \wRegInTop_1_1[11] , 
        \wRegInTop_1_1[10] , \wRegInTop_1_1[9] , \wRegInTop_1_1[8] , 
        \wRegInTop_1_1[7] , \wRegInTop_1_1[6] , \wRegInTop_1_1[5] , 
        \wRegInTop_1_1[4] , \wRegInTop_1_1[3] , \wRegInTop_1_1[2] , 
        \wRegInTop_1_1[1] , \wRegInTop_1_1[0] }), .In2({\wRegInBot_1_1[31] , 
        \wRegInBot_1_1[30] , \wRegInBot_1_1[29] , \wRegInBot_1_1[28] , 
        \wRegInBot_1_1[27] , \wRegInBot_1_1[26] , \wRegInBot_1_1[25] , 
        \wRegInBot_1_1[24] , \wRegInBot_1_1[23] , \wRegInBot_1_1[22] , 
        \wRegInBot_1_1[21] , \wRegInBot_1_1[20] , \wRegInBot_1_1[19] , 
        \wRegInBot_1_1[18] , \wRegInBot_1_1[17] , \wRegInBot_1_1[16] , 
        \wRegInBot_1_1[15] , \wRegInBot_1_1[14] , \wRegInBot_1_1[13] , 
        \wRegInBot_1_1[12] , \wRegInBot_1_1[11] , \wRegInBot_1_1[10] , 
        \wRegInBot_1_1[9] , \wRegInBot_1_1[8] , \wRegInBot_1_1[7] , 
        \wRegInBot_1_1[6] , \wRegInBot_1_1[5] , \wRegInBot_1_1[4] , 
        \wRegInBot_1_1[3] , \wRegInBot_1_1[2] , \wRegInBot_1_1[1] , 
        \wRegInBot_1_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_2_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink6[31] , \ScanLink6[30] , \ScanLink6[29] , 
        \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , \ScanLink6[25] , 
        \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , \ScanLink6[21] , 
        \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , \ScanLink6[17] , 
        \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , \ScanLink6[13] , 
        \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , \ScanLink6[9] , 
        \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , \ScanLink6[5] , 
        \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , \ScanLink6[1] , 
        \ScanLink6[0] }), .ScanOut({\ScanLink5[31] , \ScanLink5[30] , 
        \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , 
        \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , 
        \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , 
        \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , 
        \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , 
        \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_2_2[31] , \wRegOut_2_2[30] , \wRegOut_2_2[29] , 
        \wRegOut_2_2[28] , \wRegOut_2_2[27] , \wRegOut_2_2[26] , 
        \wRegOut_2_2[25] , \wRegOut_2_2[24] , \wRegOut_2_2[23] , 
        \wRegOut_2_2[22] , \wRegOut_2_2[21] , \wRegOut_2_2[20] , 
        \wRegOut_2_2[19] , \wRegOut_2_2[18] , \wRegOut_2_2[17] , 
        \wRegOut_2_2[16] , \wRegOut_2_2[15] , \wRegOut_2_2[14] , 
        \wRegOut_2_2[13] , \wRegOut_2_2[12] , \wRegOut_2_2[11] , 
        \wRegOut_2_2[10] , \wRegOut_2_2[9] , \wRegOut_2_2[8] , 
        \wRegOut_2_2[7] , \wRegOut_2_2[6] , \wRegOut_2_2[5] , \wRegOut_2_2[4] , 
        \wRegOut_2_2[3] , \wRegOut_2_2[2] , \wRegOut_2_2[1] , \wRegOut_2_2[0] 
        }), .Enable1(\wRegEnTop_2_2[0] ), .Enable2(\wRegEnBot_2_2[0] ), .In1({
        \wRegInTop_2_2[31] , \wRegInTop_2_2[30] , \wRegInTop_2_2[29] , 
        \wRegInTop_2_2[28] , \wRegInTop_2_2[27] , \wRegInTop_2_2[26] , 
        \wRegInTop_2_2[25] , \wRegInTop_2_2[24] , \wRegInTop_2_2[23] , 
        \wRegInTop_2_2[22] , \wRegInTop_2_2[21] , \wRegInTop_2_2[20] , 
        \wRegInTop_2_2[19] , \wRegInTop_2_2[18] , \wRegInTop_2_2[17] , 
        \wRegInTop_2_2[16] , \wRegInTop_2_2[15] , \wRegInTop_2_2[14] , 
        \wRegInTop_2_2[13] , \wRegInTop_2_2[12] , \wRegInTop_2_2[11] , 
        \wRegInTop_2_2[10] , \wRegInTop_2_2[9] , \wRegInTop_2_2[8] , 
        \wRegInTop_2_2[7] , \wRegInTop_2_2[6] , \wRegInTop_2_2[5] , 
        \wRegInTop_2_2[4] , \wRegInTop_2_2[3] , \wRegInTop_2_2[2] , 
        \wRegInTop_2_2[1] , \wRegInTop_2_2[0] }), .In2({\wRegInBot_2_2[31] , 
        \wRegInBot_2_2[30] , \wRegInBot_2_2[29] , \wRegInBot_2_2[28] , 
        \wRegInBot_2_2[27] , \wRegInBot_2_2[26] , \wRegInBot_2_2[25] , 
        \wRegInBot_2_2[24] , \wRegInBot_2_2[23] , \wRegInBot_2_2[22] , 
        \wRegInBot_2_2[21] , \wRegInBot_2_2[20] , \wRegInBot_2_2[19] , 
        \wRegInBot_2_2[18] , \wRegInBot_2_2[17] , \wRegInBot_2_2[16] , 
        \wRegInBot_2_2[15] , \wRegInBot_2_2[14] , \wRegInBot_2_2[13] , 
        \wRegInBot_2_2[12] , \wRegInBot_2_2[11] , \wRegInBot_2_2[10] , 
        \wRegInBot_2_2[9] , \wRegInBot_2_2[8] , \wRegInBot_2_2[7] , 
        \wRegInBot_2_2[6] , \wRegInBot_2_2[5] , \wRegInBot_2_2[4] , 
        \wRegInBot_2_2[3] , \wRegInBot_2_2[2] , \wRegInBot_2_2[1] , 
        \wRegInBot_2_2[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink10[31] , \ScanLink10[30] , \ScanLink10[29] , 
        \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , \ScanLink10[25] , 
        \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , \ScanLink10[21] , 
        \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , \ScanLink10[17] , 
        \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , \ScanLink10[13] , 
        \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , \ScanLink10[9] , 
        \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , \ScanLink10[5] , 
        \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , \ScanLink10[1] , 
        \ScanLink10[0] }), .ScanOut({\ScanLink9[31] , \ScanLink9[30] , 
        \ScanLink9[29] , \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , 
        \ScanLink9[25] , \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , 
        \ScanLink9[21] , \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , 
        \ScanLink9[17] , \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , 
        \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , 
        \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , 
        \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , 
        \ScanLink9[1] , \ScanLink9[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_2[31] , \wRegOut_3_2[30] , \wRegOut_3_2[29] , 
        \wRegOut_3_2[28] , \wRegOut_3_2[27] , \wRegOut_3_2[26] , 
        \wRegOut_3_2[25] , \wRegOut_3_2[24] , \wRegOut_3_2[23] , 
        \wRegOut_3_2[22] , \wRegOut_3_2[21] , \wRegOut_3_2[20] , 
        \wRegOut_3_2[19] , \wRegOut_3_2[18] , \wRegOut_3_2[17] , 
        \wRegOut_3_2[16] , \wRegOut_3_2[15] , \wRegOut_3_2[14] , 
        \wRegOut_3_2[13] , \wRegOut_3_2[12] , \wRegOut_3_2[11] , 
        \wRegOut_3_2[10] , \wRegOut_3_2[9] , \wRegOut_3_2[8] , 
        \wRegOut_3_2[7] , \wRegOut_3_2[6] , \wRegOut_3_2[5] , \wRegOut_3_2[4] , 
        \wRegOut_3_2[3] , \wRegOut_3_2[2] , \wRegOut_3_2[1] , \wRegOut_3_2[0] 
        }), .Enable1(\wRegEnTop_3_2[0] ), .Enable2(\wRegEnBot_3_2[0] ), .In1({
        \wRegInTop_3_2[31] , \wRegInTop_3_2[30] , \wRegInTop_3_2[29] , 
        \wRegInTop_3_2[28] , \wRegInTop_3_2[27] , \wRegInTop_3_2[26] , 
        \wRegInTop_3_2[25] , \wRegInTop_3_2[24] , \wRegInTop_3_2[23] , 
        \wRegInTop_3_2[22] , \wRegInTop_3_2[21] , \wRegInTop_3_2[20] , 
        \wRegInTop_3_2[19] , \wRegInTop_3_2[18] , \wRegInTop_3_2[17] , 
        \wRegInTop_3_2[16] , \wRegInTop_3_2[15] , \wRegInTop_3_2[14] , 
        \wRegInTop_3_2[13] , \wRegInTop_3_2[12] , \wRegInTop_3_2[11] , 
        \wRegInTop_3_2[10] , \wRegInTop_3_2[9] , \wRegInTop_3_2[8] , 
        \wRegInTop_3_2[7] , \wRegInTop_3_2[6] , \wRegInTop_3_2[5] , 
        \wRegInTop_3_2[4] , \wRegInTop_3_2[3] , \wRegInTop_3_2[2] , 
        \wRegInTop_3_2[1] , \wRegInTop_3_2[0] }), .In2({\wRegInBot_3_2[31] , 
        \wRegInBot_3_2[30] , \wRegInBot_3_2[29] , \wRegInBot_3_2[28] , 
        \wRegInBot_3_2[27] , \wRegInBot_3_2[26] , \wRegInBot_3_2[25] , 
        \wRegInBot_3_2[24] , \wRegInBot_3_2[23] , \wRegInBot_3_2[22] , 
        \wRegInBot_3_2[21] , \wRegInBot_3_2[20] , \wRegInBot_3_2[19] , 
        \wRegInBot_3_2[18] , \wRegInBot_3_2[17] , \wRegInBot_3_2[16] , 
        \wRegInBot_3_2[15] , \wRegInBot_3_2[14] , \wRegInBot_3_2[13] , 
        \wRegInBot_3_2[12] , \wRegInBot_3_2[11] , \wRegInBot_3_2[10] , 
        \wRegInBot_3_2[9] , \wRegInBot_3_2[8] , \wRegInBot_3_2[7] , 
        \wRegInBot_3_2[6] , \wRegInBot_3_2[5] , \wRegInBot_3_2[4] , 
        \wRegInBot_3_2[3] , \wRegInBot_3_2[2] , \wRegInBot_3_2[1] , 
        \wRegInBot_3_2[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink17[31] , \ScanLink17[30] , \ScanLink17[29] , 
        \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , \ScanLink17[25] , 
        \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , \ScanLink17[21] , 
        \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , \ScanLink17[17] , 
        \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , \ScanLink17[13] , 
        \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , \ScanLink17[9] , 
        \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , \ScanLink17[5] , 
        \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , \ScanLink17[1] , 
        \ScanLink17[0] }), .ScanOut({\ScanLink16[31] , \ScanLink16[30] , 
        \ScanLink16[29] , \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , 
        \ScanLink16[25] , \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , 
        \ScanLink16[21] , \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , 
        \ScanLink16[17] , \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , 
        \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , 
        \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , 
        \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , 
        \ScanLink16[1] , \ScanLink16[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_1[31] , \wRegOut_4_1[30] , \wRegOut_4_1[29] , 
        \wRegOut_4_1[28] , \wRegOut_4_1[27] , \wRegOut_4_1[26] , 
        \wRegOut_4_1[25] , \wRegOut_4_1[24] , \wRegOut_4_1[23] , 
        \wRegOut_4_1[22] , \wRegOut_4_1[21] , \wRegOut_4_1[20] , 
        \wRegOut_4_1[19] , \wRegOut_4_1[18] , \wRegOut_4_1[17] , 
        \wRegOut_4_1[16] , \wRegOut_4_1[15] , \wRegOut_4_1[14] , 
        \wRegOut_4_1[13] , \wRegOut_4_1[12] , \wRegOut_4_1[11] , 
        \wRegOut_4_1[10] , \wRegOut_4_1[9] , \wRegOut_4_1[8] , 
        \wRegOut_4_1[7] , \wRegOut_4_1[6] , \wRegOut_4_1[5] , \wRegOut_4_1[4] , 
        \wRegOut_4_1[3] , \wRegOut_4_1[2] , \wRegOut_4_1[1] , \wRegOut_4_1[0] 
        }), .Enable1(\wRegEnTop_4_1[0] ), .Enable2(\wRegEnBot_4_1[0] ), .In1({
        \wRegInTop_4_1[31] , \wRegInTop_4_1[30] , \wRegInTop_4_1[29] , 
        \wRegInTop_4_1[28] , \wRegInTop_4_1[27] , \wRegInTop_4_1[26] , 
        \wRegInTop_4_1[25] , \wRegInTop_4_1[24] , \wRegInTop_4_1[23] , 
        \wRegInTop_4_1[22] , \wRegInTop_4_1[21] , \wRegInTop_4_1[20] , 
        \wRegInTop_4_1[19] , \wRegInTop_4_1[18] , \wRegInTop_4_1[17] , 
        \wRegInTop_4_1[16] , \wRegInTop_4_1[15] , \wRegInTop_4_1[14] , 
        \wRegInTop_4_1[13] , \wRegInTop_4_1[12] , \wRegInTop_4_1[11] , 
        \wRegInTop_4_1[10] , \wRegInTop_4_1[9] , \wRegInTop_4_1[8] , 
        \wRegInTop_4_1[7] , \wRegInTop_4_1[6] , \wRegInTop_4_1[5] , 
        \wRegInTop_4_1[4] , \wRegInTop_4_1[3] , \wRegInTop_4_1[2] , 
        \wRegInTop_4_1[1] , \wRegInTop_4_1[0] }), .In2({\wRegInBot_4_1[31] , 
        \wRegInBot_4_1[30] , \wRegInBot_4_1[29] , \wRegInBot_4_1[28] , 
        \wRegInBot_4_1[27] , \wRegInBot_4_1[26] , \wRegInBot_4_1[25] , 
        \wRegInBot_4_1[24] , \wRegInBot_4_1[23] , \wRegInBot_4_1[22] , 
        \wRegInBot_4_1[21] , \wRegInBot_4_1[20] , \wRegInBot_4_1[19] , 
        \wRegInBot_4_1[18] , \wRegInBot_4_1[17] , \wRegInBot_4_1[16] , 
        \wRegInBot_4_1[15] , \wRegInBot_4_1[14] , \wRegInBot_4_1[13] , 
        \wRegInBot_4_1[12] , \wRegInBot_4_1[11] , \wRegInBot_4_1[10] , 
        \wRegInBot_4_1[9] , \wRegInBot_4_1[8] , \wRegInBot_4_1[7] , 
        \wRegInBot_4_1[6] , \wRegInBot_4_1[5] , \wRegInBot_4_1[4] , 
        \wRegInBot_4_1[3] , \wRegInBot_4_1[2] , \wRegInBot_4_1[1] , 
        \wRegInBot_4_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink46[31] , \ScanLink46[30] , \ScanLink46[29] , 
        \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , \ScanLink46[25] , 
        \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , \ScanLink46[21] , 
        \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , \ScanLink46[17] , 
        \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , \ScanLink46[13] , 
        \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , \ScanLink46[9] , 
        \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , \ScanLink46[5] , 
        \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , \ScanLink46[1] , 
        \ScanLink46[0] }), .ScanOut({\ScanLink45[31] , \ScanLink45[30] , 
        \ScanLink45[29] , \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , 
        \ScanLink45[25] , \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , 
        \ScanLink45[21] , \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , 
        \ScanLink45[17] , \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , 
        \ScanLink45[13] , \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , 
        \ScanLink45[9] , \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , 
        \ScanLink45[5] , \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , 
        \ScanLink45[1] , \ScanLink45[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_14[31] , \wRegOut_5_14[30] , 
        \wRegOut_5_14[29] , \wRegOut_5_14[28] , \wRegOut_5_14[27] , 
        \wRegOut_5_14[26] , \wRegOut_5_14[25] , \wRegOut_5_14[24] , 
        \wRegOut_5_14[23] , \wRegOut_5_14[22] , \wRegOut_5_14[21] , 
        \wRegOut_5_14[20] , \wRegOut_5_14[19] , \wRegOut_5_14[18] , 
        \wRegOut_5_14[17] , \wRegOut_5_14[16] , \wRegOut_5_14[15] , 
        \wRegOut_5_14[14] , \wRegOut_5_14[13] , \wRegOut_5_14[12] , 
        \wRegOut_5_14[11] , \wRegOut_5_14[10] , \wRegOut_5_14[9] , 
        \wRegOut_5_14[8] , \wRegOut_5_14[7] , \wRegOut_5_14[6] , 
        \wRegOut_5_14[5] , \wRegOut_5_14[4] , \wRegOut_5_14[3] , 
        \wRegOut_5_14[2] , \wRegOut_5_14[1] , \wRegOut_5_14[0] }), .Enable1(
        \wRegEnTop_5_14[0] ), .Enable2(\wRegEnBot_5_14[0] ), .In1({
        \wRegInTop_5_14[31] , \wRegInTop_5_14[30] , \wRegInTop_5_14[29] , 
        \wRegInTop_5_14[28] , \wRegInTop_5_14[27] , \wRegInTop_5_14[26] , 
        \wRegInTop_5_14[25] , \wRegInTop_5_14[24] , \wRegInTop_5_14[23] , 
        \wRegInTop_5_14[22] , \wRegInTop_5_14[21] , \wRegInTop_5_14[20] , 
        \wRegInTop_5_14[19] , \wRegInTop_5_14[18] , \wRegInTop_5_14[17] , 
        \wRegInTop_5_14[16] , \wRegInTop_5_14[15] , \wRegInTop_5_14[14] , 
        \wRegInTop_5_14[13] , \wRegInTop_5_14[12] , \wRegInTop_5_14[11] , 
        \wRegInTop_5_14[10] , \wRegInTop_5_14[9] , \wRegInTop_5_14[8] , 
        \wRegInTop_5_14[7] , \wRegInTop_5_14[6] , \wRegInTop_5_14[5] , 
        \wRegInTop_5_14[4] , \wRegInTop_5_14[3] , \wRegInTop_5_14[2] , 
        \wRegInTop_5_14[1] , \wRegInTop_5_14[0] }), .In2({\wRegInBot_5_14[31] , 
        \wRegInBot_5_14[30] , \wRegInBot_5_14[29] , \wRegInBot_5_14[28] , 
        \wRegInBot_5_14[27] , \wRegInBot_5_14[26] , \wRegInBot_5_14[25] , 
        \wRegInBot_5_14[24] , \wRegInBot_5_14[23] , \wRegInBot_5_14[22] , 
        \wRegInBot_5_14[21] , \wRegInBot_5_14[20] , \wRegInBot_5_14[19] , 
        \wRegInBot_5_14[18] , \wRegInBot_5_14[17] , \wRegInBot_5_14[16] , 
        \wRegInBot_5_14[15] , \wRegInBot_5_14[14] , \wRegInBot_5_14[13] , 
        \wRegInBot_5_14[12] , \wRegInBot_5_14[11] , \wRegInBot_5_14[10] , 
        \wRegInBot_5_14[9] , \wRegInBot_5_14[8] , \wRegInBot_5_14[7] , 
        \wRegInBot_5_14[6] , \wRegInBot_5_14[5] , \wRegInBot_5_14[4] , 
        \wRegInBot_5_14[3] , \wRegInBot_5_14[2] , \wRegInBot_5_14[1] , 
        \wRegInBot_5_14[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_50 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink178[31] , \ScanLink178[30] , \ScanLink178[29] , 
        \ScanLink178[28] , \ScanLink178[27] , \ScanLink178[26] , 
        \ScanLink178[25] , \ScanLink178[24] , \ScanLink178[23] , 
        \ScanLink178[22] , \ScanLink178[21] , \ScanLink178[20] , 
        \ScanLink178[19] , \ScanLink178[18] , \ScanLink178[17] , 
        \ScanLink178[16] , \ScanLink178[15] , \ScanLink178[14] , 
        \ScanLink178[13] , \ScanLink178[12] , \ScanLink178[11] , 
        \ScanLink178[10] , \ScanLink178[9] , \ScanLink178[8] , 
        \ScanLink178[7] , \ScanLink178[6] , \ScanLink178[5] , \ScanLink178[4] , 
        \ScanLink178[3] , \ScanLink178[2] , \ScanLink178[1] , \ScanLink178[0] 
        }), .ScanOut({\ScanLink177[31] , \ScanLink177[30] , \ScanLink177[29] , 
        \ScanLink177[28] , \ScanLink177[27] , \ScanLink177[26] , 
        \ScanLink177[25] , \ScanLink177[24] , \ScanLink177[23] , 
        \ScanLink177[22] , \ScanLink177[21] , \ScanLink177[20] , 
        \ScanLink177[19] , \ScanLink177[18] , \ScanLink177[17] , 
        \ScanLink177[16] , \ScanLink177[15] , \ScanLink177[14] , 
        \ScanLink177[13] , \ScanLink177[12] , \ScanLink177[11] , 
        \ScanLink177[10] , \ScanLink177[9] , \ScanLink177[8] , 
        \ScanLink177[7] , \ScanLink177[6] , \ScanLink177[5] , \ScanLink177[4] , 
        \ScanLink177[3] , \ScanLink177[2] , \ScanLink177[1] , \ScanLink177[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_50[31] , 
        \wRegOut_7_50[30] , \wRegOut_7_50[29] , \wRegOut_7_50[28] , 
        \wRegOut_7_50[27] , \wRegOut_7_50[26] , \wRegOut_7_50[25] , 
        \wRegOut_7_50[24] , \wRegOut_7_50[23] , \wRegOut_7_50[22] , 
        \wRegOut_7_50[21] , \wRegOut_7_50[20] , \wRegOut_7_50[19] , 
        \wRegOut_7_50[18] , \wRegOut_7_50[17] , \wRegOut_7_50[16] , 
        \wRegOut_7_50[15] , \wRegOut_7_50[14] , \wRegOut_7_50[13] , 
        \wRegOut_7_50[12] , \wRegOut_7_50[11] , \wRegOut_7_50[10] , 
        \wRegOut_7_50[9] , \wRegOut_7_50[8] , \wRegOut_7_50[7] , 
        \wRegOut_7_50[6] , \wRegOut_7_50[5] , \wRegOut_7_50[4] , 
        \wRegOut_7_50[3] , \wRegOut_7_50[2] , \wRegOut_7_50[1] , 
        \wRegOut_7_50[0] }), .Enable1(\wRegEnTop_7_50[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_50[31] , \wRegInTop_7_50[30] , \wRegInTop_7_50[29] , 
        \wRegInTop_7_50[28] , \wRegInTop_7_50[27] , \wRegInTop_7_50[26] , 
        \wRegInTop_7_50[25] , \wRegInTop_7_50[24] , \wRegInTop_7_50[23] , 
        \wRegInTop_7_50[22] , \wRegInTop_7_50[21] , \wRegInTop_7_50[20] , 
        \wRegInTop_7_50[19] , \wRegInTop_7_50[18] , \wRegInTop_7_50[17] , 
        \wRegInTop_7_50[16] , \wRegInTop_7_50[15] , \wRegInTop_7_50[14] , 
        \wRegInTop_7_50[13] , \wRegInTop_7_50[12] , \wRegInTop_7_50[11] , 
        \wRegInTop_7_50[10] , \wRegInTop_7_50[9] , \wRegInTop_7_50[8] , 
        \wRegInTop_7_50[7] , \wRegInTop_7_50[6] , \wRegInTop_7_50[5] , 
        \wRegInTop_7_50[4] , \wRegInTop_7_50[3] , \wRegInTop_7_50[2] , 
        \wRegInTop_7_50[1] , \wRegInTop_7_50[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_57 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink185[31] , \ScanLink185[30] , \ScanLink185[29] , 
        \ScanLink185[28] , \ScanLink185[27] , \ScanLink185[26] , 
        \ScanLink185[25] , \ScanLink185[24] , \ScanLink185[23] , 
        \ScanLink185[22] , \ScanLink185[21] , \ScanLink185[20] , 
        \ScanLink185[19] , \ScanLink185[18] , \ScanLink185[17] , 
        \ScanLink185[16] , \ScanLink185[15] , \ScanLink185[14] , 
        \ScanLink185[13] , \ScanLink185[12] , \ScanLink185[11] , 
        \ScanLink185[10] , \ScanLink185[9] , \ScanLink185[8] , 
        \ScanLink185[7] , \ScanLink185[6] , \ScanLink185[5] , \ScanLink185[4] , 
        \ScanLink185[3] , \ScanLink185[2] , \ScanLink185[1] , \ScanLink185[0] 
        }), .ScanOut({\ScanLink184[31] , \ScanLink184[30] , \ScanLink184[29] , 
        \ScanLink184[28] , \ScanLink184[27] , \ScanLink184[26] , 
        \ScanLink184[25] , \ScanLink184[24] , \ScanLink184[23] , 
        \ScanLink184[22] , \ScanLink184[21] , \ScanLink184[20] , 
        \ScanLink184[19] , \ScanLink184[18] , \ScanLink184[17] , 
        \ScanLink184[16] , \ScanLink184[15] , \ScanLink184[14] , 
        \ScanLink184[13] , \ScanLink184[12] , \ScanLink184[11] , 
        \ScanLink184[10] , \ScanLink184[9] , \ScanLink184[8] , 
        \ScanLink184[7] , \ScanLink184[6] , \ScanLink184[5] , \ScanLink184[4] , 
        \ScanLink184[3] , \ScanLink184[2] , \ScanLink184[1] , \ScanLink184[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_57[31] , 
        \wRegOut_7_57[30] , \wRegOut_7_57[29] , \wRegOut_7_57[28] , 
        \wRegOut_7_57[27] , \wRegOut_7_57[26] , \wRegOut_7_57[25] , 
        \wRegOut_7_57[24] , \wRegOut_7_57[23] , \wRegOut_7_57[22] , 
        \wRegOut_7_57[21] , \wRegOut_7_57[20] , \wRegOut_7_57[19] , 
        \wRegOut_7_57[18] , \wRegOut_7_57[17] , \wRegOut_7_57[16] , 
        \wRegOut_7_57[15] , \wRegOut_7_57[14] , \wRegOut_7_57[13] , 
        \wRegOut_7_57[12] , \wRegOut_7_57[11] , \wRegOut_7_57[10] , 
        \wRegOut_7_57[9] , \wRegOut_7_57[8] , \wRegOut_7_57[7] , 
        \wRegOut_7_57[6] , \wRegOut_7_57[5] , \wRegOut_7_57[4] , 
        \wRegOut_7_57[3] , \wRegOut_7_57[2] , \wRegOut_7_57[1] , 
        \wRegOut_7_57[0] }), .Enable1(\wRegEnTop_7_57[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_57[31] , \wRegInTop_7_57[30] , \wRegInTop_7_57[29] , 
        \wRegInTop_7_57[28] , \wRegInTop_7_57[27] , \wRegInTop_7_57[26] , 
        \wRegInTop_7_57[25] , \wRegInTop_7_57[24] , \wRegInTop_7_57[23] , 
        \wRegInTop_7_57[22] , \wRegInTop_7_57[21] , \wRegInTop_7_57[20] , 
        \wRegInTop_7_57[19] , \wRegInTop_7_57[18] , \wRegInTop_7_57[17] , 
        \wRegInTop_7_57[16] , \wRegInTop_7_57[15] , \wRegInTop_7_57[14] , 
        \wRegInTop_7_57[13] , \wRegInTop_7_57[12] , \wRegInTop_7_57[11] , 
        \wRegInTop_7_57[10] , \wRegInTop_7_57[9] , \wRegInTop_7_57[8] , 
        \wRegInTop_7_57[7] , \wRegInTop_7_57[6] , \wRegInTop_7_57[5] , 
        \wRegInTop_7_57[4] , \wRegInTop_7_57[3] , \wRegInTop_7_57[2] , 
        \wRegInTop_7_57[1] , \wRegInTop_7_57[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_24 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink88[31] , \ScanLink88[30] , \ScanLink88[29] , 
        \ScanLink88[28] , \ScanLink88[27] , \ScanLink88[26] , \ScanLink88[25] , 
        \ScanLink88[24] , \ScanLink88[23] , \ScanLink88[22] , \ScanLink88[21] , 
        \ScanLink88[20] , \ScanLink88[19] , \ScanLink88[18] , \ScanLink88[17] , 
        \ScanLink88[16] , \ScanLink88[15] , \ScanLink88[14] , \ScanLink88[13] , 
        \ScanLink88[12] , \ScanLink88[11] , \ScanLink88[10] , \ScanLink88[9] , 
        \ScanLink88[8] , \ScanLink88[7] , \ScanLink88[6] , \ScanLink88[5] , 
        \ScanLink88[4] , \ScanLink88[3] , \ScanLink88[2] , \ScanLink88[1] , 
        \ScanLink88[0] }), .ScanOut({\ScanLink87[31] , \ScanLink87[30] , 
        \ScanLink87[29] , \ScanLink87[28] , \ScanLink87[27] , \ScanLink87[26] , 
        \ScanLink87[25] , \ScanLink87[24] , \ScanLink87[23] , \ScanLink87[22] , 
        \ScanLink87[21] , \ScanLink87[20] , \ScanLink87[19] , \ScanLink87[18] , 
        \ScanLink87[17] , \ScanLink87[16] , \ScanLink87[15] , \ScanLink87[14] , 
        \ScanLink87[13] , \ScanLink87[12] , \ScanLink87[11] , \ScanLink87[10] , 
        \ScanLink87[9] , \ScanLink87[8] , \ScanLink87[7] , \ScanLink87[6] , 
        \ScanLink87[5] , \ScanLink87[4] , \ScanLink87[3] , \ScanLink87[2] , 
        \ScanLink87[1] , \ScanLink87[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_24[31] , \wRegOut_6_24[30] , 
        \wRegOut_6_24[29] , \wRegOut_6_24[28] , \wRegOut_6_24[27] , 
        \wRegOut_6_24[26] , \wRegOut_6_24[25] , \wRegOut_6_24[24] , 
        \wRegOut_6_24[23] , \wRegOut_6_24[22] , \wRegOut_6_24[21] , 
        \wRegOut_6_24[20] , \wRegOut_6_24[19] , \wRegOut_6_24[18] , 
        \wRegOut_6_24[17] , \wRegOut_6_24[16] , \wRegOut_6_24[15] , 
        \wRegOut_6_24[14] , \wRegOut_6_24[13] , \wRegOut_6_24[12] , 
        \wRegOut_6_24[11] , \wRegOut_6_24[10] , \wRegOut_6_24[9] , 
        \wRegOut_6_24[8] , \wRegOut_6_24[7] , \wRegOut_6_24[6] , 
        \wRegOut_6_24[5] , \wRegOut_6_24[4] , \wRegOut_6_24[3] , 
        \wRegOut_6_24[2] , \wRegOut_6_24[1] , \wRegOut_6_24[0] }), .Enable1(
        \wRegEnTop_6_24[0] ), .Enable2(\wRegEnBot_6_24[0] ), .In1({
        \wRegInTop_6_24[31] , \wRegInTop_6_24[30] , \wRegInTop_6_24[29] , 
        \wRegInTop_6_24[28] , \wRegInTop_6_24[27] , \wRegInTop_6_24[26] , 
        \wRegInTop_6_24[25] , \wRegInTop_6_24[24] , \wRegInTop_6_24[23] , 
        \wRegInTop_6_24[22] , \wRegInTop_6_24[21] , \wRegInTop_6_24[20] , 
        \wRegInTop_6_24[19] , \wRegInTop_6_24[18] , \wRegInTop_6_24[17] , 
        \wRegInTop_6_24[16] , \wRegInTop_6_24[15] , \wRegInTop_6_24[14] , 
        \wRegInTop_6_24[13] , \wRegInTop_6_24[12] , \wRegInTop_6_24[11] , 
        \wRegInTop_6_24[10] , \wRegInTop_6_24[9] , \wRegInTop_6_24[8] , 
        \wRegInTop_6_24[7] , \wRegInTop_6_24[6] , \wRegInTop_6_24[5] , 
        \wRegInTop_6_24[4] , \wRegInTop_6_24[3] , \wRegInTop_6_24[2] , 
        \wRegInTop_6_24[1] , \wRegInTop_6_24[0] }), .In2({\wRegInBot_6_24[31] , 
        \wRegInBot_6_24[30] , \wRegInBot_6_24[29] , \wRegInBot_6_24[28] , 
        \wRegInBot_6_24[27] , \wRegInBot_6_24[26] , \wRegInBot_6_24[25] , 
        \wRegInBot_6_24[24] , \wRegInBot_6_24[23] , \wRegInBot_6_24[22] , 
        \wRegInBot_6_24[21] , \wRegInBot_6_24[20] , \wRegInBot_6_24[19] , 
        \wRegInBot_6_24[18] , \wRegInBot_6_24[17] , \wRegInBot_6_24[16] , 
        \wRegInBot_6_24[15] , \wRegInBot_6_24[14] , \wRegInBot_6_24[13] , 
        \wRegInBot_6_24[12] , \wRegInBot_6_24[11] , \wRegInBot_6_24[10] , 
        \wRegInBot_6_24[9] , \wRegInBot_6_24[8] , \wRegInBot_6_24[7] , 
        \wRegInBot_6_24[6] , \wRegInBot_6_24[5] , \wRegInBot_6_24[4] , 
        \wRegInBot_6_24[3] , \wRegInBot_6_24[2] , \wRegInBot_6_24[1] , 
        \wRegInBot_6_24[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink31[31] , \ScanLink31[30] , \ScanLink31[29] , 
        \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , \ScanLink31[25] , 
        \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , \ScanLink31[21] , 
        \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , \ScanLink31[17] , 
        \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , \ScanLink31[13] , 
        \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , \ScanLink31[9] , 
        \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , \ScanLink31[5] , 
        \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , \ScanLink31[1] , 
        \ScanLink31[0] }), .ScanOut({\ScanLink30[31] , \ScanLink30[30] , 
        \ScanLink30[29] , \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , 
        \ScanLink30[25] , \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , 
        \ScanLink30[21] , \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , 
        \ScanLink30[17] , \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , 
        \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , 
        \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , 
        \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , 
        \ScanLink30[1] , \ScanLink30[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_15[31] , \wRegOut_4_15[30] , 
        \wRegOut_4_15[29] , \wRegOut_4_15[28] , \wRegOut_4_15[27] , 
        \wRegOut_4_15[26] , \wRegOut_4_15[25] , \wRegOut_4_15[24] , 
        \wRegOut_4_15[23] , \wRegOut_4_15[22] , \wRegOut_4_15[21] , 
        \wRegOut_4_15[20] , \wRegOut_4_15[19] , \wRegOut_4_15[18] , 
        \wRegOut_4_15[17] , \wRegOut_4_15[16] , \wRegOut_4_15[15] , 
        \wRegOut_4_15[14] , \wRegOut_4_15[13] , \wRegOut_4_15[12] , 
        \wRegOut_4_15[11] , \wRegOut_4_15[10] , \wRegOut_4_15[9] , 
        \wRegOut_4_15[8] , \wRegOut_4_15[7] , \wRegOut_4_15[6] , 
        \wRegOut_4_15[5] , \wRegOut_4_15[4] , \wRegOut_4_15[3] , 
        \wRegOut_4_15[2] , \wRegOut_4_15[1] , \wRegOut_4_15[0] }), .Enable1(
        \wRegEnTop_4_15[0] ), .Enable2(\wRegEnBot_4_15[0] ), .In1({
        \wRegInTop_4_15[31] , \wRegInTop_4_15[30] , \wRegInTop_4_15[29] , 
        \wRegInTop_4_15[28] , \wRegInTop_4_15[27] , \wRegInTop_4_15[26] , 
        \wRegInTop_4_15[25] , \wRegInTop_4_15[24] , \wRegInTop_4_15[23] , 
        \wRegInTop_4_15[22] , \wRegInTop_4_15[21] , \wRegInTop_4_15[20] , 
        \wRegInTop_4_15[19] , \wRegInTop_4_15[18] , \wRegInTop_4_15[17] , 
        \wRegInTop_4_15[16] , \wRegInTop_4_15[15] , \wRegInTop_4_15[14] , 
        \wRegInTop_4_15[13] , \wRegInTop_4_15[12] , \wRegInTop_4_15[11] , 
        \wRegInTop_4_15[10] , \wRegInTop_4_15[9] , \wRegInTop_4_15[8] , 
        \wRegInTop_4_15[7] , \wRegInTop_4_15[6] , \wRegInTop_4_15[5] , 
        \wRegInTop_4_15[4] , \wRegInTop_4_15[3] , \wRegInTop_4_15[2] , 
        \wRegInTop_4_15[1] , \wRegInTop_4_15[0] }), .In2({\wRegInBot_4_15[31] , 
        \wRegInBot_4_15[30] , \wRegInBot_4_15[29] , \wRegInBot_4_15[28] , 
        \wRegInBot_4_15[27] , \wRegInBot_4_15[26] , \wRegInBot_4_15[25] , 
        \wRegInBot_4_15[24] , \wRegInBot_4_15[23] , \wRegInBot_4_15[22] , 
        \wRegInBot_4_15[21] , \wRegInBot_4_15[20] , \wRegInBot_4_15[19] , 
        \wRegInBot_4_15[18] , \wRegInBot_4_15[17] , \wRegInBot_4_15[16] , 
        \wRegInBot_4_15[15] , \wRegInBot_4_15[14] , \wRegInBot_4_15[13] , 
        \wRegInBot_4_15[12] , \wRegInBot_4_15[11] , \wRegInBot_4_15[10] , 
        \wRegInBot_4_15[9] , \wRegInBot_4_15[8] , \wRegInBot_4_15[7] , 
        \wRegInBot_4_15[6] , \wRegInBot_4_15[5] , \wRegInBot_4_15[4] , 
        \wRegInBot_4_15[3] , \wRegInBot_4_15[2] , \wRegInBot_4_15[1] , 
        \wRegInBot_4_15[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_51 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink115[31] , \ScanLink115[30] , \ScanLink115[29] , 
        \ScanLink115[28] , \ScanLink115[27] , \ScanLink115[26] , 
        \ScanLink115[25] , \ScanLink115[24] , \ScanLink115[23] , 
        \ScanLink115[22] , \ScanLink115[21] , \ScanLink115[20] , 
        \ScanLink115[19] , \ScanLink115[18] , \ScanLink115[17] , 
        \ScanLink115[16] , \ScanLink115[15] , \ScanLink115[14] , 
        \ScanLink115[13] , \ScanLink115[12] , \ScanLink115[11] , 
        \ScanLink115[10] , \ScanLink115[9] , \ScanLink115[8] , 
        \ScanLink115[7] , \ScanLink115[6] , \ScanLink115[5] , \ScanLink115[4] , 
        \ScanLink115[3] , \ScanLink115[2] , \ScanLink115[1] , \ScanLink115[0] 
        }), .ScanOut({\ScanLink114[31] , \ScanLink114[30] , \ScanLink114[29] , 
        \ScanLink114[28] , \ScanLink114[27] , \ScanLink114[26] , 
        \ScanLink114[25] , \ScanLink114[24] , \ScanLink114[23] , 
        \ScanLink114[22] , \ScanLink114[21] , \ScanLink114[20] , 
        \ScanLink114[19] , \ScanLink114[18] , \ScanLink114[17] , 
        \ScanLink114[16] , \ScanLink114[15] , \ScanLink114[14] , 
        \ScanLink114[13] , \ScanLink114[12] , \ScanLink114[11] , 
        \ScanLink114[10] , \ScanLink114[9] , \ScanLink114[8] , 
        \ScanLink114[7] , \ScanLink114[6] , \ScanLink114[5] , \ScanLink114[4] , 
        \ScanLink114[3] , \ScanLink114[2] , \ScanLink114[1] , \ScanLink114[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_51[31] , 
        \wRegOut_6_51[30] , \wRegOut_6_51[29] , \wRegOut_6_51[28] , 
        \wRegOut_6_51[27] , \wRegOut_6_51[26] , \wRegOut_6_51[25] , 
        \wRegOut_6_51[24] , \wRegOut_6_51[23] , \wRegOut_6_51[22] , 
        \wRegOut_6_51[21] , \wRegOut_6_51[20] , \wRegOut_6_51[19] , 
        \wRegOut_6_51[18] , \wRegOut_6_51[17] , \wRegOut_6_51[16] , 
        \wRegOut_6_51[15] , \wRegOut_6_51[14] , \wRegOut_6_51[13] , 
        \wRegOut_6_51[12] , \wRegOut_6_51[11] , \wRegOut_6_51[10] , 
        \wRegOut_6_51[9] , \wRegOut_6_51[8] , \wRegOut_6_51[7] , 
        \wRegOut_6_51[6] , \wRegOut_6_51[5] , \wRegOut_6_51[4] , 
        \wRegOut_6_51[3] , \wRegOut_6_51[2] , \wRegOut_6_51[1] , 
        \wRegOut_6_51[0] }), .Enable1(\wRegEnTop_6_51[0] ), .Enable2(
        \wRegEnBot_6_51[0] ), .In1({\wRegInTop_6_51[31] , \wRegInTop_6_51[30] , 
        \wRegInTop_6_51[29] , \wRegInTop_6_51[28] , \wRegInTop_6_51[27] , 
        \wRegInTop_6_51[26] , \wRegInTop_6_51[25] , \wRegInTop_6_51[24] , 
        \wRegInTop_6_51[23] , \wRegInTop_6_51[22] , \wRegInTop_6_51[21] , 
        \wRegInTop_6_51[20] , \wRegInTop_6_51[19] , \wRegInTop_6_51[18] , 
        \wRegInTop_6_51[17] , \wRegInTop_6_51[16] , \wRegInTop_6_51[15] , 
        \wRegInTop_6_51[14] , \wRegInTop_6_51[13] , \wRegInTop_6_51[12] , 
        \wRegInTop_6_51[11] , \wRegInTop_6_51[10] , \wRegInTop_6_51[9] , 
        \wRegInTop_6_51[8] , \wRegInTop_6_51[7] , \wRegInTop_6_51[6] , 
        \wRegInTop_6_51[5] , \wRegInTop_6_51[4] , \wRegInTop_6_51[3] , 
        \wRegInTop_6_51[2] , \wRegInTop_6_51[1] , \wRegInTop_6_51[0] }), .In2(
        {\wRegInBot_6_51[31] , \wRegInBot_6_51[30] , \wRegInBot_6_51[29] , 
        \wRegInBot_6_51[28] , \wRegInBot_6_51[27] , \wRegInBot_6_51[26] , 
        \wRegInBot_6_51[25] , \wRegInBot_6_51[24] , \wRegInBot_6_51[23] , 
        \wRegInBot_6_51[22] , \wRegInBot_6_51[21] , \wRegInBot_6_51[20] , 
        \wRegInBot_6_51[19] , \wRegInBot_6_51[18] , \wRegInBot_6_51[17] , 
        \wRegInBot_6_51[16] , \wRegInBot_6_51[15] , \wRegInBot_6_51[14] , 
        \wRegInBot_6_51[13] , \wRegInBot_6_51[12] , \wRegInBot_6_51[11] , 
        \wRegInBot_6_51[10] , \wRegInBot_6_51[9] , \wRegInBot_6_51[8] , 
        \wRegInBot_6_51[7] , \wRegInBot_6_51[6] , \wRegInBot_6_51[5] , 
        \wRegInBot_6_51[4] , \wRegInBot_6_51[3] , \wRegInBot_6_51[2] , 
        \wRegInBot_6_51[1] , \wRegInBot_6_51[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_19 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink147[31] , \ScanLink147[30] , \ScanLink147[29] , 
        \ScanLink147[28] , \ScanLink147[27] , \ScanLink147[26] , 
        \ScanLink147[25] , \ScanLink147[24] , \ScanLink147[23] , 
        \ScanLink147[22] , \ScanLink147[21] , \ScanLink147[20] , 
        \ScanLink147[19] , \ScanLink147[18] , \ScanLink147[17] , 
        \ScanLink147[16] , \ScanLink147[15] , \ScanLink147[14] , 
        \ScanLink147[13] , \ScanLink147[12] , \ScanLink147[11] , 
        \ScanLink147[10] , \ScanLink147[9] , \ScanLink147[8] , 
        \ScanLink147[7] , \ScanLink147[6] , \ScanLink147[5] , \ScanLink147[4] , 
        \ScanLink147[3] , \ScanLink147[2] , \ScanLink147[1] , \ScanLink147[0] 
        }), .ScanOut({\ScanLink146[31] , \ScanLink146[30] , \ScanLink146[29] , 
        \ScanLink146[28] , \ScanLink146[27] , \ScanLink146[26] , 
        \ScanLink146[25] , \ScanLink146[24] , \ScanLink146[23] , 
        \ScanLink146[22] , \ScanLink146[21] , \ScanLink146[20] , 
        \ScanLink146[19] , \ScanLink146[18] , \ScanLink146[17] , 
        \ScanLink146[16] , \ScanLink146[15] , \ScanLink146[14] , 
        \ScanLink146[13] , \ScanLink146[12] , \ScanLink146[11] , 
        \ScanLink146[10] , \ScanLink146[9] , \ScanLink146[8] , 
        \ScanLink146[7] , \ScanLink146[6] , \ScanLink146[5] , \ScanLink146[4] , 
        \ScanLink146[3] , \ScanLink146[2] , \ScanLink146[1] , \ScanLink146[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_19[31] , 
        \wRegOut_7_19[30] , \wRegOut_7_19[29] , \wRegOut_7_19[28] , 
        \wRegOut_7_19[27] , \wRegOut_7_19[26] , \wRegOut_7_19[25] , 
        \wRegOut_7_19[24] , \wRegOut_7_19[23] , \wRegOut_7_19[22] , 
        \wRegOut_7_19[21] , \wRegOut_7_19[20] , \wRegOut_7_19[19] , 
        \wRegOut_7_19[18] , \wRegOut_7_19[17] , \wRegOut_7_19[16] , 
        \wRegOut_7_19[15] , \wRegOut_7_19[14] , \wRegOut_7_19[13] , 
        \wRegOut_7_19[12] , \wRegOut_7_19[11] , \wRegOut_7_19[10] , 
        \wRegOut_7_19[9] , \wRegOut_7_19[8] , \wRegOut_7_19[7] , 
        \wRegOut_7_19[6] , \wRegOut_7_19[5] , \wRegOut_7_19[4] , 
        \wRegOut_7_19[3] , \wRegOut_7_19[2] , \wRegOut_7_19[1] , 
        \wRegOut_7_19[0] }), .Enable1(\wRegEnTop_7_19[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_19[31] , \wRegInTop_7_19[30] , \wRegInTop_7_19[29] , 
        \wRegInTop_7_19[28] , \wRegInTop_7_19[27] , \wRegInTop_7_19[26] , 
        \wRegInTop_7_19[25] , \wRegInTop_7_19[24] , \wRegInTop_7_19[23] , 
        \wRegInTop_7_19[22] , \wRegInTop_7_19[21] , \wRegInTop_7_19[20] , 
        \wRegInTop_7_19[19] , \wRegInTop_7_19[18] , \wRegInTop_7_19[17] , 
        \wRegInTop_7_19[16] , \wRegInTop_7_19[15] , \wRegInTop_7_19[14] , 
        \wRegInTop_7_19[13] , \wRegInTop_7_19[12] , \wRegInTop_7_19[11] , 
        \wRegInTop_7_19[10] , \wRegInTop_7_19[9] , \wRegInTop_7_19[8] , 
        \wRegInTop_7_19[7] , \wRegInTop_7_19[6] , \wRegInTop_7_19[5] , 
        \wRegInTop_7_19[4] , \wRegInTop_7_19[3] , \wRegInTop_7_19[2] , 
        \wRegInTop_7_19[1] , \wRegInTop_7_19[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_77 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink205[31] , \ScanLink205[30] , \ScanLink205[29] , 
        \ScanLink205[28] , \ScanLink205[27] , \ScanLink205[26] , 
        \ScanLink205[25] , \ScanLink205[24] , \ScanLink205[23] , 
        \ScanLink205[22] , \ScanLink205[21] , \ScanLink205[20] , 
        \ScanLink205[19] , \ScanLink205[18] , \ScanLink205[17] , 
        \ScanLink205[16] , \ScanLink205[15] , \ScanLink205[14] , 
        \ScanLink205[13] , \ScanLink205[12] , \ScanLink205[11] , 
        \ScanLink205[10] , \ScanLink205[9] , \ScanLink205[8] , 
        \ScanLink205[7] , \ScanLink205[6] , \ScanLink205[5] , \ScanLink205[4] , 
        \ScanLink205[3] , \ScanLink205[2] , \ScanLink205[1] , \ScanLink205[0] 
        }), .ScanOut({\ScanLink204[31] , \ScanLink204[30] , \ScanLink204[29] , 
        \ScanLink204[28] , \ScanLink204[27] , \ScanLink204[26] , 
        \ScanLink204[25] , \ScanLink204[24] , \ScanLink204[23] , 
        \ScanLink204[22] , \ScanLink204[21] , \ScanLink204[20] , 
        \ScanLink204[19] , \ScanLink204[18] , \ScanLink204[17] , 
        \ScanLink204[16] , \ScanLink204[15] , \ScanLink204[14] , 
        \ScanLink204[13] , \ScanLink204[12] , \ScanLink204[11] , 
        \ScanLink204[10] , \ScanLink204[9] , \ScanLink204[8] , 
        \ScanLink204[7] , \ScanLink204[6] , \ScanLink204[5] , \ScanLink204[4] , 
        \ScanLink204[3] , \ScanLink204[2] , \ScanLink204[1] , \ScanLink204[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_77[31] , 
        \wRegOut_7_77[30] , \wRegOut_7_77[29] , \wRegOut_7_77[28] , 
        \wRegOut_7_77[27] , \wRegOut_7_77[26] , \wRegOut_7_77[25] , 
        \wRegOut_7_77[24] , \wRegOut_7_77[23] , \wRegOut_7_77[22] , 
        \wRegOut_7_77[21] , \wRegOut_7_77[20] , \wRegOut_7_77[19] , 
        \wRegOut_7_77[18] , \wRegOut_7_77[17] , \wRegOut_7_77[16] , 
        \wRegOut_7_77[15] , \wRegOut_7_77[14] , \wRegOut_7_77[13] , 
        \wRegOut_7_77[12] , \wRegOut_7_77[11] , \wRegOut_7_77[10] , 
        \wRegOut_7_77[9] , \wRegOut_7_77[8] , \wRegOut_7_77[7] , 
        \wRegOut_7_77[6] , \wRegOut_7_77[5] , \wRegOut_7_77[4] , 
        \wRegOut_7_77[3] , \wRegOut_7_77[2] , \wRegOut_7_77[1] , 
        \wRegOut_7_77[0] }), .Enable1(\wRegEnTop_7_77[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_77[31] , \wRegInTop_7_77[30] , \wRegInTop_7_77[29] , 
        \wRegInTop_7_77[28] , \wRegInTop_7_77[27] , \wRegInTop_7_77[26] , 
        \wRegInTop_7_77[25] , \wRegInTop_7_77[24] , \wRegInTop_7_77[23] , 
        \wRegInTop_7_77[22] , \wRegInTop_7_77[21] , \wRegInTop_7_77[20] , 
        \wRegInTop_7_77[19] , \wRegInTop_7_77[18] , \wRegInTop_7_77[17] , 
        \wRegInTop_7_77[16] , \wRegInTop_7_77[15] , \wRegInTop_7_77[14] , 
        \wRegInTop_7_77[13] , \wRegInTop_7_77[12] , \wRegInTop_7_77[11] , 
        \wRegInTop_7_77[10] , \wRegInTop_7_77[9] , \wRegInTop_7_77[8] , 
        \wRegInTop_7_77[7] , \wRegInTop_7_77[6] , \wRegInTop_7_77[5] , 
        \wRegInTop_7_77[4] , \wRegInTop_7_77[3] , \wRegInTop_7_77[2] , 
        \wRegInTop_7_77[1] , \wRegInTop_7_77[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_45[0] ), .P_In({\wRegOut_6_45[31] , 
        \wRegOut_6_45[30] , \wRegOut_6_45[29] , \wRegOut_6_45[28] , 
        \wRegOut_6_45[27] , \wRegOut_6_45[26] , \wRegOut_6_45[25] , 
        \wRegOut_6_45[24] , \wRegOut_6_45[23] , \wRegOut_6_45[22] , 
        \wRegOut_6_45[21] , \wRegOut_6_45[20] , \wRegOut_6_45[19] , 
        \wRegOut_6_45[18] , \wRegOut_6_45[17] , \wRegOut_6_45[16] , 
        \wRegOut_6_45[15] , \wRegOut_6_45[14] , \wRegOut_6_45[13] , 
        \wRegOut_6_45[12] , \wRegOut_6_45[11] , \wRegOut_6_45[10] , 
        \wRegOut_6_45[9] , \wRegOut_6_45[8] , \wRegOut_6_45[7] , 
        \wRegOut_6_45[6] , \wRegOut_6_45[5] , \wRegOut_6_45[4] , 
        \wRegOut_6_45[3] , \wRegOut_6_45[2] , \wRegOut_6_45[1] , 
        \wRegOut_6_45[0] }), .P_Out({\wRegInBot_6_45[31] , 
        \wRegInBot_6_45[30] , \wRegInBot_6_45[29] , \wRegInBot_6_45[28] , 
        \wRegInBot_6_45[27] , \wRegInBot_6_45[26] , \wRegInBot_6_45[25] , 
        \wRegInBot_6_45[24] , \wRegInBot_6_45[23] , \wRegInBot_6_45[22] , 
        \wRegInBot_6_45[21] , \wRegInBot_6_45[20] , \wRegInBot_6_45[19] , 
        \wRegInBot_6_45[18] , \wRegInBot_6_45[17] , \wRegInBot_6_45[16] , 
        \wRegInBot_6_45[15] , \wRegInBot_6_45[14] , \wRegInBot_6_45[13] , 
        \wRegInBot_6_45[12] , \wRegInBot_6_45[11] , \wRegInBot_6_45[10] , 
        \wRegInBot_6_45[9] , \wRegInBot_6_45[8] , \wRegInBot_6_45[7] , 
        \wRegInBot_6_45[6] , \wRegInBot_6_45[5] , \wRegInBot_6_45[4] , 
        \wRegInBot_6_45[3] , \wRegInBot_6_45[2] , \wRegInBot_6_45[1] , 
        \wRegInBot_6_45[0] }), .L_WR(\wRegEnTop_7_90[0] ), .L_In({
        \wRegOut_7_90[31] , \wRegOut_7_90[30] , \wRegOut_7_90[29] , 
        \wRegOut_7_90[28] , \wRegOut_7_90[27] , \wRegOut_7_90[26] , 
        \wRegOut_7_90[25] , \wRegOut_7_90[24] , \wRegOut_7_90[23] , 
        \wRegOut_7_90[22] , \wRegOut_7_90[21] , \wRegOut_7_90[20] , 
        \wRegOut_7_90[19] , \wRegOut_7_90[18] , \wRegOut_7_90[17] , 
        \wRegOut_7_90[16] , \wRegOut_7_90[15] , \wRegOut_7_90[14] , 
        \wRegOut_7_90[13] , \wRegOut_7_90[12] , \wRegOut_7_90[11] , 
        \wRegOut_7_90[10] , \wRegOut_7_90[9] , \wRegOut_7_90[8] , 
        \wRegOut_7_90[7] , \wRegOut_7_90[6] , \wRegOut_7_90[5] , 
        \wRegOut_7_90[4] , \wRegOut_7_90[3] , \wRegOut_7_90[2] , 
        \wRegOut_7_90[1] , \wRegOut_7_90[0] }), .L_Out({\wRegInTop_7_90[31] , 
        \wRegInTop_7_90[30] , \wRegInTop_7_90[29] , \wRegInTop_7_90[28] , 
        \wRegInTop_7_90[27] , \wRegInTop_7_90[26] , \wRegInTop_7_90[25] , 
        \wRegInTop_7_90[24] , \wRegInTop_7_90[23] , \wRegInTop_7_90[22] , 
        \wRegInTop_7_90[21] , \wRegInTop_7_90[20] , \wRegInTop_7_90[19] , 
        \wRegInTop_7_90[18] , \wRegInTop_7_90[17] , \wRegInTop_7_90[16] , 
        \wRegInTop_7_90[15] , \wRegInTop_7_90[14] , \wRegInTop_7_90[13] , 
        \wRegInTop_7_90[12] , \wRegInTop_7_90[11] , \wRegInTop_7_90[10] , 
        \wRegInTop_7_90[9] , \wRegInTop_7_90[8] , \wRegInTop_7_90[7] , 
        \wRegInTop_7_90[6] , \wRegInTop_7_90[5] , \wRegInTop_7_90[4] , 
        \wRegInTop_7_90[3] , \wRegInTop_7_90[2] , \wRegInTop_7_90[1] , 
        \wRegInTop_7_90[0] }), .R_WR(\wRegEnTop_7_91[0] ), .R_In({
        \wRegOut_7_91[31] , \wRegOut_7_91[30] , \wRegOut_7_91[29] , 
        \wRegOut_7_91[28] , \wRegOut_7_91[27] , \wRegOut_7_91[26] , 
        \wRegOut_7_91[25] , \wRegOut_7_91[24] , \wRegOut_7_91[23] , 
        \wRegOut_7_91[22] , \wRegOut_7_91[21] , \wRegOut_7_91[20] , 
        \wRegOut_7_91[19] , \wRegOut_7_91[18] , \wRegOut_7_91[17] , 
        \wRegOut_7_91[16] , \wRegOut_7_91[15] , \wRegOut_7_91[14] , 
        \wRegOut_7_91[13] , \wRegOut_7_91[12] , \wRegOut_7_91[11] , 
        \wRegOut_7_91[10] , \wRegOut_7_91[9] , \wRegOut_7_91[8] , 
        \wRegOut_7_91[7] , \wRegOut_7_91[6] , \wRegOut_7_91[5] , 
        \wRegOut_7_91[4] , \wRegOut_7_91[3] , \wRegOut_7_91[2] , 
        \wRegOut_7_91[1] , \wRegOut_7_91[0] }), .R_Out({\wRegInTop_7_91[31] , 
        \wRegInTop_7_91[30] , \wRegInTop_7_91[29] , \wRegInTop_7_91[28] , 
        \wRegInTop_7_91[27] , \wRegInTop_7_91[26] , \wRegInTop_7_91[25] , 
        \wRegInTop_7_91[24] , \wRegInTop_7_91[23] , \wRegInTop_7_91[22] , 
        \wRegInTop_7_91[21] , \wRegInTop_7_91[20] , \wRegInTop_7_91[19] , 
        \wRegInTop_7_91[18] , \wRegInTop_7_91[17] , \wRegInTop_7_91[16] , 
        \wRegInTop_7_91[15] , \wRegInTop_7_91[14] , \wRegInTop_7_91[13] , 
        \wRegInTop_7_91[12] , \wRegInTop_7_91[11] , \wRegInTop_7_91[10] , 
        \wRegInTop_7_91[9] , \wRegInTop_7_91[8] , \wRegInTop_7_91[7] , 
        \wRegInTop_7_91[6] , \wRegInTop_7_91[5] , \wRegInTop_7_91[4] , 
        \wRegInTop_7_91[3] , \wRegInTop_7_91[2] , \wRegInTop_7_91[1] , 
        \wRegInTop_7_91[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_89 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink217[31] , \ScanLink217[30] , \ScanLink217[29] , 
        \ScanLink217[28] , \ScanLink217[27] , \ScanLink217[26] , 
        \ScanLink217[25] , \ScanLink217[24] , \ScanLink217[23] , 
        \ScanLink217[22] , \ScanLink217[21] , \ScanLink217[20] , 
        \ScanLink217[19] , \ScanLink217[18] , \ScanLink217[17] , 
        \ScanLink217[16] , \ScanLink217[15] , \ScanLink217[14] , 
        \ScanLink217[13] , \ScanLink217[12] , \ScanLink217[11] , 
        \ScanLink217[10] , \ScanLink217[9] , \ScanLink217[8] , 
        \ScanLink217[7] , \ScanLink217[6] , \ScanLink217[5] , \ScanLink217[4] , 
        \ScanLink217[3] , \ScanLink217[2] , \ScanLink217[1] , \ScanLink217[0] 
        }), .ScanOut({\ScanLink216[31] , \ScanLink216[30] , \ScanLink216[29] , 
        \ScanLink216[28] , \ScanLink216[27] , \ScanLink216[26] , 
        \ScanLink216[25] , \ScanLink216[24] , \ScanLink216[23] , 
        \ScanLink216[22] , \ScanLink216[21] , \ScanLink216[20] , 
        \ScanLink216[19] , \ScanLink216[18] , \ScanLink216[17] , 
        \ScanLink216[16] , \ScanLink216[15] , \ScanLink216[14] , 
        \ScanLink216[13] , \ScanLink216[12] , \ScanLink216[11] , 
        \ScanLink216[10] , \ScanLink216[9] , \ScanLink216[8] , 
        \ScanLink216[7] , \ScanLink216[6] , \ScanLink216[5] , \ScanLink216[4] , 
        \ScanLink216[3] , \ScanLink216[2] , \ScanLink216[1] , \ScanLink216[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_89[31] , 
        \wRegOut_7_89[30] , \wRegOut_7_89[29] , \wRegOut_7_89[28] , 
        \wRegOut_7_89[27] , \wRegOut_7_89[26] , \wRegOut_7_89[25] , 
        \wRegOut_7_89[24] , \wRegOut_7_89[23] , \wRegOut_7_89[22] , 
        \wRegOut_7_89[21] , \wRegOut_7_89[20] , \wRegOut_7_89[19] , 
        \wRegOut_7_89[18] , \wRegOut_7_89[17] , \wRegOut_7_89[16] , 
        \wRegOut_7_89[15] , \wRegOut_7_89[14] , \wRegOut_7_89[13] , 
        \wRegOut_7_89[12] , \wRegOut_7_89[11] , \wRegOut_7_89[10] , 
        \wRegOut_7_89[9] , \wRegOut_7_89[8] , \wRegOut_7_89[7] , 
        \wRegOut_7_89[6] , \wRegOut_7_89[5] , \wRegOut_7_89[4] , 
        \wRegOut_7_89[3] , \wRegOut_7_89[2] , \wRegOut_7_89[1] , 
        \wRegOut_7_89[0] }), .Enable1(\wRegEnTop_7_89[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_89[31] , \wRegInTop_7_89[30] , \wRegInTop_7_89[29] , 
        \wRegInTop_7_89[28] , \wRegInTop_7_89[27] , \wRegInTop_7_89[26] , 
        \wRegInTop_7_89[25] , \wRegInTop_7_89[24] , \wRegInTop_7_89[23] , 
        \wRegInTop_7_89[22] , \wRegInTop_7_89[21] , \wRegInTop_7_89[20] , 
        \wRegInTop_7_89[19] , \wRegInTop_7_89[18] , \wRegInTop_7_89[17] , 
        \wRegInTop_7_89[16] , \wRegInTop_7_89[15] , \wRegInTop_7_89[14] , 
        \wRegInTop_7_89[13] , \wRegInTop_7_89[12] , \wRegInTop_7_89[11] , 
        \wRegInTop_7_89[10] , \wRegInTop_7_89[9] , \wRegInTop_7_89[8] , 
        \wRegInTop_7_89[7] , \wRegInTop_7_89[6] , \wRegInTop_7_89[5] , 
        \wRegInTop_7_89[4] , \wRegInTop_7_89[3] , \wRegInTop_7_89[2] , 
        \wRegInTop_7_89[1] , \wRegInTop_7_89[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_92 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink220[31] , \ScanLink220[30] , \ScanLink220[29] , 
        \ScanLink220[28] , \ScanLink220[27] , \ScanLink220[26] , 
        \ScanLink220[25] , \ScanLink220[24] , \ScanLink220[23] , 
        \ScanLink220[22] , \ScanLink220[21] , \ScanLink220[20] , 
        \ScanLink220[19] , \ScanLink220[18] , \ScanLink220[17] , 
        \ScanLink220[16] , \ScanLink220[15] , \ScanLink220[14] , 
        \ScanLink220[13] , \ScanLink220[12] , \ScanLink220[11] , 
        \ScanLink220[10] , \ScanLink220[9] , \ScanLink220[8] , 
        \ScanLink220[7] , \ScanLink220[6] , \ScanLink220[5] , \ScanLink220[4] , 
        \ScanLink220[3] , \ScanLink220[2] , \ScanLink220[1] , \ScanLink220[0] 
        }), .ScanOut({\ScanLink219[31] , \ScanLink219[30] , \ScanLink219[29] , 
        \ScanLink219[28] , \ScanLink219[27] , \ScanLink219[26] , 
        \ScanLink219[25] , \ScanLink219[24] , \ScanLink219[23] , 
        \ScanLink219[22] , \ScanLink219[21] , \ScanLink219[20] , 
        \ScanLink219[19] , \ScanLink219[18] , \ScanLink219[17] , 
        \ScanLink219[16] , \ScanLink219[15] , \ScanLink219[14] , 
        \ScanLink219[13] , \ScanLink219[12] , \ScanLink219[11] , 
        \ScanLink219[10] , \ScanLink219[9] , \ScanLink219[8] , 
        \ScanLink219[7] , \ScanLink219[6] , \ScanLink219[5] , \ScanLink219[4] , 
        \ScanLink219[3] , \ScanLink219[2] , \ScanLink219[1] , \ScanLink219[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_92[31] , 
        \wRegOut_7_92[30] , \wRegOut_7_92[29] , \wRegOut_7_92[28] , 
        \wRegOut_7_92[27] , \wRegOut_7_92[26] , \wRegOut_7_92[25] , 
        \wRegOut_7_92[24] , \wRegOut_7_92[23] , \wRegOut_7_92[22] , 
        \wRegOut_7_92[21] , \wRegOut_7_92[20] , \wRegOut_7_92[19] , 
        \wRegOut_7_92[18] , \wRegOut_7_92[17] , \wRegOut_7_92[16] , 
        \wRegOut_7_92[15] , \wRegOut_7_92[14] , \wRegOut_7_92[13] , 
        \wRegOut_7_92[12] , \wRegOut_7_92[11] , \wRegOut_7_92[10] , 
        \wRegOut_7_92[9] , \wRegOut_7_92[8] , \wRegOut_7_92[7] , 
        \wRegOut_7_92[6] , \wRegOut_7_92[5] , \wRegOut_7_92[4] , 
        \wRegOut_7_92[3] , \wRegOut_7_92[2] , \wRegOut_7_92[1] , 
        \wRegOut_7_92[0] }), .Enable1(\wRegEnTop_7_92[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_92[31] , \wRegInTop_7_92[30] , \wRegInTop_7_92[29] , 
        \wRegInTop_7_92[28] , \wRegInTop_7_92[27] , \wRegInTop_7_92[26] , 
        \wRegInTop_7_92[25] , \wRegInTop_7_92[24] , \wRegInTop_7_92[23] , 
        \wRegInTop_7_92[22] , \wRegInTop_7_92[21] , \wRegInTop_7_92[20] , 
        \wRegInTop_7_92[19] , \wRegInTop_7_92[18] , \wRegInTop_7_92[17] , 
        \wRegInTop_7_92[16] , \wRegInTop_7_92[15] , \wRegInTop_7_92[14] , 
        \wRegInTop_7_92[13] , \wRegInTop_7_92[12] , \wRegInTop_7_92[11] , 
        \wRegInTop_7_92[10] , \wRegInTop_7_92[9] , \wRegInTop_7_92[8] , 
        \wRegInTop_7_92[7] , \wRegInTop_7_92[6] , \wRegInTop_7_92[5] , 
        \wRegInTop_7_92[4] , \wRegInTop_7_92[3] , \wRegInTop_7_92[2] , 
        \wRegInTop_7_92[1] , \wRegInTop_7_92[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_3[0] ), .P_In({\wRegOut_5_3[31] , 
        \wRegOut_5_3[30] , \wRegOut_5_3[29] , \wRegOut_5_3[28] , 
        \wRegOut_5_3[27] , \wRegOut_5_3[26] , \wRegOut_5_3[25] , 
        \wRegOut_5_3[24] , \wRegOut_5_3[23] , \wRegOut_5_3[22] , 
        \wRegOut_5_3[21] , \wRegOut_5_3[20] , \wRegOut_5_3[19] , 
        \wRegOut_5_3[18] , \wRegOut_5_3[17] , \wRegOut_5_3[16] , 
        \wRegOut_5_3[15] , \wRegOut_5_3[14] , \wRegOut_5_3[13] , 
        \wRegOut_5_3[12] , \wRegOut_5_3[11] , \wRegOut_5_3[10] , 
        \wRegOut_5_3[9] , \wRegOut_5_3[8] , \wRegOut_5_3[7] , \wRegOut_5_3[6] , 
        \wRegOut_5_3[5] , \wRegOut_5_3[4] , \wRegOut_5_3[3] , \wRegOut_5_3[2] , 
        \wRegOut_5_3[1] , \wRegOut_5_3[0] }), .P_Out({\wRegInBot_5_3[31] , 
        \wRegInBot_5_3[30] , \wRegInBot_5_3[29] , \wRegInBot_5_3[28] , 
        \wRegInBot_5_3[27] , \wRegInBot_5_3[26] , \wRegInBot_5_3[25] , 
        \wRegInBot_5_3[24] , \wRegInBot_5_3[23] , \wRegInBot_5_3[22] , 
        \wRegInBot_5_3[21] , \wRegInBot_5_3[20] , \wRegInBot_5_3[19] , 
        \wRegInBot_5_3[18] , \wRegInBot_5_3[17] , \wRegInBot_5_3[16] , 
        \wRegInBot_5_3[15] , \wRegInBot_5_3[14] , \wRegInBot_5_3[13] , 
        \wRegInBot_5_3[12] , \wRegInBot_5_3[11] , \wRegInBot_5_3[10] , 
        \wRegInBot_5_3[9] , \wRegInBot_5_3[8] , \wRegInBot_5_3[7] , 
        \wRegInBot_5_3[6] , \wRegInBot_5_3[5] , \wRegInBot_5_3[4] , 
        \wRegInBot_5_3[3] , \wRegInBot_5_3[2] , \wRegInBot_5_3[1] , 
        \wRegInBot_5_3[0] }), .L_WR(\wRegEnTop_6_6[0] ), .L_In({
        \wRegOut_6_6[31] , \wRegOut_6_6[30] , \wRegOut_6_6[29] , 
        \wRegOut_6_6[28] , \wRegOut_6_6[27] , \wRegOut_6_6[26] , 
        \wRegOut_6_6[25] , \wRegOut_6_6[24] , \wRegOut_6_6[23] , 
        \wRegOut_6_6[22] , \wRegOut_6_6[21] , \wRegOut_6_6[20] , 
        \wRegOut_6_6[19] , \wRegOut_6_6[18] , \wRegOut_6_6[17] , 
        \wRegOut_6_6[16] , \wRegOut_6_6[15] , \wRegOut_6_6[14] , 
        \wRegOut_6_6[13] , \wRegOut_6_6[12] , \wRegOut_6_6[11] , 
        \wRegOut_6_6[10] , \wRegOut_6_6[9] , \wRegOut_6_6[8] , 
        \wRegOut_6_6[7] , \wRegOut_6_6[6] , \wRegOut_6_6[5] , \wRegOut_6_6[4] , 
        \wRegOut_6_6[3] , \wRegOut_6_6[2] , \wRegOut_6_6[1] , \wRegOut_6_6[0] 
        }), .L_Out({\wRegInTop_6_6[31] , \wRegInTop_6_6[30] , 
        \wRegInTop_6_6[29] , \wRegInTop_6_6[28] , \wRegInTop_6_6[27] , 
        \wRegInTop_6_6[26] , \wRegInTop_6_6[25] , \wRegInTop_6_6[24] , 
        \wRegInTop_6_6[23] , \wRegInTop_6_6[22] , \wRegInTop_6_6[21] , 
        \wRegInTop_6_6[20] , \wRegInTop_6_6[19] , \wRegInTop_6_6[18] , 
        \wRegInTop_6_6[17] , \wRegInTop_6_6[16] , \wRegInTop_6_6[15] , 
        \wRegInTop_6_6[14] , \wRegInTop_6_6[13] , \wRegInTop_6_6[12] , 
        \wRegInTop_6_6[11] , \wRegInTop_6_6[10] , \wRegInTop_6_6[9] , 
        \wRegInTop_6_6[8] , \wRegInTop_6_6[7] , \wRegInTop_6_6[6] , 
        \wRegInTop_6_6[5] , \wRegInTop_6_6[4] , \wRegInTop_6_6[3] , 
        \wRegInTop_6_6[2] , \wRegInTop_6_6[1] , \wRegInTop_6_6[0] }), .R_WR(
        \wRegEnTop_6_7[0] ), .R_In({\wRegOut_6_7[31] , \wRegOut_6_7[30] , 
        \wRegOut_6_7[29] , \wRegOut_6_7[28] , \wRegOut_6_7[27] , 
        \wRegOut_6_7[26] , \wRegOut_6_7[25] , \wRegOut_6_7[24] , 
        \wRegOut_6_7[23] , \wRegOut_6_7[22] , \wRegOut_6_7[21] , 
        \wRegOut_6_7[20] , \wRegOut_6_7[19] , \wRegOut_6_7[18] , 
        \wRegOut_6_7[17] , \wRegOut_6_7[16] , \wRegOut_6_7[15] , 
        \wRegOut_6_7[14] , \wRegOut_6_7[13] , \wRegOut_6_7[12] , 
        \wRegOut_6_7[11] , \wRegOut_6_7[10] , \wRegOut_6_7[9] , 
        \wRegOut_6_7[8] , \wRegOut_6_7[7] , \wRegOut_6_7[6] , \wRegOut_6_7[5] , 
        \wRegOut_6_7[4] , \wRegOut_6_7[3] , \wRegOut_6_7[2] , \wRegOut_6_7[1] , 
        \wRegOut_6_7[0] }), .R_Out({\wRegInTop_6_7[31] , \wRegInTop_6_7[30] , 
        \wRegInTop_6_7[29] , \wRegInTop_6_7[28] , \wRegInTop_6_7[27] , 
        \wRegInTop_6_7[26] , \wRegInTop_6_7[25] , \wRegInTop_6_7[24] , 
        \wRegInTop_6_7[23] , \wRegInTop_6_7[22] , \wRegInTop_6_7[21] , 
        \wRegInTop_6_7[20] , \wRegInTop_6_7[19] , \wRegInTop_6_7[18] , 
        \wRegInTop_6_7[17] , \wRegInTop_6_7[16] , \wRegInTop_6_7[15] , 
        \wRegInTop_6_7[14] , \wRegInTop_6_7[13] , \wRegInTop_6_7[12] , 
        \wRegInTop_6_7[11] , \wRegInTop_6_7[10] , \wRegInTop_6_7[9] , 
        \wRegInTop_6_7[8] , \wRegInTop_6_7[7] , \wRegInTop_6_7[6] , 
        \wRegInTop_6_7[5] , \wRegInTop_6_7[4] , \wRegInTop_6_7[3] , 
        \wRegInTop_6_7[2] , \wRegInTop_6_7[1] , \wRegInTop_6_7[0] }) );
    BHeap_Node_WIDTH32 BHN_6_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_62[0] ), .P_In({\wRegOut_6_62[31] , 
        \wRegOut_6_62[30] , \wRegOut_6_62[29] , \wRegOut_6_62[28] , 
        \wRegOut_6_62[27] , \wRegOut_6_62[26] , \wRegOut_6_62[25] , 
        \wRegOut_6_62[24] , \wRegOut_6_62[23] , \wRegOut_6_62[22] , 
        \wRegOut_6_62[21] , \wRegOut_6_62[20] , \wRegOut_6_62[19] , 
        \wRegOut_6_62[18] , \wRegOut_6_62[17] , \wRegOut_6_62[16] , 
        \wRegOut_6_62[15] , \wRegOut_6_62[14] , \wRegOut_6_62[13] , 
        \wRegOut_6_62[12] , \wRegOut_6_62[11] , \wRegOut_6_62[10] , 
        \wRegOut_6_62[9] , \wRegOut_6_62[8] , \wRegOut_6_62[7] , 
        \wRegOut_6_62[6] , \wRegOut_6_62[5] , \wRegOut_6_62[4] , 
        \wRegOut_6_62[3] , \wRegOut_6_62[2] , \wRegOut_6_62[1] , 
        \wRegOut_6_62[0] }), .P_Out({\wRegInBot_6_62[31] , 
        \wRegInBot_6_62[30] , \wRegInBot_6_62[29] , \wRegInBot_6_62[28] , 
        \wRegInBot_6_62[27] , \wRegInBot_6_62[26] , \wRegInBot_6_62[25] , 
        \wRegInBot_6_62[24] , \wRegInBot_6_62[23] , \wRegInBot_6_62[22] , 
        \wRegInBot_6_62[21] , \wRegInBot_6_62[20] , \wRegInBot_6_62[19] , 
        \wRegInBot_6_62[18] , \wRegInBot_6_62[17] , \wRegInBot_6_62[16] , 
        \wRegInBot_6_62[15] , \wRegInBot_6_62[14] , \wRegInBot_6_62[13] , 
        \wRegInBot_6_62[12] , \wRegInBot_6_62[11] , \wRegInBot_6_62[10] , 
        \wRegInBot_6_62[9] , \wRegInBot_6_62[8] , \wRegInBot_6_62[7] , 
        \wRegInBot_6_62[6] , \wRegInBot_6_62[5] , \wRegInBot_6_62[4] , 
        \wRegInBot_6_62[3] , \wRegInBot_6_62[2] , \wRegInBot_6_62[1] , 
        \wRegInBot_6_62[0] }), .L_WR(\wRegEnTop_7_124[0] ), .L_In({
        \wRegOut_7_124[31] , \wRegOut_7_124[30] , \wRegOut_7_124[29] , 
        \wRegOut_7_124[28] , \wRegOut_7_124[27] , \wRegOut_7_124[26] , 
        \wRegOut_7_124[25] , \wRegOut_7_124[24] , \wRegOut_7_124[23] , 
        \wRegOut_7_124[22] , \wRegOut_7_124[21] , \wRegOut_7_124[20] , 
        \wRegOut_7_124[19] , \wRegOut_7_124[18] , \wRegOut_7_124[17] , 
        \wRegOut_7_124[16] , \wRegOut_7_124[15] , \wRegOut_7_124[14] , 
        \wRegOut_7_124[13] , \wRegOut_7_124[12] , \wRegOut_7_124[11] , 
        \wRegOut_7_124[10] , \wRegOut_7_124[9] , \wRegOut_7_124[8] , 
        \wRegOut_7_124[7] , \wRegOut_7_124[6] , \wRegOut_7_124[5] , 
        \wRegOut_7_124[4] , \wRegOut_7_124[3] , \wRegOut_7_124[2] , 
        \wRegOut_7_124[1] , \wRegOut_7_124[0] }), .L_Out({
        \wRegInTop_7_124[31] , \wRegInTop_7_124[30] , \wRegInTop_7_124[29] , 
        \wRegInTop_7_124[28] , \wRegInTop_7_124[27] , \wRegInTop_7_124[26] , 
        \wRegInTop_7_124[25] , \wRegInTop_7_124[24] , \wRegInTop_7_124[23] , 
        \wRegInTop_7_124[22] , \wRegInTop_7_124[21] , \wRegInTop_7_124[20] , 
        \wRegInTop_7_124[19] , \wRegInTop_7_124[18] , \wRegInTop_7_124[17] , 
        \wRegInTop_7_124[16] , \wRegInTop_7_124[15] , \wRegInTop_7_124[14] , 
        \wRegInTop_7_124[13] , \wRegInTop_7_124[12] , \wRegInTop_7_124[11] , 
        \wRegInTop_7_124[10] , \wRegInTop_7_124[9] , \wRegInTop_7_124[8] , 
        \wRegInTop_7_124[7] , \wRegInTop_7_124[6] , \wRegInTop_7_124[5] , 
        \wRegInTop_7_124[4] , \wRegInTop_7_124[3] , \wRegInTop_7_124[2] , 
        \wRegInTop_7_124[1] , \wRegInTop_7_124[0] }), .R_WR(
        \wRegEnTop_7_125[0] ), .R_In({\wRegOut_7_125[31] , \wRegOut_7_125[30] , 
        \wRegOut_7_125[29] , \wRegOut_7_125[28] , \wRegOut_7_125[27] , 
        \wRegOut_7_125[26] , \wRegOut_7_125[25] , \wRegOut_7_125[24] , 
        \wRegOut_7_125[23] , \wRegOut_7_125[22] , \wRegOut_7_125[21] , 
        \wRegOut_7_125[20] , \wRegOut_7_125[19] , \wRegOut_7_125[18] , 
        \wRegOut_7_125[17] , \wRegOut_7_125[16] , \wRegOut_7_125[15] , 
        \wRegOut_7_125[14] , \wRegOut_7_125[13] , \wRegOut_7_125[12] , 
        \wRegOut_7_125[11] , \wRegOut_7_125[10] , \wRegOut_7_125[9] , 
        \wRegOut_7_125[8] , \wRegOut_7_125[7] , \wRegOut_7_125[6] , 
        \wRegOut_7_125[5] , \wRegOut_7_125[4] , \wRegOut_7_125[3] , 
        \wRegOut_7_125[2] , \wRegOut_7_125[1] , \wRegOut_7_125[0] }), .R_Out({
        \wRegInTop_7_125[31] , \wRegInTop_7_125[30] , \wRegInTop_7_125[29] , 
        \wRegInTop_7_125[28] , \wRegInTop_7_125[27] , \wRegInTop_7_125[26] , 
        \wRegInTop_7_125[25] , \wRegInTop_7_125[24] , \wRegInTop_7_125[23] , 
        \wRegInTop_7_125[22] , \wRegInTop_7_125[21] , \wRegInTop_7_125[20] , 
        \wRegInTop_7_125[19] , \wRegInTop_7_125[18] , \wRegInTop_7_125[17] , 
        \wRegInTop_7_125[16] , \wRegInTop_7_125[15] , \wRegInTop_7_125[14] , 
        \wRegInTop_7_125[13] , \wRegInTop_7_125[12] , \wRegInTop_7_125[11] , 
        \wRegInTop_7_125[10] , \wRegInTop_7_125[9] , \wRegInTop_7_125[8] , 
        \wRegInTop_7_125[7] , \wRegInTop_7_125[6] , \wRegInTop_7_125[5] , 
        \wRegInTop_7_125[4] , \wRegInTop_7_125[3] , \wRegInTop_7_125[2] , 
        \wRegInTop_7_125[1] , \wRegInTop_7_125[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink33[31] , \ScanLink33[30] , \ScanLink33[29] , 
        \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , \ScanLink33[25] , 
        \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , \ScanLink33[21] , 
        \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , \ScanLink33[17] , 
        \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , \ScanLink33[13] , 
        \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , \ScanLink33[9] , 
        \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , \ScanLink33[5] , 
        \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , \ScanLink33[1] , 
        \ScanLink33[0] }), .ScanOut({\ScanLink32[31] , \ScanLink32[30] , 
        \ScanLink32[29] , \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , 
        \ScanLink32[25] , \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , 
        \ScanLink32[21] , \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , 
        \ScanLink32[17] , \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , 
        \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , 
        \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , 
        \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , 
        \ScanLink32[1] , \ScanLink32[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_1[31] , \wRegOut_5_1[30] , \wRegOut_5_1[29] , 
        \wRegOut_5_1[28] , \wRegOut_5_1[27] , \wRegOut_5_1[26] , 
        \wRegOut_5_1[25] , \wRegOut_5_1[24] , \wRegOut_5_1[23] , 
        \wRegOut_5_1[22] , \wRegOut_5_1[21] , \wRegOut_5_1[20] , 
        \wRegOut_5_1[19] , \wRegOut_5_1[18] , \wRegOut_5_1[17] , 
        \wRegOut_5_1[16] , \wRegOut_5_1[15] , \wRegOut_5_1[14] , 
        \wRegOut_5_1[13] , \wRegOut_5_1[12] , \wRegOut_5_1[11] , 
        \wRegOut_5_1[10] , \wRegOut_5_1[9] , \wRegOut_5_1[8] , 
        \wRegOut_5_1[7] , \wRegOut_5_1[6] , \wRegOut_5_1[5] , \wRegOut_5_1[4] , 
        \wRegOut_5_1[3] , \wRegOut_5_1[2] , \wRegOut_5_1[1] , \wRegOut_5_1[0] 
        }), .Enable1(\wRegEnTop_5_1[0] ), .Enable2(\wRegEnBot_5_1[0] ), .In1({
        \wRegInTop_5_1[31] , \wRegInTop_5_1[30] , \wRegInTop_5_1[29] , 
        \wRegInTop_5_1[28] , \wRegInTop_5_1[27] , \wRegInTop_5_1[26] , 
        \wRegInTop_5_1[25] , \wRegInTop_5_1[24] , \wRegInTop_5_1[23] , 
        \wRegInTop_5_1[22] , \wRegInTop_5_1[21] , \wRegInTop_5_1[20] , 
        \wRegInTop_5_1[19] , \wRegInTop_5_1[18] , \wRegInTop_5_1[17] , 
        \wRegInTop_5_1[16] , \wRegInTop_5_1[15] , \wRegInTop_5_1[14] , 
        \wRegInTop_5_1[13] , \wRegInTop_5_1[12] , \wRegInTop_5_1[11] , 
        \wRegInTop_5_1[10] , \wRegInTop_5_1[9] , \wRegInTop_5_1[8] , 
        \wRegInTop_5_1[7] , \wRegInTop_5_1[6] , \wRegInTop_5_1[5] , 
        \wRegInTop_5_1[4] , \wRegInTop_5_1[3] , \wRegInTop_5_1[2] , 
        \wRegInTop_5_1[1] , \wRegInTop_5_1[0] }), .In2({\wRegInBot_5_1[31] , 
        \wRegInBot_5_1[30] , \wRegInBot_5_1[29] , \wRegInBot_5_1[28] , 
        \wRegInBot_5_1[27] , \wRegInBot_5_1[26] , \wRegInBot_5_1[25] , 
        \wRegInBot_5_1[24] , \wRegInBot_5_1[23] , \wRegInBot_5_1[22] , 
        \wRegInBot_5_1[21] , \wRegInBot_5_1[20] , \wRegInBot_5_1[19] , 
        \wRegInBot_5_1[18] , \wRegInBot_5_1[17] , \wRegInBot_5_1[16] , 
        \wRegInBot_5_1[15] , \wRegInBot_5_1[14] , \wRegInBot_5_1[13] , 
        \wRegInBot_5_1[12] , \wRegInBot_5_1[11] , \wRegInBot_5_1[10] , 
        \wRegInBot_5_1[9] , \wRegInBot_5_1[8] , \wRegInBot_5_1[7] , 
        \wRegInBot_5_1[6] , \wRegInBot_5_1[5] , \wRegInBot_5_1[4] , 
        \wRegInBot_5_1[3] , \wRegInBot_5_1[2] , \wRegInBot_5_1[1] , 
        \wRegInBot_5_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_28 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink60[31] , \ScanLink60[30] , \ScanLink60[29] , 
        \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , \ScanLink60[25] , 
        \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , \ScanLink60[21] , 
        \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , \ScanLink60[17] , 
        \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , \ScanLink60[13] , 
        \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , \ScanLink60[9] , 
        \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , \ScanLink60[5] , 
        \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , \ScanLink60[1] , 
        \ScanLink60[0] }), .ScanOut({\ScanLink59[31] , \ScanLink59[30] , 
        \ScanLink59[29] , \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , 
        \ScanLink59[25] , \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , 
        \ScanLink59[21] , \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , 
        \ScanLink59[17] , \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , 
        \ScanLink59[13] , \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , 
        \ScanLink59[9] , \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , 
        \ScanLink59[5] , \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , 
        \ScanLink59[1] , \ScanLink59[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_28[31] , \wRegOut_5_28[30] , 
        \wRegOut_5_28[29] , \wRegOut_5_28[28] , \wRegOut_5_28[27] , 
        \wRegOut_5_28[26] , \wRegOut_5_28[25] , \wRegOut_5_28[24] , 
        \wRegOut_5_28[23] , \wRegOut_5_28[22] , \wRegOut_5_28[21] , 
        \wRegOut_5_28[20] , \wRegOut_5_28[19] , \wRegOut_5_28[18] , 
        \wRegOut_5_28[17] , \wRegOut_5_28[16] , \wRegOut_5_28[15] , 
        \wRegOut_5_28[14] , \wRegOut_5_28[13] , \wRegOut_5_28[12] , 
        \wRegOut_5_28[11] , \wRegOut_5_28[10] , \wRegOut_5_28[9] , 
        \wRegOut_5_28[8] , \wRegOut_5_28[7] , \wRegOut_5_28[6] , 
        \wRegOut_5_28[5] , \wRegOut_5_28[4] , \wRegOut_5_28[3] , 
        \wRegOut_5_28[2] , \wRegOut_5_28[1] , \wRegOut_5_28[0] }), .Enable1(
        \wRegEnTop_5_28[0] ), .Enable2(\wRegEnBot_5_28[0] ), .In1({
        \wRegInTop_5_28[31] , \wRegInTop_5_28[30] , \wRegInTop_5_28[29] , 
        \wRegInTop_5_28[28] , \wRegInTop_5_28[27] , \wRegInTop_5_28[26] , 
        \wRegInTop_5_28[25] , \wRegInTop_5_28[24] , \wRegInTop_5_28[23] , 
        \wRegInTop_5_28[22] , \wRegInTop_5_28[21] , \wRegInTop_5_28[20] , 
        \wRegInTop_5_28[19] , \wRegInTop_5_28[18] , \wRegInTop_5_28[17] , 
        \wRegInTop_5_28[16] , \wRegInTop_5_28[15] , \wRegInTop_5_28[14] , 
        \wRegInTop_5_28[13] , \wRegInTop_5_28[12] , \wRegInTop_5_28[11] , 
        \wRegInTop_5_28[10] , \wRegInTop_5_28[9] , \wRegInTop_5_28[8] , 
        \wRegInTop_5_28[7] , \wRegInTop_5_28[6] , \wRegInTop_5_28[5] , 
        \wRegInTop_5_28[4] , \wRegInTop_5_28[3] , \wRegInTop_5_28[2] , 
        \wRegInTop_5_28[1] , \wRegInTop_5_28[0] }), .In2({\wRegInBot_5_28[31] , 
        \wRegInBot_5_28[30] , \wRegInBot_5_28[29] , \wRegInBot_5_28[28] , 
        \wRegInBot_5_28[27] , \wRegInBot_5_28[26] , \wRegInBot_5_28[25] , 
        \wRegInBot_5_28[24] , \wRegInBot_5_28[23] , \wRegInBot_5_28[22] , 
        \wRegInBot_5_28[21] , \wRegInBot_5_28[20] , \wRegInBot_5_28[19] , 
        \wRegInBot_5_28[18] , \wRegInBot_5_28[17] , \wRegInBot_5_28[16] , 
        \wRegInBot_5_28[15] , \wRegInBot_5_28[14] , \wRegInBot_5_28[13] , 
        \wRegInBot_5_28[12] , \wRegInBot_5_28[11] , \wRegInBot_5_28[10] , 
        \wRegInBot_5_28[9] , \wRegInBot_5_28[8] , \wRegInBot_5_28[7] , 
        \wRegInBot_5_28[6] , \wRegInBot_5_28[5] , \wRegInBot_5_28[4] , 
        \wRegInBot_5_28[3] , \wRegInBot_5_28[2] , \wRegInBot_5_28[1] , 
        \wRegInBot_5_28[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_18 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink82[31] , \ScanLink82[30] , \ScanLink82[29] , 
        \ScanLink82[28] , \ScanLink82[27] , \ScanLink82[26] , \ScanLink82[25] , 
        \ScanLink82[24] , \ScanLink82[23] , \ScanLink82[22] , \ScanLink82[21] , 
        \ScanLink82[20] , \ScanLink82[19] , \ScanLink82[18] , \ScanLink82[17] , 
        \ScanLink82[16] , \ScanLink82[15] , \ScanLink82[14] , \ScanLink82[13] , 
        \ScanLink82[12] , \ScanLink82[11] , \ScanLink82[10] , \ScanLink82[9] , 
        \ScanLink82[8] , \ScanLink82[7] , \ScanLink82[6] , \ScanLink82[5] , 
        \ScanLink82[4] , \ScanLink82[3] , \ScanLink82[2] , \ScanLink82[1] , 
        \ScanLink82[0] }), .ScanOut({\ScanLink81[31] , \ScanLink81[30] , 
        \ScanLink81[29] , \ScanLink81[28] , \ScanLink81[27] , \ScanLink81[26] , 
        \ScanLink81[25] , \ScanLink81[24] , \ScanLink81[23] , \ScanLink81[22] , 
        \ScanLink81[21] , \ScanLink81[20] , \ScanLink81[19] , \ScanLink81[18] , 
        \ScanLink81[17] , \ScanLink81[16] , \ScanLink81[15] , \ScanLink81[14] , 
        \ScanLink81[13] , \ScanLink81[12] , \ScanLink81[11] , \ScanLink81[10] , 
        \ScanLink81[9] , \ScanLink81[8] , \ScanLink81[7] , \ScanLink81[6] , 
        \ScanLink81[5] , \ScanLink81[4] , \ScanLink81[3] , \ScanLink81[2] , 
        \ScanLink81[1] , \ScanLink81[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_18[31] , \wRegOut_6_18[30] , 
        \wRegOut_6_18[29] , \wRegOut_6_18[28] , \wRegOut_6_18[27] , 
        \wRegOut_6_18[26] , \wRegOut_6_18[25] , \wRegOut_6_18[24] , 
        \wRegOut_6_18[23] , \wRegOut_6_18[22] , \wRegOut_6_18[21] , 
        \wRegOut_6_18[20] , \wRegOut_6_18[19] , \wRegOut_6_18[18] , 
        \wRegOut_6_18[17] , \wRegOut_6_18[16] , \wRegOut_6_18[15] , 
        \wRegOut_6_18[14] , \wRegOut_6_18[13] , \wRegOut_6_18[12] , 
        \wRegOut_6_18[11] , \wRegOut_6_18[10] , \wRegOut_6_18[9] , 
        \wRegOut_6_18[8] , \wRegOut_6_18[7] , \wRegOut_6_18[6] , 
        \wRegOut_6_18[5] , \wRegOut_6_18[4] , \wRegOut_6_18[3] , 
        \wRegOut_6_18[2] , \wRegOut_6_18[1] , \wRegOut_6_18[0] }), .Enable1(
        \wRegEnTop_6_18[0] ), .Enable2(\wRegEnBot_6_18[0] ), .In1({
        \wRegInTop_6_18[31] , \wRegInTop_6_18[30] , \wRegInTop_6_18[29] , 
        \wRegInTop_6_18[28] , \wRegInTop_6_18[27] , \wRegInTop_6_18[26] , 
        \wRegInTop_6_18[25] , \wRegInTop_6_18[24] , \wRegInTop_6_18[23] , 
        \wRegInTop_6_18[22] , \wRegInTop_6_18[21] , \wRegInTop_6_18[20] , 
        \wRegInTop_6_18[19] , \wRegInTop_6_18[18] , \wRegInTop_6_18[17] , 
        \wRegInTop_6_18[16] , \wRegInTop_6_18[15] , \wRegInTop_6_18[14] , 
        \wRegInTop_6_18[13] , \wRegInTop_6_18[12] , \wRegInTop_6_18[11] , 
        \wRegInTop_6_18[10] , \wRegInTop_6_18[9] , \wRegInTop_6_18[8] , 
        \wRegInTop_6_18[7] , \wRegInTop_6_18[6] , \wRegInTop_6_18[5] , 
        \wRegInTop_6_18[4] , \wRegInTop_6_18[3] , \wRegInTop_6_18[2] , 
        \wRegInTop_6_18[1] , \wRegInTop_6_18[0] }), .In2({\wRegInBot_6_18[31] , 
        \wRegInBot_6_18[30] , \wRegInBot_6_18[29] , \wRegInBot_6_18[28] , 
        \wRegInBot_6_18[27] , \wRegInBot_6_18[26] , \wRegInBot_6_18[25] , 
        \wRegInBot_6_18[24] , \wRegInBot_6_18[23] , \wRegInBot_6_18[22] , 
        \wRegInBot_6_18[21] , \wRegInBot_6_18[20] , \wRegInBot_6_18[19] , 
        \wRegInBot_6_18[18] , \wRegInBot_6_18[17] , \wRegInBot_6_18[16] , 
        \wRegInBot_6_18[15] , \wRegInBot_6_18[14] , \wRegInBot_6_18[13] , 
        \wRegInBot_6_18[12] , \wRegInBot_6_18[11] , \wRegInBot_6_18[10] , 
        \wRegInBot_6_18[9] , \wRegInBot_6_18[8] , \wRegInBot_6_18[7] , 
        \wRegInBot_6_18[6] , \wRegInBot_6_18[5] , \wRegInBot_6_18[4] , 
        \wRegInBot_6_18[3] , \wRegInBot_6_18[2] , \wRegInBot_6_18[1] , 
        \wRegInBot_6_18[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_25 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink153[31] , \ScanLink153[30] , \ScanLink153[29] , 
        \ScanLink153[28] , \ScanLink153[27] , \ScanLink153[26] , 
        \ScanLink153[25] , \ScanLink153[24] , \ScanLink153[23] , 
        \ScanLink153[22] , \ScanLink153[21] , \ScanLink153[20] , 
        \ScanLink153[19] , \ScanLink153[18] , \ScanLink153[17] , 
        \ScanLink153[16] , \ScanLink153[15] , \ScanLink153[14] , 
        \ScanLink153[13] , \ScanLink153[12] , \ScanLink153[11] , 
        \ScanLink153[10] , \ScanLink153[9] , \ScanLink153[8] , 
        \ScanLink153[7] , \ScanLink153[6] , \ScanLink153[5] , \ScanLink153[4] , 
        \ScanLink153[3] , \ScanLink153[2] , \ScanLink153[1] , \ScanLink153[0] 
        }), .ScanOut({\ScanLink152[31] , \ScanLink152[30] , \ScanLink152[29] , 
        \ScanLink152[28] , \ScanLink152[27] , \ScanLink152[26] , 
        \ScanLink152[25] , \ScanLink152[24] , \ScanLink152[23] , 
        \ScanLink152[22] , \ScanLink152[21] , \ScanLink152[20] , 
        \ScanLink152[19] , \ScanLink152[18] , \ScanLink152[17] , 
        \ScanLink152[16] , \ScanLink152[15] , \ScanLink152[14] , 
        \ScanLink152[13] , \ScanLink152[12] , \ScanLink152[11] , 
        \ScanLink152[10] , \ScanLink152[9] , \ScanLink152[8] , 
        \ScanLink152[7] , \ScanLink152[6] , \ScanLink152[5] , \ScanLink152[4] , 
        \ScanLink152[3] , \ScanLink152[2] , \ScanLink152[1] , \ScanLink152[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_25[31] , 
        \wRegOut_7_25[30] , \wRegOut_7_25[29] , \wRegOut_7_25[28] , 
        \wRegOut_7_25[27] , \wRegOut_7_25[26] , \wRegOut_7_25[25] , 
        \wRegOut_7_25[24] , \wRegOut_7_25[23] , \wRegOut_7_25[22] , 
        \wRegOut_7_25[21] , \wRegOut_7_25[20] , \wRegOut_7_25[19] , 
        \wRegOut_7_25[18] , \wRegOut_7_25[17] , \wRegOut_7_25[16] , 
        \wRegOut_7_25[15] , \wRegOut_7_25[14] , \wRegOut_7_25[13] , 
        \wRegOut_7_25[12] , \wRegOut_7_25[11] , \wRegOut_7_25[10] , 
        \wRegOut_7_25[9] , \wRegOut_7_25[8] , \wRegOut_7_25[7] , 
        \wRegOut_7_25[6] , \wRegOut_7_25[5] , \wRegOut_7_25[4] , 
        \wRegOut_7_25[3] , \wRegOut_7_25[2] , \wRegOut_7_25[1] , 
        \wRegOut_7_25[0] }), .Enable1(\wRegEnTop_7_25[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_25[31] , \wRegInTop_7_25[30] , \wRegInTop_7_25[29] , 
        \wRegInTop_7_25[28] , \wRegInTop_7_25[27] , \wRegInTop_7_25[26] , 
        \wRegInTop_7_25[25] , \wRegInTop_7_25[24] , \wRegInTop_7_25[23] , 
        \wRegInTop_7_25[22] , \wRegInTop_7_25[21] , \wRegInTop_7_25[20] , 
        \wRegInTop_7_25[19] , \wRegInTop_7_25[18] , \wRegInTop_7_25[17] , 
        \wRegInTop_7_25[16] , \wRegInTop_7_25[15] , \wRegInTop_7_25[14] , 
        \wRegInTop_7_25[13] , \wRegInTop_7_25[12] , \wRegInTop_7_25[11] , 
        \wRegInTop_7_25[10] , \wRegInTop_7_25[9] , \wRegInTop_7_25[8] , 
        \wRegInTop_7_25[7] , \wRegInTop_7_25[6] , \wRegInTop_7_25[5] , 
        \wRegInTop_7_25[4] , \wRegInTop_7_25[3] , \wRegInTop_7_25[2] , 
        \wRegInTop_7_25[1] , \wRegInTop_7_25[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_116 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink244[31] , \ScanLink244[30] , \ScanLink244[29] , 
        \ScanLink244[28] , \ScanLink244[27] , \ScanLink244[26] , 
        \ScanLink244[25] , \ScanLink244[24] , \ScanLink244[23] , 
        \ScanLink244[22] , \ScanLink244[21] , \ScanLink244[20] , 
        \ScanLink244[19] , \ScanLink244[18] , \ScanLink244[17] , 
        \ScanLink244[16] , \ScanLink244[15] , \ScanLink244[14] , 
        \ScanLink244[13] , \ScanLink244[12] , \ScanLink244[11] , 
        \ScanLink244[10] , \ScanLink244[9] , \ScanLink244[8] , 
        \ScanLink244[7] , \ScanLink244[6] , \ScanLink244[5] , \ScanLink244[4] , 
        \ScanLink244[3] , \ScanLink244[2] , \ScanLink244[1] , \ScanLink244[0] 
        }), .ScanOut({\ScanLink243[31] , \ScanLink243[30] , \ScanLink243[29] , 
        \ScanLink243[28] , \ScanLink243[27] , \ScanLink243[26] , 
        \ScanLink243[25] , \ScanLink243[24] , \ScanLink243[23] , 
        \ScanLink243[22] , \ScanLink243[21] , \ScanLink243[20] , 
        \ScanLink243[19] , \ScanLink243[18] , \ScanLink243[17] , 
        \ScanLink243[16] , \ScanLink243[15] , \ScanLink243[14] , 
        \ScanLink243[13] , \ScanLink243[12] , \ScanLink243[11] , 
        \ScanLink243[10] , \ScanLink243[9] , \ScanLink243[8] , 
        \ScanLink243[7] , \ScanLink243[6] , \ScanLink243[5] , \ScanLink243[4] , 
        \ScanLink243[3] , \ScanLink243[2] , \ScanLink243[1] , \ScanLink243[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_116[31] , 
        \wRegOut_7_116[30] , \wRegOut_7_116[29] , \wRegOut_7_116[28] , 
        \wRegOut_7_116[27] , \wRegOut_7_116[26] , \wRegOut_7_116[25] , 
        \wRegOut_7_116[24] , \wRegOut_7_116[23] , \wRegOut_7_116[22] , 
        \wRegOut_7_116[21] , \wRegOut_7_116[20] , \wRegOut_7_116[19] , 
        \wRegOut_7_116[18] , \wRegOut_7_116[17] , \wRegOut_7_116[16] , 
        \wRegOut_7_116[15] , \wRegOut_7_116[14] , \wRegOut_7_116[13] , 
        \wRegOut_7_116[12] , \wRegOut_7_116[11] , \wRegOut_7_116[10] , 
        \wRegOut_7_116[9] , \wRegOut_7_116[8] , \wRegOut_7_116[7] , 
        \wRegOut_7_116[6] , \wRegOut_7_116[5] , \wRegOut_7_116[4] , 
        \wRegOut_7_116[3] , \wRegOut_7_116[2] , \wRegOut_7_116[1] , 
        \wRegOut_7_116[0] }), .Enable1(\wRegEnTop_7_116[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_116[31] , \wRegInTop_7_116[30] , 
        \wRegInTop_7_116[29] , \wRegInTop_7_116[28] , \wRegInTop_7_116[27] , 
        \wRegInTop_7_116[26] , \wRegInTop_7_116[25] , \wRegInTop_7_116[24] , 
        \wRegInTop_7_116[23] , \wRegInTop_7_116[22] , \wRegInTop_7_116[21] , 
        \wRegInTop_7_116[20] , \wRegInTop_7_116[19] , \wRegInTop_7_116[18] , 
        \wRegInTop_7_116[17] , \wRegInTop_7_116[16] , \wRegInTop_7_116[15] , 
        \wRegInTop_7_116[14] , \wRegInTop_7_116[13] , \wRegInTop_7_116[12] , 
        \wRegInTop_7_116[11] , \wRegInTop_7_116[10] , \wRegInTop_7_116[9] , 
        \wRegInTop_7_116[8] , \wRegInTop_7_116[7] , \wRegInTop_7_116[6] , 
        \wRegInTop_7_116[5] , \wRegInTop_7_116[4] , \wRegInTop_7_116[3] , 
        \wRegInTop_7_116[2] , \wRegInTop_7_116[1] , \wRegInTop_7_116[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_3[0] ), .P_In({\wRegOut_4_3[31] , 
        \wRegOut_4_3[30] , \wRegOut_4_3[29] , \wRegOut_4_3[28] , 
        \wRegOut_4_3[27] , \wRegOut_4_3[26] , \wRegOut_4_3[25] , 
        \wRegOut_4_3[24] , \wRegOut_4_3[23] , \wRegOut_4_3[22] , 
        \wRegOut_4_3[21] , \wRegOut_4_3[20] , \wRegOut_4_3[19] , 
        \wRegOut_4_3[18] , \wRegOut_4_3[17] , \wRegOut_4_3[16] , 
        \wRegOut_4_3[15] , \wRegOut_4_3[14] , \wRegOut_4_3[13] , 
        \wRegOut_4_3[12] , \wRegOut_4_3[11] , \wRegOut_4_3[10] , 
        \wRegOut_4_3[9] , \wRegOut_4_3[8] , \wRegOut_4_3[7] , \wRegOut_4_3[6] , 
        \wRegOut_4_3[5] , \wRegOut_4_3[4] , \wRegOut_4_3[3] , \wRegOut_4_3[2] , 
        \wRegOut_4_3[1] , \wRegOut_4_3[0] }), .P_Out({\wRegInBot_4_3[31] , 
        \wRegInBot_4_3[30] , \wRegInBot_4_3[29] , \wRegInBot_4_3[28] , 
        \wRegInBot_4_3[27] , \wRegInBot_4_3[26] , \wRegInBot_4_3[25] , 
        \wRegInBot_4_3[24] , \wRegInBot_4_3[23] , \wRegInBot_4_3[22] , 
        \wRegInBot_4_3[21] , \wRegInBot_4_3[20] , \wRegInBot_4_3[19] , 
        \wRegInBot_4_3[18] , \wRegInBot_4_3[17] , \wRegInBot_4_3[16] , 
        \wRegInBot_4_3[15] , \wRegInBot_4_3[14] , \wRegInBot_4_3[13] , 
        \wRegInBot_4_3[12] , \wRegInBot_4_3[11] , \wRegInBot_4_3[10] , 
        \wRegInBot_4_3[9] , \wRegInBot_4_3[8] , \wRegInBot_4_3[7] , 
        \wRegInBot_4_3[6] , \wRegInBot_4_3[5] , \wRegInBot_4_3[4] , 
        \wRegInBot_4_3[3] , \wRegInBot_4_3[2] , \wRegInBot_4_3[1] , 
        \wRegInBot_4_3[0] }), .L_WR(\wRegEnTop_5_6[0] ), .L_In({
        \wRegOut_5_6[31] , \wRegOut_5_6[30] , \wRegOut_5_6[29] , 
        \wRegOut_5_6[28] , \wRegOut_5_6[27] , \wRegOut_5_6[26] , 
        \wRegOut_5_6[25] , \wRegOut_5_6[24] , \wRegOut_5_6[23] , 
        \wRegOut_5_6[22] , \wRegOut_5_6[21] , \wRegOut_5_6[20] , 
        \wRegOut_5_6[19] , \wRegOut_5_6[18] , \wRegOut_5_6[17] , 
        \wRegOut_5_6[16] , \wRegOut_5_6[15] , \wRegOut_5_6[14] , 
        \wRegOut_5_6[13] , \wRegOut_5_6[12] , \wRegOut_5_6[11] , 
        \wRegOut_5_6[10] , \wRegOut_5_6[9] , \wRegOut_5_6[8] , 
        \wRegOut_5_6[7] , \wRegOut_5_6[6] , \wRegOut_5_6[5] , \wRegOut_5_6[4] , 
        \wRegOut_5_6[3] , \wRegOut_5_6[2] , \wRegOut_5_6[1] , \wRegOut_5_6[0] 
        }), .L_Out({\wRegInTop_5_6[31] , \wRegInTop_5_6[30] , 
        \wRegInTop_5_6[29] , \wRegInTop_5_6[28] , \wRegInTop_5_6[27] , 
        \wRegInTop_5_6[26] , \wRegInTop_5_6[25] , \wRegInTop_5_6[24] , 
        \wRegInTop_5_6[23] , \wRegInTop_5_6[22] , \wRegInTop_5_6[21] , 
        \wRegInTop_5_6[20] , \wRegInTop_5_6[19] , \wRegInTop_5_6[18] , 
        \wRegInTop_5_6[17] , \wRegInTop_5_6[16] , \wRegInTop_5_6[15] , 
        \wRegInTop_5_6[14] , \wRegInTop_5_6[13] , \wRegInTop_5_6[12] , 
        \wRegInTop_5_6[11] , \wRegInTop_5_6[10] , \wRegInTop_5_6[9] , 
        \wRegInTop_5_6[8] , \wRegInTop_5_6[7] , \wRegInTop_5_6[6] , 
        \wRegInTop_5_6[5] , \wRegInTop_5_6[4] , \wRegInTop_5_6[3] , 
        \wRegInTop_5_6[2] , \wRegInTop_5_6[1] , \wRegInTop_5_6[0] }), .R_WR(
        \wRegEnTop_5_7[0] ), .R_In({\wRegOut_5_7[31] , \wRegOut_5_7[30] , 
        \wRegOut_5_7[29] , \wRegOut_5_7[28] , \wRegOut_5_7[27] , 
        \wRegOut_5_7[26] , \wRegOut_5_7[25] , \wRegOut_5_7[24] , 
        \wRegOut_5_7[23] , \wRegOut_5_7[22] , \wRegOut_5_7[21] , 
        \wRegOut_5_7[20] , \wRegOut_5_7[19] , \wRegOut_5_7[18] , 
        \wRegOut_5_7[17] , \wRegOut_5_7[16] , \wRegOut_5_7[15] , 
        \wRegOut_5_7[14] , \wRegOut_5_7[13] , \wRegOut_5_7[12] , 
        \wRegOut_5_7[11] , \wRegOut_5_7[10] , \wRegOut_5_7[9] , 
        \wRegOut_5_7[8] , \wRegOut_5_7[7] , \wRegOut_5_7[6] , \wRegOut_5_7[5] , 
        \wRegOut_5_7[4] , \wRegOut_5_7[3] , \wRegOut_5_7[2] , \wRegOut_5_7[1] , 
        \wRegOut_5_7[0] }), .R_Out({\wRegInTop_5_7[31] , \wRegInTop_5_7[30] , 
        \wRegInTop_5_7[29] , \wRegInTop_5_7[28] , \wRegInTop_5_7[27] , 
        \wRegInTop_5_7[26] , \wRegInTop_5_7[25] , \wRegInTop_5_7[24] , 
        \wRegInTop_5_7[23] , \wRegInTop_5_7[22] , \wRegInTop_5_7[21] , 
        \wRegInTop_5_7[20] , \wRegInTop_5_7[19] , \wRegInTop_5_7[18] , 
        \wRegInTop_5_7[17] , \wRegInTop_5_7[16] , \wRegInTop_5_7[15] , 
        \wRegInTop_5_7[14] , \wRegInTop_5_7[13] , \wRegInTop_5_7[12] , 
        \wRegInTop_5_7[11] , \wRegInTop_5_7[10] , \wRegInTop_5_7[9] , 
        \wRegInTop_5_7[8] , \wRegInTop_5_7[7] , \wRegInTop_5_7[6] , 
        \wRegInTop_5_7[5] , \wRegInTop_5_7[4] , \wRegInTop_5_7[3] , 
        \wRegInTop_5_7[2] , \wRegInTop_5_7[1] , \wRegInTop_5_7[0] }) );
    BHeap_Node_WIDTH32 BHN_5_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_27[0] ), .P_In({\wRegOut_5_27[31] , 
        \wRegOut_5_27[30] , \wRegOut_5_27[29] , \wRegOut_5_27[28] , 
        \wRegOut_5_27[27] , \wRegOut_5_27[26] , \wRegOut_5_27[25] , 
        \wRegOut_5_27[24] , \wRegOut_5_27[23] , \wRegOut_5_27[22] , 
        \wRegOut_5_27[21] , \wRegOut_5_27[20] , \wRegOut_5_27[19] , 
        \wRegOut_5_27[18] , \wRegOut_5_27[17] , \wRegOut_5_27[16] , 
        \wRegOut_5_27[15] , \wRegOut_5_27[14] , \wRegOut_5_27[13] , 
        \wRegOut_5_27[12] , \wRegOut_5_27[11] , \wRegOut_5_27[10] , 
        \wRegOut_5_27[9] , \wRegOut_5_27[8] , \wRegOut_5_27[7] , 
        \wRegOut_5_27[6] , \wRegOut_5_27[5] , \wRegOut_5_27[4] , 
        \wRegOut_5_27[3] , \wRegOut_5_27[2] , \wRegOut_5_27[1] , 
        \wRegOut_5_27[0] }), .P_Out({\wRegInBot_5_27[31] , 
        \wRegInBot_5_27[30] , \wRegInBot_5_27[29] , \wRegInBot_5_27[28] , 
        \wRegInBot_5_27[27] , \wRegInBot_5_27[26] , \wRegInBot_5_27[25] , 
        \wRegInBot_5_27[24] , \wRegInBot_5_27[23] , \wRegInBot_5_27[22] , 
        \wRegInBot_5_27[21] , \wRegInBot_5_27[20] , \wRegInBot_5_27[19] , 
        \wRegInBot_5_27[18] , \wRegInBot_5_27[17] , \wRegInBot_5_27[16] , 
        \wRegInBot_5_27[15] , \wRegInBot_5_27[14] , \wRegInBot_5_27[13] , 
        \wRegInBot_5_27[12] , \wRegInBot_5_27[11] , \wRegInBot_5_27[10] , 
        \wRegInBot_5_27[9] , \wRegInBot_5_27[8] , \wRegInBot_5_27[7] , 
        \wRegInBot_5_27[6] , \wRegInBot_5_27[5] , \wRegInBot_5_27[4] , 
        \wRegInBot_5_27[3] , \wRegInBot_5_27[2] , \wRegInBot_5_27[1] , 
        \wRegInBot_5_27[0] }), .L_WR(\wRegEnTop_6_54[0] ), .L_In({
        \wRegOut_6_54[31] , \wRegOut_6_54[30] , \wRegOut_6_54[29] , 
        \wRegOut_6_54[28] , \wRegOut_6_54[27] , \wRegOut_6_54[26] , 
        \wRegOut_6_54[25] , \wRegOut_6_54[24] , \wRegOut_6_54[23] , 
        \wRegOut_6_54[22] , \wRegOut_6_54[21] , \wRegOut_6_54[20] , 
        \wRegOut_6_54[19] , \wRegOut_6_54[18] , \wRegOut_6_54[17] , 
        \wRegOut_6_54[16] , \wRegOut_6_54[15] , \wRegOut_6_54[14] , 
        \wRegOut_6_54[13] , \wRegOut_6_54[12] , \wRegOut_6_54[11] , 
        \wRegOut_6_54[10] , \wRegOut_6_54[9] , \wRegOut_6_54[8] , 
        \wRegOut_6_54[7] , \wRegOut_6_54[6] , \wRegOut_6_54[5] , 
        \wRegOut_6_54[4] , \wRegOut_6_54[3] , \wRegOut_6_54[2] , 
        \wRegOut_6_54[1] , \wRegOut_6_54[0] }), .L_Out({\wRegInTop_6_54[31] , 
        \wRegInTop_6_54[30] , \wRegInTop_6_54[29] , \wRegInTop_6_54[28] , 
        \wRegInTop_6_54[27] , \wRegInTop_6_54[26] , \wRegInTop_6_54[25] , 
        \wRegInTop_6_54[24] , \wRegInTop_6_54[23] , \wRegInTop_6_54[22] , 
        \wRegInTop_6_54[21] , \wRegInTop_6_54[20] , \wRegInTop_6_54[19] , 
        \wRegInTop_6_54[18] , \wRegInTop_6_54[17] , \wRegInTop_6_54[16] , 
        \wRegInTop_6_54[15] , \wRegInTop_6_54[14] , \wRegInTop_6_54[13] , 
        \wRegInTop_6_54[12] , \wRegInTop_6_54[11] , \wRegInTop_6_54[10] , 
        \wRegInTop_6_54[9] , \wRegInTop_6_54[8] , \wRegInTop_6_54[7] , 
        \wRegInTop_6_54[6] , \wRegInTop_6_54[5] , \wRegInTop_6_54[4] , 
        \wRegInTop_6_54[3] , \wRegInTop_6_54[2] , \wRegInTop_6_54[1] , 
        \wRegInTop_6_54[0] }), .R_WR(\wRegEnTop_6_55[0] ), .R_In({
        \wRegOut_6_55[31] , \wRegOut_6_55[30] , \wRegOut_6_55[29] , 
        \wRegOut_6_55[28] , \wRegOut_6_55[27] , \wRegOut_6_55[26] , 
        \wRegOut_6_55[25] , \wRegOut_6_55[24] , \wRegOut_6_55[23] , 
        \wRegOut_6_55[22] , \wRegOut_6_55[21] , \wRegOut_6_55[20] , 
        \wRegOut_6_55[19] , \wRegOut_6_55[18] , \wRegOut_6_55[17] , 
        \wRegOut_6_55[16] , \wRegOut_6_55[15] , \wRegOut_6_55[14] , 
        \wRegOut_6_55[13] , \wRegOut_6_55[12] , \wRegOut_6_55[11] , 
        \wRegOut_6_55[10] , \wRegOut_6_55[9] , \wRegOut_6_55[8] , 
        \wRegOut_6_55[7] , \wRegOut_6_55[6] , \wRegOut_6_55[5] , 
        \wRegOut_6_55[4] , \wRegOut_6_55[3] , \wRegOut_6_55[2] , 
        \wRegOut_6_55[1] , \wRegOut_6_55[0] }), .R_Out({\wRegInTop_6_55[31] , 
        \wRegInTop_6_55[30] , \wRegInTop_6_55[29] , \wRegInTop_6_55[28] , 
        \wRegInTop_6_55[27] , \wRegInTop_6_55[26] , \wRegInTop_6_55[25] , 
        \wRegInTop_6_55[24] , \wRegInTop_6_55[23] , \wRegInTop_6_55[22] , 
        \wRegInTop_6_55[21] , \wRegInTop_6_55[20] , \wRegInTop_6_55[19] , 
        \wRegInTop_6_55[18] , \wRegInTop_6_55[17] , \wRegInTop_6_55[16] , 
        \wRegInTop_6_55[15] , \wRegInTop_6_55[14] , \wRegInTop_6_55[13] , 
        \wRegInTop_6_55[12] , \wRegInTop_6_55[11] , \wRegInTop_6_55[10] , 
        \wRegInTop_6_55[9] , \wRegInTop_6_55[8] , \wRegInTop_6_55[7] , 
        \wRegInTop_6_55[6] , \wRegInTop_6_55[5] , \wRegInTop_6_55[4] , 
        \wRegInTop_6_55[3] , \wRegInTop_6_55[2] , \wRegInTop_6_55[1] , 
        \wRegInTop_6_55[0] }) );
    BHeap_Node_WIDTH32 BHN_6_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_30[0] ), .P_In({\wRegOut_6_30[31] , 
        \wRegOut_6_30[30] , \wRegOut_6_30[29] , \wRegOut_6_30[28] , 
        \wRegOut_6_30[27] , \wRegOut_6_30[26] , \wRegOut_6_30[25] , 
        \wRegOut_6_30[24] , \wRegOut_6_30[23] , \wRegOut_6_30[22] , 
        \wRegOut_6_30[21] , \wRegOut_6_30[20] , \wRegOut_6_30[19] , 
        \wRegOut_6_30[18] , \wRegOut_6_30[17] , \wRegOut_6_30[16] , 
        \wRegOut_6_30[15] , \wRegOut_6_30[14] , \wRegOut_6_30[13] , 
        \wRegOut_6_30[12] , \wRegOut_6_30[11] , \wRegOut_6_30[10] , 
        \wRegOut_6_30[9] , \wRegOut_6_30[8] , \wRegOut_6_30[7] , 
        \wRegOut_6_30[6] , \wRegOut_6_30[5] , \wRegOut_6_30[4] , 
        \wRegOut_6_30[3] , \wRegOut_6_30[2] , \wRegOut_6_30[1] , 
        \wRegOut_6_30[0] }), .P_Out({\wRegInBot_6_30[31] , 
        \wRegInBot_6_30[30] , \wRegInBot_6_30[29] , \wRegInBot_6_30[28] , 
        \wRegInBot_6_30[27] , \wRegInBot_6_30[26] , \wRegInBot_6_30[25] , 
        \wRegInBot_6_30[24] , \wRegInBot_6_30[23] , \wRegInBot_6_30[22] , 
        \wRegInBot_6_30[21] , \wRegInBot_6_30[20] , \wRegInBot_6_30[19] , 
        \wRegInBot_6_30[18] , \wRegInBot_6_30[17] , \wRegInBot_6_30[16] , 
        \wRegInBot_6_30[15] , \wRegInBot_6_30[14] , \wRegInBot_6_30[13] , 
        \wRegInBot_6_30[12] , \wRegInBot_6_30[11] , \wRegInBot_6_30[10] , 
        \wRegInBot_6_30[9] , \wRegInBot_6_30[8] , \wRegInBot_6_30[7] , 
        \wRegInBot_6_30[6] , \wRegInBot_6_30[5] , \wRegInBot_6_30[4] , 
        \wRegInBot_6_30[3] , \wRegInBot_6_30[2] , \wRegInBot_6_30[1] , 
        \wRegInBot_6_30[0] }), .L_WR(\wRegEnTop_7_60[0] ), .L_In({
        \wRegOut_7_60[31] , \wRegOut_7_60[30] , \wRegOut_7_60[29] , 
        \wRegOut_7_60[28] , \wRegOut_7_60[27] , \wRegOut_7_60[26] , 
        \wRegOut_7_60[25] , \wRegOut_7_60[24] , \wRegOut_7_60[23] , 
        \wRegOut_7_60[22] , \wRegOut_7_60[21] , \wRegOut_7_60[20] , 
        \wRegOut_7_60[19] , \wRegOut_7_60[18] , \wRegOut_7_60[17] , 
        \wRegOut_7_60[16] , \wRegOut_7_60[15] , \wRegOut_7_60[14] , 
        \wRegOut_7_60[13] , \wRegOut_7_60[12] , \wRegOut_7_60[11] , 
        \wRegOut_7_60[10] , \wRegOut_7_60[9] , \wRegOut_7_60[8] , 
        \wRegOut_7_60[7] , \wRegOut_7_60[6] , \wRegOut_7_60[5] , 
        \wRegOut_7_60[4] , \wRegOut_7_60[3] , \wRegOut_7_60[2] , 
        \wRegOut_7_60[1] , \wRegOut_7_60[0] }), .L_Out({\wRegInTop_7_60[31] , 
        \wRegInTop_7_60[30] , \wRegInTop_7_60[29] , \wRegInTop_7_60[28] , 
        \wRegInTop_7_60[27] , \wRegInTop_7_60[26] , \wRegInTop_7_60[25] , 
        \wRegInTop_7_60[24] , \wRegInTop_7_60[23] , \wRegInTop_7_60[22] , 
        \wRegInTop_7_60[21] , \wRegInTop_7_60[20] , \wRegInTop_7_60[19] , 
        \wRegInTop_7_60[18] , \wRegInTop_7_60[17] , \wRegInTop_7_60[16] , 
        \wRegInTop_7_60[15] , \wRegInTop_7_60[14] , \wRegInTop_7_60[13] , 
        \wRegInTop_7_60[12] , \wRegInTop_7_60[11] , \wRegInTop_7_60[10] , 
        \wRegInTop_7_60[9] , \wRegInTop_7_60[8] , \wRegInTop_7_60[7] , 
        \wRegInTop_7_60[6] , \wRegInTop_7_60[5] , \wRegInTop_7_60[4] , 
        \wRegInTop_7_60[3] , \wRegInTop_7_60[2] , \wRegInTop_7_60[1] , 
        \wRegInTop_7_60[0] }), .R_WR(\wRegEnTop_7_61[0] ), .R_In({
        \wRegOut_7_61[31] , \wRegOut_7_61[30] , \wRegOut_7_61[29] , 
        \wRegOut_7_61[28] , \wRegOut_7_61[27] , \wRegOut_7_61[26] , 
        \wRegOut_7_61[25] , \wRegOut_7_61[24] , \wRegOut_7_61[23] , 
        \wRegOut_7_61[22] , \wRegOut_7_61[21] , \wRegOut_7_61[20] , 
        \wRegOut_7_61[19] , \wRegOut_7_61[18] , \wRegOut_7_61[17] , 
        \wRegOut_7_61[16] , \wRegOut_7_61[15] , \wRegOut_7_61[14] , 
        \wRegOut_7_61[13] , \wRegOut_7_61[12] , \wRegOut_7_61[11] , 
        \wRegOut_7_61[10] , \wRegOut_7_61[9] , \wRegOut_7_61[8] , 
        \wRegOut_7_61[7] , \wRegOut_7_61[6] , \wRegOut_7_61[5] , 
        \wRegOut_7_61[4] , \wRegOut_7_61[3] , \wRegOut_7_61[2] , 
        \wRegOut_7_61[1] , \wRegOut_7_61[0] }), .R_Out({\wRegInTop_7_61[31] , 
        \wRegInTop_7_61[30] , \wRegInTop_7_61[29] , \wRegInTop_7_61[28] , 
        \wRegInTop_7_61[27] , \wRegInTop_7_61[26] , \wRegInTop_7_61[25] , 
        \wRegInTop_7_61[24] , \wRegInTop_7_61[23] , \wRegInTop_7_61[22] , 
        \wRegInTop_7_61[21] , \wRegInTop_7_61[20] , \wRegInTop_7_61[19] , 
        \wRegInTop_7_61[18] , \wRegInTop_7_61[17] , \wRegInTop_7_61[16] , 
        \wRegInTop_7_61[15] , \wRegInTop_7_61[14] , \wRegInTop_7_61[13] , 
        \wRegInTop_7_61[12] , \wRegInTop_7_61[11] , \wRegInTop_7_61[10] , 
        \wRegInTop_7_61[9] , \wRegInTop_7_61[8] , \wRegInTop_7_61[7] , 
        \wRegInTop_7_61[6] , \wRegInTop_7_61[5] , \wRegInTop_7_61[4] , 
        \wRegInTop_7_61[3] , \wRegInTop_7_61[2] , \wRegInTop_7_61[1] , 
        \wRegInTop_7_61[0] }) );
    BHeap_Node_WIDTH32 BHN_6_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_17[0] ), .P_In({\wRegOut_6_17[31] , 
        \wRegOut_6_17[30] , \wRegOut_6_17[29] , \wRegOut_6_17[28] , 
        \wRegOut_6_17[27] , \wRegOut_6_17[26] , \wRegOut_6_17[25] , 
        \wRegOut_6_17[24] , \wRegOut_6_17[23] , \wRegOut_6_17[22] , 
        \wRegOut_6_17[21] , \wRegOut_6_17[20] , \wRegOut_6_17[19] , 
        \wRegOut_6_17[18] , \wRegOut_6_17[17] , \wRegOut_6_17[16] , 
        \wRegOut_6_17[15] , \wRegOut_6_17[14] , \wRegOut_6_17[13] , 
        \wRegOut_6_17[12] , \wRegOut_6_17[11] , \wRegOut_6_17[10] , 
        \wRegOut_6_17[9] , \wRegOut_6_17[8] , \wRegOut_6_17[7] , 
        \wRegOut_6_17[6] , \wRegOut_6_17[5] , \wRegOut_6_17[4] , 
        \wRegOut_6_17[3] , \wRegOut_6_17[2] , \wRegOut_6_17[1] , 
        \wRegOut_6_17[0] }), .P_Out({\wRegInBot_6_17[31] , 
        \wRegInBot_6_17[30] , \wRegInBot_6_17[29] , \wRegInBot_6_17[28] , 
        \wRegInBot_6_17[27] , \wRegInBot_6_17[26] , \wRegInBot_6_17[25] , 
        \wRegInBot_6_17[24] , \wRegInBot_6_17[23] , \wRegInBot_6_17[22] , 
        \wRegInBot_6_17[21] , \wRegInBot_6_17[20] , \wRegInBot_6_17[19] , 
        \wRegInBot_6_17[18] , \wRegInBot_6_17[17] , \wRegInBot_6_17[16] , 
        \wRegInBot_6_17[15] , \wRegInBot_6_17[14] , \wRegInBot_6_17[13] , 
        \wRegInBot_6_17[12] , \wRegInBot_6_17[11] , \wRegInBot_6_17[10] , 
        \wRegInBot_6_17[9] , \wRegInBot_6_17[8] , \wRegInBot_6_17[7] , 
        \wRegInBot_6_17[6] , \wRegInBot_6_17[5] , \wRegInBot_6_17[4] , 
        \wRegInBot_6_17[3] , \wRegInBot_6_17[2] , \wRegInBot_6_17[1] , 
        \wRegInBot_6_17[0] }), .L_WR(\wRegEnTop_7_34[0] ), .L_In({
        \wRegOut_7_34[31] , \wRegOut_7_34[30] , \wRegOut_7_34[29] , 
        \wRegOut_7_34[28] , \wRegOut_7_34[27] , \wRegOut_7_34[26] , 
        \wRegOut_7_34[25] , \wRegOut_7_34[24] , \wRegOut_7_34[23] , 
        \wRegOut_7_34[22] , \wRegOut_7_34[21] , \wRegOut_7_34[20] , 
        \wRegOut_7_34[19] , \wRegOut_7_34[18] , \wRegOut_7_34[17] , 
        \wRegOut_7_34[16] , \wRegOut_7_34[15] , \wRegOut_7_34[14] , 
        \wRegOut_7_34[13] , \wRegOut_7_34[12] , \wRegOut_7_34[11] , 
        \wRegOut_7_34[10] , \wRegOut_7_34[9] , \wRegOut_7_34[8] , 
        \wRegOut_7_34[7] , \wRegOut_7_34[6] , \wRegOut_7_34[5] , 
        \wRegOut_7_34[4] , \wRegOut_7_34[3] , \wRegOut_7_34[2] , 
        \wRegOut_7_34[1] , \wRegOut_7_34[0] }), .L_Out({\wRegInTop_7_34[31] , 
        \wRegInTop_7_34[30] , \wRegInTop_7_34[29] , \wRegInTop_7_34[28] , 
        \wRegInTop_7_34[27] , \wRegInTop_7_34[26] , \wRegInTop_7_34[25] , 
        \wRegInTop_7_34[24] , \wRegInTop_7_34[23] , \wRegInTop_7_34[22] , 
        \wRegInTop_7_34[21] , \wRegInTop_7_34[20] , \wRegInTop_7_34[19] , 
        \wRegInTop_7_34[18] , \wRegInTop_7_34[17] , \wRegInTop_7_34[16] , 
        \wRegInTop_7_34[15] , \wRegInTop_7_34[14] , \wRegInTop_7_34[13] , 
        \wRegInTop_7_34[12] , \wRegInTop_7_34[11] , \wRegInTop_7_34[10] , 
        \wRegInTop_7_34[9] , \wRegInTop_7_34[8] , \wRegInTop_7_34[7] , 
        \wRegInTop_7_34[6] , \wRegInTop_7_34[5] , \wRegInTop_7_34[4] , 
        \wRegInTop_7_34[3] , \wRegInTop_7_34[2] , \wRegInTop_7_34[1] , 
        \wRegInTop_7_34[0] }), .R_WR(\wRegEnTop_7_35[0] ), .R_In({
        \wRegOut_7_35[31] , \wRegOut_7_35[30] , \wRegOut_7_35[29] , 
        \wRegOut_7_35[28] , \wRegOut_7_35[27] , \wRegOut_7_35[26] , 
        \wRegOut_7_35[25] , \wRegOut_7_35[24] , \wRegOut_7_35[23] , 
        \wRegOut_7_35[22] , \wRegOut_7_35[21] , \wRegOut_7_35[20] , 
        \wRegOut_7_35[19] , \wRegOut_7_35[18] , \wRegOut_7_35[17] , 
        \wRegOut_7_35[16] , \wRegOut_7_35[15] , \wRegOut_7_35[14] , 
        \wRegOut_7_35[13] , \wRegOut_7_35[12] , \wRegOut_7_35[11] , 
        \wRegOut_7_35[10] , \wRegOut_7_35[9] , \wRegOut_7_35[8] , 
        \wRegOut_7_35[7] , \wRegOut_7_35[6] , \wRegOut_7_35[5] , 
        \wRegOut_7_35[4] , \wRegOut_7_35[3] , \wRegOut_7_35[2] , 
        \wRegOut_7_35[1] , \wRegOut_7_35[0] }), .R_Out({\wRegInTop_7_35[31] , 
        \wRegInTop_7_35[30] , \wRegInTop_7_35[29] , \wRegInTop_7_35[28] , 
        \wRegInTop_7_35[27] , \wRegInTop_7_35[26] , \wRegInTop_7_35[25] , 
        \wRegInTop_7_35[24] , \wRegInTop_7_35[23] , \wRegInTop_7_35[22] , 
        \wRegInTop_7_35[21] , \wRegInTop_7_35[20] , \wRegInTop_7_35[19] , 
        \wRegInTop_7_35[18] , \wRegInTop_7_35[17] , \wRegInTop_7_35[16] , 
        \wRegInTop_7_35[15] , \wRegInTop_7_35[14] , \wRegInTop_7_35[13] , 
        \wRegInTop_7_35[12] , \wRegInTop_7_35[11] , \wRegInTop_7_35[10] , 
        \wRegInTop_7_35[9] , \wRegInTop_7_35[8] , \wRegInTop_7_35[7] , 
        \wRegInTop_7_35[6] , \wRegInTop_7_35[5] , \wRegInTop_7_35[4] , 
        \wRegInTop_7_35[3] , \wRegInTop_7_35[2] , \wRegInTop_7_35[1] , 
        \wRegInTop_7_35[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink24[31] , \ScanLink24[30] , \ScanLink24[29] , 
        \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , \ScanLink24[25] , 
        \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , \ScanLink24[21] , 
        \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , \ScanLink24[17] , 
        \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , \ScanLink24[13] , 
        \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , \ScanLink24[9] , 
        \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , \ScanLink24[5] , 
        \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , \ScanLink24[1] , 
        \ScanLink24[0] }), .ScanOut({\ScanLink23[31] , \ScanLink23[30] , 
        \ScanLink23[29] , \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , 
        \ScanLink23[25] , \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , 
        \ScanLink23[21] , \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , 
        \ScanLink23[17] , \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , 
        \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , 
        \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , 
        \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , 
        \ScanLink23[1] , \ScanLink23[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_8[31] , \wRegOut_4_8[30] , \wRegOut_4_8[29] , 
        \wRegOut_4_8[28] , \wRegOut_4_8[27] , \wRegOut_4_8[26] , 
        \wRegOut_4_8[25] , \wRegOut_4_8[24] , \wRegOut_4_8[23] , 
        \wRegOut_4_8[22] , \wRegOut_4_8[21] , \wRegOut_4_8[20] , 
        \wRegOut_4_8[19] , \wRegOut_4_8[18] , \wRegOut_4_8[17] , 
        \wRegOut_4_8[16] , \wRegOut_4_8[15] , \wRegOut_4_8[14] , 
        \wRegOut_4_8[13] , \wRegOut_4_8[12] , \wRegOut_4_8[11] , 
        \wRegOut_4_8[10] , \wRegOut_4_8[9] , \wRegOut_4_8[8] , 
        \wRegOut_4_8[7] , \wRegOut_4_8[6] , \wRegOut_4_8[5] , \wRegOut_4_8[4] , 
        \wRegOut_4_8[3] , \wRegOut_4_8[2] , \wRegOut_4_8[1] , \wRegOut_4_8[0] 
        }), .Enable1(\wRegEnTop_4_8[0] ), .Enable2(\wRegEnBot_4_8[0] ), .In1({
        \wRegInTop_4_8[31] , \wRegInTop_4_8[30] , \wRegInTop_4_8[29] , 
        \wRegInTop_4_8[28] , \wRegInTop_4_8[27] , \wRegInTop_4_8[26] , 
        \wRegInTop_4_8[25] , \wRegInTop_4_8[24] , \wRegInTop_4_8[23] , 
        \wRegInTop_4_8[22] , \wRegInTop_4_8[21] , \wRegInTop_4_8[20] , 
        \wRegInTop_4_8[19] , \wRegInTop_4_8[18] , \wRegInTop_4_8[17] , 
        \wRegInTop_4_8[16] , \wRegInTop_4_8[15] , \wRegInTop_4_8[14] , 
        \wRegInTop_4_8[13] , \wRegInTop_4_8[12] , \wRegInTop_4_8[11] , 
        \wRegInTop_4_8[10] , \wRegInTop_4_8[9] , \wRegInTop_4_8[8] , 
        \wRegInTop_4_8[7] , \wRegInTop_4_8[6] , \wRegInTop_4_8[5] , 
        \wRegInTop_4_8[4] , \wRegInTop_4_8[3] , \wRegInTop_4_8[2] , 
        \wRegInTop_4_8[1] , \wRegInTop_4_8[0] }), .In2({\wRegInBot_4_8[31] , 
        \wRegInBot_4_8[30] , \wRegInBot_4_8[29] , \wRegInBot_4_8[28] , 
        \wRegInBot_4_8[27] , \wRegInBot_4_8[26] , \wRegInBot_4_8[25] , 
        \wRegInBot_4_8[24] , \wRegInBot_4_8[23] , \wRegInBot_4_8[22] , 
        \wRegInBot_4_8[21] , \wRegInBot_4_8[20] , \wRegInBot_4_8[19] , 
        \wRegInBot_4_8[18] , \wRegInBot_4_8[17] , \wRegInBot_4_8[16] , 
        \wRegInBot_4_8[15] , \wRegInBot_4_8[14] , \wRegInBot_4_8[13] , 
        \wRegInBot_4_8[12] , \wRegInBot_4_8[11] , \wRegInBot_4_8[10] , 
        \wRegInBot_4_8[9] , \wRegInBot_4_8[8] , \wRegInBot_4_8[7] , 
        \wRegInBot_4_8[6] , \wRegInBot_4_8[5] , \wRegInBot_4_8[4] , 
        \wRegInBot_4_8[3] , \wRegInBot_4_8[2] , \wRegInBot_4_8[1] , 
        \wRegInBot_4_8[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink68[31] , \ScanLink68[30] , \ScanLink68[29] , 
        \ScanLink68[28] , \ScanLink68[27] , \ScanLink68[26] , \ScanLink68[25] , 
        \ScanLink68[24] , \ScanLink68[23] , \ScanLink68[22] , \ScanLink68[21] , 
        \ScanLink68[20] , \ScanLink68[19] , \ScanLink68[18] , \ScanLink68[17] , 
        \ScanLink68[16] , \ScanLink68[15] , \ScanLink68[14] , \ScanLink68[13] , 
        \ScanLink68[12] , \ScanLink68[11] , \ScanLink68[10] , \ScanLink68[9] , 
        \ScanLink68[8] , \ScanLink68[7] , \ScanLink68[6] , \ScanLink68[5] , 
        \ScanLink68[4] , \ScanLink68[3] , \ScanLink68[2] , \ScanLink68[1] , 
        \ScanLink68[0] }), .ScanOut({\ScanLink67[31] , \ScanLink67[30] , 
        \ScanLink67[29] , \ScanLink67[28] , \ScanLink67[27] , \ScanLink67[26] , 
        \ScanLink67[25] , \ScanLink67[24] , \ScanLink67[23] , \ScanLink67[22] , 
        \ScanLink67[21] , \ScanLink67[20] , \ScanLink67[19] , \ScanLink67[18] , 
        \ScanLink67[17] , \ScanLink67[16] , \ScanLink67[15] , \ScanLink67[14] , 
        \ScanLink67[13] , \ScanLink67[12] , \ScanLink67[11] , \ScanLink67[10] , 
        \ScanLink67[9] , \ScanLink67[8] , \ScanLink67[7] , \ScanLink67[6] , 
        \ScanLink67[5] , \ScanLink67[4] , \ScanLink67[3] , \ScanLink67[2] , 
        \ScanLink67[1] , \ScanLink67[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_4[31] , \wRegOut_6_4[30] , \wRegOut_6_4[29] , 
        \wRegOut_6_4[28] , \wRegOut_6_4[27] , \wRegOut_6_4[26] , 
        \wRegOut_6_4[25] , \wRegOut_6_4[24] , \wRegOut_6_4[23] , 
        \wRegOut_6_4[22] , \wRegOut_6_4[21] , \wRegOut_6_4[20] , 
        \wRegOut_6_4[19] , \wRegOut_6_4[18] , \wRegOut_6_4[17] , 
        \wRegOut_6_4[16] , \wRegOut_6_4[15] , \wRegOut_6_4[14] , 
        \wRegOut_6_4[13] , \wRegOut_6_4[12] , \wRegOut_6_4[11] , 
        \wRegOut_6_4[10] , \wRegOut_6_4[9] , \wRegOut_6_4[8] , 
        \wRegOut_6_4[7] , \wRegOut_6_4[6] , \wRegOut_6_4[5] , \wRegOut_6_4[4] , 
        \wRegOut_6_4[3] , \wRegOut_6_4[2] , \wRegOut_6_4[1] , \wRegOut_6_4[0] 
        }), .Enable1(\wRegEnTop_6_4[0] ), .Enable2(\wRegEnBot_6_4[0] ), .In1({
        \wRegInTop_6_4[31] , \wRegInTop_6_4[30] , \wRegInTop_6_4[29] , 
        \wRegInTop_6_4[28] , \wRegInTop_6_4[27] , \wRegInTop_6_4[26] , 
        \wRegInTop_6_4[25] , \wRegInTop_6_4[24] , \wRegInTop_6_4[23] , 
        \wRegInTop_6_4[22] , \wRegInTop_6_4[21] , \wRegInTop_6_4[20] , 
        \wRegInTop_6_4[19] , \wRegInTop_6_4[18] , \wRegInTop_6_4[17] , 
        \wRegInTop_6_4[16] , \wRegInTop_6_4[15] , \wRegInTop_6_4[14] , 
        \wRegInTop_6_4[13] , \wRegInTop_6_4[12] , \wRegInTop_6_4[11] , 
        \wRegInTop_6_4[10] , \wRegInTop_6_4[9] , \wRegInTop_6_4[8] , 
        \wRegInTop_6_4[7] , \wRegInTop_6_4[6] , \wRegInTop_6_4[5] , 
        \wRegInTop_6_4[4] , \wRegInTop_6_4[3] , \wRegInTop_6_4[2] , 
        \wRegInTop_6_4[1] , \wRegInTop_6_4[0] }), .In2({\wRegInBot_6_4[31] , 
        \wRegInBot_6_4[30] , \wRegInBot_6_4[29] , \wRegInBot_6_4[28] , 
        \wRegInBot_6_4[27] , \wRegInBot_6_4[26] , \wRegInBot_6_4[25] , 
        \wRegInBot_6_4[24] , \wRegInBot_6_4[23] , \wRegInBot_6_4[22] , 
        \wRegInBot_6_4[21] , \wRegInBot_6_4[20] , \wRegInBot_6_4[19] , 
        \wRegInBot_6_4[18] , \wRegInBot_6_4[17] , \wRegInBot_6_4[16] , 
        \wRegInBot_6_4[15] , \wRegInBot_6_4[14] , \wRegInBot_6_4[13] , 
        \wRegInBot_6_4[12] , \wRegInBot_6_4[11] , \wRegInBot_6_4[10] , 
        \wRegInBot_6_4[9] , \wRegInBot_6_4[8] , \wRegInBot_6_4[7] , 
        \wRegInBot_6_4[6] , \wRegInBot_6_4[5] , \wRegInBot_6_4[4] , 
        \wRegInBot_6_4[3] , \wRegInBot_6_4[2] , \wRegInBot_6_4[1] , 
        \wRegInBot_6_4[0] }) );
    BHeap_Node_WIDTH32 BHN_5_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_12[0] ), .P_In({\wRegOut_5_12[31] , 
        \wRegOut_5_12[30] , \wRegOut_5_12[29] , \wRegOut_5_12[28] , 
        \wRegOut_5_12[27] , \wRegOut_5_12[26] , \wRegOut_5_12[25] , 
        \wRegOut_5_12[24] , \wRegOut_5_12[23] , \wRegOut_5_12[22] , 
        \wRegOut_5_12[21] , \wRegOut_5_12[20] , \wRegOut_5_12[19] , 
        \wRegOut_5_12[18] , \wRegOut_5_12[17] , \wRegOut_5_12[16] , 
        \wRegOut_5_12[15] , \wRegOut_5_12[14] , \wRegOut_5_12[13] , 
        \wRegOut_5_12[12] , \wRegOut_5_12[11] , \wRegOut_5_12[10] , 
        \wRegOut_5_12[9] , \wRegOut_5_12[8] , \wRegOut_5_12[7] , 
        \wRegOut_5_12[6] , \wRegOut_5_12[5] , \wRegOut_5_12[4] , 
        \wRegOut_5_12[3] , \wRegOut_5_12[2] , \wRegOut_5_12[1] , 
        \wRegOut_5_12[0] }), .P_Out({\wRegInBot_5_12[31] , 
        \wRegInBot_5_12[30] , \wRegInBot_5_12[29] , \wRegInBot_5_12[28] , 
        \wRegInBot_5_12[27] , \wRegInBot_5_12[26] , \wRegInBot_5_12[25] , 
        \wRegInBot_5_12[24] , \wRegInBot_5_12[23] , \wRegInBot_5_12[22] , 
        \wRegInBot_5_12[21] , \wRegInBot_5_12[20] , \wRegInBot_5_12[19] , 
        \wRegInBot_5_12[18] , \wRegInBot_5_12[17] , \wRegInBot_5_12[16] , 
        \wRegInBot_5_12[15] , \wRegInBot_5_12[14] , \wRegInBot_5_12[13] , 
        \wRegInBot_5_12[12] , \wRegInBot_5_12[11] , \wRegInBot_5_12[10] , 
        \wRegInBot_5_12[9] , \wRegInBot_5_12[8] , \wRegInBot_5_12[7] , 
        \wRegInBot_5_12[6] , \wRegInBot_5_12[5] , \wRegInBot_5_12[4] , 
        \wRegInBot_5_12[3] , \wRegInBot_5_12[2] , \wRegInBot_5_12[1] , 
        \wRegInBot_5_12[0] }), .L_WR(\wRegEnTop_6_24[0] ), .L_In({
        \wRegOut_6_24[31] , \wRegOut_6_24[30] , \wRegOut_6_24[29] , 
        \wRegOut_6_24[28] , \wRegOut_6_24[27] , \wRegOut_6_24[26] , 
        \wRegOut_6_24[25] , \wRegOut_6_24[24] , \wRegOut_6_24[23] , 
        \wRegOut_6_24[22] , \wRegOut_6_24[21] , \wRegOut_6_24[20] , 
        \wRegOut_6_24[19] , \wRegOut_6_24[18] , \wRegOut_6_24[17] , 
        \wRegOut_6_24[16] , \wRegOut_6_24[15] , \wRegOut_6_24[14] , 
        \wRegOut_6_24[13] , \wRegOut_6_24[12] , \wRegOut_6_24[11] , 
        \wRegOut_6_24[10] , \wRegOut_6_24[9] , \wRegOut_6_24[8] , 
        \wRegOut_6_24[7] , \wRegOut_6_24[6] , \wRegOut_6_24[5] , 
        \wRegOut_6_24[4] , \wRegOut_6_24[3] , \wRegOut_6_24[2] , 
        \wRegOut_6_24[1] , \wRegOut_6_24[0] }), .L_Out({\wRegInTop_6_24[31] , 
        \wRegInTop_6_24[30] , \wRegInTop_6_24[29] , \wRegInTop_6_24[28] , 
        \wRegInTop_6_24[27] , \wRegInTop_6_24[26] , \wRegInTop_6_24[25] , 
        \wRegInTop_6_24[24] , \wRegInTop_6_24[23] , \wRegInTop_6_24[22] , 
        \wRegInTop_6_24[21] , \wRegInTop_6_24[20] , \wRegInTop_6_24[19] , 
        \wRegInTop_6_24[18] , \wRegInTop_6_24[17] , \wRegInTop_6_24[16] , 
        \wRegInTop_6_24[15] , \wRegInTop_6_24[14] , \wRegInTop_6_24[13] , 
        \wRegInTop_6_24[12] , \wRegInTop_6_24[11] , \wRegInTop_6_24[10] , 
        \wRegInTop_6_24[9] , \wRegInTop_6_24[8] , \wRegInTop_6_24[7] , 
        \wRegInTop_6_24[6] , \wRegInTop_6_24[5] , \wRegInTop_6_24[4] , 
        \wRegInTop_6_24[3] , \wRegInTop_6_24[2] , \wRegInTop_6_24[1] , 
        \wRegInTop_6_24[0] }), .R_WR(\wRegEnTop_6_25[0] ), .R_In({
        \wRegOut_6_25[31] , \wRegOut_6_25[30] , \wRegOut_6_25[29] , 
        \wRegOut_6_25[28] , \wRegOut_6_25[27] , \wRegOut_6_25[26] , 
        \wRegOut_6_25[25] , \wRegOut_6_25[24] , \wRegOut_6_25[23] , 
        \wRegOut_6_25[22] , \wRegOut_6_25[21] , \wRegOut_6_25[20] , 
        \wRegOut_6_25[19] , \wRegOut_6_25[18] , \wRegOut_6_25[17] , 
        \wRegOut_6_25[16] , \wRegOut_6_25[15] , \wRegOut_6_25[14] , 
        \wRegOut_6_25[13] , \wRegOut_6_25[12] , \wRegOut_6_25[11] , 
        \wRegOut_6_25[10] , \wRegOut_6_25[9] , \wRegOut_6_25[8] , 
        \wRegOut_6_25[7] , \wRegOut_6_25[6] , \wRegOut_6_25[5] , 
        \wRegOut_6_25[4] , \wRegOut_6_25[3] , \wRegOut_6_25[2] , 
        \wRegOut_6_25[1] , \wRegOut_6_25[0] }), .R_Out({\wRegInTop_6_25[31] , 
        \wRegInTop_6_25[30] , \wRegInTop_6_25[29] , \wRegInTop_6_25[28] , 
        \wRegInTop_6_25[27] , \wRegInTop_6_25[26] , \wRegInTop_6_25[25] , 
        \wRegInTop_6_25[24] , \wRegInTop_6_25[23] , \wRegInTop_6_25[22] , 
        \wRegInTop_6_25[21] , \wRegInTop_6_25[20] , \wRegInTop_6_25[19] , 
        \wRegInTop_6_25[18] , \wRegInTop_6_25[17] , \wRegInTop_6_25[16] , 
        \wRegInTop_6_25[15] , \wRegInTop_6_25[14] , \wRegInTop_6_25[13] , 
        \wRegInTop_6_25[12] , \wRegInTop_6_25[11] , \wRegInTop_6_25[10] , 
        \wRegInTop_6_25[9] , \wRegInTop_6_25[8] , \wRegInTop_6_25[7] , 
        \wRegInTop_6_25[6] , \wRegInTop_6_25[5] , \wRegInTop_6_25[4] , 
        \wRegInTop_6_25[3] , \wRegInTop_6_25[2] , \wRegInTop_6_25[1] , 
        \wRegInTop_6_25[0] }) );
    BHeap_Node_WIDTH32 BHN_6_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_22[0] ), .P_In({\wRegOut_6_22[31] , 
        \wRegOut_6_22[30] , \wRegOut_6_22[29] , \wRegOut_6_22[28] , 
        \wRegOut_6_22[27] , \wRegOut_6_22[26] , \wRegOut_6_22[25] , 
        \wRegOut_6_22[24] , \wRegOut_6_22[23] , \wRegOut_6_22[22] , 
        \wRegOut_6_22[21] , \wRegOut_6_22[20] , \wRegOut_6_22[19] , 
        \wRegOut_6_22[18] , \wRegOut_6_22[17] , \wRegOut_6_22[16] , 
        \wRegOut_6_22[15] , \wRegOut_6_22[14] , \wRegOut_6_22[13] , 
        \wRegOut_6_22[12] , \wRegOut_6_22[11] , \wRegOut_6_22[10] , 
        \wRegOut_6_22[9] , \wRegOut_6_22[8] , \wRegOut_6_22[7] , 
        \wRegOut_6_22[6] , \wRegOut_6_22[5] , \wRegOut_6_22[4] , 
        \wRegOut_6_22[3] , \wRegOut_6_22[2] , \wRegOut_6_22[1] , 
        \wRegOut_6_22[0] }), .P_Out({\wRegInBot_6_22[31] , 
        \wRegInBot_6_22[30] , \wRegInBot_6_22[29] , \wRegInBot_6_22[28] , 
        \wRegInBot_6_22[27] , \wRegInBot_6_22[26] , \wRegInBot_6_22[25] , 
        \wRegInBot_6_22[24] , \wRegInBot_6_22[23] , \wRegInBot_6_22[22] , 
        \wRegInBot_6_22[21] , \wRegInBot_6_22[20] , \wRegInBot_6_22[19] , 
        \wRegInBot_6_22[18] , \wRegInBot_6_22[17] , \wRegInBot_6_22[16] , 
        \wRegInBot_6_22[15] , \wRegInBot_6_22[14] , \wRegInBot_6_22[13] , 
        \wRegInBot_6_22[12] , \wRegInBot_6_22[11] , \wRegInBot_6_22[10] , 
        \wRegInBot_6_22[9] , \wRegInBot_6_22[8] , \wRegInBot_6_22[7] , 
        \wRegInBot_6_22[6] , \wRegInBot_6_22[5] , \wRegInBot_6_22[4] , 
        \wRegInBot_6_22[3] , \wRegInBot_6_22[2] , \wRegInBot_6_22[1] , 
        \wRegInBot_6_22[0] }), .L_WR(\wRegEnTop_7_44[0] ), .L_In({
        \wRegOut_7_44[31] , \wRegOut_7_44[30] , \wRegOut_7_44[29] , 
        \wRegOut_7_44[28] , \wRegOut_7_44[27] , \wRegOut_7_44[26] , 
        \wRegOut_7_44[25] , \wRegOut_7_44[24] , \wRegOut_7_44[23] , 
        \wRegOut_7_44[22] , \wRegOut_7_44[21] , \wRegOut_7_44[20] , 
        \wRegOut_7_44[19] , \wRegOut_7_44[18] , \wRegOut_7_44[17] , 
        \wRegOut_7_44[16] , \wRegOut_7_44[15] , \wRegOut_7_44[14] , 
        \wRegOut_7_44[13] , \wRegOut_7_44[12] , \wRegOut_7_44[11] , 
        \wRegOut_7_44[10] , \wRegOut_7_44[9] , \wRegOut_7_44[8] , 
        \wRegOut_7_44[7] , \wRegOut_7_44[6] , \wRegOut_7_44[5] , 
        \wRegOut_7_44[4] , \wRegOut_7_44[3] , \wRegOut_7_44[2] , 
        \wRegOut_7_44[1] , \wRegOut_7_44[0] }), .L_Out({\wRegInTop_7_44[31] , 
        \wRegInTop_7_44[30] , \wRegInTop_7_44[29] , \wRegInTop_7_44[28] , 
        \wRegInTop_7_44[27] , \wRegInTop_7_44[26] , \wRegInTop_7_44[25] , 
        \wRegInTop_7_44[24] , \wRegInTop_7_44[23] , \wRegInTop_7_44[22] , 
        \wRegInTop_7_44[21] , \wRegInTop_7_44[20] , \wRegInTop_7_44[19] , 
        \wRegInTop_7_44[18] , \wRegInTop_7_44[17] , \wRegInTop_7_44[16] , 
        \wRegInTop_7_44[15] , \wRegInTop_7_44[14] , \wRegInTop_7_44[13] , 
        \wRegInTop_7_44[12] , \wRegInTop_7_44[11] , \wRegInTop_7_44[10] , 
        \wRegInTop_7_44[9] , \wRegInTop_7_44[8] , \wRegInTop_7_44[7] , 
        \wRegInTop_7_44[6] , \wRegInTop_7_44[5] , \wRegInTop_7_44[4] , 
        \wRegInTop_7_44[3] , \wRegInTop_7_44[2] , \wRegInTop_7_44[1] , 
        \wRegInTop_7_44[0] }), .R_WR(\wRegEnTop_7_45[0] ), .R_In({
        \wRegOut_7_45[31] , \wRegOut_7_45[30] , \wRegOut_7_45[29] , 
        \wRegOut_7_45[28] , \wRegOut_7_45[27] , \wRegOut_7_45[26] , 
        \wRegOut_7_45[25] , \wRegOut_7_45[24] , \wRegOut_7_45[23] , 
        \wRegOut_7_45[22] , \wRegOut_7_45[21] , \wRegOut_7_45[20] , 
        \wRegOut_7_45[19] , \wRegOut_7_45[18] , \wRegOut_7_45[17] , 
        \wRegOut_7_45[16] , \wRegOut_7_45[15] , \wRegOut_7_45[14] , 
        \wRegOut_7_45[13] , \wRegOut_7_45[12] , \wRegOut_7_45[11] , 
        \wRegOut_7_45[10] , \wRegOut_7_45[9] , \wRegOut_7_45[8] , 
        \wRegOut_7_45[7] , \wRegOut_7_45[6] , \wRegOut_7_45[5] , 
        \wRegOut_7_45[4] , \wRegOut_7_45[3] , \wRegOut_7_45[2] , 
        \wRegOut_7_45[1] , \wRegOut_7_45[0] }), .R_Out({\wRegInTop_7_45[31] , 
        \wRegInTop_7_45[30] , \wRegInTop_7_45[29] , \wRegInTop_7_45[28] , 
        \wRegInTop_7_45[27] , \wRegInTop_7_45[26] , \wRegInTop_7_45[25] , 
        \wRegInTop_7_45[24] , \wRegInTop_7_45[23] , \wRegInTop_7_45[22] , 
        \wRegInTop_7_45[21] , \wRegInTop_7_45[20] , \wRegInTop_7_45[19] , 
        \wRegInTop_7_45[18] , \wRegInTop_7_45[17] , \wRegInTop_7_45[16] , 
        \wRegInTop_7_45[15] , \wRegInTop_7_45[14] , \wRegInTop_7_45[13] , 
        \wRegInTop_7_45[12] , \wRegInTop_7_45[11] , \wRegInTop_7_45[10] , 
        \wRegInTop_7_45[9] , \wRegInTop_7_45[8] , \wRegInTop_7_45[7] , 
        \wRegInTop_7_45[6] , \wRegInTop_7_45[5] , \wRegInTop_7_45[4] , 
        \wRegInTop_7_45[3] , \wRegInTop_7_45[2] , \wRegInTop_7_45[1] , 
        \wRegInTop_7_45[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_36 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink100[31] , \ScanLink100[30] , \ScanLink100[29] , 
        \ScanLink100[28] , \ScanLink100[27] , \ScanLink100[26] , 
        \ScanLink100[25] , \ScanLink100[24] , \ScanLink100[23] , 
        \ScanLink100[22] , \ScanLink100[21] , \ScanLink100[20] , 
        \ScanLink100[19] , \ScanLink100[18] , \ScanLink100[17] , 
        \ScanLink100[16] , \ScanLink100[15] , \ScanLink100[14] , 
        \ScanLink100[13] , \ScanLink100[12] , \ScanLink100[11] , 
        \ScanLink100[10] , \ScanLink100[9] , \ScanLink100[8] , 
        \ScanLink100[7] , \ScanLink100[6] , \ScanLink100[5] , \ScanLink100[4] , 
        \ScanLink100[3] , \ScanLink100[2] , \ScanLink100[1] , \ScanLink100[0] 
        }), .ScanOut({\ScanLink99[31] , \ScanLink99[30] , \ScanLink99[29] , 
        \ScanLink99[28] , \ScanLink99[27] , \ScanLink99[26] , \ScanLink99[25] , 
        \ScanLink99[24] , \ScanLink99[23] , \ScanLink99[22] , \ScanLink99[21] , 
        \ScanLink99[20] , \ScanLink99[19] , \ScanLink99[18] , \ScanLink99[17] , 
        \ScanLink99[16] , \ScanLink99[15] , \ScanLink99[14] , \ScanLink99[13] , 
        \ScanLink99[12] , \ScanLink99[11] , \ScanLink99[10] , \ScanLink99[9] , 
        \ScanLink99[8] , \ScanLink99[7] , \ScanLink99[6] , \ScanLink99[5] , 
        \ScanLink99[4] , \ScanLink99[3] , \ScanLink99[2] , \ScanLink99[1] , 
        \ScanLink99[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({
        \wRegOut_6_36[31] , \wRegOut_6_36[30] , \wRegOut_6_36[29] , 
        \wRegOut_6_36[28] , \wRegOut_6_36[27] , \wRegOut_6_36[26] , 
        \wRegOut_6_36[25] , \wRegOut_6_36[24] , \wRegOut_6_36[23] , 
        \wRegOut_6_36[22] , \wRegOut_6_36[21] , \wRegOut_6_36[20] , 
        \wRegOut_6_36[19] , \wRegOut_6_36[18] , \wRegOut_6_36[17] , 
        \wRegOut_6_36[16] , \wRegOut_6_36[15] , \wRegOut_6_36[14] , 
        \wRegOut_6_36[13] , \wRegOut_6_36[12] , \wRegOut_6_36[11] , 
        \wRegOut_6_36[10] , \wRegOut_6_36[9] , \wRegOut_6_36[8] , 
        \wRegOut_6_36[7] , \wRegOut_6_36[6] , \wRegOut_6_36[5] , 
        \wRegOut_6_36[4] , \wRegOut_6_36[3] , \wRegOut_6_36[2] , 
        \wRegOut_6_36[1] , \wRegOut_6_36[0] }), .Enable1(\wRegEnTop_6_36[0] ), 
        .Enable2(\wRegEnBot_6_36[0] ), .In1({\wRegInTop_6_36[31] , 
        \wRegInTop_6_36[30] , \wRegInTop_6_36[29] , \wRegInTop_6_36[28] , 
        \wRegInTop_6_36[27] , \wRegInTop_6_36[26] , \wRegInTop_6_36[25] , 
        \wRegInTop_6_36[24] , \wRegInTop_6_36[23] , \wRegInTop_6_36[22] , 
        \wRegInTop_6_36[21] , \wRegInTop_6_36[20] , \wRegInTop_6_36[19] , 
        \wRegInTop_6_36[18] , \wRegInTop_6_36[17] , \wRegInTop_6_36[16] , 
        \wRegInTop_6_36[15] , \wRegInTop_6_36[14] , \wRegInTop_6_36[13] , 
        \wRegInTop_6_36[12] , \wRegInTop_6_36[11] , \wRegInTop_6_36[10] , 
        \wRegInTop_6_36[9] , \wRegInTop_6_36[8] , \wRegInTop_6_36[7] , 
        \wRegInTop_6_36[6] , \wRegInTop_6_36[5] , \wRegInTop_6_36[4] , 
        \wRegInTop_6_36[3] , \wRegInTop_6_36[2] , \wRegInTop_6_36[1] , 
        \wRegInTop_6_36[0] }), .In2({\wRegInBot_6_36[31] , 
        \wRegInBot_6_36[30] , \wRegInBot_6_36[29] , \wRegInBot_6_36[28] , 
        \wRegInBot_6_36[27] , \wRegInBot_6_36[26] , \wRegInBot_6_36[25] , 
        \wRegInBot_6_36[24] , \wRegInBot_6_36[23] , \wRegInBot_6_36[22] , 
        \wRegInBot_6_36[21] , \wRegInBot_6_36[20] , \wRegInBot_6_36[19] , 
        \wRegInBot_6_36[18] , \wRegInBot_6_36[17] , \wRegInBot_6_36[16] , 
        \wRegInBot_6_36[15] , \wRegInBot_6_36[14] , \wRegInBot_6_36[13] , 
        \wRegInBot_6_36[12] , \wRegInBot_6_36[11] , \wRegInBot_6_36[10] , 
        \wRegInBot_6_36[9] , \wRegInBot_6_36[8] , \wRegInBot_6_36[7] , 
        \wRegInBot_6_36[6] , \wRegInBot_6_36[5] , \wRegInBot_6_36[4] , 
        \wRegInBot_6_36[3] , \wRegInBot_6_36[2] , \wRegInBot_6_36[1] , 
        \wRegInBot_6_36[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_43 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink107[31] , \ScanLink107[30] , \ScanLink107[29] , 
        \ScanLink107[28] , \ScanLink107[27] , \ScanLink107[26] , 
        \ScanLink107[25] , \ScanLink107[24] , \ScanLink107[23] , 
        \ScanLink107[22] , \ScanLink107[21] , \ScanLink107[20] , 
        \ScanLink107[19] , \ScanLink107[18] , \ScanLink107[17] , 
        \ScanLink107[16] , \ScanLink107[15] , \ScanLink107[14] , 
        \ScanLink107[13] , \ScanLink107[12] , \ScanLink107[11] , 
        \ScanLink107[10] , \ScanLink107[9] , \ScanLink107[8] , 
        \ScanLink107[7] , \ScanLink107[6] , \ScanLink107[5] , \ScanLink107[4] , 
        \ScanLink107[3] , \ScanLink107[2] , \ScanLink107[1] , \ScanLink107[0] 
        }), .ScanOut({\ScanLink106[31] , \ScanLink106[30] , \ScanLink106[29] , 
        \ScanLink106[28] , \ScanLink106[27] , \ScanLink106[26] , 
        \ScanLink106[25] , \ScanLink106[24] , \ScanLink106[23] , 
        \ScanLink106[22] , \ScanLink106[21] , \ScanLink106[20] , 
        \ScanLink106[19] , \ScanLink106[18] , \ScanLink106[17] , 
        \ScanLink106[16] , \ScanLink106[15] , \ScanLink106[14] , 
        \ScanLink106[13] , \ScanLink106[12] , \ScanLink106[11] , 
        \ScanLink106[10] , \ScanLink106[9] , \ScanLink106[8] , 
        \ScanLink106[7] , \ScanLink106[6] , \ScanLink106[5] , \ScanLink106[4] , 
        \ScanLink106[3] , \ScanLink106[2] , \ScanLink106[1] , \ScanLink106[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_43[31] , 
        \wRegOut_6_43[30] , \wRegOut_6_43[29] , \wRegOut_6_43[28] , 
        \wRegOut_6_43[27] , \wRegOut_6_43[26] , \wRegOut_6_43[25] , 
        \wRegOut_6_43[24] , \wRegOut_6_43[23] , \wRegOut_6_43[22] , 
        \wRegOut_6_43[21] , \wRegOut_6_43[20] , \wRegOut_6_43[19] , 
        \wRegOut_6_43[18] , \wRegOut_6_43[17] , \wRegOut_6_43[16] , 
        \wRegOut_6_43[15] , \wRegOut_6_43[14] , \wRegOut_6_43[13] , 
        \wRegOut_6_43[12] , \wRegOut_6_43[11] , \wRegOut_6_43[10] , 
        \wRegOut_6_43[9] , \wRegOut_6_43[8] , \wRegOut_6_43[7] , 
        \wRegOut_6_43[6] , \wRegOut_6_43[5] , \wRegOut_6_43[4] , 
        \wRegOut_6_43[3] , \wRegOut_6_43[2] , \wRegOut_6_43[1] , 
        \wRegOut_6_43[0] }), .Enable1(\wRegEnTop_6_43[0] ), .Enable2(
        \wRegEnBot_6_43[0] ), .In1({\wRegInTop_6_43[31] , \wRegInTop_6_43[30] , 
        \wRegInTop_6_43[29] , \wRegInTop_6_43[28] , \wRegInTop_6_43[27] , 
        \wRegInTop_6_43[26] , \wRegInTop_6_43[25] , \wRegInTop_6_43[24] , 
        \wRegInTop_6_43[23] , \wRegInTop_6_43[22] , \wRegInTop_6_43[21] , 
        \wRegInTop_6_43[20] , \wRegInTop_6_43[19] , \wRegInTop_6_43[18] , 
        \wRegInTop_6_43[17] , \wRegInTop_6_43[16] , \wRegInTop_6_43[15] , 
        \wRegInTop_6_43[14] , \wRegInTop_6_43[13] , \wRegInTop_6_43[12] , 
        \wRegInTop_6_43[11] , \wRegInTop_6_43[10] , \wRegInTop_6_43[9] , 
        \wRegInTop_6_43[8] , \wRegInTop_6_43[7] , \wRegInTop_6_43[6] , 
        \wRegInTop_6_43[5] , \wRegInTop_6_43[4] , \wRegInTop_6_43[3] , 
        \wRegInTop_6_43[2] , \wRegInTop_6_43[1] , \wRegInTop_6_43[0] }), .In2(
        {\wRegInBot_6_43[31] , \wRegInBot_6_43[30] , \wRegInBot_6_43[29] , 
        \wRegInBot_6_43[28] , \wRegInBot_6_43[27] , \wRegInBot_6_43[26] , 
        \wRegInBot_6_43[25] , \wRegInBot_6_43[24] , \wRegInBot_6_43[23] , 
        \wRegInBot_6_43[22] , \wRegInBot_6_43[21] , \wRegInBot_6_43[20] , 
        \wRegInBot_6_43[19] , \wRegInBot_6_43[18] , \wRegInBot_6_43[17] , 
        \wRegInBot_6_43[16] , \wRegInBot_6_43[15] , \wRegInBot_6_43[14] , 
        \wRegInBot_6_43[13] , \wRegInBot_6_43[12] , \wRegInBot_6_43[11] , 
        \wRegInBot_6_43[10] , \wRegInBot_6_43[9] , \wRegInBot_6_43[8] , 
        \wRegInBot_6_43[7] , \wRegInBot_6_43[6] , \wRegInBot_6_43[5] , 
        \wRegInBot_6_43[4] , \wRegInBot_6_43[3] , \wRegInBot_6_43[2] , 
        \wRegInBot_6_43[1] , \wRegInBot_6_43[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_59 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink187[31] , \ScanLink187[30] , \ScanLink187[29] , 
        \ScanLink187[28] , \ScanLink187[27] , \ScanLink187[26] , 
        \ScanLink187[25] , \ScanLink187[24] , \ScanLink187[23] , 
        \ScanLink187[22] , \ScanLink187[21] , \ScanLink187[20] , 
        \ScanLink187[19] , \ScanLink187[18] , \ScanLink187[17] , 
        \ScanLink187[16] , \ScanLink187[15] , \ScanLink187[14] , 
        \ScanLink187[13] , \ScanLink187[12] , \ScanLink187[11] , 
        \ScanLink187[10] , \ScanLink187[9] , \ScanLink187[8] , 
        \ScanLink187[7] , \ScanLink187[6] , \ScanLink187[5] , \ScanLink187[4] , 
        \ScanLink187[3] , \ScanLink187[2] , \ScanLink187[1] , \ScanLink187[0] 
        }), .ScanOut({\ScanLink186[31] , \ScanLink186[30] , \ScanLink186[29] , 
        \ScanLink186[28] , \ScanLink186[27] , \ScanLink186[26] , 
        \ScanLink186[25] , \ScanLink186[24] , \ScanLink186[23] , 
        \ScanLink186[22] , \ScanLink186[21] , \ScanLink186[20] , 
        \ScanLink186[19] , \ScanLink186[18] , \ScanLink186[17] , 
        \ScanLink186[16] , \ScanLink186[15] , \ScanLink186[14] , 
        \ScanLink186[13] , \ScanLink186[12] , \ScanLink186[11] , 
        \ScanLink186[10] , \ScanLink186[9] , \ScanLink186[8] , 
        \ScanLink186[7] , \ScanLink186[6] , \ScanLink186[5] , \ScanLink186[4] , 
        \ScanLink186[3] , \ScanLink186[2] , \ScanLink186[1] , \ScanLink186[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_59[31] , 
        \wRegOut_7_59[30] , \wRegOut_7_59[29] , \wRegOut_7_59[28] , 
        \wRegOut_7_59[27] , \wRegOut_7_59[26] , \wRegOut_7_59[25] , 
        \wRegOut_7_59[24] , \wRegOut_7_59[23] , \wRegOut_7_59[22] , 
        \wRegOut_7_59[21] , \wRegOut_7_59[20] , \wRegOut_7_59[19] , 
        \wRegOut_7_59[18] , \wRegOut_7_59[17] , \wRegOut_7_59[16] , 
        \wRegOut_7_59[15] , \wRegOut_7_59[14] , \wRegOut_7_59[13] , 
        \wRegOut_7_59[12] , \wRegOut_7_59[11] , \wRegOut_7_59[10] , 
        \wRegOut_7_59[9] , \wRegOut_7_59[8] , \wRegOut_7_59[7] , 
        \wRegOut_7_59[6] , \wRegOut_7_59[5] , \wRegOut_7_59[4] , 
        \wRegOut_7_59[3] , \wRegOut_7_59[2] , \wRegOut_7_59[1] , 
        \wRegOut_7_59[0] }), .Enable1(\wRegEnTop_7_59[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_59[31] , \wRegInTop_7_59[30] , \wRegInTop_7_59[29] , 
        \wRegInTop_7_59[28] , \wRegInTop_7_59[27] , \wRegInTop_7_59[26] , 
        \wRegInTop_7_59[25] , \wRegInTop_7_59[24] , \wRegInTop_7_59[23] , 
        \wRegInTop_7_59[22] , \wRegInTop_7_59[21] , \wRegInTop_7_59[20] , 
        \wRegInTop_7_59[19] , \wRegInTop_7_59[18] , \wRegInTop_7_59[17] , 
        \wRegInTop_7_59[16] , \wRegInTop_7_59[15] , \wRegInTop_7_59[14] , 
        \wRegInTop_7_59[13] , \wRegInTop_7_59[12] , \wRegInTop_7_59[11] , 
        \wRegInTop_7_59[10] , \wRegInTop_7_59[9] , \wRegInTop_7_59[8] , 
        \wRegInTop_7_59[7] , \wRegInTop_7_59[6] , \wRegInTop_7_59[5] , 
        \wRegInTop_7_59[4] , \wRegInTop_7_59[3] , \wRegInTop_7_59[2] , 
        \wRegInTop_7_59[1] , \wRegInTop_7_59[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_58 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink122[31] , \ScanLink122[30] , \ScanLink122[29] , 
        \ScanLink122[28] , \ScanLink122[27] , \ScanLink122[26] , 
        \ScanLink122[25] , \ScanLink122[24] , \ScanLink122[23] , 
        \ScanLink122[22] , \ScanLink122[21] , \ScanLink122[20] , 
        \ScanLink122[19] , \ScanLink122[18] , \ScanLink122[17] , 
        \ScanLink122[16] , \ScanLink122[15] , \ScanLink122[14] , 
        \ScanLink122[13] , \ScanLink122[12] , \ScanLink122[11] , 
        \ScanLink122[10] , \ScanLink122[9] , \ScanLink122[8] , 
        \ScanLink122[7] , \ScanLink122[6] , \ScanLink122[5] , \ScanLink122[4] , 
        \ScanLink122[3] , \ScanLink122[2] , \ScanLink122[1] , \ScanLink122[0] 
        }), .ScanOut({\ScanLink121[31] , \ScanLink121[30] , \ScanLink121[29] , 
        \ScanLink121[28] , \ScanLink121[27] , \ScanLink121[26] , 
        \ScanLink121[25] , \ScanLink121[24] , \ScanLink121[23] , 
        \ScanLink121[22] , \ScanLink121[21] , \ScanLink121[20] , 
        \ScanLink121[19] , \ScanLink121[18] , \ScanLink121[17] , 
        \ScanLink121[16] , \ScanLink121[15] , \ScanLink121[14] , 
        \ScanLink121[13] , \ScanLink121[12] , \ScanLink121[11] , 
        \ScanLink121[10] , \ScanLink121[9] , \ScanLink121[8] , 
        \ScanLink121[7] , \ScanLink121[6] , \ScanLink121[5] , \ScanLink121[4] , 
        \ScanLink121[3] , \ScanLink121[2] , \ScanLink121[1] , \ScanLink121[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_58[31] , 
        \wRegOut_6_58[30] , \wRegOut_6_58[29] , \wRegOut_6_58[28] , 
        \wRegOut_6_58[27] , \wRegOut_6_58[26] , \wRegOut_6_58[25] , 
        \wRegOut_6_58[24] , \wRegOut_6_58[23] , \wRegOut_6_58[22] , 
        \wRegOut_6_58[21] , \wRegOut_6_58[20] , \wRegOut_6_58[19] , 
        \wRegOut_6_58[18] , \wRegOut_6_58[17] , \wRegOut_6_58[16] , 
        \wRegOut_6_58[15] , \wRegOut_6_58[14] , \wRegOut_6_58[13] , 
        \wRegOut_6_58[12] , \wRegOut_6_58[11] , \wRegOut_6_58[10] , 
        \wRegOut_6_58[9] , \wRegOut_6_58[8] , \wRegOut_6_58[7] , 
        \wRegOut_6_58[6] , \wRegOut_6_58[5] , \wRegOut_6_58[4] , 
        \wRegOut_6_58[3] , \wRegOut_6_58[2] , \wRegOut_6_58[1] , 
        \wRegOut_6_58[0] }), .Enable1(\wRegEnTop_6_58[0] ), .Enable2(
        \wRegEnBot_6_58[0] ), .In1({\wRegInTop_6_58[31] , \wRegInTop_6_58[30] , 
        \wRegInTop_6_58[29] , \wRegInTop_6_58[28] , \wRegInTop_6_58[27] , 
        \wRegInTop_6_58[26] , \wRegInTop_6_58[25] , \wRegInTop_6_58[24] , 
        \wRegInTop_6_58[23] , \wRegInTop_6_58[22] , \wRegInTop_6_58[21] , 
        \wRegInTop_6_58[20] , \wRegInTop_6_58[19] , \wRegInTop_6_58[18] , 
        \wRegInTop_6_58[17] , \wRegInTop_6_58[16] , \wRegInTop_6_58[15] , 
        \wRegInTop_6_58[14] , \wRegInTop_6_58[13] , \wRegInTop_6_58[12] , 
        \wRegInTop_6_58[11] , \wRegInTop_6_58[10] , \wRegInTop_6_58[9] , 
        \wRegInTop_6_58[8] , \wRegInTop_6_58[7] , \wRegInTop_6_58[6] , 
        \wRegInTop_6_58[5] , \wRegInTop_6_58[4] , \wRegInTop_6_58[3] , 
        \wRegInTop_6_58[2] , \wRegInTop_6_58[1] , \wRegInTop_6_58[0] }), .In2(
        {\wRegInBot_6_58[31] , \wRegInBot_6_58[30] , \wRegInBot_6_58[29] , 
        \wRegInBot_6_58[28] , \wRegInBot_6_58[27] , \wRegInBot_6_58[26] , 
        \wRegInBot_6_58[25] , \wRegInBot_6_58[24] , \wRegInBot_6_58[23] , 
        \wRegInBot_6_58[22] , \wRegInBot_6_58[21] , \wRegInBot_6_58[20] , 
        \wRegInBot_6_58[19] , \wRegInBot_6_58[18] , \wRegInBot_6_58[17] , 
        \wRegInBot_6_58[16] , \wRegInBot_6_58[15] , \wRegInBot_6_58[14] , 
        \wRegInBot_6_58[13] , \wRegInBot_6_58[12] , \wRegInBot_6_58[11] , 
        \wRegInBot_6_58[10] , \wRegInBot_6_58[9] , \wRegInBot_6_58[8] , 
        \wRegInBot_6_58[7] , \wRegInBot_6_58[6] , \wRegInBot_6_58[5] , 
        \wRegInBot_6_58[4] , \wRegInBot_6_58[3] , \wRegInBot_6_58[2] , 
        \wRegInBot_6_58[1] , \wRegInBot_6_58[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink138[31] , \ScanLink138[30] , \ScanLink138[29] , 
        \ScanLink138[28] , \ScanLink138[27] , \ScanLink138[26] , 
        \ScanLink138[25] , \ScanLink138[24] , \ScanLink138[23] , 
        \ScanLink138[22] , \ScanLink138[21] , \ScanLink138[20] , 
        \ScanLink138[19] , \ScanLink138[18] , \ScanLink138[17] , 
        \ScanLink138[16] , \ScanLink138[15] , \ScanLink138[14] , 
        \ScanLink138[13] , \ScanLink138[12] , \ScanLink138[11] , 
        \ScanLink138[10] , \ScanLink138[9] , \ScanLink138[8] , 
        \ScanLink138[7] , \ScanLink138[6] , \ScanLink138[5] , \ScanLink138[4] , 
        \ScanLink138[3] , \ScanLink138[2] , \ScanLink138[1] , \ScanLink138[0] 
        }), .ScanOut({\ScanLink137[31] , \ScanLink137[30] , \ScanLink137[29] , 
        \ScanLink137[28] , \ScanLink137[27] , \ScanLink137[26] , 
        \ScanLink137[25] , \ScanLink137[24] , \ScanLink137[23] , 
        \ScanLink137[22] , \ScanLink137[21] , \ScanLink137[20] , 
        \ScanLink137[19] , \ScanLink137[18] , \ScanLink137[17] , 
        \ScanLink137[16] , \ScanLink137[15] , \ScanLink137[14] , 
        \ScanLink137[13] , \ScanLink137[12] , \ScanLink137[11] , 
        \ScanLink137[10] , \ScanLink137[9] , \ScanLink137[8] , 
        \ScanLink137[7] , \ScanLink137[6] , \ScanLink137[5] , \ScanLink137[4] , 
        \ScanLink137[3] , \ScanLink137[2] , \ScanLink137[1] , \ScanLink137[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_10[31] , 
        \wRegOut_7_10[30] , \wRegOut_7_10[29] , \wRegOut_7_10[28] , 
        \wRegOut_7_10[27] , \wRegOut_7_10[26] , \wRegOut_7_10[25] , 
        \wRegOut_7_10[24] , \wRegOut_7_10[23] , \wRegOut_7_10[22] , 
        \wRegOut_7_10[21] , \wRegOut_7_10[20] , \wRegOut_7_10[19] , 
        \wRegOut_7_10[18] , \wRegOut_7_10[17] , \wRegOut_7_10[16] , 
        \wRegOut_7_10[15] , \wRegOut_7_10[14] , \wRegOut_7_10[13] , 
        \wRegOut_7_10[12] , \wRegOut_7_10[11] , \wRegOut_7_10[10] , 
        \wRegOut_7_10[9] , \wRegOut_7_10[8] , \wRegOut_7_10[7] , 
        \wRegOut_7_10[6] , \wRegOut_7_10[5] , \wRegOut_7_10[4] , 
        \wRegOut_7_10[3] , \wRegOut_7_10[2] , \wRegOut_7_10[1] , 
        \wRegOut_7_10[0] }), .Enable1(\wRegEnTop_7_10[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_10[31] , \wRegInTop_7_10[30] , \wRegInTop_7_10[29] , 
        \wRegInTop_7_10[28] , \wRegInTop_7_10[27] , \wRegInTop_7_10[26] , 
        \wRegInTop_7_10[25] , \wRegInTop_7_10[24] , \wRegInTop_7_10[23] , 
        \wRegInTop_7_10[22] , \wRegInTop_7_10[21] , \wRegInTop_7_10[20] , 
        \wRegInTop_7_10[19] , \wRegInTop_7_10[18] , \wRegInTop_7_10[17] , 
        \wRegInTop_7_10[16] , \wRegInTop_7_10[15] , \wRegInTop_7_10[14] , 
        \wRegInTop_7_10[13] , \wRegInTop_7_10[12] , \wRegInTop_7_10[11] , 
        \wRegInTop_7_10[10] , \wRegInTop_7_10[9] , \wRegInTop_7_10[8] , 
        \wRegInTop_7_10[7] , \wRegInTop_7_10[6] , \wRegInTop_7_10[5] , 
        \wRegInTop_7_10[4] , \wRegInTop_7_10[3] , \wRegInTop_7_10[2] , 
        \wRegInTop_7_10[1] , \wRegInTop_7_10[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_37 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink165[31] , \ScanLink165[30] , \ScanLink165[29] , 
        \ScanLink165[28] , \ScanLink165[27] , \ScanLink165[26] , 
        \ScanLink165[25] , \ScanLink165[24] , \ScanLink165[23] , 
        \ScanLink165[22] , \ScanLink165[21] , \ScanLink165[20] , 
        \ScanLink165[19] , \ScanLink165[18] , \ScanLink165[17] , 
        \ScanLink165[16] , \ScanLink165[15] , \ScanLink165[14] , 
        \ScanLink165[13] , \ScanLink165[12] , \ScanLink165[11] , 
        \ScanLink165[10] , \ScanLink165[9] , \ScanLink165[8] , 
        \ScanLink165[7] , \ScanLink165[6] , \ScanLink165[5] , \ScanLink165[4] , 
        \ScanLink165[3] , \ScanLink165[2] , \ScanLink165[1] , \ScanLink165[0] 
        }), .ScanOut({\ScanLink164[31] , \ScanLink164[30] , \ScanLink164[29] , 
        \ScanLink164[28] , \ScanLink164[27] , \ScanLink164[26] , 
        \ScanLink164[25] , \ScanLink164[24] , \ScanLink164[23] , 
        \ScanLink164[22] , \ScanLink164[21] , \ScanLink164[20] , 
        \ScanLink164[19] , \ScanLink164[18] , \ScanLink164[17] , 
        \ScanLink164[16] , \ScanLink164[15] , \ScanLink164[14] , 
        \ScanLink164[13] , \ScanLink164[12] , \ScanLink164[11] , 
        \ScanLink164[10] , \ScanLink164[9] , \ScanLink164[8] , 
        \ScanLink164[7] , \ScanLink164[6] , \ScanLink164[5] , \ScanLink164[4] , 
        \ScanLink164[3] , \ScanLink164[2] , \ScanLink164[1] , \ScanLink164[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_37[31] , 
        \wRegOut_7_37[30] , \wRegOut_7_37[29] , \wRegOut_7_37[28] , 
        \wRegOut_7_37[27] , \wRegOut_7_37[26] , \wRegOut_7_37[25] , 
        \wRegOut_7_37[24] , \wRegOut_7_37[23] , \wRegOut_7_37[22] , 
        \wRegOut_7_37[21] , \wRegOut_7_37[20] , \wRegOut_7_37[19] , 
        \wRegOut_7_37[18] , \wRegOut_7_37[17] , \wRegOut_7_37[16] , 
        \wRegOut_7_37[15] , \wRegOut_7_37[14] , \wRegOut_7_37[13] , 
        \wRegOut_7_37[12] , \wRegOut_7_37[11] , \wRegOut_7_37[10] , 
        \wRegOut_7_37[9] , \wRegOut_7_37[8] , \wRegOut_7_37[7] , 
        \wRegOut_7_37[6] , \wRegOut_7_37[5] , \wRegOut_7_37[4] , 
        \wRegOut_7_37[3] , \wRegOut_7_37[2] , \wRegOut_7_37[1] , 
        \wRegOut_7_37[0] }), .Enable1(\wRegEnTop_7_37[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_37[31] , \wRegInTop_7_37[30] , \wRegInTop_7_37[29] , 
        \wRegInTop_7_37[28] , \wRegInTop_7_37[27] , \wRegInTop_7_37[26] , 
        \wRegInTop_7_37[25] , \wRegInTop_7_37[24] , \wRegInTop_7_37[23] , 
        \wRegInTop_7_37[22] , \wRegInTop_7_37[21] , \wRegInTop_7_37[20] , 
        \wRegInTop_7_37[19] , \wRegInTop_7_37[18] , \wRegInTop_7_37[17] , 
        \wRegInTop_7_37[16] , \wRegInTop_7_37[15] , \wRegInTop_7_37[14] , 
        \wRegInTop_7_37[13] , \wRegInTop_7_37[12] , \wRegInTop_7_37[11] , 
        \wRegInTop_7_37[10] , \wRegInTop_7_37[9] , \wRegInTop_7_37[8] , 
        \wRegInTop_7_37[7] , \wRegInTop_7_37[6] , \wRegInTop_7_37[5] , 
        \wRegInTop_7_37[4] , \wRegInTop_7_37[3] , \wRegInTop_7_37[2] , 
        \wRegInTop_7_37[1] , \wRegInTop_7_37[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_123 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink251[31] , \ScanLink251[30] , \ScanLink251[29] , 
        \ScanLink251[28] , \ScanLink251[27] , \ScanLink251[26] , 
        \ScanLink251[25] , \ScanLink251[24] , \ScanLink251[23] , 
        \ScanLink251[22] , \ScanLink251[21] , \ScanLink251[20] , 
        \ScanLink251[19] , \ScanLink251[18] , \ScanLink251[17] , 
        \ScanLink251[16] , \ScanLink251[15] , \ScanLink251[14] , 
        \ScanLink251[13] , \ScanLink251[12] , \ScanLink251[11] , 
        \ScanLink251[10] , \ScanLink251[9] , \ScanLink251[8] , 
        \ScanLink251[7] , \ScanLink251[6] , \ScanLink251[5] , \ScanLink251[4] , 
        \ScanLink251[3] , \ScanLink251[2] , \ScanLink251[1] , \ScanLink251[0] 
        }), .ScanOut({\ScanLink250[31] , \ScanLink250[30] , \ScanLink250[29] , 
        \ScanLink250[28] , \ScanLink250[27] , \ScanLink250[26] , 
        \ScanLink250[25] , \ScanLink250[24] , \ScanLink250[23] , 
        \ScanLink250[22] , \ScanLink250[21] , \ScanLink250[20] , 
        \ScanLink250[19] , \ScanLink250[18] , \ScanLink250[17] , 
        \ScanLink250[16] , \ScanLink250[15] , \ScanLink250[14] , 
        \ScanLink250[13] , \ScanLink250[12] , \ScanLink250[11] , 
        \ScanLink250[10] , \ScanLink250[9] , \ScanLink250[8] , 
        \ScanLink250[7] , \ScanLink250[6] , \ScanLink250[5] , \ScanLink250[4] , 
        \ScanLink250[3] , \ScanLink250[2] , \ScanLink250[1] , \ScanLink250[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_123[31] , 
        \wRegOut_7_123[30] , \wRegOut_7_123[29] , \wRegOut_7_123[28] , 
        \wRegOut_7_123[27] , \wRegOut_7_123[26] , \wRegOut_7_123[25] , 
        \wRegOut_7_123[24] , \wRegOut_7_123[23] , \wRegOut_7_123[22] , 
        \wRegOut_7_123[21] , \wRegOut_7_123[20] , \wRegOut_7_123[19] , 
        \wRegOut_7_123[18] , \wRegOut_7_123[17] , \wRegOut_7_123[16] , 
        \wRegOut_7_123[15] , \wRegOut_7_123[14] , \wRegOut_7_123[13] , 
        \wRegOut_7_123[12] , \wRegOut_7_123[11] , \wRegOut_7_123[10] , 
        \wRegOut_7_123[9] , \wRegOut_7_123[8] , \wRegOut_7_123[7] , 
        \wRegOut_7_123[6] , \wRegOut_7_123[5] , \wRegOut_7_123[4] , 
        \wRegOut_7_123[3] , \wRegOut_7_123[2] , \wRegOut_7_123[1] , 
        \wRegOut_7_123[0] }), .Enable1(\wRegEnTop_7_123[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_123[31] , \wRegInTop_7_123[30] , 
        \wRegInTop_7_123[29] , \wRegInTop_7_123[28] , \wRegInTop_7_123[27] , 
        \wRegInTop_7_123[26] , \wRegInTop_7_123[25] , \wRegInTop_7_123[24] , 
        \wRegInTop_7_123[23] , \wRegInTop_7_123[22] , \wRegInTop_7_123[21] , 
        \wRegInTop_7_123[20] , \wRegInTop_7_123[19] , \wRegInTop_7_123[18] , 
        \wRegInTop_7_123[17] , \wRegInTop_7_123[16] , \wRegInTop_7_123[15] , 
        \wRegInTop_7_123[14] , \wRegInTop_7_123[13] , \wRegInTop_7_123[12] , 
        \wRegInTop_7_123[11] , \wRegInTop_7_123[10] , \wRegInTop_7_123[9] , 
        \wRegInTop_7_123[8] , \wRegInTop_7_123[7] , \wRegInTop_7_123[6] , 
        \wRegInTop_7_123[5] , \wRegInTop_7_123[4] , \wRegInTop_7_123[3] , 
        \wRegInTop_7_123[2] , \wRegInTop_7_123[1] , \wRegInTop_7_123[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_104 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink232[31] , \ScanLink232[30] , \ScanLink232[29] , 
        \ScanLink232[28] , \ScanLink232[27] , \ScanLink232[26] , 
        \ScanLink232[25] , \ScanLink232[24] , \ScanLink232[23] , 
        \ScanLink232[22] , \ScanLink232[21] , \ScanLink232[20] , 
        \ScanLink232[19] , \ScanLink232[18] , \ScanLink232[17] , 
        \ScanLink232[16] , \ScanLink232[15] , \ScanLink232[14] , 
        \ScanLink232[13] , \ScanLink232[12] , \ScanLink232[11] , 
        \ScanLink232[10] , \ScanLink232[9] , \ScanLink232[8] , 
        \ScanLink232[7] , \ScanLink232[6] , \ScanLink232[5] , \ScanLink232[4] , 
        \ScanLink232[3] , \ScanLink232[2] , \ScanLink232[1] , \ScanLink232[0] 
        }), .ScanOut({\ScanLink231[31] , \ScanLink231[30] , \ScanLink231[29] , 
        \ScanLink231[28] , \ScanLink231[27] , \ScanLink231[26] , 
        \ScanLink231[25] , \ScanLink231[24] , \ScanLink231[23] , 
        \ScanLink231[22] , \ScanLink231[21] , \ScanLink231[20] , 
        \ScanLink231[19] , \ScanLink231[18] , \ScanLink231[17] , 
        \ScanLink231[16] , \ScanLink231[15] , \ScanLink231[14] , 
        \ScanLink231[13] , \ScanLink231[12] , \ScanLink231[11] , 
        \ScanLink231[10] , \ScanLink231[9] , \ScanLink231[8] , 
        \ScanLink231[7] , \ScanLink231[6] , \ScanLink231[5] , \ScanLink231[4] , 
        \ScanLink231[3] , \ScanLink231[2] , \ScanLink231[1] , \ScanLink231[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_104[31] , 
        \wRegOut_7_104[30] , \wRegOut_7_104[29] , \wRegOut_7_104[28] , 
        \wRegOut_7_104[27] , \wRegOut_7_104[26] , \wRegOut_7_104[25] , 
        \wRegOut_7_104[24] , \wRegOut_7_104[23] , \wRegOut_7_104[22] , 
        \wRegOut_7_104[21] , \wRegOut_7_104[20] , \wRegOut_7_104[19] , 
        \wRegOut_7_104[18] , \wRegOut_7_104[17] , \wRegOut_7_104[16] , 
        \wRegOut_7_104[15] , \wRegOut_7_104[14] , \wRegOut_7_104[13] , 
        \wRegOut_7_104[12] , \wRegOut_7_104[11] , \wRegOut_7_104[10] , 
        \wRegOut_7_104[9] , \wRegOut_7_104[8] , \wRegOut_7_104[7] , 
        \wRegOut_7_104[6] , \wRegOut_7_104[5] , \wRegOut_7_104[4] , 
        \wRegOut_7_104[3] , \wRegOut_7_104[2] , \wRegOut_7_104[1] , 
        \wRegOut_7_104[0] }), .Enable1(\wRegEnTop_7_104[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_104[31] , \wRegInTop_7_104[30] , 
        \wRegInTop_7_104[29] , \wRegInTop_7_104[28] , \wRegInTop_7_104[27] , 
        \wRegInTop_7_104[26] , \wRegInTop_7_104[25] , \wRegInTop_7_104[24] , 
        \wRegInTop_7_104[23] , \wRegInTop_7_104[22] , \wRegInTop_7_104[21] , 
        \wRegInTop_7_104[20] , \wRegInTop_7_104[19] , \wRegInTop_7_104[18] , 
        \wRegInTop_7_104[17] , \wRegInTop_7_104[16] , \wRegInTop_7_104[15] , 
        \wRegInTop_7_104[14] , \wRegInTop_7_104[13] , \wRegInTop_7_104[12] , 
        \wRegInTop_7_104[11] , \wRegInTop_7_104[10] , \wRegInTop_7_104[9] , 
        \wRegInTop_7_104[8] , \wRegInTop_7_104[7] , \wRegInTop_7_104[6] , 
        \wRegInTop_7_104[5] , \wRegInTop_7_104[4] , \wRegInTop_7_104[3] , 
        \wRegInTop_7_104[2] , \wRegInTop_7_104[1] , \wRegInTop_7_104[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_CtrlReg_WIDTH32 BHCR_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_5[0] ), 
        .Out(\wCtrlOut_4[0] ), .Enable(\wEnable_4[0] ) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_80 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink208[31] , \ScanLink208[30] , \ScanLink208[29] , 
        \ScanLink208[28] , \ScanLink208[27] , \ScanLink208[26] , 
        \ScanLink208[25] , \ScanLink208[24] , \ScanLink208[23] , 
        \ScanLink208[22] , \ScanLink208[21] , \ScanLink208[20] , 
        \ScanLink208[19] , \ScanLink208[18] , \ScanLink208[17] , 
        \ScanLink208[16] , \ScanLink208[15] , \ScanLink208[14] , 
        \ScanLink208[13] , \ScanLink208[12] , \ScanLink208[11] , 
        \ScanLink208[10] , \ScanLink208[9] , \ScanLink208[8] , 
        \ScanLink208[7] , \ScanLink208[6] , \ScanLink208[5] , \ScanLink208[4] , 
        \ScanLink208[3] , \ScanLink208[2] , \ScanLink208[1] , \ScanLink208[0] 
        }), .ScanOut({\ScanLink207[31] , \ScanLink207[30] , \ScanLink207[29] , 
        \ScanLink207[28] , \ScanLink207[27] , \ScanLink207[26] , 
        \ScanLink207[25] , \ScanLink207[24] , \ScanLink207[23] , 
        \ScanLink207[22] , \ScanLink207[21] , \ScanLink207[20] , 
        \ScanLink207[19] , \ScanLink207[18] , \ScanLink207[17] , 
        \ScanLink207[16] , \ScanLink207[15] , \ScanLink207[14] , 
        \ScanLink207[13] , \ScanLink207[12] , \ScanLink207[11] , 
        \ScanLink207[10] , \ScanLink207[9] , \ScanLink207[8] , 
        \ScanLink207[7] , \ScanLink207[6] , \ScanLink207[5] , \ScanLink207[4] , 
        \ScanLink207[3] , \ScanLink207[2] , \ScanLink207[1] , \ScanLink207[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_80[31] , 
        \wRegOut_7_80[30] , \wRegOut_7_80[29] , \wRegOut_7_80[28] , 
        \wRegOut_7_80[27] , \wRegOut_7_80[26] , \wRegOut_7_80[25] , 
        \wRegOut_7_80[24] , \wRegOut_7_80[23] , \wRegOut_7_80[22] , 
        \wRegOut_7_80[21] , \wRegOut_7_80[20] , \wRegOut_7_80[19] , 
        \wRegOut_7_80[18] , \wRegOut_7_80[17] , \wRegOut_7_80[16] , 
        \wRegOut_7_80[15] , \wRegOut_7_80[14] , \wRegOut_7_80[13] , 
        \wRegOut_7_80[12] , \wRegOut_7_80[11] , \wRegOut_7_80[10] , 
        \wRegOut_7_80[9] , \wRegOut_7_80[8] , \wRegOut_7_80[7] , 
        \wRegOut_7_80[6] , \wRegOut_7_80[5] , \wRegOut_7_80[4] , 
        \wRegOut_7_80[3] , \wRegOut_7_80[2] , \wRegOut_7_80[1] , 
        \wRegOut_7_80[0] }), .Enable1(\wRegEnTop_7_80[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_80[31] , \wRegInTop_7_80[30] , \wRegInTop_7_80[29] , 
        \wRegInTop_7_80[28] , \wRegInTop_7_80[27] , \wRegInTop_7_80[26] , 
        \wRegInTop_7_80[25] , \wRegInTop_7_80[24] , \wRegInTop_7_80[23] , 
        \wRegInTop_7_80[22] , \wRegInTop_7_80[21] , \wRegInTop_7_80[20] , 
        \wRegInTop_7_80[19] , \wRegInTop_7_80[18] , \wRegInTop_7_80[17] , 
        \wRegInTop_7_80[16] , \wRegInTop_7_80[15] , \wRegInTop_7_80[14] , 
        \wRegInTop_7_80[13] , \wRegInTop_7_80[12] , \wRegInTop_7_80[11] , 
        \wRegInTop_7_80[10] , \wRegInTop_7_80[9] , \wRegInTop_7_80[8] , 
        \wRegInTop_7_80[7] , \wRegInTop_7_80[6] , \wRegInTop_7_80[5] , 
        \wRegInTop_7_80[4] , \wRegInTop_7_80[3] , \wRegInTop_7_80[2] , 
        \wRegInTop_7_80[1] , \wRegInTop_7_80[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_2[0] ), .P_WR(\wRegEnBot_2_0[0] ), .P_In({\wRegOut_2_0[31] , 
        \wRegOut_2_0[30] , \wRegOut_2_0[29] , \wRegOut_2_0[28] , 
        \wRegOut_2_0[27] , \wRegOut_2_0[26] , \wRegOut_2_0[25] , 
        \wRegOut_2_0[24] , \wRegOut_2_0[23] , \wRegOut_2_0[22] , 
        \wRegOut_2_0[21] , \wRegOut_2_0[20] , \wRegOut_2_0[19] , 
        \wRegOut_2_0[18] , \wRegOut_2_0[17] , \wRegOut_2_0[16] , 
        \wRegOut_2_0[15] , \wRegOut_2_0[14] , \wRegOut_2_0[13] , 
        \wRegOut_2_0[12] , \wRegOut_2_0[11] , \wRegOut_2_0[10] , 
        \wRegOut_2_0[9] , \wRegOut_2_0[8] , \wRegOut_2_0[7] , \wRegOut_2_0[6] , 
        \wRegOut_2_0[5] , \wRegOut_2_0[4] , \wRegOut_2_0[3] , \wRegOut_2_0[2] , 
        \wRegOut_2_0[1] , \wRegOut_2_0[0] }), .P_Out({\wRegInBot_2_0[31] , 
        \wRegInBot_2_0[30] , \wRegInBot_2_0[29] , \wRegInBot_2_0[28] , 
        \wRegInBot_2_0[27] , \wRegInBot_2_0[26] , \wRegInBot_2_0[25] , 
        \wRegInBot_2_0[24] , \wRegInBot_2_0[23] , \wRegInBot_2_0[22] , 
        \wRegInBot_2_0[21] , \wRegInBot_2_0[20] , \wRegInBot_2_0[19] , 
        \wRegInBot_2_0[18] , \wRegInBot_2_0[17] , \wRegInBot_2_0[16] , 
        \wRegInBot_2_0[15] , \wRegInBot_2_0[14] , \wRegInBot_2_0[13] , 
        \wRegInBot_2_0[12] , \wRegInBot_2_0[11] , \wRegInBot_2_0[10] , 
        \wRegInBot_2_0[9] , \wRegInBot_2_0[8] , \wRegInBot_2_0[7] , 
        \wRegInBot_2_0[6] , \wRegInBot_2_0[5] , \wRegInBot_2_0[4] , 
        \wRegInBot_2_0[3] , \wRegInBot_2_0[2] , \wRegInBot_2_0[1] , 
        \wRegInBot_2_0[0] }), .L_WR(\wRegEnTop_3_0[0] ), .L_In({
        \wRegOut_3_0[31] , \wRegOut_3_0[30] , \wRegOut_3_0[29] , 
        \wRegOut_3_0[28] , \wRegOut_3_0[27] , \wRegOut_3_0[26] , 
        \wRegOut_3_0[25] , \wRegOut_3_0[24] , \wRegOut_3_0[23] , 
        \wRegOut_3_0[22] , \wRegOut_3_0[21] , \wRegOut_3_0[20] , 
        \wRegOut_3_0[19] , \wRegOut_3_0[18] , \wRegOut_3_0[17] , 
        \wRegOut_3_0[16] , \wRegOut_3_0[15] , \wRegOut_3_0[14] , 
        \wRegOut_3_0[13] , \wRegOut_3_0[12] , \wRegOut_3_0[11] , 
        \wRegOut_3_0[10] , \wRegOut_3_0[9] , \wRegOut_3_0[8] , 
        \wRegOut_3_0[7] , \wRegOut_3_0[6] , \wRegOut_3_0[5] , \wRegOut_3_0[4] , 
        \wRegOut_3_0[3] , \wRegOut_3_0[2] , \wRegOut_3_0[1] , \wRegOut_3_0[0] 
        }), .L_Out({\wRegInTop_3_0[31] , \wRegInTop_3_0[30] , 
        \wRegInTop_3_0[29] , \wRegInTop_3_0[28] , \wRegInTop_3_0[27] , 
        \wRegInTop_3_0[26] , \wRegInTop_3_0[25] , \wRegInTop_3_0[24] , 
        \wRegInTop_3_0[23] , \wRegInTop_3_0[22] , \wRegInTop_3_0[21] , 
        \wRegInTop_3_0[20] , \wRegInTop_3_0[19] , \wRegInTop_3_0[18] , 
        \wRegInTop_3_0[17] , \wRegInTop_3_0[16] , \wRegInTop_3_0[15] , 
        \wRegInTop_3_0[14] , \wRegInTop_3_0[13] , \wRegInTop_3_0[12] , 
        \wRegInTop_3_0[11] , \wRegInTop_3_0[10] , \wRegInTop_3_0[9] , 
        \wRegInTop_3_0[8] , \wRegInTop_3_0[7] , \wRegInTop_3_0[6] , 
        \wRegInTop_3_0[5] , \wRegInTop_3_0[4] , \wRegInTop_3_0[3] , 
        \wRegInTop_3_0[2] , \wRegInTop_3_0[1] , \wRegInTop_3_0[0] }), .R_WR(
        \wRegEnTop_3_1[0] ), .R_In({\wRegOut_3_1[31] , \wRegOut_3_1[30] , 
        \wRegOut_3_1[29] , \wRegOut_3_1[28] , \wRegOut_3_1[27] , 
        \wRegOut_3_1[26] , \wRegOut_3_1[25] , \wRegOut_3_1[24] , 
        \wRegOut_3_1[23] , \wRegOut_3_1[22] , \wRegOut_3_1[21] , 
        \wRegOut_3_1[20] , \wRegOut_3_1[19] , \wRegOut_3_1[18] , 
        \wRegOut_3_1[17] , \wRegOut_3_1[16] , \wRegOut_3_1[15] , 
        \wRegOut_3_1[14] , \wRegOut_3_1[13] , \wRegOut_3_1[12] , 
        \wRegOut_3_1[11] , \wRegOut_3_1[10] , \wRegOut_3_1[9] , 
        \wRegOut_3_1[8] , \wRegOut_3_1[7] , \wRegOut_3_1[6] , \wRegOut_3_1[5] , 
        \wRegOut_3_1[4] , \wRegOut_3_1[3] , \wRegOut_3_1[2] , \wRegOut_3_1[1] , 
        \wRegOut_3_1[0] }), .R_Out({\wRegInTop_3_1[31] , \wRegInTop_3_1[30] , 
        \wRegInTop_3_1[29] , \wRegInTop_3_1[28] , \wRegInTop_3_1[27] , 
        \wRegInTop_3_1[26] , \wRegInTop_3_1[25] , \wRegInTop_3_1[24] , 
        \wRegInTop_3_1[23] , \wRegInTop_3_1[22] , \wRegInTop_3_1[21] , 
        \wRegInTop_3_1[20] , \wRegInTop_3_1[19] , \wRegInTop_3_1[18] , 
        \wRegInTop_3_1[17] , \wRegInTop_3_1[16] , \wRegInTop_3_1[15] , 
        \wRegInTop_3_1[14] , \wRegInTop_3_1[13] , \wRegInTop_3_1[12] , 
        \wRegInTop_3_1[11] , \wRegInTop_3_1[10] , \wRegInTop_3_1[9] , 
        \wRegInTop_3_1[8] , \wRegInTop_3_1[7] , \wRegInTop_3_1[6] , 
        \wRegInTop_3_1[5] , \wRegInTop_3_1[4] , \wRegInTop_3_1[3] , 
        \wRegInTop_3_1[2] , \wRegInTop_3_1[1] , \wRegInTop_3_1[0] }) );
    BHeap_Node_WIDTH32 BHN_3_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_0[0] ), .P_In({\wRegOut_3_0[31] , 
        \wRegOut_3_0[30] , \wRegOut_3_0[29] , \wRegOut_3_0[28] , 
        \wRegOut_3_0[27] , \wRegOut_3_0[26] , \wRegOut_3_0[25] , 
        \wRegOut_3_0[24] , \wRegOut_3_0[23] , \wRegOut_3_0[22] , 
        \wRegOut_3_0[21] , \wRegOut_3_0[20] , \wRegOut_3_0[19] , 
        \wRegOut_3_0[18] , \wRegOut_3_0[17] , \wRegOut_3_0[16] , 
        \wRegOut_3_0[15] , \wRegOut_3_0[14] , \wRegOut_3_0[13] , 
        \wRegOut_3_0[12] , \wRegOut_3_0[11] , \wRegOut_3_0[10] , 
        \wRegOut_3_0[9] , \wRegOut_3_0[8] , \wRegOut_3_0[7] , \wRegOut_3_0[6] , 
        \wRegOut_3_0[5] , \wRegOut_3_0[4] , \wRegOut_3_0[3] , \wRegOut_3_0[2] , 
        \wRegOut_3_0[1] , \wRegOut_3_0[0] }), .P_Out({\wRegInBot_3_0[31] , 
        \wRegInBot_3_0[30] , \wRegInBot_3_0[29] , \wRegInBot_3_0[28] , 
        \wRegInBot_3_0[27] , \wRegInBot_3_0[26] , \wRegInBot_3_0[25] , 
        \wRegInBot_3_0[24] , \wRegInBot_3_0[23] , \wRegInBot_3_0[22] , 
        \wRegInBot_3_0[21] , \wRegInBot_3_0[20] , \wRegInBot_3_0[19] , 
        \wRegInBot_3_0[18] , \wRegInBot_3_0[17] , \wRegInBot_3_0[16] , 
        \wRegInBot_3_0[15] , \wRegInBot_3_0[14] , \wRegInBot_3_0[13] , 
        \wRegInBot_3_0[12] , \wRegInBot_3_0[11] , \wRegInBot_3_0[10] , 
        \wRegInBot_3_0[9] , \wRegInBot_3_0[8] , \wRegInBot_3_0[7] , 
        \wRegInBot_3_0[6] , \wRegInBot_3_0[5] , \wRegInBot_3_0[4] , 
        \wRegInBot_3_0[3] , \wRegInBot_3_0[2] , \wRegInBot_3_0[1] , 
        \wRegInBot_3_0[0] }), .L_WR(\wRegEnTop_4_0[0] ), .L_In({
        \wRegOut_4_0[31] , \wRegOut_4_0[30] , \wRegOut_4_0[29] , 
        \wRegOut_4_0[28] , \wRegOut_4_0[27] , \wRegOut_4_0[26] , 
        \wRegOut_4_0[25] , \wRegOut_4_0[24] , \wRegOut_4_0[23] , 
        \wRegOut_4_0[22] , \wRegOut_4_0[21] , \wRegOut_4_0[20] , 
        \wRegOut_4_0[19] , \wRegOut_4_0[18] , \wRegOut_4_0[17] , 
        \wRegOut_4_0[16] , \wRegOut_4_0[15] , \wRegOut_4_0[14] , 
        \wRegOut_4_0[13] , \wRegOut_4_0[12] , \wRegOut_4_0[11] , 
        \wRegOut_4_0[10] , \wRegOut_4_0[9] , \wRegOut_4_0[8] , 
        \wRegOut_4_0[7] , \wRegOut_4_0[6] , \wRegOut_4_0[5] , \wRegOut_4_0[4] , 
        \wRegOut_4_0[3] , \wRegOut_4_0[2] , \wRegOut_4_0[1] , \wRegOut_4_0[0] 
        }), .L_Out({\wRegInTop_4_0[31] , \wRegInTop_4_0[30] , 
        \wRegInTop_4_0[29] , \wRegInTop_4_0[28] , \wRegInTop_4_0[27] , 
        \wRegInTop_4_0[26] , \wRegInTop_4_0[25] , \wRegInTop_4_0[24] , 
        \wRegInTop_4_0[23] , \wRegInTop_4_0[22] , \wRegInTop_4_0[21] , 
        \wRegInTop_4_0[20] , \wRegInTop_4_0[19] , \wRegInTop_4_0[18] , 
        \wRegInTop_4_0[17] , \wRegInTop_4_0[16] , \wRegInTop_4_0[15] , 
        \wRegInTop_4_0[14] , \wRegInTop_4_0[13] , \wRegInTop_4_0[12] , 
        \wRegInTop_4_0[11] , \wRegInTop_4_0[10] , \wRegInTop_4_0[9] , 
        \wRegInTop_4_0[8] , \wRegInTop_4_0[7] , \wRegInTop_4_0[6] , 
        \wRegInTop_4_0[5] , \wRegInTop_4_0[4] , \wRegInTop_4_0[3] , 
        \wRegInTop_4_0[2] , \wRegInTop_4_0[1] , \wRegInTop_4_0[0] }), .R_WR(
        \wRegEnTop_4_1[0] ), .R_In({\wRegOut_4_1[31] , \wRegOut_4_1[30] , 
        \wRegOut_4_1[29] , \wRegOut_4_1[28] , \wRegOut_4_1[27] , 
        \wRegOut_4_1[26] , \wRegOut_4_1[25] , \wRegOut_4_1[24] , 
        \wRegOut_4_1[23] , \wRegOut_4_1[22] , \wRegOut_4_1[21] , 
        \wRegOut_4_1[20] , \wRegOut_4_1[19] , \wRegOut_4_1[18] , 
        \wRegOut_4_1[17] , \wRegOut_4_1[16] , \wRegOut_4_1[15] , 
        \wRegOut_4_1[14] , \wRegOut_4_1[13] , \wRegOut_4_1[12] , 
        \wRegOut_4_1[11] , \wRegOut_4_1[10] , \wRegOut_4_1[9] , 
        \wRegOut_4_1[8] , \wRegOut_4_1[7] , \wRegOut_4_1[6] , \wRegOut_4_1[5] , 
        \wRegOut_4_1[4] , \wRegOut_4_1[3] , \wRegOut_4_1[2] , \wRegOut_4_1[1] , 
        \wRegOut_4_1[0] }), .R_Out({\wRegInTop_4_1[31] , \wRegInTop_4_1[30] , 
        \wRegInTop_4_1[29] , \wRegInTop_4_1[28] , \wRegInTop_4_1[27] , 
        \wRegInTop_4_1[26] , \wRegInTop_4_1[25] , \wRegInTop_4_1[24] , 
        \wRegInTop_4_1[23] , \wRegInTop_4_1[22] , \wRegInTop_4_1[21] , 
        \wRegInTop_4_1[20] , \wRegInTop_4_1[19] , \wRegInTop_4_1[18] , 
        \wRegInTop_4_1[17] , \wRegInTop_4_1[16] , \wRegInTop_4_1[15] , 
        \wRegInTop_4_1[14] , \wRegInTop_4_1[13] , \wRegInTop_4_1[12] , 
        \wRegInTop_4_1[11] , \wRegInTop_4_1[10] , \wRegInTop_4_1[9] , 
        \wRegInTop_4_1[8] , \wRegInTop_4_1[7] , \wRegInTop_4_1[6] , 
        \wRegInTop_4_1[5] , \wRegInTop_4_1[4] , \wRegInTop_4_1[3] , 
        \wRegInTop_4_1[2] , \wRegInTop_4_1[1] , \wRegInTop_4_1[0] }) );
    BHeap_Node_WIDTH32 BHN_4_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_13[0] ), .P_In({\wRegOut_4_13[31] , 
        \wRegOut_4_13[30] , \wRegOut_4_13[29] , \wRegOut_4_13[28] , 
        \wRegOut_4_13[27] , \wRegOut_4_13[26] , \wRegOut_4_13[25] , 
        \wRegOut_4_13[24] , \wRegOut_4_13[23] , \wRegOut_4_13[22] , 
        \wRegOut_4_13[21] , \wRegOut_4_13[20] , \wRegOut_4_13[19] , 
        \wRegOut_4_13[18] , \wRegOut_4_13[17] , \wRegOut_4_13[16] , 
        \wRegOut_4_13[15] , \wRegOut_4_13[14] , \wRegOut_4_13[13] , 
        \wRegOut_4_13[12] , \wRegOut_4_13[11] , \wRegOut_4_13[10] , 
        \wRegOut_4_13[9] , \wRegOut_4_13[8] , \wRegOut_4_13[7] , 
        \wRegOut_4_13[6] , \wRegOut_4_13[5] , \wRegOut_4_13[4] , 
        \wRegOut_4_13[3] , \wRegOut_4_13[2] , \wRegOut_4_13[1] , 
        \wRegOut_4_13[0] }), .P_Out({\wRegInBot_4_13[31] , 
        \wRegInBot_4_13[30] , \wRegInBot_4_13[29] , \wRegInBot_4_13[28] , 
        \wRegInBot_4_13[27] , \wRegInBot_4_13[26] , \wRegInBot_4_13[25] , 
        \wRegInBot_4_13[24] , \wRegInBot_4_13[23] , \wRegInBot_4_13[22] , 
        \wRegInBot_4_13[21] , \wRegInBot_4_13[20] , \wRegInBot_4_13[19] , 
        \wRegInBot_4_13[18] , \wRegInBot_4_13[17] , \wRegInBot_4_13[16] , 
        \wRegInBot_4_13[15] , \wRegInBot_4_13[14] , \wRegInBot_4_13[13] , 
        \wRegInBot_4_13[12] , \wRegInBot_4_13[11] , \wRegInBot_4_13[10] , 
        \wRegInBot_4_13[9] , \wRegInBot_4_13[8] , \wRegInBot_4_13[7] , 
        \wRegInBot_4_13[6] , \wRegInBot_4_13[5] , \wRegInBot_4_13[4] , 
        \wRegInBot_4_13[3] , \wRegInBot_4_13[2] , \wRegInBot_4_13[1] , 
        \wRegInBot_4_13[0] }), .L_WR(\wRegEnTop_5_26[0] ), .L_In({
        \wRegOut_5_26[31] , \wRegOut_5_26[30] , \wRegOut_5_26[29] , 
        \wRegOut_5_26[28] , \wRegOut_5_26[27] , \wRegOut_5_26[26] , 
        \wRegOut_5_26[25] , \wRegOut_5_26[24] , \wRegOut_5_26[23] , 
        \wRegOut_5_26[22] , \wRegOut_5_26[21] , \wRegOut_5_26[20] , 
        \wRegOut_5_26[19] , \wRegOut_5_26[18] , \wRegOut_5_26[17] , 
        \wRegOut_5_26[16] , \wRegOut_5_26[15] , \wRegOut_5_26[14] , 
        \wRegOut_5_26[13] , \wRegOut_5_26[12] , \wRegOut_5_26[11] , 
        \wRegOut_5_26[10] , \wRegOut_5_26[9] , \wRegOut_5_26[8] , 
        \wRegOut_5_26[7] , \wRegOut_5_26[6] , \wRegOut_5_26[5] , 
        \wRegOut_5_26[4] , \wRegOut_5_26[3] , \wRegOut_5_26[2] , 
        \wRegOut_5_26[1] , \wRegOut_5_26[0] }), .L_Out({\wRegInTop_5_26[31] , 
        \wRegInTop_5_26[30] , \wRegInTop_5_26[29] , \wRegInTop_5_26[28] , 
        \wRegInTop_5_26[27] , \wRegInTop_5_26[26] , \wRegInTop_5_26[25] , 
        \wRegInTop_5_26[24] , \wRegInTop_5_26[23] , \wRegInTop_5_26[22] , 
        \wRegInTop_5_26[21] , \wRegInTop_5_26[20] , \wRegInTop_5_26[19] , 
        \wRegInTop_5_26[18] , \wRegInTop_5_26[17] , \wRegInTop_5_26[16] , 
        \wRegInTop_5_26[15] , \wRegInTop_5_26[14] , \wRegInTop_5_26[13] , 
        \wRegInTop_5_26[12] , \wRegInTop_5_26[11] , \wRegInTop_5_26[10] , 
        \wRegInTop_5_26[9] , \wRegInTop_5_26[8] , \wRegInTop_5_26[7] , 
        \wRegInTop_5_26[6] , \wRegInTop_5_26[5] , \wRegInTop_5_26[4] , 
        \wRegInTop_5_26[3] , \wRegInTop_5_26[2] , \wRegInTop_5_26[1] , 
        \wRegInTop_5_26[0] }), .R_WR(\wRegEnTop_5_27[0] ), .R_In({
        \wRegOut_5_27[31] , \wRegOut_5_27[30] , \wRegOut_5_27[29] , 
        \wRegOut_5_27[28] , \wRegOut_5_27[27] , \wRegOut_5_27[26] , 
        \wRegOut_5_27[25] , \wRegOut_5_27[24] , \wRegOut_5_27[23] , 
        \wRegOut_5_27[22] , \wRegOut_5_27[21] , \wRegOut_5_27[20] , 
        \wRegOut_5_27[19] , \wRegOut_5_27[18] , \wRegOut_5_27[17] , 
        \wRegOut_5_27[16] , \wRegOut_5_27[15] , \wRegOut_5_27[14] , 
        \wRegOut_5_27[13] , \wRegOut_5_27[12] , \wRegOut_5_27[11] , 
        \wRegOut_5_27[10] , \wRegOut_5_27[9] , \wRegOut_5_27[8] , 
        \wRegOut_5_27[7] , \wRegOut_5_27[6] , \wRegOut_5_27[5] , 
        \wRegOut_5_27[4] , \wRegOut_5_27[3] , \wRegOut_5_27[2] , 
        \wRegOut_5_27[1] , \wRegOut_5_27[0] }), .R_Out({\wRegInTop_5_27[31] , 
        \wRegInTop_5_27[30] , \wRegInTop_5_27[29] , \wRegInTop_5_27[28] , 
        \wRegInTop_5_27[27] , \wRegInTop_5_27[26] , \wRegInTop_5_27[25] , 
        \wRegInTop_5_27[24] , \wRegInTop_5_27[23] , \wRegInTop_5_27[22] , 
        \wRegInTop_5_27[21] , \wRegInTop_5_27[20] , \wRegInTop_5_27[19] , 
        \wRegInTop_5_27[18] , \wRegInTop_5_27[17] , \wRegInTop_5_27[16] , 
        \wRegInTop_5_27[15] , \wRegInTop_5_27[14] , \wRegInTop_5_27[13] , 
        \wRegInTop_5_27[12] , \wRegInTop_5_27[11] , \wRegInTop_5_27[10] , 
        \wRegInTop_5_27[9] , \wRegInTop_5_27[8] , \wRegInTop_5_27[7] , 
        \wRegInTop_5_27[6] , \wRegInTop_5_27[5] , \wRegInTop_5_27[4] , 
        \wRegInTop_5_27[3] , \wRegInTop_5_27[2] , \wRegInTop_5_27[1] , 
        \wRegInTop_5_27[0] }) );
    BHeap_Node_WIDTH32 BHN_6_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_6[0] ), .P_In({\wRegOut_6_6[31] , 
        \wRegOut_6_6[30] , \wRegOut_6_6[29] , \wRegOut_6_6[28] , 
        \wRegOut_6_6[27] , \wRegOut_6_6[26] , \wRegOut_6_6[25] , 
        \wRegOut_6_6[24] , \wRegOut_6_6[23] , \wRegOut_6_6[22] , 
        \wRegOut_6_6[21] , \wRegOut_6_6[20] , \wRegOut_6_6[19] , 
        \wRegOut_6_6[18] , \wRegOut_6_6[17] , \wRegOut_6_6[16] , 
        \wRegOut_6_6[15] , \wRegOut_6_6[14] , \wRegOut_6_6[13] , 
        \wRegOut_6_6[12] , \wRegOut_6_6[11] , \wRegOut_6_6[10] , 
        \wRegOut_6_6[9] , \wRegOut_6_6[8] , \wRegOut_6_6[7] , \wRegOut_6_6[6] , 
        \wRegOut_6_6[5] , \wRegOut_6_6[4] , \wRegOut_6_6[3] , \wRegOut_6_6[2] , 
        \wRegOut_6_6[1] , \wRegOut_6_6[0] }), .P_Out({\wRegInBot_6_6[31] , 
        \wRegInBot_6_6[30] , \wRegInBot_6_6[29] , \wRegInBot_6_6[28] , 
        \wRegInBot_6_6[27] , \wRegInBot_6_6[26] , \wRegInBot_6_6[25] , 
        \wRegInBot_6_6[24] , \wRegInBot_6_6[23] , \wRegInBot_6_6[22] , 
        \wRegInBot_6_6[21] , \wRegInBot_6_6[20] , \wRegInBot_6_6[19] , 
        \wRegInBot_6_6[18] , \wRegInBot_6_6[17] , \wRegInBot_6_6[16] , 
        \wRegInBot_6_6[15] , \wRegInBot_6_6[14] , \wRegInBot_6_6[13] , 
        \wRegInBot_6_6[12] , \wRegInBot_6_6[11] , \wRegInBot_6_6[10] , 
        \wRegInBot_6_6[9] , \wRegInBot_6_6[8] , \wRegInBot_6_6[7] , 
        \wRegInBot_6_6[6] , \wRegInBot_6_6[5] , \wRegInBot_6_6[4] , 
        \wRegInBot_6_6[3] , \wRegInBot_6_6[2] , \wRegInBot_6_6[1] , 
        \wRegInBot_6_6[0] }), .L_WR(\wRegEnTop_7_12[0] ), .L_In({
        \wRegOut_7_12[31] , \wRegOut_7_12[30] , \wRegOut_7_12[29] , 
        \wRegOut_7_12[28] , \wRegOut_7_12[27] , \wRegOut_7_12[26] , 
        \wRegOut_7_12[25] , \wRegOut_7_12[24] , \wRegOut_7_12[23] , 
        \wRegOut_7_12[22] , \wRegOut_7_12[21] , \wRegOut_7_12[20] , 
        \wRegOut_7_12[19] , \wRegOut_7_12[18] , \wRegOut_7_12[17] , 
        \wRegOut_7_12[16] , \wRegOut_7_12[15] , \wRegOut_7_12[14] , 
        \wRegOut_7_12[13] , \wRegOut_7_12[12] , \wRegOut_7_12[11] , 
        \wRegOut_7_12[10] , \wRegOut_7_12[9] , \wRegOut_7_12[8] , 
        \wRegOut_7_12[7] , \wRegOut_7_12[6] , \wRegOut_7_12[5] , 
        \wRegOut_7_12[4] , \wRegOut_7_12[3] , \wRegOut_7_12[2] , 
        \wRegOut_7_12[1] , \wRegOut_7_12[0] }), .L_Out({\wRegInTop_7_12[31] , 
        \wRegInTop_7_12[30] , \wRegInTop_7_12[29] , \wRegInTop_7_12[28] , 
        \wRegInTop_7_12[27] , \wRegInTop_7_12[26] , \wRegInTop_7_12[25] , 
        \wRegInTop_7_12[24] , \wRegInTop_7_12[23] , \wRegInTop_7_12[22] , 
        \wRegInTop_7_12[21] , \wRegInTop_7_12[20] , \wRegInTop_7_12[19] , 
        \wRegInTop_7_12[18] , \wRegInTop_7_12[17] , \wRegInTop_7_12[16] , 
        \wRegInTop_7_12[15] , \wRegInTop_7_12[14] , \wRegInTop_7_12[13] , 
        \wRegInTop_7_12[12] , \wRegInTop_7_12[11] , \wRegInTop_7_12[10] , 
        \wRegInTop_7_12[9] , \wRegInTop_7_12[8] , \wRegInTop_7_12[7] , 
        \wRegInTop_7_12[6] , \wRegInTop_7_12[5] , \wRegInTop_7_12[4] , 
        \wRegInTop_7_12[3] , \wRegInTop_7_12[2] , \wRegInTop_7_12[1] , 
        \wRegInTop_7_12[0] }), .R_WR(\wRegEnTop_7_13[0] ), .R_In({
        \wRegOut_7_13[31] , \wRegOut_7_13[30] , \wRegOut_7_13[29] , 
        \wRegOut_7_13[28] , \wRegOut_7_13[27] , \wRegOut_7_13[26] , 
        \wRegOut_7_13[25] , \wRegOut_7_13[24] , \wRegOut_7_13[23] , 
        \wRegOut_7_13[22] , \wRegOut_7_13[21] , \wRegOut_7_13[20] , 
        \wRegOut_7_13[19] , \wRegOut_7_13[18] , \wRegOut_7_13[17] , 
        \wRegOut_7_13[16] , \wRegOut_7_13[15] , \wRegOut_7_13[14] , 
        \wRegOut_7_13[13] , \wRegOut_7_13[12] , \wRegOut_7_13[11] , 
        \wRegOut_7_13[10] , \wRegOut_7_13[9] , \wRegOut_7_13[8] , 
        \wRegOut_7_13[7] , \wRegOut_7_13[6] , \wRegOut_7_13[5] , 
        \wRegOut_7_13[4] , \wRegOut_7_13[3] , \wRegOut_7_13[2] , 
        \wRegOut_7_13[1] , \wRegOut_7_13[0] }), .R_Out({\wRegInTop_7_13[31] , 
        \wRegInTop_7_13[30] , \wRegInTop_7_13[29] , \wRegInTop_7_13[28] , 
        \wRegInTop_7_13[27] , \wRegInTop_7_13[26] , \wRegInTop_7_13[25] , 
        \wRegInTop_7_13[24] , \wRegInTop_7_13[23] , \wRegInTop_7_13[22] , 
        \wRegInTop_7_13[21] , \wRegInTop_7_13[20] , \wRegInTop_7_13[19] , 
        \wRegInTop_7_13[18] , \wRegInTop_7_13[17] , \wRegInTop_7_13[16] , 
        \wRegInTop_7_13[15] , \wRegInTop_7_13[14] , \wRegInTop_7_13[13] , 
        \wRegInTop_7_13[12] , \wRegInTop_7_13[11] , \wRegInTop_7_13[10] , 
        \wRegInTop_7_13[9] , \wRegInTop_7_13[8] , \wRegInTop_7_13[7] , 
        \wRegInTop_7_13[6] , \wRegInTop_7_13[5] , \wRegInTop_7_13[4] , 
        \wRegInTop_7_13[3] , \wRegInTop_7_13[2] , \wRegInTop_7_13[1] , 
        \wRegInTop_7_13[0] }) );
    BHeap_Node_WIDTH32 BHN_6_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_57[0] ), .P_In({\wRegOut_6_57[31] , 
        \wRegOut_6_57[30] , \wRegOut_6_57[29] , \wRegOut_6_57[28] , 
        \wRegOut_6_57[27] , \wRegOut_6_57[26] , \wRegOut_6_57[25] , 
        \wRegOut_6_57[24] , \wRegOut_6_57[23] , \wRegOut_6_57[22] , 
        \wRegOut_6_57[21] , \wRegOut_6_57[20] , \wRegOut_6_57[19] , 
        \wRegOut_6_57[18] , \wRegOut_6_57[17] , \wRegOut_6_57[16] , 
        \wRegOut_6_57[15] , \wRegOut_6_57[14] , \wRegOut_6_57[13] , 
        \wRegOut_6_57[12] , \wRegOut_6_57[11] , \wRegOut_6_57[10] , 
        \wRegOut_6_57[9] , \wRegOut_6_57[8] , \wRegOut_6_57[7] , 
        \wRegOut_6_57[6] , \wRegOut_6_57[5] , \wRegOut_6_57[4] , 
        \wRegOut_6_57[3] , \wRegOut_6_57[2] , \wRegOut_6_57[1] , 
        \wRegOut_6_57[0] }), .P_Out({\wRegInBot_6_57[31] , 
        \wRegInBot_6_57[30] , \wRegInBot_6_57[29] , \wRegInBot_6_57[28] , 
        \wRegInBot_6_57[27] , \wRegInBot_6_57[26] , \wRegInBot_6_57[25] , 
        \wRegInBot_6_57[24] , \wRegInBot_6_57[23] , \wRegInBot_6_57[22] , 
        \wRegInBot_6_57[21] , \wRegInBot_6_57[20] , \wRegInBot_6_57[19] , 
        \wRegInBot_6_57[18] , \wRegInBot_6_57[17] , \wRegInBot_6_57[16] , 
        \wRegInBot_6_57[15] , \wRegInBot_6_57[14] , \wRegInBot_6_57[13] , 
        \wRegInBot_6_57[12] , \wRegInBot_6_57[11] , \wRegInBot_6_57[10] , 
        \wRegInBot_6_57[9] , \wRegInBot_6_57[8] , \wRegInBot_6_57[7] , 
        \wRegInBot_6_57[6] , \wRegInBot_6_57[5] , \wRegInBot_6_57[4] , 
        \wRegInBot_6_57[3] , \wRegInBot_6_57[2] , \wRegInBot_6_57[1] , 
        \wRegInBot_6_57[0] }), .L_WR(\wRegEnTop_7_114[0] ), .L_In({
        \wRegOut_7_114[31] , \wRegOut_7_114[30] , \wRegOut_7_114[29] , 
        \wRegOut_7_114[28] , \wRegOut_7_114[27] , \wRegOut_7_114[26] , 
        \wRegOut_7_114[25] , \wRegOut_7_114[24] , \wRegOut_7_114[23] , 
        \wRegOut_7_114[22] , \wRegOut_7_114[21] , \wRegOut_7_114[20] , 
        \wRegOut_7_114[19] , \wRegOut_7_114[18] , \wRegOut_7_114[17] , 
        \wRegOut_7_114[16] , \wRegOut_7_114[15] , \wRegOut_7_114[14] , 
        \wRegOut_7_114[13] , \wRegOut_7_114[12] , \wRegOut_7_114[11] , 
        \wRegOut_7_114[10] , \wRegOut_7_114[9] , \wRegOut_7_114[8] , 
        \wRegOut_7_114[7] , \wRegOut_7_114[6] , \wRegOut_7_114[5] , 
        \wRegOut_7_114[4] , \wRegOut_7_114[3] , \wRegOut_7_114[2] , 
        \wRegOut_7_114[1] , \wRegOut_7_114[0] }), .L_Out({
        \wRegInTop_7_114[31] , \wRegInTop_7_114[30] , \wRegInTop_7_114[29] , 
        \wRegInTop_7_114[28] , \wRegInTop_7_114[27] , \wRegInTop_7_114[26] , 
        \wRegInTop_7_114[25] , \wRegInTop_7_114[24] , \wRegInTop_7_114[23] , 
        \wRegInTop_7_114[22] , \wRegInTop_7_114[21] , \wRegInTop_7_114[20] , 
        \wRegInTop_7_114[19] , \wRegInTop_7_114[18] , \wRegInTop_7_114[17] , 
        \wRegInTop_7_114[16] , \wRegInTop_7_114[15] , \wRegInTop_7_114[14] , 
        \wRegInTop_7_114[13] , \wRegInTop_7_114[12] , \wRegInTop_7_114[11] , 
        \wRegInTop_7_114[10] , \wRegInTop_7_114[9] , \wRegInTop_7_114[8] , 
        \wRegInTop_7_114[7] , \wRegInTop_7_114[6] , \wRegInTop_7_114[5] , 
        \wRegInTop_7_114[4] , \wRegInTop_7_114[3] , \wRegInTop_7_114[2] , 
        \wRegInTop_7_114[1] , \wRegInTop_7_114[0] }), .R_WR(
        \wRegEnTop_7_115[0] ), .R_In({\wRegOut_7_115[31] , \wRegOut_7_115[30] , 
        \wRegOut_7_115[29] , \wRegOut_7_115[28] , \wRegOut_7_115[27] , 
        \wRegOut_7_115[26] , \wRegOut_7_115[25] , \wRegOut_7_115[24] , 
        \wRegOut_7_115[23] , \wRegOut_7_115[22] , \wRegOut_7_115[21] , 
        \wRegOut_7_115[20] , \wRegOut_7_115[19] , \wRegOut_7_115[18] , 
        \wRegOut_7_115[17] , \wRegOut_7_115[16] , \wRegOut_7_115[15] , 
        \wRegOut_7_115[14] , \wRegOut_7_115[13] , \wRegOut_7_115[12] , 
        \wRegOut_7_115[11] , \wRegOut_7_115[10] , \wRegOut_7_115[9] , 
        \wRegOut_7_115[8] , \wRegOut_7_115[7] , \wRegOut_7_115[6] , 
        \wRegOut_7_115[5] , \wRegOut_7_115[4] , \wRegOut_7_115[3] , 
        \wRegOut_7_115[2] , \wRegOut_7_115[1] , \wRegOut_7_115[0] }), .R_Out({
        \wRegInTop_7_115[31] , \wRegInTop_7_115[30] , \wRegInTop_7_115[29] , 
        \wRegInTop_7_115[28] , \wRegInTop_7_115[27] , \wRegInTop_7_115[26] , 
        \wRegInTop_7_115[25] , \wRegInTop_7_115[24] , \wRegInTop_7_115[23] , 
        \wRegInTop_7_115[22] , \wRegInTop_7_115[21] , \wRegInTop_7_115[20] , 
        \wRegInTop_7_115[19] , \wRegInTop_7_115[18] , \wRegInTop_7_115[17] , 
        \wRegInTop_7_115[16] , \wRegInTop_7_115[15] , \wRegInTop_7_115[14] , 
        \wRegInTop_7_115[13] , \wRegInTop_7_115[12] , \wRegInTop_7_115[11] , 
        \wRegInTop_7_115[10] , \wRegInTop_7_115[9] , \wRegInTop_7_115[8] , 
        \wRegInTop_7_115[7] , \wRegInTop_7_115[6] , \wRegInTop_7_115[5] , 
        \wRegInTop_7_115[4] , \wRegInTop_7_115[3] , \wRegInTop_7_115[2] , 
        \wRegInTop_7_115[1] , \wRegInTop_7_115[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink132[31] , \ScanLink132[30] , \ScanLink132[29] , 
        \ScanLink132[28] , \ScanLink132[27] , \ScanLink132[26] , 
        \ScanLink132[25] , \ScanLink132[24] , \ScanLink132[23] , 
        \ScanLink132[22] , \ScanLink132[21] , \ScanLink132[20] , 
        \ScanLink132[19] , \ScanLink132[18] , \ScanLink132[17] , 
        \ScanLink132[16] , \ScanLink132[15] , \ScanLink132[14] , 
        \ScanLink132[13] , \ScanLink132[12] , \ScanLink132[11] , 
        \ScanLink132[10] , \ScanLink132[9] , \ScanLink132[8] , 
        \ScanLink132[7] , \ScanLink132[6] , \ScanLink132[5] , \ScanLink132[4] , 
        \ScanLink132[3] , \ScanLink132[2] , \ScanLink132[1] , \ScanLink132[0] 
        }), .ScanOut({\ScanLink131[31] , \ScanLink131[30] , \ScanLink131[29] , 
        \ScanLink131[28] , \ScanLink131[27] , \ScanLink131[26] , 
        \ScanLink131[25] , \ScanLink131[24] , \ScanLink131[23] , 
        \ScanLink131[22] , \ScanLink131[21] , \ScanLink131[20] , 
        \ScanLink131[19] , \ScanLink131[18] , \ScanLink131[17] , 
        \ScanLink131[16] , \ScanLink131[15] , \ScanLink131[14] , 
        \ScanLink131[13] , \ScanLink131[12] , \ScanLink131[11] , 
        \ScanLink131[10] , \ScanLink131[9] , \ScanLink131[8] , 
        \ScanLink131[7] , \ScanLink131[6] , \ScanLink131[5] , \ScanLink131[4] , 
        \ScanLink131[3] , \ScanLink131[2] , \ScanLink131[1] , \ScanLink131[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_4[31] , 
        \wRegOut_7_4[30] , \wRegOut_7_4[29] , \wRegOut_7_4[28] , 
        \wRegOut_7_4[27] , \wRegOut_7_4[26] , \wRegOut_7_4[25] , 
        \wRegOut_7_4[24] , \wRegOut_7_4[23] , \wRegOut_7_4[22] , 
        \wRegOut_7_4[21] , \wRegOut_7_4[20] , \wRegOut_7_4[19] , 
        \wRegOut_7_4[18] , \wRegOut_7_4[17] , \wRegOut_7_4[16] , 
        \wRegOut_7_4[15] , \wRegOut_7_4[14] , \wRegOut_7_4[13] , 
        \wRegOut_7_4[12] , \wRegOut_7_4[11] , \wRegOut_7_4[10] , 
        \wRegOut_7_4[9] , \wRegOut_7_4[8] , \wRegOut_7_4[7] , \wRegOut_7_4[6] , 
        \wRegOut_7_4[5] , \wRegOut_7_4[4] , \wRegOut_7_4[3] , \wRegOut_7_4[2] , 
        \wRegOut_7_4[1] , \wRegOut_7_4[0] }), .Enable1(\wRegEnTop_7_4[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_4[31] , \wRegInTop_7_4[30] , 
        \wRegInTop_7_4[29] , \wRegInTop_7_4[28] , \wRegInTop_7_4[27] , 
        \wRegInTop_7_4[26] , \wRegInTop_7_4[25] , \wRegInTop_7_4[24] , 
        \wRegInTop_7_4[23] , \wRegInTop_7_4[22] , \wRegInTop_7_4[21] , 
        \wRegInTop_7_4[20] , \wRegInTop_7_4[19] , \wRegInTop_7_4[18] , 
        \wRegInTop_7_4[17] , \wRegInTop_7_4[16] , \wRegInTop_7_4[15] , 
        \wRegInTop_7_4[14] , \wRegInTop_7_4[13] , \wRegInTop_7_4[12] , 
        \wRegInTop_7_4[11] , \wRegInTop_7_4[10] , \wRegInTop_7_4[9] , 
        \wRegInTop_7_4[8] , \wRegInTop_7_4[7] , \wRegInTop_7_4[6] , 
        \wRegInTop_7_4[5] , \wRegInTop_7_4[4] , \wRegInTop_7_4[3] , 
        \wRegInTop_7_4[2] , \wRegInTop_7_4[1] , \wRegInTop_7_4[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_42 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink170[31] , \ScanLink170[30] , \ScanLink170[29] , 
        \ScanLink170[28] , \ScanLink170[27] , \ScanLink170[26] , 
        \ScanLink170[25] , \ScanLink170[24] , \ScanLink170[23] , 
        \ScanLink170[22] , \ScanLink170[21] , \ScanLink170[20] , 
        \ScanLink170[19] , \ScanLink170[18] , \ScanLink170[17] , 
        \ScanLink170[16] , \ScanLink170[15] , \ScanLink170[14] , 
        \ScanLink170[13] , \ScanLink170[12] , \ScanLink170[11] , 
        \ScanLink170[10] , \ScanLink170[9] , \ScanLink170[8] , 
        \ScanLink170[7] , \ScanLink170[6] , \ScanLink170[5] , \ScanLink170[4] , 
        \ScanLink170[3] , \ScanLink170[2] , \ScanLink170[1] , \ScanLink170[0] 
        }), .ScanOut({\ScanLink169[31] , \ScanLink169[30] , \ScanLink169[29] , 
        \ScanLink169[28] , \ScanLink169[27] , \ScanLink169[26] , 
        \ScanLink169[25] , \ScanLink169[24] , \ScanLink169[23] , 
        \ScanLink169[22] , \ScanLink169[21] , \ScanLink169[20] , 
        \ScanLink169[19] , \ScanLink169[18] , \ScanLink169[17] , 
        \ScanLink169[16] , \ScanLink169[15] , \ScanLink169[14] , 
        \ScanLink169[13] , \ScanLink169[12] , \ScanLink169[11] , 
        \ScanLink169[10] , \ScanLink169[9] , \ScanLink169[8] , 
        \ScanLink169[7] , \ScanLink169[6] , \ScanLink169[5] , \ScanLink169[4] , 
        \ScanLink169[3] , \ScanLink169[2] , \ScanLink169[1] , \ScanLink169[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_42[31] , 
        \wRegOut_7_42[30] , \wRegOut_7_42[29] , \wRegOut_7_42[28] , 
        \wRegOut_7_42[27] , \wRegOut_7_42[26] , \wRegOut_7_42[25] , 
        \wRegOut_7_42[24] , \wRegOut_7_42[23] , \wRegOut_7_42[22] , 
        \wRegOut_7_42[21] , \wRegOut_7_42[20] , \wRegOut_7_42[19] , 
        \wRegOut_7_42[18] , \wRegOut_7_42[17] , \wRegOut_7_42[16] , 
        \wRegOut_7_42[15] , \wRegOut_7_42[14] , \wRegOut_7_42[13] , 
        \wRegOut_7_42[12] , \wRegOut_7_42[11] , \wRegOut_7_42[10] , 
        \wRegOut_7_42[9] , \wRegOut_7_42[8] , \wRegOut_7_42[7] , 
        \wRegOut_7_42[6] , \wRegOut_7_42[5] , \wRegOut_7_42[4] , 
        \wRegOut_7_42[3] , \wRegOut_7_42[2] , \wRegOut_7_42[1] , 
        \wRegOut_7_42[0] }), .Enable1(\wRegEnTop_7_42[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_42[31] , \wRegInTop_7_42[30] , \wRegInTop_7_42[29] , 
        \wRegInTop_7_42[28] , \wRegInTop_7_42[27] , \wRegInTop_7_42[26] , 
        \wRegInTop_7_42[25] , \wRegInTop_7_42[24] , \wRegInTop_7_42[23] , 
        \wRegInTop_7_42[22] , \wRegInTop_7_42[21] , \wRegInTop_7_42[20] , 
        \wRegInTop_7_42[19] , \wRegInTop_7_42[18] , \wRegInTop_7_42[17] , 
        \wRegInTop_7_42[16] , \wRegInTop_7_42[15] , \wRegInTop_7_42[14] , 
        \wRegInTop_7_42[13] , \wRegInTop_7_42[12] , \wRegInTop_7_42[11] , 
        \wRegInTop_7_42[10] , \wRegInTop_7_42[9] , \wRegInTop_7_42[8] , 
        \wRegInTop_7_42[7] , \wRegInTop_7_42[6] , \wRegInTop_7_42[5] , 
        \wRegInTop_7_42[4] , \wRegInTop_7_42[3] , \wRegInTop_7_42[2] , 
        \wRegInTop_7_42[1] , \wRegInTop_7_42[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_2_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink7[31] , \ScanLink7[30] , \ScanLink7[29] , 
        \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , \ScanLink7[25] , 
        \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , \ScanLink7[21] , 
        \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , \ScanLink7[17] , 
        \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , \ScanLink7[13] , 
        \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , \ScanLink7[9] , 
        \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , \ScanLink7[5] , 
        \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , \ScanLink7[1] , 
        \ScanLink7[0] }), .ScanOut({\ScanLink6[31] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , 
        \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , 
        \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , 
        \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , 
        \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , 
        \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_2_3[31] , \wRegOut_2_3[30] , \wRegOut_2_3[29] , 
        \wRegOut_2_3[28] , \wRegOut_2_3[27] , \wRegOut_2_3[26] , 
        \wRegOut_2_3[25] , \wRegOut_2_3[24] , \wRegOut_2_3[23] , 
        \wRegOut_2_3[22] , \wRegOut_2_3[21] , \wRegOut_2_3[20] , 
        \wRegOut_2_3[19] , \wRegOut_2_3[18] , \wRegOut_2_3[17] , 
        \wRegOut_2_3[16] , \wRegOut_2_3[15] , \wRegOut_2_3[14] , 
        \wRegOut_2_3[13] , \wRegOut_2_3[12] , \wRegOut_2_3[11] , 
        \wRegOut_2_3[10] , \wRegOut_2_3[9] , \wRegOut_2_3[8] , 
        \wRegOut_2_3[7] , \wRegOut_2_3[6] , \wRegOut_2_3[5] , \wRegOut_2_3[4] , 
        \wRegOut_2_3[3] , \wRegOut_2_3[2] , \wRegOut_2_3[1] , \wRegOut_2_3[0] 
        }), .Enable1(\wRegEnTop_2_3[0] ), .Enable2(\wRegEnBot_2_3[0] ), .In1({
        \wRegInTop_2_3[31] , \wRegInTop_2_3[30] , \wRegInTop_2_3[29] , 
        \wRegInTop_2_3[28] , \wRegInTop_2_3[27] , \wRegInTop_2_3[26] , 
        \wRegInTop_2_3[25] , \wRegInTop_2_3[24] , \wRegInTop_2_3[23] , 
        \wRegInTop_2_3[22] , \wRegInTop_2_3[21] , \wRegInTop_2_3[20] , 
        \wRegInTop_2_3[19] , \wRegInTop_2_3[18] , \wRegInTop_2_3[17] , 
        \wRegInTop_2_3[16] , \wRegInTop_2_3[15] , \wRegInTop_2_3[14] , 
        \wRegInTop_2_3[13] , \wRegInTop_2_3[12] , \wRegInTop_2_3[11] , 
        \wRegInTop_2_3[10] , \wRegInTop_2_3[9] , \wRegInTop_2_3[8] , 
        \wRegInTop_2_3[7] , \wRegInTop_2_3[6] , \wRegInTop_2_3[5] , 
        \wRegInTop_2_3[4] , \wRegInTop_2_3[3] , \wRegInTop_2_3[2] , 
        \wRegInTop_2_3[1] , \wRegInTop_2_3[0] }), .In2({\wRegInBot_2_3[31] , 
        \wRegInBot_2_3[30] , \wRegInBot_2_3[29] , \wRegInBot_2_3[28] , 
        \wRegInBot_2_3[27] , \wRegInBot_2_3[26] , \wRegInBot_2_3[25] , 
        \wRegInBot_2_3[24] , \wRegInBot_2_3[23] , \wRegInBot_2_3[22] , 
        \wRegInBot_2_3[21] , \wRegInBot_2_3[20] , \wRegInBot_2_3[19] , 
        \wRegInBot_2_3[18] , \wRegInBot_2_3[17] , \wRegInBot_2_3[16] , 
        \wRegInBot_2_3[15] , \wRegInBot_2_3[14] , \wRegInBot_2_3[13] , 
        \wRegInBot_2_3[12] , \wRegInBot_2_3[11] , \wRegInBot_2_3[10] , 
        \wRegInBot_2_3[9] , \wRegInBot_2_3[8] , \wRegInBot_2_3[7] , 
        \wRegInBot_2_3[6] , \wRegInBot_2_3[5] , \wRegInBot_2_3[4] , 
        \wRegInBot_2_3[3] , \wRegInBot_2_3[2] , \wRegInBot_2_3[1] , 
        \wRegInBot_2_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink16[31] , \ScanLink16[30] , \ScanLink16[29] , 
        \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , \ScanLink16[25] , 
        \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , \ScanLink16[21] , 
        \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , \ScanLink16[17] , 
        \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , \ScanLink16[13] , 
        \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , \ScanLink16[9] , 
        \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , \ScanLink16[5] , 
        \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , \ScanLink16[1] , 
        \ScanLink16[0] }), .ScanOut({\ScanLink15[31] , \ScanLink15[30] , 
        \ScanLink15[29] , \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , 
        \ScanLink15[25] , \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , 
        \ScanLink15[21] , \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , 
        \ScanLink15[17] , \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , 
        \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , 
        \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , 
        \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , 
        \ScanLink15[1] , \ScanLink15[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_0[31] , \wRegOut_4_0[30] , \wRegOut_4_0[29] , 
        \wRegOut_4_0[28] , \wRegOut_4_0[27] , \wRegOut_4_0[26] , 
        \wRegOut_4_0[25] , \wRegOut_4_0[24] , \wRegOut_4_0[23] , 
        \wRegOut_4_0[22] , \wRegOut_4_0[21] , \wRegOut_4_0[20] , 
        \wRegOut_4_0[19] , \wRegOut_4_0[18] , \wRegOut_4_0[17] , 
        \wRegOut_4_0[16] , \wRegOut_4_0[15] , \wRegOut_4_0[14] , 
        \wRegOut_4_0[13] , \wRegOut_4_0[12] , \wRegOut_4_0[11] , 
        \wRegOut_4_0[10] , \wRegOut_4_0[9] , \wRegOut_4_0[8] , 
        \wRegOut_4_0[7] , \wRegOut_4_0[6] , \wRegOut_4_0[5] , \wRegOut_4_0[4] , 
        \wRegOut_4_0[3] , \wRegOut_4_0[2] , \wRegOut_4_0[1] , \wRegOut_4_0[0] 
        }), .Enable1(\wRegEnTop_4_0[0] ), .Enable2(\wRegEnBot_4_0[0] ), .In1({
        \wRegInTop_4_0[31] , \wRegInTop_4_0[30] , \wRegInTop_4_0[29] , 
        \wRegInTop_4_0[28] , \wRegInTop_4_0[27] , \wRegInTop_4_0[26] , 
        \wRegInTop_4_0[25] , \wRegInTop_4_0[24] , \wRegInTop_4_0[23] , 
        \wRegInTop_4_0[22] , \wRegInTop_4_0[21] , \wRegInTop_4_0[20] , 
        \wRegInTop_4_0[19] , \wRegInTop_4_0[18] , \wRegInTop_4_0[17] , 
        \wRegInTop_4_0[16] , \wRegInTop_4_0[15] , \wRegInTop_4_0[14] , 
        \wRegInTop_4_0[13] , \wRegInTop_4_0[12] , \wRegInTop_4_0[11] , 
        \wRegInTop_4_0[10] , \wRegInTop_4_0[9] , \wRegInTop_4_0[8] , 
        \wRegInTop_4_0[7] , \wRegInTop_4_0[6] , \wRegInTop_4_0[5] , 
        \wRegInTop_4_0[4] , \wRegInTop_4_0[3] , \wRegInTop_4_0[2] , 
        \wRegInTop_4_0[1] , \wRegInTop_4_0[0] }), .In2({\wRegInBot_4_0[31] , 
        \wRegInBot_4_0[30] , \wRegInBot_4_0[29] , \wRegInBot_4_0[28] , 
        \wRegInBot_4_0[27] , \wRegInBot_4_0[26] , \wRegInBot_4_0[25] , 
        \wRegInBot_4_0[24] , \wRegInBot_4_0[23] , \wRegInBot_4_0[22] , 
        \wRegInBot_4_0[21] , \wRegInBot_4_0[20] , \wRegInBot_4_0[19] , 
        \wRegInBot_4_0[18] , \wRegInBot_4_0[17] , \wRegInBot_4_0[16] , 
        \wRegInBot_4_0[15] , \wRegInBot_4_0[14] , \wRegInBot_4_0[13] , 
        \wRegInBot_4_0[12] , \wRegInBot_4_0[11] , \wRegInBot_4_0[10] , 
        \wRegInBot_4_0[9] , \wRegInBot_4_0[8] , \wRegInBot_4_0[7] , 
        \wRegInBot_4_0[6] , \wRegInBot_4_0[5] , \wRegInBot_4_0[4] , 
        \wRegInBot_4_0[3] , \wRegInBot_4_0[2] , \wRegInBot_4_0[1] , 
        \wRegInBot_4_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink30[31] , \ScanLink30[30] , \ScanLink30[29] , 
        \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , \ScanLink30[25] , 
        \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , \ScanLink30[21] , 
        \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , \ScanLink30[17] , 
        \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , \ScanLink30[13] , 
        \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , \ScanLink30[9] , 
        \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , \ScanLink30[5] , 
        \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , \ScanLink30[1] , 
        \ScanLink30[0] }), .ScanOut({\ScanLink29[31] , \ScanLink29[30] , 
        \ScanLink29[29] , \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , 
        \ScanLink29[25] , \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , 
        \ScanLink29[21] , \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , 
        \ScanLink29[17] , \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , 
        \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , 
        \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , 
        \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , 
        \ScanLink29[1] , \ScanLink29[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_14[31] , \wRegOut_4_14[30] , 
        \wRegOut_4_14[29] , \wRegOut_4_14[28] , \wRegOut_4_14[27] , 
        \wRegOut_4_14[26] , \wRegOut_4_14[25] , \wRegOut_4_14[24] , 
        \wRegOut_4_14[23] , \wRegOut_4_14[22] , \wRegOut_4_14[21] , 
        \wRegOut_4_14[20] , \wRegOut_4_14[19] , \wRegOut_4_14[18] , 
        \wRegOut_4_14[17] , \wRegOut_4_14[16] , \wRegOut_4_14[15] , 
        \wRegOut_4_14[14] , \wRegOut_4_14[13] , \wRegOut_4_14[12] , 
        \wRegOut_4_14[11] , \wRegOut_4_14[10] , \wRegOut_4_14[9] , 
        \wRegOut_4_14[8] , \wRegOut_4_14[7] , \wRegOut_4_14[6] , 
        \wRegOut_4_14[5] , \wRegOut_4_14[4] , \wRegOut_4_14[3] , 
        \wRegOut_4_14[2] , \wRegOut_4_14[1] , \wRegOut_4_14[0] }), .Enable1(
        \wRegEnTop_4_14[0] ), .Enable2(\wRegEnBot_4_14[0] ), .In1({
        \wRegInTop_4_14[31] , \wRegInTop_4_14[30] , \wRegInTop_4_14[29] , 
        \wRegInTop_4_14[28] , \wRegInTop_4_14[27] , \wRegInTop_4_14[26] , 
        \wRegInTop_4_14[25] , \wRegInTop_4_14[24] , \wRegInTop_4_14[23] , 
        \wRegInTop_4_14[22] , \wRegInTop_4_14[21] , \wRegInTop_4_14[20] , 
        \wRegInTop_4_14[19] , \wRegInTop_4_14[18] , \wRegInTop_4_14[17] , 
        \wRegInTop_4_14[16] , \wRegInTop_4_14[15] , \wRegInTop_4_14[14] , 
        \wRegInTop_4_14[13] , \wRegInTop_4_14[12] , \wRegInTop_4_14[11] , 
        \wRegInTop_4_14[10] , \wRegInTop_4_14[9] , \wRegInTop_4_14[8] , 
        \wRegInTop_4_14[7] , \wRegInTop_4_14[6] , \wRegInTop_4_14[5] , 
        \wRegInTop_4_14[4] , \wRegInTop_4_14[3] , \wRegInTop_4_14[2] , 
        \wRegInTop_4_14[1] , \wRegInTop_4_14[0] }), .In2({\wRegInBot_4_14[31] , 
        \wRegInBot_4_14[30] , \wRegInBot_4_14[29] , \wRegInBot_4_14[28] , 
        \wRegInBot_4_14[27] , \wRegInBot_4_14[26] , \wRegInBot_4_14[25] , 
        \wRegInBot_4_14[24] , \wRegInBot_4_14[23] , \wRegInBot_4_14[22] , 
        \wRegInBot_4_14[21] , \wRegInBot_4_14[20] , \wRegInBot_4_14[19] , 
        \wRegInBot_4_14[18] , \wRegInBot_4_14[17] , \wRegInBot_4_14[16] , 
        \wRegInBot_4_14[15] , \wRegInBot_4_14[14] , \wRegInBot_4_14[13] , 
        \wRegInBot_4_14[12] , \wRegInBot_4_14[11] , \wRegInBot_4_14[10] , 
        \wRegInBot_4_14[9] , \wRegInBot_4_14[8] , \wRegInBot_4_14[7] , 
        \wRegInBot_4_14[6] , \wRegInBot_4_14[5] , \wRegInBot_4_14[4] , 
        \wRegInBot_4_14[3] , \wRegInBot_4_14[2] , \wRegInBot_4_14[1] , 
        \wRegInBot_4_14[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink32[31] , \ScanLink32[30] , \ScanLink32[29] , 
        \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , \ScanLink32[25] , 
        \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , \ScanLink32[21] , 
        \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , \ScanLink32[17] , 
        \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , \ScanLink32[13] , 
        \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , \ScanLink32[9] , 
        \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , \ScanLink32[5] , 
        \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , \ScanLink32[1] , 
        \ScanLink32[0] }), .ScanOut({\ScanLink31[31] , \ScanLink31[30] , 
        \ScanLink31[29] , \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , 
        \ScanLink31[25] , \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , 
        \ScanLink31[21] , \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , 
        \ScanLink31[17] , \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , 
        \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , 
        \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , 
        \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , 
        \ScanLink31[1] , \ScanLink31[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_0[31] , \wRegOut_5_0[30] , \wRegOut_5_0[29] , 
        \wRegOut_5_0[28] , \wRegOut_5_0[27] , \wRegOut_5_0[26] , 
        \wRegOut_5_0[25] , \wRegOut_5_0[24] , \wRegOut_5_0[23] , 
        \wRegOut_5_0[22] , \wRegOut_5_0[21] , \wRegOut_5_0[20] , 
        \wRegOut_5_0[19] , \wRegOut_5_0[18] , \wRegOut_5_0[17] , 
        \wRegOut_5_0[16] , \wRegOut_5_0[15] , \wRegOut_5_0[14] , 
        \wRegOut_5_0[13] , \wRegOut_5_0[12] , \wRegOut_5_0[11] , 
        \wRegOut_5_0[10] , \wRegOut_5_0[9] , \wRegOut_5_0[8] , 
        \wRegOut_5_0[7] , \wRegOut_5_0[6] , \wRegOut_5_0[5] , \wRegOut_5_0[4] , 
        \wRegOut_5_0[3] , \wRegOut_5_0[2] , \wRegOut_5_0[1] , \wRegOut_5_0[0] 
        }), .Enable1(\wRegEnTop_5_0[0] ), .Enable2(\wRegEnBot_5_0[0] ), .In1({
        \wRegInTop_5_0[31] , \wRegInTop_5_0[30] , \wRegInTop_5_0[29] , 
        \wRegInTop_5_0[28] , \wRegInTop_5_0[27] , \wRegInTop_5_0[26] , 
        \wRegInTop_5_0[25] , \wRegInTop_5_0[24] , \wRegInTop_5_0[23] , 
        \wRegInTop_5_0[22] , \wRegInTop_5_0[21] , \wRegInTop_5_0[20] , 
        \wRegInTop_5_0[19] , \wRegInTop_5_0[18] , \wRegInTop_5_0[17] , 
        \wRegInTop_5_0[16] , \wRegInTop_5_0[15] , \wRegInTop_5_0[14] , 
        \wRegInTop_5_0[13] , \wRegInTop_5_0[12] , \wRegInTop_5_0[11] , 
        \wRegInTop_5_0[10] , \wRegInTop_5_0[9] , \wRegInTop_5_0[8] , 
        \wRegInTop_5_0[7] , \wRegInTop_5_0[6] , \wRegInTop_5_0[5] , 
        \wRegInTop_5_0[4] , \wRegInTop_5_0[3] , \wRegInTop_5_0[2] , 
        \wRegInTop_5_0[1] , \wRegInTop_5_0[0] }), .In2({\wRegInBot_5_0[31] , 
        \wRegInBot_5_0[30] , \wRegInBot_5_0[29] , \wRegInBot_5_0[28] , 
        \wRegInBot_5_0[27] , \wRegInBot_5_0[26] , \wRegInBot_5_0[25] , 
        \wRegInBot_5_0[24] , \wRegInBot_5_0[23] , \wRegInBot_5_0[22] , 
        \wRegInBot_5_0[21] , \wRegInBot_5_0[20] , \wRegInBot_5_0[19] , 
        \wRegInBot_5_0[18] , \wRegInBot_5_0[17] , \wRegInBot_5_0[16] , 
        \wRegInBot_5_0[15] , \wRegInBot_5_0[14] , \wRegInBot_5_0[13] , 
        \wRegInBot_5_0[12] , \wRegInBot_5_0[11] , \wRegInBot_5_0[10] , 
        \wRegInBot_5_0[9] , \wRegInBot_5_0[8] , \wRegInBot_5_0[7] , 
        \wRegInBot_5_0[6] , \wRegInBot_5_0[5] , \wRegInBot_5_0[4] , 
        \wRegInBot_5_0[3] , \wRegInBot_5_0[2] , \wRegInBot_5_0[1] , 
        \wRegInBot_5_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink40[31] , \ScanLink40[30] , \ScanLink40[29] , 
        \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , \ScanLink40[25] , 
        \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , \ScanLink40[21] , 
        \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , \ScanLink40[17] , 
        \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , \ScanLink40[13] , 
        \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , \ScanLink40[9] , 
        \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , \ScanLink40[5] , 
        \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , \ScanLink40[1] , 
        \ScanLink40[0] }), .ScanOut({\ScanLink39[31] , \ScanLink39[30] , 
        \ScanLink39[29] , \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , 
        \ScanLink39[25] , \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , 
        \ScanLink39[21] , \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , 
        \ScanLink39[17] , \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , 
        \ScanLink39[13] , \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , 
        \ScanLink39[9] , \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , 
        \ScanLink39[5] , \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , 
        \ScanLink39[1] , \ScanLink39[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_8[31] , \wRegOut_5_8[30] , \wRegOut_5_8[29] , 
        \wRegOut_5_8[28] , \wRegOut_5_8[27] , \wRegOut_5_8[26] , 
        \wRegOut_5_8[25] , \wRegOut_5_8[24] , \wRegOut_5_8[23] , 
        \wRegOut_5_8[22] , \wRegOut_5_8[21] , \wRegOut_5_8[20] , 
        \wRegOut_5_8[19] , \wRegOut_5_8[18] , \wRegOut_5_8[17] , 
        \wRegOut_5_8[16] , \wRegOut_5_8[15] , \wRegOut_5_8[14] , 
        \wRegOut_5_8[13] , \wRegOut_5_8[12] , \wRegOut_5_8[11] , 
        \wRegOut_5_8[10] , \wRegOut_5_8[9] , \wRegOut_5_8[8] , 
        \wRegOut_5_8[7] , \wRegOut_5_8[6] , \wRegOut_5_8[5] , \wRegOut_5_8[4] , 
        \wRegOut_5_8[3] , \wRegOut_5_8[2] , \wRegOut_5_8[1] , \wRegOut_5_8[0] 
        }), .Enable1(\wRegEnTop_5_8[0] ), .Enable2(\wRegEnBot_5_8[0] ), .In1({
        \wRegInTop_5_8[31] , \wRegInTop_5_8[30] , \wRegInTop_5_8[29] , 
        \wRegInTop_5_8[28] , \wRegInTop_5_8[27] , \wRegInTop_5_8[26] , 
        \wRegInTop_5_8[25] , \wRegInTop_5_8[24] , \wRegInTop_5_8[23] , 
        \wRegInTop_5_8[22] , \wRegInTop_5_8[21] , \wRegInTop_5_8[20] , 
        \wRegInTop_5_8[19] , \wRegInTop_5_8[18] , \wRegInTop_5_8[17] , 
        \wRegInTop_5_8[16] , \wRegInTop_5_8[15] , \wRegInTop_5_8[14] , 
        \wRegInTop_5_8[13] , \wRegInTop_5_8[12] , \wRegInTop_5_8[11] , 
        \wRegInTop_5_8[10] , \wRegInTop_5_8[9] , \wRegInTop_5_8[8] , 
        \wRegInTop_5_8[7] , \wRegInTop_5_8[6] , \wRegInTop_5_8[5] , 
        \wRegInTop_5_8[4] , \wRegInTop_5_8[3] , \wRegInTop_5_8[2] , 
        \wRegInTop_5_8[1] , \wRegInTop_5_8[0] }), .In2({\wRegInBot_5_8[31] , 
        \wRegInBot_5_8[30] , \wRegInBot_5_8[29] , \wRegInBot_5_8[28] , 
        \wRegInBot_5_8[27] , \wRegInBot_5_8[26] , \wRegInBot_5_8[25] , 
        \wRegInBot_5_8[24] , \wRegInBot_5_8[23] , \wRegInBot_5_8[22] , 
        \wRegInBot_5_8[21] , \wRegInBot_5_8[20] , \wRegInBot_5_8[19] , 
        \wRegInBot_5_8[18] , \wRegInBot_5_8[17] , \wRegInBot_5_8[16] , 
        \wRegInBot_5_8[15] , \wRegInBot_5_8[14] , \wRegInBot_5_8[13] , 
        \wRegInBot_5_8[12] , \wRegInBot_5_8[11] , \wRegInBot_5_8[10] , 
        \wRegInBot_5_8[9] , \wRegInBot_5_8[8] , \wRegInBot_5_8[7] , 
        \wRegInBot_5_8[6] , \wRegInBot_5_8[5] , \wRegInBot_5_8[4] , 
        \wRegInBot_5_8[3] , \wRegInBot_5_8[2] , \wRegInBot_5_8[1] , 
        \wRegInBot_5_8[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_21 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink53[31] , \ScanLink53[30] , \ScanLink53[29] , 
        \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , \ScanLink53[25] , 
        \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , \ScanLink53[21] , 
        \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , \ScanLink53[17] , 
        \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , \ScanLink53[13] , 
        \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , \ScanLink53[9] , 
        \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , \ScanLink53[5] , 
        \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , \ScanLink53[1] , 
        \ScanLink53[0] }), .ScanOut({\ScanLink52[31] , \ScanLink52[30] , 
        \ScanLink52[29] , \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , 
        \ScanLink52[25] , \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , 
        \ScanLink52[21] , \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , 
        \ScanLink52[17] , \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , 
        \ScanLink52[13] , \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , 
        \ScanLink52[9] , \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , 
        \ScanLink52[5] , \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , 
        \ScanLink52[1] , \ScanLink52[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_21[31] , \wRegOut_5_21[30] , 
        \wRegOut_5_21[29] , \wRegOut_5_21[28] , \wRegOut_5_21[27] , 
        \wRegOut_5_21[26] , \wRegOut_5_21[25] , \wRegOut_5_21[24] , 
        \wRegOut_5_21[23] , \wRegOut_5_21[22] , \wRegOut_5_21[21] , 
        \wRegOut_5_21[20] , \wRegOut_5_21[19] , \wRegOut_5_21[18] , 
        \wRegOut_5_21[17] , \wRegOut_5_21[16] , \wRegOut_5_21[15] , 
        \wRegOut_5_21[14] , \wRegOut_5_21[13] , \wRegOut_5_21[12] , 
        \wRegOut_5_21[11] , \wRegOut_5_21[10] , \wRegOut_5_21[9] , 
        \wRegOut_5_21[8] , \wRegOut_5_21[7] , \wRegOut_5_21[6] , 
        \wRegOut_5_21[5] , \wRegOut_5_21[4] , \wRegOut_5_21[3] , 
        \wRegOut_5_21[2] , \wRegOut_5_21[1] , \wRegOut_5_21[0] }), .Enable1(
        \wRegEnTop_5_21[0] ), .Enable2(\wRegEnBot_5_21[0] ), .In1({
        \wRegInTop_5_21[31] , \wRegInTop_5_21[30] , \wRegInTop_5_21[29] , 
        \wRegInTop_5_21[28] , \wRegInTop_5_21[27] , \wRegInTop_5_21[26] , 
        \wRegInTop_5_21[25] , \wRegInTop_5_21[24] , \wRegInTop_5_21[23] , 
        \wRegInTop_5_21[22] , \wRegInTop_5_21[21] , \wRegInTop_5_21[20] , 
        \wRegInTop_5_21[19] , \wRegInTop_5_21[18] , \wRegInTop_5_21[17] , 
        \wRegInTop_5_21[16] , \wRegInTop_5_21[15] , \wRegInTop_5_21[14] , 
        \wRegInTop_5_21[13] , \wRegInTop_5_21[12] , \wRegInTop_5_21[11] , 
        \wRegInTop_5_21[10] , \wRegInTop_5_21[9] , \wRegInTop_5_21[8] , 
        \wRegInTop_5_21[7] , \wRegInTop_5_21[6] , \wRegInTop_5_21[5] , 
        \wRegInTop_5_21[4] , \wRegInTop_5_21[3] , \wRegInTop_5_21[2] , 
        \wRegInTop_5_21[1] , \wRegInTop_5_21[0] }), .In2({\wRegInBot_5_21[31] , 
        \wRegInBot_5_21[30] , \wRegInBot_5_21[29] , \wRegInBot_5_21[28] , 
        \wRegInBot_5_21[27] , \wRegInBot_5_21[26] , \wRegInBot_5_21[25] , 
        \wRegInBot_5_21[24] , \wRegInBot_5_21[23] , \wRegInBot_5_21[22] , 
        \wRegInBot_5_21[21] , \wRegInBot_5_21[20] , \wRegInBot_5_21[19] , 
        \wRegInBot_5_21[18] , \wRegInBot_5_21[17] , \wRegInBot_5_21[16] , 
        \wRegInBot_5_21[15] , \wRegInBot_5_21[14] , \wRegInBot_5_21[13] , 
        \wRegInBot_5_21[12] , \wRegInBot_5_21[11] , \wRegInBot_5_21[10] , 
        \wRegInBot_5_21[9] , \wRegInBot_5_21[8] , \wRegInBot_5_21[7] , 
        \wRegInBot_5_21[6] , \wRegInBot_5_21[5] , \wRegInBot_5_21[4] , 
        \wRegInBot_5_21[3] , \wRegInBot_5_21[2] , \wRegInBot_5_21[1] , 
        \wRegInBot_5_21[0] }) );
    BHeap_Node_WIDTH32 BHN_6_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_39[0] ), .P_In({\wRegOut_6_39[31] , 
        \wRegOut_6_39[30] , \wRegOut_6_39[29] , \wRegOut_6_39[28] , 
        \wRegOut_6_39[27] , \wRegOut_6_39[26] , \wRegOut_6_39[25] , 
        \wRegOut_6_39[24] , \wRegOut_6_39[23] , \wRegOut_6_39[22] , 
        \wRegOut_6_39[21] , \wRegOut_6_39[20] , \wRegOut_6_39[19] , 
        \wRegOut_6_39[18] , \wRegOut_6_39[17] , \wRegOut_6_39[16] , 
        \wRegOut_6_39[15] , \wRegOut_6_39[14] , \wRegOut_6_39[13] , 
        \wRegOut_6_39[12] , \wRegOut_6_39[11] , \wRegOut_6_39[10] , 
        \wRegOut_6_39[9] , \wRegOut_6_39[8] , \wRegOut_6_39[7] , 
        \wRegOut_6_39[6] , \wRegOut_6_39[5] , \wRegOut_6_39[4] , 
        \wRegOut_6_39[3] , \wRegOut_6_39[2] , \wRegOut_6_39[1] , 
        \wRegOut_6_39[0] }), .P_Out({\wRegInBot_6_39[31] , 
        \wRegInBot_6_39[30] , \wRegInBot_6_39[29] , \wRegInBot_6_39[28] , 
        \wRegInBot_6_39[27] , \wRegInBot_6_39[26] , \wRegInBot_6_39[25] , 
        \wRegInBot_6_39[24] , \wRegInBot_6_39[23] , \wRegInBot_6_39[22] , 
        \wRegInBot_6_39[21] , \wRegInBot_6_39[20] , \wRegInBot_6_39[19] , 
        \wRegInBot_6_39[18] , \wRegInBot_6_39[17] , \wRegInBot_6_39[16] , 
        \wRegInBot_6_39[15] , \wRegInBot_6_39[14] , \wRegInBot_6_39[13] , 
        \wRegInBot_6_39[12] , \wRegInBot_6_39[11] , \wRegInBot_6_39[10] , 
        \wRegInBot_6_39[9] , \wRegInBot_6_39[8] , \wRegInBot_6_39[7] , 
        \wRegInBot_6_39[6] , \wRegInBot_6_39[5] , \wRegInBot_6_39[4] , 
        \wRegInBot_6_39[3] , \wRegInBot_6_39[2] , \wRegInBot_6_39[1] , 
        \wRegInBot_6_39[0] }), .L_WR(\wRegEnTop_7_78[0] ), .L_In({
        \wRegOut_7_78[31] , \wRegOut_7_78[30] , \wRegOut_7_78[29] , 
        \wRegOut_7_78[28] , \wRegOut_7_78[27] , \wRegOut_7_78[26] , 
        \wRegOut_7_78[25] , \wRegOut_7_78[24] , \wRegOut_7_78[23] , 
        \wRegOut_7_78[22] , \wRegOut_7_78[21] , \wRegOut_7_78[20] , 
        \wRegOut_7_78[19] , \wRegOut_7_78[18] , \wRegOut_7_78[17] , 
        \wRegOut_7_78[16] , \wRegOut_7_78[15] , \wRegOut_7_78[14] , 
        \wRegOut_7_78[13] , \wRegOut_7_78[12] , \wRegOut_7_78[11] , 
        \wRegOut_7_78[10] , \wRegOut_7_78[9] , \wRegOut_7_78[8] , 
        \wRegOut_7_78[7] , \wRegOut_7_78[6] , \wRegOut_7_78[5] , 
        \wRegOut_7_78[4] , \wRegOut_7_78[3] , \wRegOut_7_78[2] , 
        \wRegOut_7_78[1] , \wRegOut_7_78[0] }), .L_Out({\wRegInTop_7_78[31] , 
        \wRegInTop_7_78[30] , \wRegInTop_7_78[29] , \wRegInTop_7_78[28] , 
        \wRegInTop_7_78[27] , \wRegInTop_7_78[26] , \wRegInTop_7_78[25] , 
        \wRegInTop_7_78[24] , \wRegInTop_7_78[23] , \wRegInTop_7_78[22] , 
        \wRegInTop_7_78[21] , \wRegInTop_7_78[20] , \wRegInTop_7_78[19] , 
        \wRegInTop_7_78[18] , \wRegInTop_7_78[17] , \wRegInTop_7_78[16] , 
        \wRegInTop_7_78[15] , \wRegInTop_7_78[14] , \wRegInTop_7_78[13] , 
        \wRegInTop_7_78[12] , \wRegInTop_7_78[11] , \wRegInTop_7_78[10] , 
        \wRegInTop_7_78[9] , \wRegInTop_7_78[8] , \wRegInTop_7_78[7] , 
        \wRegInTop_7_78[6] , \wRegInTop_7_78[5] , \wRegInTop_7_78[4] , 
        \wRegInTop_7_78[3] , \wRegInTop_7_78[2] , \wRegInTop_7_78[1] , 
        \wRegInTop_7_78[0] }), .R_WR(\wRegEnTop_7_79[0] ), .R_In({
        \wRegOut_7_79[31] , \wRegOut_7_79[30] , \wRegOut_7_79[29] , 
        \wRegOut_7_79[28] , \wRegOut_7_79[27] , \wRegOut_7_79[26] , 
        \wRegOut_7_79[25] , \wRegOut_7_79[24] , \wRegOut_7_79[23] , 
        \wRegOut_7_79[22] , \wRegOut_7_79[21] , \wRegOut_7_79[20] , 
        \wRegOut_7_79[19] , \wRegOut_7_79[18] , \wRegOut_7_79[17] , 
        \wRegOut_7_79[16] , \wRegOut_7_79[15] , \wRegOut_7_79[14] , 
        \wRegOut_7_79[13] , \wRegOut_7_79[12] , \wRegOut_7_79[11] , 
        \wRegOut_7_79[10] , \wRegOut_7_79[9] , \wRegOut_7_79[8] , 
        \wRegOut_7_79[7] , \wRegOut_7_79[6] , \wRegOut_7_79[5] , 
        \wRegOut_7_79[4] , \wRegOut_7_79[3] , \wRegOut_7_79[2] , 
        \wRegOut_7_79[1] , \wRegOut_7_79[0] }), .R_Out({\wRegInTop_7_79[31] , 
        \wRegInTop_7_79[30] , \wRegInTop_7_79[29] , \wRegInTop_7_79[28] , 
        \wRegInTop_7_79[27] , \wRegInTop_7_79[26] , \wRegInTop_7_79[25] , 
        \wRegInTop_7_79[24] , \wRegInTop_7_79[23] , \wRegInTop_7_79[22] , 
        \wRegInTop_7_79[21] , \wRegInTop_7_79[20] , \wRegInTop_7_79[19] , 
        \wRegInTop_7_79[18] , \wRegInTop_7_79[17] , \wRegInTop_7_79[16] , 
        \wRegInTop_7_79[15] , \wRegInTop_7_79[14] , \wRegInTop_7_79[13] , 
        \wRegInTop_7_79[12] , \wRegInTop_7_79[11] , \wRegInTop_7_79[10] , 
        \wRegInTop_7_79[9] , \wRegInTop_7_79[8] , \wRegInTop_7_79[7] , 
        \wRegInTop_7_79[6] , \wRegInTop_7_79[5] , \wRegInTop_7_79[4] , 
        \wRegInTop_7_79[3] , \wRegInTop_7_79[2] , \wRegInTop_7_79[1] , 
        \wRegInTop_7_79[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink75[31] , \ScanLink75[30] , \ScanLink75[29] , 
        \ScanLink75[28] , \ScanLink75[27] , \ScanLink75[26] , \ScanLink75[25] , 
        \ScanLink75[24] , \ScanLink75[23] , \ScanLink75[22] , \ScanLink75[21] , 
        \ScanLink75[20] , \ScanLink75[19] , \ScanLink75[18] , \ScanLink75[17] , 
        \ScanLink75[16] , \ScanLink75[15] , \ScanLink75[14] , \ScanLink75[13] , 
        \ScanLink75[12] , \ScanLink75[11] , \ScanLink75[10] , \ScanLink75[9] , 
        \ScanLink75[8] , \ScanLink75[7] , \ScanLink75[6] , \ScanLink75[5] , 
        \ScanLink75[4] , \ScanLink75[3] , \ScanLink75[2] , \ScanLink75[1] , 
        \ScanLink75[0] }), .ScanOut({\ScanLink74[31] , \ScanLink74[30] , 
        \ScanLink74[29] , \ScanLink74[28] , \ScanLink74[27] , \ScanLink74[26] , 
        \ScanLink74[25] , \ScanLink74[24] , \ScanLink74[23] , \ScanLink74[22] , 
        \ScanLink74[21] , \ScanLink74[20] , \ScanLink74[19] , \ScanLink74[18] , 
        \ScanLink74[17] , \ScanLink74[16] , \ScanLink74[15] , \ScanLink74[14] , 
        \ScanLink74[13] , \ScanLink74[12] , \ScanLink74[11] , \ScanLink74[10] , 
        \ScanLink74[9] , \ScanLink74[8] , \ScanLink74[7] , \ScanLink74[6] , 
        \ScanLink74[5] , \ScanLink74[4] , \ScanLink74[3] , \ScanLink74[2] , 
        \ScanLink74[1] , \ScanLink74[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_11[31] , \wRegOut_6_11[30] , 
        \wRegOut_6_11[29] , \wRegOut_6_11[28] , \wRegOut_6_11[27] , 
        \wRegOut_6_11[26] , \wRegOut_6_11[25] , \wRegOut_6_11[24] , 
        \wRegOut_6_11[23] , \wRegOut_6_11[22] , \wRegOut_6_11[21] , 
        \wRegOut_6_11[20] , \wRegOut_6_11[19] , \wRegOut_6_11[18] , 
        \wRegOut_6_11[17] , \wRegOut_6_11[16] , \wRegOut_6_11[15] , 
        \wRegOut_6_11[14] , \wRegOut_6_11[13] , \wRegOut_6_11[12] , 
        \wRegOut_6_11[11] , \wRegOut_6_11[10] , \wRegOut_6_11[9] , 
        \wRegOut_6_11[8] , \wRegOut_6_11[7] , \wRegOut_6_11[6] , 
        \wRegOut_6_11[5] , \wRegOut_6_11[4] , \wRegOut_6_11[3] , 
        \wRegOut_6_11[2] , \wRegOut_6_11[1] , \wRegOut_6_11[0] }), .Enable1(
        \wRegEnTop_6_11[0] ), .Enable2(\wRegEnBot_6_11[0] ), .In1({
        \wRegInTop_6_11[31] , \wRegInTop_6_11[30] , \wRegInTop_6_11[29] , 
        \wRegInTop_6_11[28] , \wRegInTop_6_11[27] , \wRegInTop_6_11[26] , 
        \wRegInTop_6_11[25] , \wRegInTop_6_11[24] , \wRegInTop_6_11[23] , 
        \wRegInTop_6_11[22] , \wRegInTop_6_11[21] , \wRegInTop_6_11[20] , 
        \wRegInTop_6_11[19] , \wRegInTop_6_11[18] , \wRegInTop_6_11[17] , 
        \wRegInTop_6_11[16] , \wRegInTop_6_11[15] , \wRegInTop_6_11[14] , 
        \wRegInTop_6_11[13] , \wRegInTop_6_11[12] , \wRegInTop_6_11[11] , 
        \wRegInTop_6_11[10] , \wRegInTop_6_11[9] , \wRegInTop_6_11[8] , 
        \wRegInTop_6_11[7] , \wRegInTop_6_11[6] , \wRegInTop_6_11[5] , 
        \wRegInTop_6_11[4] , \wRegInTop_6_11[3] , \wRegInTop_6_11[2] , 
        \wRegInTop_6_11[1] , \wRegInTop_6_11[0] }), .In2({\wRegInBot_6_11[31] , 
        \wRegInBot_6_11[30] , \wRegInBot_6_11[29] , \wRegInBot_6_11[28] , 
        \wRegInBot_6_11[27] , \wRegInBot_6_11[26] , \wRegInBot_6_11[25] , 
        \wRegInBot_6_11[24] , \wRegInBot_6_11[23] , \wRegInBot_6_11[22] , 
        \wRegInBot_6_11[21] , \wRegInBot_6_11[20] , \wRegInBot_6_11[19] , 
        \wRegInBot_6_11[18] , \wRegInBot_6_11[17] , \wRegInBot_6_11[16] , 
        \wRegInBot_6_11[15] , \wRegInBot_6_11[14] , \wRegInBot_6_11[13] , 
        \wRegInBot_6_11[12] , \wRegInBot_6_11[11] , \wRegInBot_6_11[10] , 
        \wRegInBot_6_11[9] , \wRegInBot_6_11[8] , \wRegInBot_6_11[7] , 
        \wRegInBot_6_11[6] , \wRegInBot_6_11[5] , \wRegInBot_6_11[4] , 
        \wRegInBot_6_11[3] , \wRegInBot_6_11[2] , \wRegInBot_6_11[1] , 
        \wRegInBot_6_11[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_65 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink193[31] , \ScanLink193[30] , \ScanLink193[29] , 
        \ScanLink193[28] , \ScanLink193[27] , \ScanLink193[26] , 
        \ScanLink193[25] , \ScanLink193[24] , \ScanLink193[23] , 
        \ScanLink193[22] , \ScanLink193[21] , \ScanLink193[20] , 
        \ScanLink193[19] , \ScanLink193[18] , \ScanLink193[17] , 
        \ScanLink193[16] , \ScanLink193[15] , \ScanLink193[14] , 
        \ScanLink193[13] , \ScanLink193[12] , \ScanLink193[11] , 
        \ScanLink193[10] , \ScanLink193[9] , \ScanLink193[8] , 
        \ScanLink193[7] , \ScanLink193[6] , \ScanLink193[5] , \ScanLink193[4] , 
        \ScanLink193[3] , \ScanLink193[2] , \ScanLink193[1] , \ScanLink193[0] 
        }), .ScanOut({\ScanLink192[31] , \ScanLink192[30] , \ScanLink192[29] , 
        \ScanLink192[28] , \ScanLink192[27] , \ScanLink192[26] , 
        \ScanLink192[25] , \ScanLink192[24] , \ScanLink192[23] , 
        \ScanLink192[22] , \ScanLink192[21] , \ScanLink192[20] , 
        \ScanLink192[19] , \ScanLink192[18] , \ScanLink192[17] , 
        \ScanLink192[16] , \ScanLink192[15] , \ScanLink192[14] , 
        \ScanLink192[13] , \ScanLink192[12] , \ScanLink192[11] , 
        \ScanLink192[10] , \ScanLink192[9] , \ScanLink192[8] , 
        \ScanLink192[7] , \ScanLink192[6] , \ScanLink192[5] , \ScanLink192[4] , 
        \ScanLink192[3] , \ScanLink192[2] , \ScanLink192[1] , \ScanLink192[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_65[31] , 
        \wRegOut_7_65[30] , \wRegOut_7_65[29] , \wRegOut_7_65[28] , 
        \wRegOut_7_65[27] , \wRegOut_7_65[26] , \wRegOut_7_65[25] , 
        \wRegOut_7_65[24] , \wRegOut_7_65[23] , \wRegOut_7_65[22] , 
        \wRegOut_7_65[21] , \wRegOut_7_65[20] , \wRegOut_7_65[19] , 
        \wRegOut_7_65[18] , \wRegOut_7_65[17] , \wRegOut_7_65[16] , 
        \wRegOut_7_65[15] , \wRegOut_7_65[14] , \wRegOut_7_65[13] , 
        \wRegOut_7_65[12] , \wRegOut_7_65[11] , \wRegOut_7_65[10] , 
        \wRegOut_7_65[9] , \wRegOut_7_65[8] , \wRegOut_7_65[7] , 
        \wRegOut_7_65[6] , \wRegOut_7_65[5] , \wRegOut_7_65[4] , 
        \wRegOut_7_65[3] , \wRegOut_7_65[2] , \wRegOut_7_65[1] , 
        \wRegOut_7_65[0] }), .Enable1(\wRegEnTop_7_65[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_65[31] , \wRegInTop_7_65[30] , \wRegInTop_7_65[29] , 
        \wRegInTop_7_65[28] , \wRegInTop_7_65[27] , \wRegInTop_7_65[26] , 
        \wRegInTop_7_65[25] , \wRegInTop_7_65[24] , \wRegInTop_7_65[23] , 
        \wRegInTop_7_65[22] , \wRegInTop_7_65[21] , \wRegInTop_7_65[20] , 
        \wRegInTop_7_65[19] , \wRegInTop_7_65[18] , \wRegInTop_7_65[17] , 
        \wRegInTop_7_65[16] , \wRegInTop_7_65[15] , \wRegInTop_7_65[14] , 
        \wRegInTop_7_65[13] , \wRegInTop_7_65[12] , \wRegInTop_7_65[11] , 
        \wRegInTop_7_65[10] , \wRegInTop_7_65[9] , \wRegInTop_7_65[8] , 
        \wRegInTop_7_65[7] , \wRegInTop_7_65[6] , \wRegInTop_7_65[5] , 
        \wRegInTop_7_65[4] , \wRegInTop_7_65[3] , \wRegInTop_7_65[2] , 
        \wRegInTop_7_65[1] , \wRegInTop_7_65[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_29 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink61[31] , \ScanLink61[30] , \ScanLink61[29] , 
        \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , \ScanLink61[25] , 
        \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , \ScanLink61[21] , 
        \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , \ScanLink61[17] , 
        \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , \ScanLink61[13] , 
        \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , \ScanLink61[9] , 
        \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , \ScanLink61[5] , 
        \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , \ScanLink61[1] , 
        \ScanLink61[0] }), .ScanOut({\ScanLink60[31] , \ScanLink60[30] , 
        \ScanLink60[29] , \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , 
        \ScanLink60[25] , \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , 
        \ScanLink60[21] , \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , 
        \ScanLink60[17] , \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , 
        \ScanLink60[13] , \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , 
        \ScanLink60[9] , \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , 
        \ScanLink60[5] , \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , 
        \ScanLink60[1] , \ScanLink60[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_29[31] , \wRegOut_5_29[30] , 
        \wRegOut_5_29[29] , \wRegOut_5_29[28] , \wRegOut_5_29[27] , 
        \wRegOut_5_29[26] , \wRegOut_5_29[25] , \wRegOut_5_29[24] , 
        \wRegOut_5_29[23] , \wRegOut_5_29[22] , \wRegOut_5_29[21] , 
        \wRegOut_5_29[20] , \wRegOut_5_29[19] , \wRegOut_5_29[18] , 
        \wRegOut_5_29[17] , \wRegOut_5_29[16] , \wRegOut_5_29[15] , 
        \wRegOut_5_29[14] , \wRegOut_5_29[13] , \wRegOut_5_29[12] , 
        \wRegOut_5_29[11] , \wRegOut_5_29[10] , \wRegOut_5_29[9] , 
        \wRegOut_5_29[8] , \wRegOut_5_29[7] , \wRegOut_5_29[6] , 
        \wRegOut_5_29[5] , \wRegOut_5_29[4] , \wRegOut_5_29[3] , 
        \wRegOut_5_29[2] , \wRegOut_5_29[1] , \wRegOut_5_29[0] }), .Enable1(
        \wRegEnTop_5_29[0] ), .Enable2(\wRegEnBot_5_29[0] ), .In1({
        \wRegInTop_5_29[31] , \wRegInTop_5_29[30] , \wRegInTop_5_29[29] , 
        \wRegInTop_5_29[28] , \wRegInTop_5_29[27] , \wRegInTop_5_29[26] , 
        \wRegInTop_5_29[25] , \wRegInTop_5_29[24] , \wRegInTop_5_29[23] , 
        \wRegInTop_5_29[22] , \wRegInTop_5_29[21] , \wRegInTop_5_29[20] , 
        \wRegInTop_5_29[19] , \wRegInTop_5_29[18] , \wRegInTop_5_29[17] , 
        \wRegInTop_5_29[16] , \wRegInTop_5_29[15] , \wRegInTop_5_29[14] , 
        \wRegInTop_5_29[13] , \wRegInTop_5_29[12] , \wRegInTop_5_29[11] , 
        \wRegInTop_5_29[10] , \wRegInTop_5_29[9] , \wRegInTop_5_29[8] , 
        \wRegInTop_5_29[7] , \wRegInTop_5_29[6] , \wRegInTop_5_29[5] , 
        \wRegInTop_5_29[4] , \wRegInTop_5_29[3] , \wRegInTop_5_29[2] , 
        \wRegInTop_5_29[1] , \wRegInTop_5_29[0] }), .In2({\wRegInBot_5_29[31] , 
        \wRegInBot_5_29[30] , \wRegInBot_5_29[29] , \wRegInBot_5_29[28] , 
        \wRegInBot_5_29[27] , \wRegInBot_5_29[26] , \wRegInBot_5_29[25] , 
        \wRegInBot_5_29[24] , \wRegInBot_5_29[23] , \wRegInBot_5_29[22] , 
        \wRegInBot_5_29[21] , \wRegInBot_5_29[20] , \wRegInBot_5_29[19] , 
        \wRegInBot_5_29[18] , \wRegInBot_5_29[17] , \wRegInBot_5_29[16] , 
        \wRegInBot_5_29[15] , \wRegInBot_5_29[14] , \wRegInBot_5_29[13] , 
        \wRegInBot_5_29[12] , \wRegInBot_5_29[11] , \wRegInBot_5_29[10] , 
        \wRegInBot_5_29[9] , \wRegInBot_5_29[8] , \wRegInBot_5_29[7] , 
        \wRegInBot_5_29[6] , \wRegInBot_5_29[5] , \wRegInBot_5_29[4] , 
        \wRegInBot_5_29[3] , \wRegInBot_5_29[2] , \wRegInBot_5_29[1] , 
        \wRegInBot_5_29[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_19 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink83[31] , \ScanLink83[30] , \ScanLink83[29] , 
        \ScanLink83[28] , \ScanLink83[27] , \ScanLink83[26] , \ScanLink83[25] , 
        \ScanLink83[24] , \ScanLink83[23] , \ScanLink83[22] , \ScanLink83[21] , 
        \ScanLink83[20] , \ScanLink83[19] , \ScanLink83[18] , \ScanLink83[17] , 
        \ScanLink83[16] , \ScanLink83[15] , \ScanLink83[14] , \ScanLink83[13] , 
        \ScanLink83[12] , \ScanLink83[11] , \ScanLink83[10] , \ScanLink83[9] , 
        \ScanLink83[8] , \ScanLink83[7] , \ScanLink83[6] , \ScanLink83[5] , 
        \ScanLink83[4] , \ScanLink83[3] , \ScanLink83[2] , \ScanLink83[1] , 
        \ScanLink83[0] }), .ScanOut({\ScanLink82[31] , \ScanLink82[30] , 
        \ScanLink82[29] , \ScanLink82[28] , \ScanLink82[27] , \ScanLink82[26] , 
        \ScanLink82[25] , \ScanLink82[24] , \ScanLink82[23] , \ScanLink82[22] , 
        \ScanLink82[21] , \ScanLink82[20] , \ScanLink82[19] , \ScanLink82[18] , 
        \ScanLink82[17] , \ScanLink82[16] , \ScanLink82[15] , \ScanLink82[14] , 
        \ScanLink82[13] , \ScanLink82[12] , \ScanLink82[11] , \ScanLink82[10] , 
        \ScanLink82[9] , \ScanLink82[8] , \ScanLink82[7] , \ScanLink82[6] , 
        \ScanLink82[5] , \ScanLink82[4] , \ScanLink82[3] , \ScanLink82[2] , 
        \ScanLink82[1] , \ScanLink82[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_19[31] , \wRegOut_6_19[30] , 
        \wRegOut_6_19[29] , \wRegOut_6_19[28] , \wRegOut_6_19[27] , 
        \wRegOut_6_19[26] , \wRegOut_6_19[25] , \wRegOut_6_19[24] , 
        \wRegOut_6_19[23] , \wRegOut_6_19[22] , \wRegOut_6_19[21] , 
        \wRegOut_6_19[20] , \wRegOut_6_19[19] , \wRegOut_6_19[18] , 
        \wRegOut_6_19[17] , \wRegOut_6_19[16] , \wRegOut_6_19[15] , 
        \wRegOut_6_19[14] , \wRegOut_6_19[13] , \wRegOut_6_19[12] , 
        \wRegOut_6_19[11] , \wRegOut_6_19[10] , \wRegOut_6_19[9] , 
        \wRegOut_6_19[8] , \wRegOut_6_19[7] , \wRegOut_6_19[6] , 
        \wRegOut_6_19[5] , \wRegOut_6_19[4] , \wRegOut_6_19[3] , 
        \wRegOut_6_19[2] , \wRegOut_6_19[1] , \wRegOut_6_19[0] }), .Enable1(
        \wRegEnTop_6_19[0] ), .Enable2(\wRegEnBot_6_19[0] ), .In1({
        \wRegInTop_6_19[31] , \wRegInTop_6_19[30] , \wRegInTop_6_19[29] , 
        \wRegInTop_6_19[28] , \wRegInTop_6_19[27] , \wRegInTop_6_19[26] , 
        \wRegInTop_6_19[25] , \wRegInTop_6_19[24] , \wRegInTop_6_19[23] , 
        \wRegInTop_6_19[22] , \wRegInTop_6_19[21] , \wRegInTop_6_19[20] , 
        \wRegInTop_6_19[19] , \wRegInTop_6_19[18] , \wRegInTop_6_19[17] , 
        \wRegInTop_6_19[16] , \wRegInTop_6_19[15] , \wRegInTop_6_19[14] , 
        \wRegInTop_6_19[13] , \wRegInTop_6_19[12] , \wRegInTop_6_19[11] , 
        \wRegInTop_6_19[10] , \wRegInTop_6_19[9] , \wRegInTop_6_19[8] , 
        \wRegInTop_6_19[7] , \wRegInTop_6_19[6] , \wRegInTop_6_19[5] , 
        \wRegInTop_6_19[4] , \wRegInTop_6_19[3] , \wRegInTop_6_19[2] , 
        \wRegInTop_6_19[1] , \wRegInTop_6_19[0] }), .In2({\wRegInBot_6_19[31] , 
        \wRegInBot_6_19[30] , \wRegInBot_6_19[29] , \wRegInBot_6_19[28] , 
        \wRegInBot_6_19[27] , \wRegInBot_6_19[26] , \wRegInBot_6_19[25] , 
        \wRegInBot_6_19[24] , \wRegInBot_6_19[23] , \wRegInBot_6_19[22] , 
        \wRegInBot_6_19[21] , \wRegInBot_6_19[20] , \wRegInBot_6_19[19] , 
        \wRegInBot_6_19[18] , \wRegInBot_6_19[17] , \wRegInBot_6_19[16] , 
        \wRegInBot_6_19[15] , \wRegInBot_6_19[14] , \wRegInBot_6_19[13] , 
        \wRegInBot_6_19[12] , \wRegInBot_6_19[11] , \wRegInBot_6_19[10] , 
        \wRegInBot_6_19[9] , \wRegInBot_6_19[8] , \wRegInBot_6_19[7] , 
        \wRegInBot_6_19[6] , \wRegInBot_6_19[5] , \wRegInBot_6_19[4] , 
        \wRegInBot_6_19[3] , \wRegInBot_6_19[2] , \wRegInBot_6_19[1] , 
        \wRegInBot_6_19[0] }) );
    BHeap_Node_WIDTH32 BHN_6_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_31[0] ), .P_In({\wRegOut_6_31[31] , 
        \wRegOut_6_31[30] , \wRegOut_6_31[29] , \wRegOut_6_31[28] , 
        \wRegOut_6_31[27] , \wRegOut_6_31[26] , \wRegOut_6_31[25] , 
        \wRegOut_6_31[24] , \wRegOut_6_31[23] , \wRegOut_6_31[22] , 
        \wRegOut_6_31[21] , \wRegOut_6_31[20] , \wRegOut_6_31[19] , 
        \wRegOut_6_31[18] , \wRegOut_6_31[17] , \wRegOut_6_31[16] , 
        \wRegOut_6_31[15] , \wRegOut_6_31[14] , \wRegOut_6_31[13] , 
        \wRegOut_6_31[12] , \wRegOut_6_31[11] , \wRegOut_6_31[10] , 
        \wRegOut_6_31[9] , \wRegOut_6_31[8] , \wRegOut_6_31[7] , 
        \wRegOut_6_31[6] , \wRegOut_6_31[5] , \wRegOut_6_31[4] , 
        \wRegOut_6_31[3] , \wRegOut_6_31[2] , \wRegOut_6_31[1] , 
        \wRegOut_6_31[0] }), .P_Out({\wRegInBot_6_31[31] , 
        \wRegInBot_6_31[30] , \wRegInBot_6_31[29] , \wRegInBot_6_31[28] , 
        \wRegInBot_6_31[27] , \wRegInBot_6_31[26] , \wRegInBot_6_31[25] , 
        \wRegInBot_6_31[24] , \wRegInBot_6_31[23] , \wRegInBot_6_31[22] , 
        \wRegInBot_6_31[21] , \wRegInBot_6_31[20] , \wRegInBot_6_31[19] , 
        \wRegInBot_6_31[18] , \wRegInBot_6_31[17] , \wRegInBot_6_31[16] , 
        \wRegInBot_6_31[15] , \wRegInBot_6_31[14] , \wRegInBot_6_31[13] , 
        \wRegInBot_6_31[12] , \wRegInBot_6_31[11] , \wRegInBot_6_31[10] , 
        \wRegInBot_6_31[9] , \wRegInBot_6_31[8] , \wRegInBot_6_31[7] , 
        \wRegInBot_6_31[6] , \wRegInBot_6_31[5] , \wRegInBot_6_31[4] , 
        \wRegInBot_6_31[3] , \wRegInBot_6_31[2] , \wRegInBot_6_31[1] , 
        \wRegInBot_6_31[0] }), .L_WR(\wRegEnTop_7_62[0] ), .L_In({
        \wRegOut_7_62[31] , \wRegOut_7_62[30] , \wRegOut_7_62[29] , 
        \wRegOut_7_62[28] , \wRegOut_7_62[27] , \wRegOut_7_62[26] , 
        \wRegOut_7_62[25] , \wRegOut_7_62[24] , \wRegOut_7_62[23] , 
        \wRegOut_7_62[22] , \wRegOut_7_62[21] , \wRegOut_7_62[20] , 
        \wRegOut_7_62[19] , \wRegOut_7_62[18] , \wRegOut_7_62[17] , 
        \wRegOut_7_62[16] , \wRegOut_7_62[15] , \wRegOut_7_62[14] , 
        \wRegOut_7_62[13] , \wRegOut_7_62[12] , \wRegOut_7_62[11] , 
        \wRegOut_7_62[10] , \wRegOut_7_62[9] , \wRegOut_7_62[8] , 
        \wRegOut_7_62[7] , \wRegOut_7_62[6] , \wRegOut_7_62[5] , 
        \wRegOut_7_62[4] , \wRegOut_7_62[3] , \wRegOut_7_62[2] , 
        \wRegOut_7_62[1] , \wRegOut_7_62[0] }), .L_Out({\wRegInTop_7_62[31] , 
        \wRegInTop_7_62[30] , \wRegInTop_7_62[29] , \wRegInTop_7_62[28] , 
        \wRegInTop_7_62[27] , \wRegInTop_7_62[26] , \wRegInTop_7_62[25] , 
        \wRegInTop_7_62[24] , \wRegInTop_7_62[23] , \wRegInTop_7_62[22] , 
        \wRegInTop_7_62[21] , \wRegInTop_7_62[20] , \wRegInTop_7_62[19] , 
        \wRegInTop_7_62[18] , \wRegInTop_7_62[17] , \wRegInTop_7_62[16] , 
        \wRegInTop_7_62[15] , \wRegInTop_7_62[14] , \wRegInTop_7_62[13] , 
        \wRegInTop_7_62[12] , \wRegInTop_7_62[11] , \wRegInTop_7_62[10] , 
        \wRegInTop_7_62[9] , \wRegInTop_7_62[8] , \wRegInTop_7_62[7] , 
        \wRegInTop_7_62[6] , \wRegInTop_7_62[5] , \wRegInTop_7_62[4] , 
        \wRegInTop_7_62[3] , \wRegInTop_7_62[2] , \wRegInTop_7_62[1] , 
        \wRegInTop_7_62[0] }), .R_WR(\wRegEnTop_7_63[0] ), .R_In({
        \wRegOut_7_63[31] , \wRegOut_7_63[30] , \wRegOut_7_63[29] , 
        \wRegOut_7_63[28] , \wRegOut_7_63[27] , \wRegOut_7_63[26] , 
        \wRegOut_7_63[25] , \wRegOut_7_63[24] , \wRegOut_7_63[23] , 
        \wRegOut_7_63[22] , \wRegOut_7_63[21] , \wRegOut_7_63[20] , 
        \wRegOut_7_63[19] , \wRegOut_7_63[18] , \wRegOut_7_63[17] , 
        \wRegOut_7_63[16] , \wRegOut_7_63[15] , \wRegOut_7_63[14] , 
        \wRegOut_7_63[13] , \wRegOut_7_63[12] , \wRegOut_7_63[11] , 
        \wRegOut_7_63[10] , \wRegOut_7_63[9] , \wRegOut_7_63[8] , 
        \wRegOut_7_63[7] , \wRegOut_7_63[6] , \wRegOut_7_63[5] , 
        \wRegOut_7_63[4] , \wRegOut_7_63[3] , \wRegOut_7_63[2] , 
        \wRegOut_7_63[1] , \wRegOut_7_63[0] }), .R_Out({\wRegInTop_7_63[31] , 
        \wRegInTop_7_63[30] , \wRegInTop_7_63[29] , \wRegInTop_7_63[28] , 
        \wRegInTop_7_63[27] , \wRegInTop_7_63[26] , \wRegInTop_7_63[25] , 
        \wRegInTop_7_63[24] , \wRegInTop_7_63[23] , \wRegInTop_7_63[22] , 
        \wRegInTop_7_63[21] , \wRegInTop_7_63[20] , \wRegInTop_7_63[19] , 
        \wRegInTop_7_63[18] , \wRegInTop_7_63[17] , \wRegInTop_7_63[16] , 
        \wRegInTop_7_63[15] , \wRegInTop_7_63[14] , \wRegInTop_7_63[13] , 
        \wRegInTop_7_63[12] , \wRegInTop_7_63[11] , \wRegInTop_7_63[10] , 
        \wRegInTop_7_63[9] , \wRegInTop_7_63[8] , \wRegInTop_7_63[7] , 
        \wRegInTop_7_63[6] , \wRegInTop_7_63[5] , \wRegInTop_7_63[4] , 
        \wRegInTop_7_63[3] , \wRegInTop_7_63[2] , \wRegInTop_7_63[1] , 
        \wRegInTop_7_63[0] }) );
    BHeap_Node_WIDTH32 BHN_5_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_26[0] ), .P_In({\wRegOut_5_26[31] , 
        \wRegOut_5_26[30] , \wRegOut_5_26[29] , \wRegOut_5_26[28] , 
        \wRegOut_5_26[27] , \wRegOut_5_26[26] , \wRegOut_5_26[25] , 
        \wRegOut_5_26[24] , \wRegOut_5_26[23] , \wRegOut_5_26[22] , 
        \wRegOut_5_26[21] , \wRegOut_5_26[20] , \wRegOut_5_26[19] , 
        \wRegOut_5_26[18] , \wRegOut_5_26[17] , \wRegOut_5_26[16] , 
        \wRegOut_5_26[15] , \wRegOut_5_26[14] , \wRegOut_5_26[13] , 
        \wRegOut_5_26[12] , \wRegOut_5_26[11] , \wRegOut_5_26[10] , 
        \wRegOut_5_26[9] , \wRegOut_5_26[8] , \wRegOut_5_26[7] , 
        \wRegOut_5_26[6] , \wRegOut_5_26[5] , \wRegOut_5_26[4] , 
        \wRegOut_5_26[3] , \wRegOut_5_26[2] , \wRegOut_5_26[1] , 
        \wRegOut_5_26[0] }), .P_Out({\wRegInBot_5_26[31] , 
        \wRegInBot_5_26[30] , \wRegInBot_5_26[29] , \wRegInBot_5_26[28] , 
        \wRegInBot_5_26[27] , \wRegInBot_5_26[26] , \wRegInBot_5_26[25] , 
        \wRegInBot_5_26[24] , \wRegInBot_5_26[23] , \wRegInBot_5_26[22] , 
        \wRegInBot_5_26[21] , \wRegInBot_5_26[20] , \wRegInBot_5_26[19] , 
        \wRegInBot_5_26[18] , \wRegInBot_5_26[17] , \wRegInBot_5_26[16] , 
        \wRegInBot_5_26[15] , \wRegInBot_5_26[14] , \wRegInBot_5_26[13] , 
        \wRegInBot_5_26[12] , \wRegInBot_5_26[11] , \wRegInBot_5_26[10] , 
        \wRegInBot_5_26[9] , \wRegInBot_5_26[8] , \wRegInBot_5_26[7] , 
        \wRegInBot_5_26[6] , \wRegInBot_5_26[5] , \wRegInBot_5_26[4] , 
        \wRegInBot_5_26[3] , \wRegInBot_5_26[2] , \wRegInBot_5_26[1] , 
        \wRegInBot_5_26[0] }), .L_WR(\wRegEnTop_6_52[0] ), .L_In({
        \wRegOut_6_52[31] , \wRegOut_6_52[30] , \wRegOut_6_52[29] , 
        \wRegOut_6_52[28] , \wRegOut_6_52[27] , \wRegOut_6_52[26] , 
        \wRegOut_6_52[25] , \wRegOut_6_52[24] , \wRegOut_6_52[23] , 
        \wRegOut_6_52[22] , \wRegOut_6_52[21] , \wRegOut_6_52[20] , 
        \wRegOut_6_52[19] , \wRegOut_6_52[18] , \wRegOut_6_52[17] , 
        \wRegOut_6_52[16] , \wRegOut_6_52[15] , \wRegOut_6_52[14] , 
        \wRegOut_6_52[13] , \wRegOut_6_52[12] , \wRegOut_6_52[11] , 
        \wRegOut_6_52[10] , \wRegOut_6_52[9] , \wRegOut_6_52[8] , 
        \wRegOut_6_52[7] , \wRegOut_6_52[6] , \wRegOut_6_52[5] , 
        \wRegOut_6_52[4] , \wRegOut_6_52[3] , \wRegOut_6_52[2] , 
        \wRegOut_6_52[1] , \wRegOut_6_52[0] }), .L_Out({\wRegInTop_6_52[31] , 
        \wRegInTop_6_52[30] , \wRegInTop_6_52[29] , \wRegInTop_6_52[28] , 
        \wRegInTop_6_52[27] , \wRegInTop_6_52[26] , \wRegInTop_6_52[25] , 
        \wRegInTop_6_52[24] , \wRegInTop_6_52[23] , \wRegInTop_6_52[22] , 
        \wRegInTop_6_52[21] , \wRegInTop_6_52[20] , \wRegInTop_6_52[19] , 
        \wRegInTop_6_52[18] , \wRegInTop_6_52[17] , \wRegInTop_6_52[16] , 
        \wRegInTop_6_52[15] , \wRegInTop_6_52[14] , \wRegInTop_6_52[13] , 
        \wRegInTop_6_52[12] , \wRegInTop_6_52[11] , \wRegInTop_6_52[10] , 
        \wRegInTop_6_52[9] , \wRegInTop_6_52[8] , \wRegInTop_6_52[7] , 
        \wRegInTop_6_52[6] , \wRegInTop_6_52[5] , \wRegInTop_6_52[4] , 
        \wRegInTop_6_52[3] , \wRegInTop_6_52[2] , \wRegInTop_6_52[1] , 
        \wRegInTop_6_52[0] }), .R_WR(\wRegEnTop_6_53[0] ), .R_In({
        \wRegOut_6_53[31] , \wRegOut_6_53[30] , \wRegOut_6_53[29] , 
        \wRegOut_6_53[28] , \wRegOut_6_53[27] , \wRegOut_6_53[26] , 
        \wRegOut_6_53[25] , \wRegOut_6_53[24] , \wRegOut_6_53[23] , 
        \wRegOut_6_53[22] , \wRegOut_6_53[21] , \wRegOut_6_53[20] , 
        \wRegOut_6_53[19] , \wRegOut_6_53[18] , \wRegOut_6_53[17] , 
        \wRegOut_6_53[16] , \wRegOut_6_53[15] , \wRegOut_6_53[14] , 
        \wRegOut_6_53[13] , \wRegOut_6_53[12] , \wRegOut_6_53[11] , 
        \wRegOut_6_53[10] , \wRegOut_6_53[9] , \wRegOut_6_53[8] , 
        \wRegOut_6_53[7] , \wRegOut_6_53[6] , \wRegOut_6_53[5] , 
        \wRegOut_6_53[4] , \wRegOut_6_53[3] , \wRegOut_6_53[2] , 
        \wRegOut_6_53[1] , \wRegOut_6_53[0] }), .R_Out({\wRegInTop_6_53[31] , 
        \wRegInTop_6_53[30] , \wRegInTop_6_53[29] , \wRegInTop_6_53[28] , 
        \wRegInTop_6_53[27] , \wRegInTop_6_53[26] , \wRegInTop_6_53[25] , 
        \wRegInTop_6_53[24] , \wRegInTop_6_53[23] , \wRegInTop_6_53[22] , 
        \wRegInTop_6_53[21] , \wRegInTop_6_53[20] , \wRegInTop_6_53[19] , 
        \wRegInTop_6_53[18] , \wRegInTop_6_53[17] , \wRegInTop_6_53[16] , 
        \wRegInTop_6_53[15] , \wRegInTop_6_53[14] , \wRegInTop_6_53[13] , 
        \wRegInTop_6_53[12] , \wRegInTop_6_53[11] , \wRegInTop_6_53[10] , 
        \wRegInTop_6_53[9] , \wRegInTop_6_53[8] , \wRegInTop_6_53[7] , 
        \wRegInTop_6_53[6] , \wRegInTop_6_53[5] , \wRegInTop_6_53[4] , 
        \wRegInTop_6_53[3] , \wRegInTop_6_53[2] , \wRegInTop_6_53[1] , 
        \wRegInTop_6_53[0] }) );
    BHeap_Node_WIDTH32 BHN_6_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_16[0] ), .P_In({\wRegOut_6_16[31] , 
        \wRegOut_6_16[30] , \wRegOut_6_16[29] , \wRegOut_6_16[28] , 
        \wRegOut_6_16[27] , \wRegOut_6_16[26] , \wRegOut_6_16[25] , 
        \wRegOut_6_16[24] , \wRegOut_6_16[23] , \wRegOut_6_16[22] , 
        \wRegOut_6_16[21] , \wRegOut_6_16[20] , \wRegOut_6_16[19] , 
        \wRegOut_6_16[18] , \wRegOut_6_16[17] , \wRegOut_6_16[16] , 
        \wRegOut_6_16[15] , \wRegOut_6_16[14] , \wRegOut_6_16[13] , 
        \wRegOut_6_16[12] , \wRegOut_6_16[11] , \wRegOut_6_16[10] , 
        \wRegOut_6_16[9] , \wRegOut_6_16[8] , \wRegOut_6_16[7] , 
        \wRegOut_6_16[6] , \wRegOut_6_16[5] , \wRegOut_6_16[4] , 
        \wRegOut_6_16[3] , \wRegOut_6_16[2] , \wRegOut_6_16[1] , 
        \wRegOut_6_16[0] }), .P_Out({\wRegInBot_6_16[31] , 
        \wRegInBot_6_16[30] , \wRegInBot_6_16[29] , \wRegInBot_6_16[28] , 
        \wRegInBot_6_16[27] , \wRegInBot_6_16[26] , \wRegInBot_6_16[25] , 
        \wRegInBot_6_16[24] , \wRegInBot_6_16[23] , \wRegInBot_6_16[22] , 
        \wRegInBot_6_16[21] , \wRegInBot_6_16[20] , \wRegInBot_6_16[19] , 
        \wRegInBot_6_16[18] , \wRegInBot_6_16[17] , \wRegInBot_6_16[16] , 
        \wRegInBot_6_16[15] , \wRegInBot_6_16[14] , \wRegInBot_6_16[13] , 
        \wRegInBot_6_16[12] , \wRegInBot_6_16[11] , \wRegInBot_6_16[10] , 
        \wRegInBot_6_16[9] , \wRegInBot_6_16[8] , \wRegInBot_6_16[7] , 
        \wRegInBot_6_16[6] , \wRegInBot_6_16[5] , \wRegInBot_6_16[4] , 
        \wRegInBot_6_16[3] , \wRegInBot_6_16[2] , \wRegInBot_6_16[1] , 
        \wRegInBot_6_16[0] }), .L_WR(\wRegEnTop_7_32[0] ), .L_In({
        \wRegOut_7_32[31] , \wRegOut_7_32[30] , \wRegOut_7_32[29] , 
        \wRegOut_7_32[28] , \wRegOut_7_32[27] , \wRegOut_7_32[26] , 
        \wRegOut_7_32[25] , \wRegOut_7_32[24] , \wRegOut_7_32[23] , 
        \wRegOut_7_32[22] , \wRegOut_7_32[21] , \wRegOut_7_32[20] , 
        \wRegOut_7_32[19] , \wRegOut_7_32[18] , \wRegOut_7_32[17] , 
        \wRegOut_7_32[16] , \wRegOut_7_32[15] , \wRegOut_7_32[14] , 
        \wRegOut_7_32[13] , \wRegOut_7_32[12] , \wRegOut_7_32[11] , 
        \wRegOut_7_32[10] , \wRegOut_7_32[9] , \wRegOut_7_32[8] , 
        \wRegOut_7_32[7] , \wRegOut_7_32[6] , \wRegOut_7_32[5] , 
        \wRegOut_7_32[4] , \wRegOut_7_32[3] , \wRegOut_7_32[2] , 
        \wRegOut_7_32[1] , \wRegOut_7_32[0] }), .L_Out({\wRegInTop_7_32[31] , 
        \wRegInTop_7_32[30] , \wRegInTop_7_32[29] , \wRegInTop_7_32[28] , 
        \wRegInTop_7_32[27] , \wRegInTop_7_32[26] , \wRegInTop_7_32[25] , 
        \wRegInTop_7_32[24] , \wRegInTop_7_32[23] , \wRegInTop_7_32[22] , 
        \wRegInTop_7_32[21] , \wRegInTop_7_32[20] , \wRegInTop_7_32[19] , 
        \wRegInTop_7_32[18] , \wRegInTop_7_32[17] , \wRegInTop_7_32[16] , 
        \wRegInTop_7_32[15] , \wRegInTop_7_32[14] , \wRegInTop_7_32[13] , 
        \wRegInTop_7_32[12] , \wRegInTop_7_32[11] , \wRegInTop_7_32[10] , 
        \wRegInTop_7_32[9] , \wRegInTop_7_32[8] , \wRegInTop_7_32[7] , 
        \wRegInTop_7_32[6] , \wRegInTop_7_32[5] , \wRegInTop_7_32[4] , 
        \wRegInTop_7_32[3] , \wRegInTop_7_32[2] , \wRegInTop_7_32[1] , 
        \wRegInTop_7_32[0] }), .R_WR(\wRegEnTop_7_33[0] ), .R_In({
        \wRegOut_7_33[31] , \wRegOut_7_33[30] , \wRegOut_7_33[29] , 
        \wRegOut_7_33[28] , \wRegOut_7_33[27] , \wRegOut_7_33[26] , 
        \wRegOut_7_33[25] , \wRegOut_7_33[24] , \wRegOut_7_33[23] , 
        \wRegOut_7_33[22] , \wRegOut_7_33[21] , \wRegOut_7_33[20] , 
        \wRegOut_7_33[19] , \wRegOut_7_33[18] , \wRegOut_7_33[17] , 
        \wRegOut_7_33[16] , \wRegOut_7_33[15] , \wRegOut_7_33[14] , 
        \wRegOut_7_33[13] , \wRegOut_7_33[12] , \wRegOut_7_33[11] , 
        \wRegOut_7_33[10] , \wRegOut_7_33[9] , \wRegOut_7_33[8] , 
        \wRegOut_7_33[7] , \wRegOut_7_33[6] , \wRegOut_7_33[5] , 
        \wRegOut_7_33[4] , \wRegOut_7_33[3] , \wRegOut_7_33[2] , 
        \wRegOut_7_33[1] , \wRegOut_7_33[0] }), .R_Out({\wRegInTop_7_33[31] , 
        \wRegInTop_7_33[30] , \wRegInTop_7_33[29] , \wRegInTop_7_33[28] , 
        \wRegInTop_7_33[27] , \wRegInTop_7_33[26] , \wRegInTop_7_33[25] , 
        \wRegInTop_7_33[24] , \wRegInTop_7_33[23] , \wRegInTop_7_33[22] , 
        \wRegInTop_7_33[21] , \wRegInTop_7_33[20] , \wRegInTop_7_33[19] , 
        \wRegInTop_7_33[18] , \wRegInTop_7_33[17] , \wRegInTop_7_33[16] , 
        \wRegInTop_7_33[15] , \wRegInTop_7_33[14] , \wRegInTop_7_33[13] , 
        \wRegInTop_7_33[12] , \wRegInTop_7_33[11] , \wRegInTop_7_33[10] , 
        \wRegInTop_7_33[9] , \wRegInTop_7_33[8] , \wRegInTop_7_33[7] , 
        \wRegInTop_7_33[6] , \wRegInTop_7_33[5] , \wRegInTop_7_33[4] , 
        \wRegInTop_7_33[3] , \wRegInTop_7_33[2] , \wRegInTop_7_33[1] , 
        \wRegInTop_7_33[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_50 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink114[31] , \ScanLink114[30] , \ScanLink114[29] , 
        \ScanLink114[28] , \ScanLink114[27] , \ScanLink114[26] , 
        \ScanLink114[25] , \ScanLink114[24] , \ScanLink114[23] , 
        \ScanLink114[22] , \ScanLink114[21] , \ScanLink114[20] , 
        \ScanLink114[19] , \ScanLink114[18] , \ScanLink114[17] , 
        \ScanLink114[16] , \ScanLink114[15] , \ScanLink114[14] , 
        \ScanLink114[13] , \ScanLink114[12] , \ScanLink114[11] , 
        \ScanLink114[10] , \ScanLink114[9] , \ScanLink114[8] , 
        \ScanLink114[7] , \ScanLink114[6] , \ScanLink114[5] , \ScanLink114[4] , 
        \ScanLink114[3] , \ScanLink114[2] , \ScanLink114[1] , \ScanLink114[0] 
        }), .ScanOut({\ScanLink113[31] , \ScanLink113[30] , \ScanLink113[29] , 
        \ScanLink113[28] , \ScanLink113[27] , \ScanLink113[26] , 
        \ScanLink113[25] , \ScanLink113[24] , \ScanLink113[23] , 
        \ScanLink113[22] , \ScanLink113[21] , \ScanLink113[20] , 
        \ScanLink113[19] , \ScanLink113[18] , \ScanLink113[17] , 
        \ScanLink113[16] , \ScanLink113[15] , \ScanLink113[14] , 
        \ScanLink113[13] , \ScanLink113[12] , \ScanLink113[11] , 
        \ScanLink113[10] , \ScanLink113[9] , \ScanLink113[8] , 
        \ScanLink113[7] , \ScanLink113[6] , \ScanLink113[5] , \ScanLink113[4] , 
        \ScanLink113[3] , \ScanLink113[2] , \ScanLink113[1] , \ScanLink113[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_50[31] , 
        \wRegOut_6_50[30] , \wRegOut_6_50[29] , \wRegOut_6_50[28] , 
        \wRegOut_6_50[27] , \wRegOut_6_50[26] , \wRegOut_6_50[25] , 
        \wRegOut_6_50[24] , \wRegOut_6_50[23] , \wRegOut_6_50[22] , 
        \wRegOut_6_50[21] , \wRegOut_6_50[20] , \wRegOut_6_50[19] , 
        \wRegOut_6_50[18] , \wRegOut_6_50[17] , \wRegOut_6_50[16] , 
        \wRegOut_6_50[15] , \wRegOut_6_50[14] , \wRegOut_6_50[13] , 
        \wRegOut_6_50[12] , \wRegOut_6_50[11] , \wRegOut_6_50[10] , 
        \wRegOut_6_50[9] , \wRegOut_6_50[8] , \wRegOut_6_50[7] , 
        \wRegOut_6_50[6] , \wRegOut_6_50[5] , \wRegOut_6_50[4] , 
        \wRegOut_6_50[3] , \wRegOut_6_50[2] , \wRegOut_6_50[1] , 
        \wRegOut_6_50[0] }), .Enable1(\wRegEnTop_6_50[0] ), .Enable2(
        \wRegEnBot_6_50[0] ), .In1({\wRegInTop_6_50[31] , \wRegInTop_6_50[30] , 
        \wRegInTop_6_50[29] , \wRegInTop_6_50[28] , \wRegInTop_6_50[27] , 
        \wRegInTop_6_50[26] , \wRegInTop_6_50[25] , \wRegInTop_6_50[24] , 
        \wRegInTop_6_50[23] , \wRegInTop_6_50[22] , \wRegInTop_6_50[21] , 
        \wRegInTop_6_50[20] , \wRegInTop_6_50[19] , \wRegInTop_6_50[18] , 
        \wRegInTop_6_50[17] , \wRegInTop_6_50[16] , \wRegInTop_6_50[15] , 
        \wRegInTop_6_50[14] , \wRegInTop_6_50[13] , \wRegInTop_6_50[12] , 
        \wRegInTop_6_50[11] , \wRegInTop_6_50[10] , \wRegInTop_6_50[9] , 
        \wRegInTop_6_50[8] , \wRegInTop_6_50[7] , \wRegInTop_6_50[6] , 
        \wRegInTop_6_50[5] , \wRegInTop_6_50[4] , \wRegInTop_6_50[3] , 
        \wRegInTop_6_50[2] , \wRegInTop_6_50[1] , \wRegInTop_6_50[0] }), .In2(
        {\wRegInBot_6_50[31] , \wRegInBot_6_50[30] , \wRegInBot_6_50[29] , 
        \wRegInBot_6_50[28] , \wRegInBot_6_50[27] , \wRegInBot_6_50[26] , 
        \wRegInBot_6_50[25] , \wRegInBot_6_50[24] , \wRegInBot_6_50[23] , 
        \wRegInBot_6_50[22] , \wRegInBot_6_50[21] , \wRegInBot_6_50[20] , 
        \wRegInBot_6_50[19] , \wRegInBot_6_50[18] , \wRegInBot_6_50[17] , 
        \wRegInBot_6_50[16] , \wRegInBot_6_50[15] , \wRegInBot_6_50[14] , 
        \wRegInBot_6_50[13] , \wRegInBot_6_50[12] , \wRegInBot_6_50[11] , 
        \wRegInBot_6_50[10] , \wRegInBot_6_50[9] , \wRegInBot_6_50[8] , 
        \wRegInBot_6_50[7] , \wRegInBot_6_50[6] , \wRegInBot_6_50[5] , 
        \wRegInBot_6_50[4] , \wRegInBot_6_50[3] , \wRegInBot_6_50[2] , 
        \wRegInBot_6_50[1] , \wRegInBot_6_50[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_24 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink152[31] , \ScanLink152[30] , \ScanLink152[29] , 
        \ScanLink152[28] , \ScanLink152[27] , \ScanLink152[26] , 
        \ScanLink152[25] , \ScanLink152[24] , \ScanLink152[23] , 
        \ScanLink152[22] , \ScanLink152[21] , \ScanLink152[20] , 
        \ScanLink152[19] , \ScanLink152[18] , \ScanLink152[17] , 
        \ScanLink152[16] , \ScanLink152[15] , \ScanLink152[14] , 
        \ScanLink152[13] , \ScanLink152[12] , \ScanLink152[11] , 
        \ScanLink152[10] , \ScanLink152[9] , \ScanLink152[8] , 
        \ScanLink152[7] , \ScanLink152[6] , \ScanLink152[5] , \ScanLink152[4] , 
        \ScanLink152[3] , \ScanLink152[2] , \ScanLink152[1] , \ScanLink152[0] 
        }), .ScanOut({\ScanLink151[31] , \ScanLink151[30] , \ScanLink151[29] , 
        \ScanLink151[28] , \ScanLink151[27] , \ScanLink151[26] , 
        \ScanLink151[25] , \ScanLink151[24] , \ScanLink151[23] , 
        \ScanLink151[22] , \ScanLink151[21] , \ScanLink151[20] , 
        \ScanLink151[19] , \ScanLink151[18] , \ScanLink151[17] , 
        \ScanLink151[16] , \ScanLink151[15] , \ScanLink151[14] , 
        \ScanLink151[13] , \ScanLink151[12] , \ScanLink151[11] , 
        \ScanLink151[10] , \ScanLink151[9] , \ScanLink151[8] , 
        \ScanLink151[7] , \ScanLink151[6] , \ScanLink151[5] , \ScanLink151[4] , 
        \ScanLink151[3] , \ScanLink151[2] , \ScanLink151[1] , \ScanLink151[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_24[31] , 
        \wRegOut_7_24[30] , \wRegOut_7_24[29] , \wRegOut_7_24[28] , 
        \wRegOut_7_24[27] , \wRegOut_7_24[26] , \wRegOut_7_24[25] , 
        \wRegOut_7_24[24] , \wRegOut_7_24[23] , \wRegOut_7_24[22] , 
        \wRegOut_7_24[21] , \wRegOut_7_24[20] , \wRegOut_7_24[19] , 
        \wRegOut_7_24[18] , \wRegOut_7_24[17] , \wRegOut_7_24[16] , 
        \wRegOut_7_24[15] , \wRegOut_7_24[14] , \wRegOut_7_24[13] , 
        \wRegOut_7_24[12] , \wRegOut_7_24[11] , \wRegOut_7_24[10] , 
        \wRegOut_7_24[9] , \wRegOut_7_24[8] , \wRegOut_7_24[7] , 
        \wRegOut_7_24[6] , \wRegOut_7_24[5] , \wRegOut_7_24[4] , 
        \wRegOut_7_24[3] , \wRegOut_7_24[2] , \wRegOut_7_24[1] , 
        \wRegOut_7_24[0] }), .Enable1(\wRegEnTop_7_24[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_24[31] , \wRegInTop_7_24[30] , \wRegInTop_7_24[29] , 
        \wRegInTop_7_24[28] , \wRegInTop_7_24[27] , \wRegInTop_7_24[26] , 
        \wRegInTop_7_24[25] , \wRegInTop_7_24[24] , \wRegInTop_7_24[23] , 
        \wRegInTop_7_24[22] , \wRegInTop_7_24[21] , \wRegInTop_7_24[20] , 
        \wRegInTop_7_24[19] , \wRegInTop_7_24[18] , \wRegInTop_7_24[17] , 
        \wRegInTop_7_24[16] , \wRegInTop_7_24[15] , \wRegInTop_7_24[14] , 
        \wRegInTop_7_24[13] , \wRegInTop_7_24[12] , \wRegInTop_7_24[11] , 
        \wRegInTop_7_24[10] , \wRegInTop_7_24[9] , \wRegInTop_7_24[8] , 
        \wRegInTop_7_24[7] , \wRegInTop_7_24[6] , \wRegInTop_7_24[5] , 
        \wRegInTop_7_24[4] , \wRegInTop_7_24[3] , \wRegInTop_7_24[2] , 
        \wRegInTop_7_24[1] , \wRegInTop_7_24[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_88 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink216[31] , \ScanLink216[30] , \ScanLink216[29] , 
        \ScanLink216[28] , \ScanLink216[27] , \ScanLink216[26] , 
        \ScanLink216[25] , \ScanLink216[24] , \ScanLink216[23] , 
        \ScanLink216[22] , \ScanLink216[21] , \ScanLink216[20] , 
        \ScanLink216[19] , \ScanLink216[18] , \ScanLink216[17] , 
        \ScanLink216[16] , \ScanLink216[15] , \ScanLink216[14] , 
        \ScanLink216[13] , \ScanLink216[12] , \ScanLink216[11] , 
        \ScanLink216[10] , \ScanLink216[9] , \ScanLink216[8] , 
        \ScanLink216[7] , \ScanLink216[6] , \ScanLink216[5] , \ScanLink216[4] , 
        \ScanLink216[3] , \ScanLink216[2] , \ScanLink216[1] , \ScanLink216[0] 
        }), .ScanOut({\ScanLink215[31] , \ScanLink215[30] , \ScanLink215[29] , 
        \ScanLink215[28] , \ScanLink215[27] , \ScanLink215[26] , 
        \ScanLink215[25] , \ScanLink215[24] , \ScanLink215[23] , 
        \ScanLink215[22] , \ScanLink215[21] , \ScanLink215[20] , 
        \ScanLink215[19] , \ScanLink215[18] , \ScanLink215[17] , 
        \ScanLink215[16] , \ScanLink215[15] , \ScanLink215[14] , 
        \ScanLink215[13] , \ScanLink215[12] , \ScanLink215[11] , 
        \ScanLink215[10] , \ScanLink215[9] , \ScanLink215[8] , 
        \ScanLink215[7] , \ScanLink215[6] , \ScanLink215[5] , \ScanLink215[4] , 
        \ScanLink215[3] , \ScanLink215[2] , \ScanLink215[1] , \ScanLink215[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_88[31] , 
        \wRegOut_7_88[30] , \wRegOut_7_88[29] , \wRegOut_7_88[28] , 
        \wRegOut_7_88[27] , \wRegOut_7_88[26] , \wRegOut_7_88[25] , 
        \wRegOut_7_88[24] , \wRegOut_7_88[23] , \wRegOut_7_88[22] , 
        \wRegOut_7_88[21] , \wRegOut_7_88[20] , \wRegOut_7_88[19] , 
        \wRegOut_7_88[18] , \wRegOut_7_88[17] , \wRegOut_7_88[16] , 
        \wRegOut_7_88[15] , \wRegOut_7_88[14] , \wRegOut_7_88[13] , 
        \wRegOut_7_88[12] , \wRegOut_7_88[11] , \wRegOut_7_88[10] , 
        \wRegOut_7_88[9] , \wRegOut_7_88[8] , \wRegOut_7_88[7] , 
        \wRegOut_7_88[6] , \wRegOut_7_88[5] , \wRegOut_7_88[4] , 
        \wRegOut_7_88[3] , \wRegOut_7_88[2] , \wRegOut_7_88[1] , 
        \wRegOut_7_88[0] }), .Enable1(\wRegEnTop_7_88[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_88[31] , \wRegInTop_7_88[30] , \wRegInTop_7_88[29] , 
        \wRegInTop_7_88[28] , \wRegInTop_7_88[27] , \wRegInTop_7_88[26] , 
        \wRegInTop_7_88[25] , \wRegInTop_7_88[24] , \wRegInTop_7_88[23] , 
        \wRegInTop_7_88[22] , \wRegInTop_7_88[21] , \wRegInTop_7_88[20] , 
        \wRegInTop_7_88[19] , \wRegInTop_7_88[18] , \wRegInTop_7_88[17] , 
        \wRegInTop_7_88[16] , \wRegInTop_7_88[15] , \wRegInTop_7_88[14] , 
        \wRegInTop_7_88[13] , \wRegInTop_7_88[12] , \wRegInTop_7_88[11] , 
        \wRegInTop_7_88[10] , \wRegInTop_7_88[9] , \wRegInTop_7_88[8] , 
        \wRegInTop_7_88[7] , \wRegInTop_7_88[6] , \wRegInTop_7_88[5] , 
        \wRegInTop_7_88[4] , \wRegInTop_7_88[3] , \wRegInTop_7_88[2] , 
        \wRegInTop_7_88[1] , \wRegInTop_7_88[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink47[31] , \ScanLink47[30] , \ScanLink47[29] , 
        \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , \ScanLink47[25] , 
        \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , \ScanLink47[21] , 
        \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , \ScanLink47[17] , 
        \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , \ScanLink47[13] , 
        \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , \ScanLink47[9] , 
        \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , \ScanLink47[5] , 
        \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , \ScanLink47[1] , 
        \ScanLink47[0] }), .ScanOut({\ScanLink46[31] , \ScanLink46[30] , 
        \ScanLink46[29] , \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , 
        \ScanLink46[25] , \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , 
        \ScanLink46[21] , \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , 
        \ScanLink46[17] , \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , 
        \ScanLink46[13] , \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , 
        \ScanLink46[9] , \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , 
        \ScanLink46[5] , \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , 
        \ScanLink46[1] , \ScanLink46[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_15[31] , \wRegOut_5_15[30] , 
        \wRegOut_5_15[29] , \wRegOut_5_15[28] , \wRegOut_5_15[27] , 
        \wRegOut_5_15[26] , \wRegOut_5_15[25] , \wRegOut_5_15[24] , 
        \wRegOut_5_15[23] , \wRegOut_5_15[22] , \wRegOut_5_15[21] , 
        \wRegOut_5_15[20] , \wRegOut_5_15[19] , \wRegOut_5_15[18] , 
        \wRegOut_5_15[17] , \wRegOut_5_15[16] , \wRegOut_5_15[15] , 
        \wRegOut_5_15[14] , \wRegOut_5_15[13] , \wRegOut_5_15[12] , 
        \wRegOut_5_15[11] , \wRegOut_5_15[10] , \wRegOut_5_15[9] , 
        \wRegOut_5_15[8] , \wRegOut_5_15[7] , \wRegOut_5_15[6] , 
        \wRegOut_5_15[5] , \wRegOut_5_15[4] , \wRegOut_5_15[3] , 
        \wRegOut_5_15[2] , \wRegOut_5_15[1] , \wRegOut_5_15[0] }), .Enable1(
        \wRegEnTop_5_15[0] ), .Enable2(\wRegEnBot_5_15[0] ), .In1({
        \wRegInTop_5_15[31] , \wRegInTop_5_15[30] , \wRegInTop_5_15[29] , 
        \wRegInTop_5_15[28] , \wRegInTop_5_15[27] , \wRegInTop_5_15[26] , 
        \wRegInTop_5_15[25] , \wRegInTop_5_15[24] , \wRegInTop_5_15[23] , 
        \wRegInTop_5_15[22] , \wRegInTop_5_15[21] , \wRegInTop_5_15[20] , 
        \wRegInTop_5_15[19] , \wRegInTop_5_15[18] , \wRegInTop_5_15[17] , 
        \wRegInTop_5_15[16] , \wRegInTop_5_15[15] , \wRegInTop_5_15[14] , 
        \wRegInTop_5_15[13] , \wRegInTop_5_15[12] , \wRegInTop_5_15[11] , 
        \wRegInTop_5_15[10] , \wRegInTop_5_15[9] , \wRegInTop_5_15[8] , 
        \wRegInTop_5_15[7] , \wRegInTop_5_15[6] , \wRegInTop_5_15[5] , 
        \wRegInTop_5_15[4] , \wRegInTop_5_15[3] , \wRegInTop_5_15[2] , 
        \wRegInTop_5_15[1] , \wRegInTop_5_15[0] }), .In2({\wRegInBot_5_15[31] , 
        \wRegInBot_5_15[30] , \wRegInBot_5_15[29] , \wRegInBot_5_15[28] , 
        \wRegInBot_5_15[27] , \wRegInBot_5_15[26] , \wRegInBot_5_15[25] , 
        \wRegInBot_5_15[24] , \wRegInBot_5_15[23] , \wRegInBot_5_15[22] , 
        \wRegInBot_5_15[21] , \wRegInBot_5_15[20] , \wRegInBot_5_15[19] , 
        \wRegInBot_5_15[18] , \wRegInBot_5_15[17] , \wRegInBot_5_15[16] , 
        \wRegInBot_5_15[15] , \wRegInBot_5_15[14] , \wRegInBot_5_15[13] , 
        \wRegInBot_5_15[12] , \wRegInBot_5_15[11] , \wRegInBot_5_15[10] , 
        \wRegInBot_5_15[9] , \wRegInBot_5_15[8] , \wRegInBot_5_15[7] , 
        \wRegInBot_5_15[6] , \wRegInBot_5_15[5] , \wRegInBot_5_15[4] , 
        \wRegInBot_5_15[3] , \wRegInBot_5_15[2] , \wRegInBot_5_15[1] , 
        \wRegInBot_5_15[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_25 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink89[31] , \ScanLink89[30] , \ScanLink89[29] , 
        \ScanLink89[28] , \ScanLink89[27] , \ScanLink89[26] , \ScanLink89[25] , 
        \ScanLink89[24] , \ScanLink89[23] , \ScanLink89[22] , \ScanLink89[21] , 
        \ScanLink89[20] , \ScanLink89[19] , \ScanLink89[18] , \ScanLink89[17] , 
        \ScanLink89[16] , \ScanLink89[15] , \ScanLink89[14] , \ScanLink89[13] , 
        \ScanLink89[12] , \ScanLink89[11] , \ScanLink89[10] , \ScanLink89[9] , 
        \ScanLink89[8] , \ScanLink89[7] , \ScanLink89[6] , \ScanLink89[5] , 
        \ScanLink89[4] , \ScanLink89[3] , \ScanLink89[2] , \ScanLink89[1] , 
        \ScanLink89[0] }), .ScanOut({\ScanLink88[31] , \ScanLink88[30] , 
        \ScanLink88[29] , \ScanLink88[28] , \ScanLink88[27] , \ScanLink88[26] , 
        \ScanLink88[25] , \ScanLink88[24] , \ScanLink88[23] , \ScanLink88[22] , 
        \ScanLink88[21] , \ScanLink88[20] , \ScanLink88[19] , \ScanLink88[18] , 
        \ScanLink88[17] , \ScanLink88[16] , \ScanLink88[15] , \ScanLink88[14] , 
        \ScanLink88[13] , \ScanLink88[12] , \ScanLink88[11] , \ScanLink88[10] , 
        \ScanLink88[9] , \ScanLink88[8] , \ScanLink88[7] , \ScanLink88[6] , 
        \ScanLink88[5] , \ScanLink88[4] , \ScanLink88[3] , \ScanLink88[2] , 
        \ScanLink88[1] , \ScanLink88[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_25[31] , \wRegOut_6_25[30] , 
        \wRegOut_6_25[29] , \wRegOut_6_25[28] , \wRegOut_6_25[27] , 
        \wRegOut_6_25[26] , \wRegOut_6_25[25] , \wRegOut_6_25[24] , 
        \wRegOut_6_25[23] , \wRegOut_6_25[22] , \wRegOut_6_25[21] , 
        \wRegOut_6_25[20] , \wRegOut_6_25[19] , \wRegOut_6_25[18] , 
        \wRegOut_6_25[17] , \wRegOut_6_25[16] , \wRegOut_6_25[15] , 
        \wRegOut_6_25[14] , \wRegOut_6_25[13] , \wRegOut_6_25[12] , 
        \wRegOut_6_25[11] , \wRegOut_6_25[10] , \wRegOut_6_25[9] , 
        \wRegOut_6_25[8] , \wRegOut_6_25[7] , \wRegOut_6_25[6] , 
        \wRegOut_6_25[5] , \wRegOut_6_25[4] , \wRegOut_6_25[3] , 
        \wRegOut_6_25[2] , \wRegOut_6_25[1] , \wRegOut_6_25[0] }), .Enable1(
        \wRegEnTop_6_25[0] ), .Enable2(\wRegEnBot_6_25[0] ), .In1({
        \wRegInTop_6_25[31] , \wRegInTop_6_25[30] , \wRegInTop_6_25[29] , 
        \wRegInTop_6_25[28] , \wRegInTop_6_25[27] , \wRegInTop_6_25[26] , 
        \wRegInTop_6_25[25] , \wRegInTop_6_25[24] , \wRegInTop_6_25[23] , 
        \wRegInTop_6_25[22] , \wRegInTop_6_25[21] , \wRegInTop_6_25[20] , 
        \wRegInTop_6_25[19] , \wRegInTop_6_25[18] , \wRegInTop_6_25[17] , 
        \wRegInTop_6_25[16] , \wRegInTop_6_25[15] , \wRegInTop_6_25[14] , 
        \wRegInTop_6_25[13] , \wRegInTop_6_25[12] , \wRegInTop_6_25[11] , 
        \wRegInTop_6_25[10] , \wRegInTop_6_25[9] , \wRegInTop_6_25[8] , 
        \wRegInTop_6_25[7] , \wRegInTop_6_25[6] , \wRegInTop_6_25[5] , 
        \wRegInTop_6_25[4] , \wRegInTop_6_25[3] , \wRegInTop_6_25[2] , 
        \wRegInTop_6_25[1] , \wRegInTop_6_25[0] }), .In2({\wRegInBot_6_25[31] , 
        \wRegInBot_6_25[30] , \wRegInBot_6_25[29] , \wRegInBot_6_25[28] , 
        \wRegInBot_6_25[27] , \wRegInBot_6_25[26] , \wRegInBot_6_25[25] , 
        \wRegInBot_6_25[24] , \wRegInBot_6_25[23] , \wRegInBot_6_25[22] , 
        \wRegInBot_6_25[21] , \wRegInBot_6_25[20] , \wRegInBot_6_25[19] , 
        \wRegInBot_6_25[18] , \wRegInBot_6_25[17] , \wRegInBot_6_25[16] , 
        \wRegInBot_6_25[15] , \wRegInBot_6_25[14] , \wRegInBot_6_25[13] , 
        \wRegInBot_6_25[12] , \wRegInBot_6_25[11] , \wRegInBot_6_25[10] , 
        \wRegInBot_6_25[9] , \wRegInBot_6_25[8] , \wRegInBot_6_25[7] , 
        \wRegInBot_6_25[6] , \wRegInBot_6_25[5] , \wRegInBot_6_25[4] , 
        \wRegInBot_6_25[3] , \wRegInBot_6_25[2] , \wRegInBot_6_25[1] , 
        \wRegInBot_6_25[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_18 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink146[31] , \ScanLink146[30] , \ScanLink146[29] , 
        \ScanLink146[28] , \ScanLink146[27] , \ScanLink146[26] , 
        \ScanLink146[25] , \ScanLink146[24] , \ScanLink146[23] , 
        \ScanLink146[22] , \ScanLink146[21] , \ScanLink146[20] , 
        \ScanLink146[19] , \ScanLink146[18] , \ScanLink146[17] , 
        \ScanLink146[16] , \ScanLink146[15] , \ScanLink146[14] , 
        \ScanLink146[13] , \ScanLink146[12] , \ScanLink146[11] , 
        \ScanLink146[10] , \ScanLink146[9] , \ScanLink146[8] , 
        \ScanLink146[7] , \ScanLink146[6] , \ScanLink146[5] , \ScanLink146[4] , 
        \ScanLink146[3] , \ScanLink146[2] , \ScanLink146[1] , \ScanLink146[0] 
        }), .ScanOut({\ScanLink145[31] , \ScanLink145[30] , \ScanLink145[29] , 
        \ScanLink145[28] , \ScanLink145[27] , \ScanLink145[26] , 
        \ScanLink145[25] , \ScanLink145[24] , \ScanLink145[23] , 
        \ScanLink145[22] , \ScanLink145[21] , \ScanLink145[20] , 
        \ScanLink145[19] , \ScanLink145[18] , \ScanLink145[17] , 
        \ScanLink145[16] , \ScanLink145[15] , \ScanLink145[14] , 
        \ScanLink145[13] , \ScanLink145[12] , \ScanLink145[11] , 
        \ScanLink145[10] , \ScanLink145[9] , \ScanLink145[8] , 
        \ScanLink145[7] , \ScanLink145[6] , \ScanLink145[5] , \ScanLink145[4] , 
        \ScanLink145[3] , \ScanLink145[2] , \ScanLink145[1] , \ScanLink145[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_18[31] , 
        \wRegOut_7_18[30] , \wRegOut_7_18[29] , \wRegOut_7_18[28] , 
        \wRegOut_7_18[27] , \wRegOut_7_18[26] , \wRegOut_7_18[25] , 
        \wRegOut_7_18[24] , \wRegOut_7_18[23] , \wRegOut_7_18[22] , 
        \wRegOut_7_18[21] , \wRegOut_7_18[20] , \wRegOut_7_18[19] , 
        \wRegOut_7_18[18] , \wRegOut_7_18[17] , \wRegOut_7_18[16] , 
        \wRegOut_7_18[15] , \wRegOut_7_18[14] , \wRegOut_7_18[13] , 
        \wRegOut_7_18[12] , \wRegOut_7_18[11] , \wRegOut_7_18[10] , 
        \wRegOut_7_18[9] , \wRegOut_7_18[8] , \wRegOut_7_18[7] , 
        \wRegOut_7_18[6] , \wRegOut_7_18[5] , \wRegOut_7_18[4] , 
        \wRegOut_7_18[3] , \wRegOut_7_18[2] , \wRegOut_7_18[1] , 
        \wRegOut_7_18[0] }), .Enable1(\wRegEnTop_7_18[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_18[31] , \wRegInTop_7_18[30] , \wRegInTop_7_18[29] , 
        \wRegInTop_7_18[28] , \wRegInTop_7_18[27] , \wRegInTop_7_18[26] , 
        \wRegInTop_7_18[25] , \wRegInTop_7_18[24] , \wRegInTop_7_18[23] , 
        \wRegInTop_7_18[22] , \wRegInTop_7_18[21] , \wRegInTop_7_18[20] , 
        \wRegInTop_7_18[19] , \wRegInTop_7_18[18] , \wRegInTop_7_18[17] , 
        \wRegInTop_7_18[16] , \wRegInTop_7_18[15] , \wRegInTop_7_18[14] , 
        \wRegInTop_7_18[13] , \wRegInTop_7_18[12] , \wRegInTop_7_18[11] , 
        \wRegInTop_7_18[10] , \wRegInTop_7_18[9] , \wRegInTop_7_18[8] , 
        \wRegInTop_7_18[7] , \wRegInTop_7_18[6] , \wRegInTop_7_18[5] , 
        \wRegInTop_7_18[4] , \wRegInTop_7_18[3] , \wRegInTop_7_18[2] , 
        \wRegInTop_7_18[1] , \wRegInTop_7_18[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_117 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink245[31] , \ScanLink245[30] , \ScanLink245[29] , 
        \ScanLink245[28] , \ScanLink245[27] , \ScanLink245[26] , 
        \ScanLink245[25] , \ScanLink245[24] , \ScanLink245[23] , 
        \ScanLink245[22] , \ScanLink245[21] , \ScanLink245[20] , 
        \ScanLink245[19] , \ScanLink245[18] , \ScanLink245[17] , 
        \ScanLink245[16] , \ScanLink245[15] , \ScanLink245[14] , 
        \ScanLink245[13] , \ScanLink245[12] , \ScanLink245[11] , 
        \ScanLink245[10] , \ScanLink245[9] , \ScanLink245[8] , 
        \ScanLink245[7] , \ScanLink245[6] , \ScanLink245[5] , \ScanLink245[4] , 
        \ScanLink245[3] , \ScanLink245[2] , \ScanLink245[1] , \ScanLink245[0] 
        }), .ScanOut({\ScanLink244[31] , \ScanLink244[30] , \ScanLink244[29] , 
        \ScanLink244[28] , \ScanLink244[27] , \ScanLink244[26] , 
        \ScanLink244[25] , \ScanLink244[24] , \ScanLink244[23] , 
        \ScanLink244[22] , \ScanLink244[21] , \ScanLink244[20] , 
        \ScanLink244[19] , \ScanLink244[18] , \ScanLink244[17] , 
        \ScanLink244[16] , \ScanLink244[15] , \ScanLink244[14] , 
        \ScanLink244[13] , \ScanLink244[12] , \ScanLink244[11] , 
        \ScanLink244[10] , \ScanLink244[9] , \ScanLink244[8] , 
        \ScanLink244[7] , \ScanLink244[6] , \ScanLink244[5] , \ScanLink244[4] , 
        \ScanLink244[3] , \ScanLink244[2] , \ScanLink244[1] , \ScanLink244[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_117[31] , 
        \wRegOut_7_117[30] , \wRegOut_7_117[29] , \wRegOut_7_117[28] , 
        \wRegOut_7_117[27] , \wRegOut_7_117[26] , \wRegOut_7_117[25] , 
        \wRegOut_7_117[24] , \wRegOut_7_117[23] , \wRegOut_7_117[22] , 
        \wRegOut_7_117[21] , \wRegOut_7_117[20] , \wRegOut_7_117[19] , 
        \wRegOut_7_117[18] , \wRegOut_7_117[17] , \wRegOut_7_117[16] , 
        \wRegOut_7_117[15] , \wRegOut_7_117[14] , \wRegOut_7_117[13] , 
        \wRegOut_7_117[12] , \wRegOut_7_117[11] , \wRegOut_7_117[10] , 
        \wRegOut_7_117[9] , \wRegOut_7_117[8] , \wRegOut_7_117[7] , 
        \wRegOut_7_117[6] , \wRegOut_7_117[5] , \wRegOut_7_117[4] , 
        \wRegOut_7_117[3] , \wRegOut_7_117[2] , \wRegOut_7_117[1] , 
        \wRegOut_7_117[0] }), .Enable1(\wRegEnTop_7_117[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_117[31] , \wRegInTop_7_117[30] , 
        \wRegInTop_7_117[29] , \wRegInTop_7_117[28] , \wRegInTop_7_117[27] , 
        \wRegInTop_7_117[26] , \wRegInTop_7_117[25] , \wRegInTop_7_117[24] , 
        \wRegInTop_7_117[23] , \wRegInTop_7_117[22] , \wRegInTop_7_117[21] , 
        \wRegInTop_7_117[20] , \wRegInTop_7_117[19] , \wRegInTop_7_117[18] , 
        \wRegInTop_7_117[17] , \wRegInTop_7_117[16] , \wRegInTop_7_117[15] , 
        \wRegInTop_7_117[14] , \wRegInTop_7_117[13] , \wRegInTop_7_117[12] , 
        \wRegInTop_7_117[11] , \wRegInTop_7_117[10] , \wRegInTop_7_117[9] , 
        \wRegInTop_7_117[8] , \wRegInTop_7_117[7] , \wRegInTop_7_117[6] , 
        \wRegInTop_7_117[5] , \wRegInTop_7_117[4] , \wRegInTop_7_117[3] , 
        \wRegInTop_7_117[2] , \wRegInTop_7_117[1] , \wRegInTop_7_117[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_2[0] ), .P_In({\wRegOut_4_2[31] , 
        \wRegOut_4_2[30] , \wRegOut_4_2[29] , \wRegOut_4_2[28] , 
        \wRegOut_4_2[27] , \wRegOut_4_2[26] , \wRegOut_4_2[25] , 
        \wRegOut_4_2[24] , \wRegOut_4_2[23] , \wRegOut_4_2[22] , 
        \wRegOut_4_2[21] , \wRegOut_4_2[20] , \wRegOut_4_2[19] , 
        \wRegOut_4_2[18] , \wRegOut_4_2[17] , \wRegOut_4_2[16] , 
        \wRegOut_4_2[15] , \wRegOut_4_2[14] , \wRegOut_4_2[13] , 
        \wRegOut_4_2[12] , \wRegOut_4_2[11] , \wRegOut_4_2[10] , 
        \wRegOut_4_2[9] , \wRegOut_4_2[8] , \wRegOut_4_2[7] , \wRegOut_4_2[6] , 
        \wRegOut_4_2[5] , \wRegOut_4_2[4] , \wRegOut_4_2[3] , \wRegOut_4_2[2] , 
        \wRegOut_4_2[1] , \wRegOut_4_2[0] }), .P_Out({\wRegInBot_4_2[31] , 
        \wRegInBot_4_2[30] , \wRegInBot_4_2[29] , \wRegInBot_4_2[28] , 
        \wRegInBot_4_2[27] , \wRegInBot_4_2[26] , \wRegInBot_4_2[25] , 
        \wRegInBot_4_2[24] , \wRegInBot_4_2[23] , \wRegInBot_4_2[22] , 
        \wRegInBot_4_2[21] , \wRegInBot_4_2[20] , \wRegInBot_4_2[19] , 
        \wRegInBot_4_2[18] , \wRegInBot_4_2[17] , \wRegInBot_4_2[16] , 
        \wRegInBot_4_2[15] , \wRegInBot_4_2[14] , \wRegInBot_4_2[13] , 
        \wRegInBot_4_2[12] , \wRegInBot_4_2[11] , \wRegInBot_4_2[10] , 
        \wRegInBot_4_2[9] , \wRegInBot_4_2[8] , \wRegInBot_4_2[7] , 
        \wRegInBot_4_2[6] , \wRegInBot_4_2[5] , \wRegInBot_4_2[4] , 
        \wRegInBot_4_2[3] , \wRegInBot_4_2[2] , \wRegInBot_4_2[1] , 
        \wRegInBot_4_2[0] }), .L_WR(\wRegEnTop_5_4[0] ), .L_In({
        \wRegOut_5_4[31] , \wRegOut_5_4[30] , \wRegOut_5_4[29] , 
        \wRegOut_5_4[28] , \wRegOut_5_4[27] , \wRegOut_5_4[26] , 
        \wRegOut_5_4[25] , \wRegOut_5_4[24] , \wRegOut_5_4[23] , 
        \wRegOut_5_4[22] , \wRegOut_5_4[21] , \wRegOut_5_4[20] , 
        \wRegOut_5_4[19] , \wRegOut_5_4[18] , \wRegOut_5_4[17] , 
        \wRegOut_5_4[16] , \wRegOut_5_4[15] , \wRegOut_5_4[14] , 
        \wRegOut_5_4[13] , \wRegOut_5_4[12] , \wRegOut_5_4[11] , 
        \wRegOut_5_4[10] , \wRegOut_5_4[9] , \wRegOut_5_4[8] , 
        \wRegOut_5_4[7] , \wRegOut_5_4[6] , \wRegOut_5_4[5] , \wRegOut_5_4[4] , 
        \wRegOut_5_4[3] , \wRegOut_5_4[2] , \wRegOut_5_4[1] , \wRegOut_5_4[0] 
        }), .L_Out({\wRegInTop_5_4[31] , \wRegInTop_5_4[30] , 
        \wRegInTop_5_4[29] , \wRegInTop_5_4[28] , \wRegInTop_5_4[27] , 
        \wRegInTop_5_4[26] , \wRegInTop_5_4[25] , \wRegInTop_5_4[24] , 
        \wRegInTop_5_4[23] , \wRegInTop_5_4[22] , \wRegInTop_5_4[21] , 
        \wRegInTop_5_4[20] , \wRegInTop_5_4[19] , \wRegInTop_5_4[18] , 
        \wRegInTop_5_4[17] , \wRegInTop_5_4[16] , \wRegInTop_5_4[15] , 
        \wRegInTop_5_4[14] , \wRegInTop_5_4[13] , \wRegInTop_5_4[12] , 
        \wRegInTop_5_4[11] , \wRegInTop_5_4[10] , \wRegInTop_5_4[9] , 
        \wRegInTop_5_4[8] , \wRegInTop_5_4[7] , \wRegInTop_5_4[6] , 
        \wRegInTop_5_4[5] , \wRegInTop_5_4[4] , \wRegInTop_5_4[3] , 
        \wRegInTop_5_4[2] , \wRegInTop_5_4[1] , \wRegInTop_5_4[0] }), .R_WR(
        \wRegEnTop_5_5[0] ), .R_In({\wRegOut_5_5[31] , \wRegOut_5_5[30] , 
        \wRegOut_5_5[29] , \wRegOut_5_5[28] , \wRegOut_5_5[27] , 
        \wRegOut_5_5[26] , \wRegOut_5_5[25] , \wRegOut_5_5[24] , 
        \wRegOut_5_5[23] , \wRegOut_5_5[22] , \wRegOut_5_5[21] , 
        \wRegOut_5_5[20] , \wRegOut_5_5[19] , \wRegOut_5_5[18] , 
        \wRegOut_5_5[17] , \wRegOut_5_5[16] , \wRegOut_5_5[15] , 
        \wRegOut_5_5[14] , \wRegOut_5_5[13] , \wRegOut_5_5[12] , 
        \wRegOut_5_5[11] , \wRegOut_5_5[10] , \wRegOut_5_5[9] , 
        \wRegOut_5_5[8] , \wRegOut_5_5[7] , \wRegOut_5_5[6] , \wRegOut_5_5[5] , 
        \wRegOut_5_5[4] , \wRegOut_5_5[3] , \wRegOut_5_5[2] , \wRegOut_5_5[1] , 
        \wRegOut_5_5[0] }), .R_Out({\wRegInTop_5_5[31] , \wRegInTop_5_5[30] , 
        \wRegInTop_5_5[29] , \wRegInTop_5_5[28] , \wRegInTop_5_5[27] , 
        \wRegInTop_5_5[26] , \wRegInTop_5_5[25] , \wRegInTop_5_5[24] , 
        \wRegInTop_5_5[23] , \wRegInTop_5_5[22] , \wRegInTop_5_5[21] , 
        \wRegInTop_5_5[20] , \wRegInTop_5_5[19] , \wRegInTop_5_5[18] , 
        \wRegInTop_5_5[17] , \wRegInTop_5_5[16] , \wRegInTop_5_5[15] , 
        \wRegInTop_5_5[14] , \wRegInTop_5_5[13] , \wRegInTop_5_5[12] , 
        \wRegInTop_5_5[11] , \wRegInTop_5_5[10] , \wRegInTop_5_5[9] , 
        \wRegInTop_5_5[8] , \wRegInTop_5_5[7] , \wRegInTop_5_5[6] , 
        \wRegInTop_5_5[5] , \wRegInTop_5_5[4] , \wRegInTop_5_5[3] , 
        \wRegInTop_5_5[2] , \wRegInTop_5_5[1] , \wRegInTop_5_5[0] }) );
    BHeap_Node_WIDTH32 BHN_6_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_44[0] ), .P_In({\wRegOut_6_44[31] , 
        \wRegOut_6_44[30] , \wRegOut_6_44[29] , \wRegOut_6_44[28] , 
        \wRegOut_6_44[27] , \wRegOut_6_44[26] , \wRegOut_6_44[25] , 
        \wRegOut_6_44[24] , \wRegOut_6_44[23] , \wRegOut_6_44[22] , 
        \wRegOut_6_44[21] , \wRegOut_6_44[20] , \wRegOut_6_44[19] , 
        \wRegOut_6_44[18] , \wRegOut_6_44[17] , \wRegOut_6_44[16] , 
        \wRegOut_6_44[15] , \wRegOut_6_44[14] , \wRegOut_6_44[13] , 
        \wRegOut_6_44[12] , \wRegOut_6_44[11] , \wRegOut_6_44[10] , 
        \wRegOut_6_44[9] , \wRegOut_6_44[8] , \wRegOut_6_44[7] , 
        \wRegOut_6_44[6] , \wRegOut_6_44[5] , \wRegOut_6_44[4] , 
        \wRegOut_6_44[3] , \wRegOut_6_44[2] , \wRegOut_6_44[1] , 
        \wRegOut_6_44[0] }), .P_Out({\wRegInBot_6_44[31] , 
        \wRegInBot_6_44[30] , \wRegInBot_6_44[29] , \wRegInBot_6_44[28] , 
        \wRegInBot_6_44[27] , \wRegInBot_6_44[26] , \wRegInBot_6_44[25] , 
        \wRegInBot_6_44[24] , \wRegInBot_6_44[23] , \wRegInBot_6_44[22] , 
        \wRegInBot_6_44[21] , \wRegInBot_6_44[20] , \wRegInBot_6_44[19] , 
        \wRegInBot_6_44[18] , \wRegInBot_6_44[17] , \wRegInBot_6_44[16] , 
        \wRegInBot_6_44[15] , \wRegInBot_6_44[14] , \wRegInBot_6_44[13] , 
        \wRegInBot_6_44[12] , \wRegInBot_6_44[11] , \wRegInBot_6_44[10] , 
        \wRegInBot_6_44[9] , \wRegInBot_6_44[8] , \wRegInBot_6_44[7] , 
        \wRegInBot_6_44[6] , \wRegInBot_6_44[5] , \wRegInBot_6_44[4] , 
        \wRegInBot_6_44[3] , \wRegInBot_6_44[2] , \wRegInBot_6_44[1] , 
        \wRegInBot_6_44[0] }), .L_WR(\wRegEnTop_7_88[0] ), .L_In({
        \wRegOut_7_88[31] , \wRegOut_7_88[30] , \wRegOut_7_88[29] , 
        \wRegOut_7_88[28] , \wRegOut_7_88[27] , \wRegOut_7_88[26] , 
        \wRegOut_7_88[25] , \wRegOut_7_88[24] , \wRegOut_7_88[23] , 
        \wRegOut_7_88[22] , \wRegOut_7_88[21] , \wRegOut_7_88[20] , 
        \wRegOut_7_88[19] , \wRegOut_7_88[18] , \wRegOut_7_88[17] , 
        \wRegOut_7_88[16] , \wRegOut_7_88[15] , \wRegOut_7_88[14] , 
        \wRegOut_7_88[13] , \wRegOut_7_88[12] , \wRegOut_7_88[11] , 
        \wRegOut_7_88[10] , \wRegOut_7_88[9] , \wRegOut_7_88[8] , 
        \wRegOut_7_88[7] , \wRegOut_7_88[6] , \wRegOut_7_88[5] , 
        \wRegOut_7_88[4] , \wRegOut_7_88[3] , \wRegOut_7_88[2] , 
        \wRegOut_7_88[1] , \wRegOut_7_88[0] }), .L_Out({\wRegInTop_7_88[31] , 
        \wRegInTop_7_88[30] , \wRegInTop_7_88[29] , \wRegInTop_7_88[28] , 
        \wRegInTop_7_88[27] , \wRegInTop_7_88[26] , \wRegInTop_7_88[25] , 
        \wRegInTop_7_88[24] , \wRegInTop_7_88[23] , \wRegInTop_7_88[22] , 
        \wRegInTop_7_88[21] , \wRegInTop_7_88[20] , \wRegInTop_7_88[19] , 
        \wRegInTop_7_88[18] , \wRegInTop_7_88[17] , \wRegInTop_7_88[16] , 
        \wRegInTop_7_88[15] , \wRegInTop_7_88[14] , \wRegInTop_7_88[13] , 
        \wRegInTop_7_88[12] , \wRegInTop_7_88[11] , \wRegInTop_7_88[10] , 
        \wRegInTop_7_88[9] , \wRegInTop_7_88[8] , \wRegInTop_7_88[7] , 
        \wRegInTop_7_88[6] , \wRegInTop_7_88[5] , \wRegInTop_7_88[4] , 
        \wRegInTop_7_88[3] , \wRegInTop_7_88[2] , \wRegInTop_7_88[1] , 
        \wRegInTop_7_88[0] }), .R_WR(\wRegEnTop_7_89[0] ), .R_In({
        \wRegOut_7_89[31] , \wRegOut_7_89[30] , \wRegOut_7_89[29] , 
        \wRegOut_7_89[28] , \wRegOut_7_89[27] , \wRegOut_7_89[26] , 
        \wRegOut_7_89[25] , \wRegOut_7_89[24] , \wRegOut_7_89[23] , 
        \wRegOut_7_89[22] , \wRegOut_7_89[21] , \wRegOut_7_89[20] , 
        \wRegOut_7_89[19] , \wRegOut_7_89[18] , \wRegOut_7_89[17] , 
        \wRegOut_7_89[16] , \wRegOut_7_89[15] , \wRegOut_7_89[14] , 
        \wRegOut_7_89[13] , \wRegOut_7_89[12] , \wRegOut_7_89[11] , 
        \wRegOut_7_89[10] , \wRegOut_7_89[9] , \wRegOut_7_89[8] , 
        \wRegOut_7_89[7] , \wRegOut_7_89[6] , \wRegOut_7_89[5] , 
        \wRegOut_7_89[4] , \wRegOut_7_89[3] , \wRegOut_7_89[2] , 
        \wRegOut_7_89[1] , \wRegOut_7_89[0] }), .R_Out({\wRegInTop_7_89[31] , 
        \wRegInTop_7_89[30] , \wRegInTop_7_89[29] , \wRegInTop_7_89[28] , 
        \wRegInTop_7_89[27] , \wRegInTop_7_89[26] , \wRegInTop_7_89[25] , 
        \wRegInTop_7_89[24] , \wRegInTop_7_89[23] , \wRegInTop_7_89[22] , 
        \wRegInTop_7_89[21] , \wRegInTop_7_89[20] , \wRegInTop_7_89[19] , 
        \wRegInTop_7_89[18] , \wRegInTop_7_89[17] , \wRegInTop_7_89[16] , 
        \wRegInTop_7_89[15] , \wRegInTop_7_89[14] , \wRegInTop_7_89[13] , 
        \wRegInTop_7_89[12] , \wRegInTop_7_89[11] , \wRegInTop_7_89[10] , 
        \wRegInTop_7_89[9] , \wRegInTop_7_89[8] , \wRegInTop_7_89[7] , 
        \wRegInTop_7_89[6] , \wRegInTop_7_89[5] , \wRegInTop_7_89[4] , 
        \wRegInTop_7_89[3] , \wRegInTop_7_89[2] , \wRegInTop_7_89[1] , 
        \wRegInTop_7_89[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_93 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink221[31] , \ScanLink221[30] , \ScanLink221[29] , 
        \ScanLink221[28] , \ScanLink221[27] , \ScanLink221[26] , 
        \ScanLink221[25] , \ScanLink221[24] , \ScanLink221[23] , 
        \ScanLink221[22] , \ScanLink221[21] , \ScanLink221[20] , 
        \ScanLink221[19] , \ScanLink221[18] , \ScanLink221[17] , 
        \ScanLink221[16] , \ScanLink221[15] , \ScanLink221[14] , 
        \ScanLink221[13] , \ScanLink221[12] , \ScanLink221[11] , 
        \ScanLink221[10] , \ScanLink221[9] , \ScanLink221[8] , 
        \ScanLink221[7] , \ScanLink221[6] , \ScanLink221[5] , \ScanLink221[4] , 
        \ScanLink221[3] , \ScanLink221[2] , \ScanLink221[1] , \ScanLink221[0] 
        }), .ScanOut({\ScanLink220[31] , \ScanLink220[30] , \ScanLink220[29] , 
        \ScanLink220[28] , \ScanLink220[27] , \ScanLink220[26] , 
        \ScanLink220[25] , \ScanLink220[24] , \ScanLink220[23] , 
        \ScanLink220[22] , \ScanLink220[21] , \ScanLink220[20] , 
        \ScanLink220[19] , \ScanLink220[18] , \ScanLink220[17] , 
        \ScanLink220[16] , \ScanLink220[15] , \ScanLink220[14] , 
        \ScanLink220[13] , \ScanLink220[12] , \ScanLink220[11] , 
        \ScanLink220[10] , \ScanLink220[9] , \ScanLink220[8] , 
        \ScanLink220[7] , \ScanLink220[6] , \ScanLink220[5] , \ScanLink220[4] , 
        \ScanLink220[3] , \ScanLink220[2] , \ScanLink220[1] , \ScanLink220[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_93[31] , 
        \wRegOut_7_93[30] , \wRegOut_7_93[29] , \wRegOut_7_93[28] , 
        \wRegOut_7_93[27] , \wRegOut_7_93[26] , \wRegOut_7_93[25] , 
        \wRegOut_7_93[24] , \wRegOut_7_93[23] , \wRegOut_7_93[22] , 
        \wRegOut_7_93[21] , \wRegOut_7_93[20] , \wRegOut_7_93[19] , 
        \wRegOut_7_93[18] , \wRegOut_7_93[17] , \wRegOut_7_93[16] , 
        \wRegOut_7_93[15] , \wRegOut_7_93[14] , \wRegOut_7_93[13] , 
        \wRegOut_7_93[12] , \wRegOut_7_93[11] , \wRegOut_7_93[10] , 
        \wRegOut_7_93[9] , \wRegOut_7_93[8] , \wRegOut_7_93[7] , 
        \wRegOut_7_93[6] , \wRegOut_7_93[5] , \wRegOut_7_93[4] , 
        \wRegOut_7_93[3] , \wRegOut_7_93[2] , \wRegOut_7_93[1] , 
        \wRegOut_7_93[0] }), .Enable1(\wRegEnTop_7_93[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_93[31] , \wRegInTop_7_93[30] , \wRegInTop_7_93[29] , 
        \wRegInTop_7_93[28] , \wRegInTop_7_93[27] , \wRegInTop_7_93[26] , 
        \wRegInTop_7_93[25] , \wRegInTop_7_93[24] , \wRegInTop_7_93[23] , 
        \wRegInTop_7_93[22] , \wRegInTop_7_93[21] , \wRegInTop_7_93[20] , 
        \wRegInTop_7_93[19] , \wRegInTop_7_93[18] , \wRegInTop_7_93[17] , 
        \wRegInTop_7_93[16] , \wRegInTop_7_93[15] , \wRegInTop_7_93[14] , 
        \wRegInTop_7_93[13] , \wRegInTop_7_93[12] , \wRegInTop_7_93[11] , 
        \wRegInTop_7_93[10] , \wRegInTop_7_93[9] , \wRegInTop_7_93[8] , 
        \wRegInTop_7_93[7] , \wRegInTop_7_93[6] , \wRegInTop_7_93[5] , 
        \wRegInTop_7_93[4] , \wRegInTop_7_93[3] , \wRegInTop_7_93[2] , 
        \wRegInTop_7_93[1] , \wRegInTop_7_93[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_2[0] ), .P_In({\wRegOut_5_2[31] , 
        \wRegOut_5_2[30] , \wRegOut_5_2[29] , \wRegOut_5_2[28] , 
        \wRegOut_5_2[27] , \wRegOut_5_2[26] , \wRegOut_5_2[25] , 
        \wRegOut_5_2[24] , \wRegOut_5_2[23] , \wRegOut_5_2[22] , 
        \wRegOut_5_2[21] , \wRegOut_5_2[20] , \wRegOut_5_2[19] , 
        \wRegOut_5_2[18] , \wRegOut_5_2[17] , \wRegOut_5_2[16] , 
        \wRegOut_5_2[15] , \wRegOut_5_2[14] , \wRegOut_5_2[13] , 
        \wRegOut_5_2[12] , \wRegOut_5_2[11] , \wRegOut_5_2[10] , 
        \wRegOut_5_2[9] , \wRegOut_5_2[8] , \wRegOut_5_2[7] , \wRegOut_5_2[6] , 
        \wRegOut_5_2[5] , \wRegOut_5_2[4] , \wRegOut_5_2[3] , \wRegOut_5_2[2] , 
        \wRegOut_5_2[1] , \wRegOut_5_2[0] }), .P_Out({\wRegInBot_5_2[31] , 
        \wRegInBot_5_2[30] , \wRegInBot_5_2[29] , \wRegInBot_5_2[28] , 
        \wRegInBot_5_2[27] , \wRegInBot_5_2[26] , \wRegInBot_5_2[25] , 
        \wRegInBot_5_2[24] , \wRegInBot_5_2[23] , \wRegInBot_5_2[22] , 
        \wRegInBot_5_2[21] , \wRegInBot_5_2[20] , \wRegInBot_5_2[19] , 
        \wRegInBot_5_2[18] , \wRegInBot_5_2[17] , \wRegInBot_5_2[16] , 
        \wRegInBot_5_2[15] , \wRegInBot_5_2[14] , \wRegInBot_5_2[13] , 
        \wRegInBot_5_2[12] , \wRegInBot_5_2[11] , \wRegInBot_5_2[10] , 
        \wRegInBot_5_2[9] , \wRegInBot_5_2[8] , \wRegInBot_5_2[7] , 
        \wRegInBot_5_2[6] , \wRegInBot_5_2[5] , \wRegInBot_5_2[4] , 
        \wRegInBot_5_2[3] , \wRegInBot_5_2[2] , \wRegInBot_5_2[1] , 
        \wRegInBot_5_2[0] }), .L_WR(\wRegEnTop_6_4[0] ), .L_In({
        \wRegOut_6_4[31] , \wRegOut_6_4[30] , \wRegOut_6_4[29] , 
        \wRegOut_6_4[28] , \wRegOut_6_4[27] , \wRegOut_6_4[26] , 
        \wRegOut_6_4[25] , \wRegOut_6_4[24] , \wRegOut_6_4[23] , 
        \wRegOut_6_4[22] , \wRegOut_6_4[21] , \wRegOut_6_4[20] , 
        \wRegOut_6_4[19] , \wRegOut_6_4[18] , \wRegOut_6_4[17] , 
        \wRegOut_6_4[16] , \wRegOut_6_4[15] , \wRegOut_6_4[14] , 
        \wRegOut_6_4[13] , \wRegOut_6_4[12] , \wRegOut_6_4[11] , 
        \wRegOut_6_4[10] , \wRegOut_6_4[9] , \wRegOut_6_4[8] , 
        \wRegOut_6_4[7] , \wRegOut_6_4[6] , \wRegOut_6_4[5] , \wRegOut_6_4[4] , 
        \wRegOut_6_4[3] , \wRegOut_6_4[2] , \wRegOut_6_4[1] , \wRegOut_6_4[0] 
        }), .L_Out({\wRegInTop_6_4[31] , \wRegInTop_6_4[30] , 
        \wRegInTop_6_4[29] , \wRegInTop_6_4[28] , \wRegInTop_6_4[27] , 
        \wRegInTop_6_4[26] , \wRegInTop_6_4[25] , \wRegInTop_6_4[24] , 
        \wRegInTop_6_4[23] , \wRegInTop_6_4[22] , \wRegInTop_6_4[21] , 
        \wRegInTop_6_4[20] , \wRegInTop_6_4[19] , \wRegInTop_6_4[18] , 
        \wRegInTop_6_4[17] , \wRegInTop_6_4[16] , \wRegInTop_6_4[15] , 
        \wRegInTop_6_4[14] , \wRegInTop_6_4[13] , \wRegInTop_6_4[12] , 
        \wRegInTop_6_4[11] , \wRegInTop_6_4[10] , \wRegInTop_6_4[9] , 
        \wRegInTop_6_4[8] , \wRegInTop_6_4[7] , \wRegInTop_6_4[6] , 
        \wRegInTop_6_4[5] , \wRegInTop_6_4[4] , \wRegInTop_6_4[3] , 
        \wRegInTop_6_4[2] , \wRegInTop_6_4[1] , \wRegInTop_6_4[0] }), .R_WR(
        \wRegEnTop_6_5[0] ), .R_In({\wRegOut_6_5[31] , \wRegOut_6_5[30] , 
        \wRegOut_6_5[29] , \wRegOut_6_5[28] , \wRegOut_6_5[27] , 
        \wRegOut_6_5[26] , \wRegOut_6_5[25] , \wRegOut_6_5[24] , 
        \wRegOut_6_5[23] , \wRegOut_6_5[22] , \wRegOut_6_5[21] , 
        \wRegOut_6_5[20] , \wRegOut_6_5[19] , \wRegOut_6_5[18] , 
        \wRegOut_6_5[17] , \wRegOut_6_5[16] , \wRegOut_6_5[15] , 
        \wRegOut_6_5[14] , \wRegOut_6_5[13] , \wRegOut_6_5[12] , 
        \wRegOut_6_5[11] , \wRegOut_6_5[10] , \wRegOut_6_5[9] , 
        \wRegOut_6_5[8] , \wRegOut_6_5[7] , \wRegOut_6_5[6] , \wRegOut_6_5[5] , 
        \wRegOut_6_5[4] , \wRegOut_6_5[3] , \wRegOut_6_5[2] , \wRegOut_6_5[1] , 
        \wRegOut_6_5[0] }), .R_Out({\wRegInTop_6_5[31] , \wRegInTop_6_5[30] , 
        \wRegInTop_6_5[29] , \wRegInTop_6_5[28] , \wRegInTop_6_5[27] , 
        \wRegInTop_6_5[26] , \wRegInTop_6_5[25] , \wRegInTop_6_5[24] , 
        \wRegInTop_6_5[23] , \wRegInTop_6_5[22] , \wRegInTop_6_5[21] , 
        \wRegInTop_6_5[20] , \wRegInTop_6_5[19] , \wRegInTop_6_5[18] , 
        \wRegInTop_6_5[17] , \wRegInTop_6_5[16] , \wRegInTop_6_5[15] , 
        \wRegInTop_6_5[14] , \wRegInTop_6_5[13] , \wRegInTop_6_5[12] , 
        \wRegInTop_6_5[11] , \wRegInTop_6_5[10] , \wRegInTop_6_5[9] , 
        \wRegInTop_6_5[8] , \wRegInTop_6_5[7] , \wRegInTop_6_5[6] , 
        \wRegInTop_6_5[5] , \wRegInTop_6_5[4] , \wRegInTop_6_5[3] , 
        \wRegInTop_6_5[2] , \wRegInTop_6_5[1] , \wRegInTop_6_5[0] }) );
    BHeap_Node_WIDTH32 BHN_6_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_63[0] ), .P_In({\wRegOut_6_63[31] , 
        \wRegOut_6_63[30] , \wRegOut_6_63[29] , \wRegOut_6_63[28] , 
        \wRegOut_6_63[27] , \wRegOut_6_63[26] , \wRegOut_6_63[25] , 
        \wRegOut_6_63[24] , \wRegOut_6_63[23] , \wRegOut_6_63[22] , 
        \wRegOut_6_63[21] , \wRegOut_6_63[20] , \wRegOut_6_63[19] , 
        \wRegOut_6_63[18] , \wRegOut_6_63[17] , \wRegOut_6_63[16] , 
        \wRegOut_6_63[15] , \wRegOut_6_63[14] , \wRegOut_6_63[13] , 
        \wRegOut_6_63[12] , \wRegOut_6_63[11] , \wRegOut_6_63[10] , 
        \wRegOut_6_63[9] , \wRegOut_6_63[8] , \wRegOut_6_63[7] , 
        \wRegOut_6_63[6] , \wRegOut_6_63[5] , \wRegOut_6_63[4] , 
        \wRegOut_6_63[3] , \wRegOut_6_63[2] , \wRegOut_6_63[1] , 
        \wRegOut_6_63[0] }), .P_Out({\wRegInBot_6_63[31] , 
        \wRegInBot_6_63[30] , \wRegInBot_6_63[29] , \wRegInBot_6_63[28] , 
        \wRegInBot_6_63[27] , \wRegInBot_6_63[26] , \wRegInBot_6_63[25] , 
        \wRegInBot_6_63[24] , \wRegInBot_6_63[23] , \wRegInBot_6_63[22] , 
        \wRegInBot_6_63[21] , \wRegInBot_6_63[20] , \wRegInBot_6_63[19] , 
        \wRegInBot_6_63[18] , \wRegInBot_6_63[17] , \wRegInBot_6_63[16] , 
        \wRegInBot_6_63[15] , \wRegInBot_6_63[14] , \wRegInBot_6_63[13] , 
        \wRegInBot_6_63[12] , \wRegInBot_6_63[11] , \wRegInBot_6_63[10] , 
        \wRegInBot_6_63[9] , \wRegInBot_6_63[8] , \wRegInBot_6_63[7] , 
        \wRegInBot_6_63[6] , \wRegInBot_6_63[5] , \wRegInBot_6_63[4] , 
        \wRegInBot_6_63[3] , \wRegInBot_6_63[2] , \wRegInBot_6_63[1] , 
        \wRegInBot_6_63[0] }), .L_WR(\wRegEnTop_7_126[0] ), .L_In({
        \wRegOut_7_126[31] , \wRegOut_7_126[30] , \wRegOut_7_126[29] , 
        \wRegOut_7_126[28] , \wRegOut_7_126[27] , \wRegOut_7_126[26] , 
        \wRegOut_7_126[25] , \wRegOut_7_126[24] , \wRegOut_7_126[23] , 
        \wRegOut_7_126[22] , \wRegOut_7_126[21] , \wRegOut_7_126[20] , 
        \wRegOut_7_126[19] , \wRegOut_7_126[18] , \wRegOut_7_126[17] , 
        \wRegOut_7_126[16] , \wRegOut_7_126[15] , \wRegOut_7_126[14] , 
        \wRegOut_7_126[13] , \wRegOut_7_126[12] , \wRegOut_7_126[11] , 
        \wRegOut_7_126[10] , \wRegOut_7_126[9] , \wRegOut_7_126[8] , 
        \wRegOut_7_126[7] , \wRegOut_7_126[6] , \wRegOut_7_126[5] , 
        \wRegOut_7_126[4] , \wRegOut_7_126[3] , \wRegOut_7_126[2] , 
        \wRegOut_7_126[1] , \wRegOut_7_126[0] }), .L_Out({
        \wRegInTop_7_126[31] , \wRegInTop_7_126[30] , \wRegInTop_7_126[29] , 
        \wRegInTop_7_126[28] , \wRegInTop_7_126[27] , \wRegInTop_7_126[26] , 
        \wRegInTop_7_126[25] , \wRegInTop_7_126[24] , \wRegInTop_7_126[23] , 
        \wRegInTop_7_126[22] , \wRegInTop_7_126[21] , \wRegInTop_7_126[20] , 
        \wRegInTop_7_126[19] , \wRegInTop_7_126[18] , \wRegInTop_7_126[17] , 
        \wRegInTop_7_126[16] , \wRegInTop_7_126[15] , \wRegInTop_7_126[14] , 
        \wRegInTop_7_126[13] , \wRegInTop_7_126[12] , \wRegInTop_7_126[11] , 
        \wRegInTop_7_126[10] , \wRegInTop_7_126[9] , \wRegInTop_7_126[8] , 
        \wRegInTop_7_126[7] , \wRegInTop_7_126[6] , \wRegInTop_7_126[5] , 
        \wRegInTop_7_126[4] , \wRegInTop_7_126[3] , \wRegInTop_7_126[2] , 
        \wRegInTop_7_126[1] , \wRegInTop_7_126[0] }), .R_WR(
        \wRegEnTop_7_127[0] ), .R_In({\wRegOut_7_127[31] , \wRegOut_7_127[30] , 
        \wRegOut_7_127[29] , \wRegOut_7_127[28] , \wRegOut_7_127[27] , 
        \wRegOut_7_127[26] , \wRegOut_7_127[25] , \wRegOut_7_127[24] , 
        \wRegOut_7_127[23] , \wRegOut_7_127[22] , \wRegOut_7_127[21] , 
        \wRegOut_7_127[20] , \wRegOut_7_127[19] , \wRegOut_7_127[18] , 
        \wRegOut_7_127[17] , \wRegOut_7_127[16] , \wRegOut_7_127[15] , 
        \wRegOut_7_127[14] , \wRegOut_7_127[13] , \wRegOut_7_127[12] , 
        \wRegOut_7_127[11] , \wRegOut_7_127[10] , \wRegOut_7_127[9] , 
        \wRegOut_7_127[8] , \wRegOut_7_127[7] , \wRegOut_7_127[6] , 
        \wRegOut_7_127[5] , \wRegOut_7_127[4] , \wRegOut_7_127[3] , 
        \wRegOut_7_127[2] , \wRegOut_7_127[1] , \wRegOut_7_127[0] }), .R_Out({
        \wRegInTop_7_127[31] , \wRegInTop_7_127[30] , \wRegInTop_7_127[29] , 
        \wRegInTop_7_127[28] , \wRegInTop_7_127[27] , \wRegInTop_7_127[26] , 
        \wRegInTop_7_127[25] , \wRegInTop_7_127[24] , \wRegInTop_7_127[23] , 
        \wRegInTop_7_127[22] , \wRegInTop_7_127[21] , \wRegInTop_7_127[20] , 
        \wRegInTop_7_127[19] , \wRegInTop_7_127[18] , \wRegInTop_7_127[17] , 
        \wRegInTop_7_127[16] , \wRegInTop_7_127[15] , \wRegInTop_7_127[14] , 
        \wRegInTop_7_127[13] , \wRegInTop_7_127[12] , \wRegInTop_7_127[11] , 
        \wRegInTop_7_127[10] , \wRegInTop_7_127[9] , \wRegInTop_7_127[8] , 
        \wRegInTop_7_127[7] , \wRegInTop_7_127[6] , \wRegInTop_7_127[5] , 
        \wRegInTop_7_127[4] , \wRegInTop_7_127[3] , \wRegInTop_7_127[2] , 
        \wRegInTop_7_127[1] , \wRegInTop_7_127[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_51 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink179[31] , \ScanLink179[30] , \ScanLink179[29] , 
        \ScanLink179[28] , \ScanLink179[27] , \ScanLink179[26] , 
        \ScanLink179[25] , \ScanLink179[24] , \ScanLink179[23] , 
        \ScanLink179[22] , \ScanLink179[21] , \ScanLink179[20] , 
        \ScanLink179[19] , \ScanLink179[18] , \ScanLink179[17] , 
        \ScanLink179[16] , \ScanLink179[15] , \ScanLink179[14] , 
        \ScanLink179[13] , \ScanLink179[12] , \ScanLink179[11] , 
        \ScanLink179[10] , \ScanLink179[9] , \ScanLink179[8] , 
        \ScanLink179[7] , \ScanLink179[6] , \ScanLink179[5] , \ScanLink179[4] , 
        \ScanLink179[3] , \ScanLink179[2] , \ScanLink179[1] , \ScanLink179[0] 
        }), .ScanOut({\ScanLink178[31] , \ScanLink178[30] , \ScanLink178[29] , 
        \ScanLink178[28] , \ScanLink178[27] , \ScanLink178[26] , 
        \ScanLink178[25] , \ScanLink178[24] , \ScanLink178[23] , 
        \ScanLink178[22] , \ScanLink178[21] , \ScanLink178[20] , 
        \ScanLink178[19] , \ScanLink178[18] , \ScanLink178[17] , 
        \ScanLink178[16] , \ScanLink178[15] , \ScanLink178[14] , 
        \ScanLink178[13] , \ScanLink178[12] , \ScanLink178[11] , 
        \ScanLink178[10] , \ScanLink178[9] , \ScanLink178[8] , 
        \ScanLink178[7] , \ScanLink178[6] , \ScanLink178[5] , \ScanLink178[4] , 
        \ScanLink178[3] , \ScanLink178[2] , \ScanLink178[1] , \ScanLink178[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_51[31] , 
        \wRegOut_7_51[30] , \wRegOut_7_51[29] , \wRegOut_7_51[28] , 
        \wRegOut_7_51[27] , \wRegOut_7_51[26] , \wRegOut_7_51[25] , 
        \wRegOut_7_51[24] , \wRegOut_7_51[23] , \wRegOut_7_51[22] , 
        \wRegOut_7_51[21] , \wRegOut_7_51[20] , \wRegOut_7_51[19] , 
        \wRegOut_7_51[18] , \wRegOut_7_51[17] , \wRegOut_7_51[16] , 
        \wRegOut_7_51[15] , \wRegOut_7_51[14] , \wRegOut_7_51[13] , 
        \wRegOut_7_51[12] , \wRegOut_7_51[11] , \wRegOut_7_51[10] , 
        \wRegOut_7_51[9] , \wRegOut_7_51[8] , \wRegOut_7_51[7] , 
        \wRegOut_7_51[6] , \wRegOut_7_51[5] , \wRegOut_7_51[4] , 
        \wRegOut_7_51[3] , \wRegOut_7_51[2] , \wRegOut_7_51[1] , 
        \wRegOut_7_51[0] }), .Enable1(\wRegEnTop_7_51[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_51[31] , \wRegInTop_7_51[30] , \wRegInTop_7_51[29] , 
        \wRegInTop_7_51[28] , \wRegInTop_7_51[27] , \wRegInTop_7_51[26] , 
        \wRegInTop_7_51[25] , \wRegInTop_7_51[24] , \wRegInTop_7_51[23] , 
        \wRegInTop_7_51[22] , \wRegInTop_7_51[21] , \wRegInTop_7_51[20] , 
        \wRegInTop_7_51[19] , \wRegInTop_7_51[18] , \wRegInTop_7_51[17] , 
        \wRegInTop_7_51[16] , \wRegInTop_7_51[15] , \wRegInTop_7_51[14] , 
        \wRegInTop_7_51[13] , \wRegInTop_7_51[12] , \wRegInTop_7_51[11] , 
        \wRegInTop_7_51[10] , \wRegInTop_7_51[9] , \wRegInTop_7_51[8] , 
        \wRegInTop_7_51[7] , \wRegInTop_7_51[6] , \wRegInTop_7_51[5] , 
        \wRegInTop_7_51[4] , \wRegInTop_7_51[3] , \wRegInTop_7_51[2] , 
        \wRegInTop_7_51[1] , \wRegInTop_7_51[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_37 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink101[31] , \ScanLink101[30] , \ScanLink101[29] , 
        \ScanLink101[28] , \ScanLink101[27] , \ScanLink101[26] , 
        \ScanLink101[25] , \ScanLink101[24] , \ScanLink101[23] , 
        \ScanLink101[22] , \ScanLink101[21] , \ScanLink101[20] , 
        \ScanLink101[19] , \ScanLink101[18] , \ScanLink101[17] , 
        \ScanLink101[16] , \ScanLink101[15] , \ScanLink101[14] , 
        \ScanLink101[13] , \ScanLink101[12] , \ScanLink101[11] , 
        \ScanLink101[10] , \ScanLink101[9] , \ScanLink101[8] , 
        \ScanLink101[7] , \ScanLink101[6] , \ScanLink101[5] , \ScanLink101[4] , 
        \ScanLink101[3] , \ScanLink101[2] , \ScanLink101[1] , \ScanLink101[0] 
        }), .ScanOut({\ScanLink100[31] , \ScanLink100[30] , \ScanLink100[29] , 
        \ScanLink100[28] , \ScanLink100[27] , \ScanLink100[26] , 
        \ScanLink100[25] , \ScanLink100[24] , \ScanLink100[23] , 
        \ScanLink100[22] , \ScanLink100[21] , \ScanLink100[20] , 
        \ScanLink100[19] , \ScanLink100[18] , \ScanLink100[17] , 
        \ScanLink100[16] , \ScanLink100[15] , \ScanLink100[14] , 
        \ScanLink100[13] , \ScanLink100[12] , \ScanLink100[11] , 
        \ScanLink100[10] , \ScanLink100[9] , \ScanLink100[8] , 
        \ScanLink100[7] , \ScanLink100[6] , \ScanLink100[5] , \ScanLink100[4] , 
        \ScanLink100[3] , \ScanLink100[2] , \ScanLink100[1] , \ScanLink100[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_37[31] , 
        \wRegOut_6_37[30] , \wRegOut_6_37[29] , \wRegOut_6_37[28] , 
        \wRegOut_6_37[27] , \wRegOut_6_37[26] , \wRegOut_6_37[25] , 
        \wRegOut_6_37[24] , \wRegOut_6_37[23] , \wRegOut_6_37[22] , 
        \wRegOut_6_37[21] , \wRegOut_6_37[20] , \wRegOut_6_37[19] , 
        \wRegOut_6_37[18] , \wRegOut_6_37[17] , \wRegOut_6_37[16] , 
        \wRegOut_6_37[15] , \wRegOut_6_37[14] , \wRegOut_6_37[13] , 
        \wRegOut_6_37[12] , \wRegOut_6_37[11] , \wRegOut_6_37[10] , 
        \wRegOut_6_37[9] , \wRegOut_6_37[8] , \wRegOut_6_37[7] , 
        \wRegOut_6_37[6] , \wRegOut_6_37[5] , \wRegOut_6_37[4] , 
        \wRegOut_6_37[3] , \wRegOut_6_37[2] , \wRegOut_6_37[1] , 
        \wRegOut_6_37[0] }), .Enable1(\wRegEnTop_6_37[0] ), .Enable2(
        \wRegEnBot_6_37[0] ), .In1({\wRegInTop_6_37[31] , \wRegInTop_6_37[30] , 
        \wRegInTop_6_37[29] , \wRegInTop_6_37[28] , \wRegInTop_6_37[27] , 
        \wRegInTop_6_37[26] , \wRegInTop_6_37[25] , \wRegInTop_6_37[24] , 
        \wRegInTop_6_37[23] , \wRegInTop_6_37[22] , \wRegInTop_6_37[21] , 
        \wRegInTop_6_37[20] , \wRegInTop_6_37[19] , \wRegInTop_6_37[18] , 
        \wRegInTop_6_37[17] , \wRegInTop_6_37[16] , \wRegInTop_6_37[15] , 
        \wRegInTop_6_37[14] , \wRegInTop_6_37[13] , \wRegInTop_6_37[12] , 
        \wRegInTop_6_37[11] , \wRegInTop_6_37[10] , \wRegInTop_6_37[9] , 
        \wRegInTop_6_37[8] , \wRegInTop_6_37[7] , \wRegInTop_6_37[6] , 
        \wRegInTop_6_37[5] , \wRegInTop_6_37[4] , \wRegInTop_6_37[3] , 
        \wRegInTop_6_37[2] , \wRegInTop_6_37[1] , \wRegInTop_6_37[0] }), .In2(
        {\wRegInBot_6_37[31] , \wRegInBot_6_37[30] , \wRegInBot_6_37[29] , 
        \wRegInBot_6_37[28] , \wRegInBot_6_37[27] , \wRegInBot_6_37[26] , 
        \wRegInBot_6_37[25] , \wRegInBot_6_37[24] , \wRegInBot_6_37[23] , 
        \wRegInBot_6_37[22] , \wRegInBot_6_37[21] , \wRegInBot_6_37[20] , 
        \wRegInBot_6_37[19] , \wRegInBot_6_37[18] , \wRegInBot_6_37[17] , 
        \wRegInBot_6_37[16] , \wRegInBot_6_37[15] , \wRegInBot_6_37[14] , 
        \wRegInBot_6_37[13] , \wRegInBot_6_37[12] , \wRegInBot_6_37[11] , 
        \wRegInBot_6_37[10] , \wRegInBot_6_37[9] , \wRegInBot_6_37[8] , 
        \wRegInBot_6_37[7] , \wRegInBot_6_37[6] , \wRegInBot_6_37[5] , 
        \wRegInBot_6_37[4] , \wRegInBot_6_37[3] , \wRegInBot_6_37[2] , 
        \wRegInBot_6_37[1] , \wRegInBot_6_37[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_76 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink204[31] , \ScanLink204[30] , \ScanLink204[29] , 
        \ScanLink204[28] , \ScanLink204[27] , \ScanLink204[26] , 
        \ScanLink204[25] , \ScanLink204[24] , \ScanLink204[23] , 
        \ScanLink204[22] , \ScanLink204[21] , \ScanLink204[20] , 
        \ScanLink204[19] , \ScanLink204[18] , \ScanLink204[17] , 
        \ScanLink204[16] , \ScanLink204[15] , \ScanLink204[14] , 
        \ScanLink204[13] , \ScanLink204[12] , \ScanLink204[11] , 
        \ScanLink204[10] , \ScanLink204[9] , \ScanLink204[8] , 
        \ScanLink204[7] , \ScanLink204[6] , \ScanLink204[5] , \ScanLink204[4] , 
        \ScanLink204[3] , \ScanLink204[2] , \ScanLink204[1] , \ScanLink204[0] 
        }), .ScanOut({\ScanLink203[31] , \ScanLink203[30] , \ScanLink203[29] , 
        \ScanLink203[28] , \ScanLink203[27] , \ScanLink203[26] , 
        \ScanLink203[25] , \ScanLink203[24] , \ScanLink203[23] , 
        \ScanLink203[22] , \ScanLink203[21] , \ScanLink203[20] , 
        \ScanLink203[19] , \ScanLink203[18] , \ScanLink203[17] , 
        \ScanLink203[16] , \ScanLink203[15] , \ScanLink203[14] , 
        \ScanLink203[13] , \ScanLink203[12] , \ScanLink203[11] , 
        \ScanLink203[10] , \ScanLink203[9] , \ScanLink203[8] , 
        \ScanLink203[7] , \ScanLink203[6] , \ScanLink203[5] , \ScanLink203[4] , 
        \ScanLink203[3] , \ScanLink203[2] , \ScanLink203[1] , \ScanLink203[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_76[31] , 
        \wRegOut_7_76[30] , \wRegOut_7_76[29] , \wRegOut_7_76[28] , 
        \wRegOut_7_76[27] , \wRegOut_7_76[26] , \wRegOut_7_76[25] , 
        \wRegOut_7_76[24] , \wRegOut_7_76[23] , \wRegOut_7_76[22] , 
        \wRegOut_7_76[21] , \wRegOut_7_76[20] , \wRegOut_7_76[19] , 
        \wRegOut_7_76[18] , \wRegOut_7_76[17] , \wRegOut_7_76[16] , 
        \wRegOut_7_76[15] , \wRegOut_7_76[14] , \wRegOut_7_76[13] , 
        \wRegOut_7_76[12] , \wRegOut_7_76[11] , \wRegOut_7_76[10] , 
        \wRegOut_7_76[9] , \wRegOut_7_76[8] , \wRegOut_7_76[7] , 
        \wRegOut_7_76[6] , \wRegOut_7_76[5] , \wRegOut_7_76[4] , 
        \wRegOut_7_76[3] , \wRegOut_7_76[2] , \wRegOut_7_76[1] , 
        \wRegOut_7_76[0] }), .Enable1(\wRegEnTop_7_76[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_76[31] , \wRegInTop_7_76[30] , \wRegInTop_7_76[29] , 
        \wRegInTop_7_76[28] , \wRegInTop_7_76[27] , \wRegInTop_7_76[26] , 
        \wRegInTop_7_76[25] , \wRegInTop_7_76[24] , \wRegInTop_7_76[23] , 
        \wRegInTop_7_76[22] , \wRegInTop_7_76[21] , \wRegInTop_7_76[20] , 
        \wRegInTop_7_76[19] , \wRegInTop_7_76[18] , \wRegInTop_7_76[17] , 
        \wRegInTop_7_76[16] , \wRegInTop_7_76[15] , \wRegInTop_7_76[14] , 
        \wRegInTop_7_76[13] , \wRegInTop_7_76[12] , \wRegInTop_7_76[11] , 
        \wRegInTop_7_76[10] , \wRegInTop_7_76[9] , \wRegInTop_7_76[8] , 
        \wRegInTop_7_76[7] , \wRegInTop_7_76[6] , \wRegInTop_7_76[5] , 
        \wRegInTop_7_76[4] , \wRegInTop_7_76[3] , \wRegInTop_7_76[2] , 
        \wRegInTop_7_76[1] , \wRegInTop_7_76[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink133[31] , \ScanLink133[30] , \ScanLink133[29] , 
        \ScanLink133[28] , \ScanLink133[27] , \ScanLink133[26] , 
        \ScanLink133[25] , \ScanLink133[24] , \ScanLink133[23] , 
        \ScanLink133[22] , \ScanLink133[21] , \ScanLink133[20] , 
        \ScanLink133[19] , \ScanLink133[18] , \ScanLink133[17] , 
        \ScanLink133[16] , \ScanLink133[15] , \ScanLink133[14] , 
        \ScanLink133[13] , \ScanLink133[12] , \ScanLink133[11] , 
        \ScanLink133[10] , \ScanLink133[9] , \ScanLink133[8] , 
        \ScanLink133[7] , \ScanLink133[6] , \ScanLink133[5] , \ScanLink133[4] , 
        \ScanLink133[3] , \ScanLink133[2] , \ScanLink133[1] , \ScanLink133[0] 
        }), .ScanOut({\ScanLink132[31] , \ScanLink132[30] , \ScanLink132[29] , 
        \ScanLink132[28] , \ScanLink132[27] , \ScanLink132[26] , 
        \ScanLink132[25] , \ScanLink132[24] , \ScanLink132[23] , 
        \ScanLink132[22] , \ScanLink132[21] , \ScanLink132[20] , 
        \ScanLink132[19] , \ScanLink132[18] , \ScanLink132[17] , 
        \ScanLink132[16] , \ScanLink132[15] , \ScanLink132[14] , 
        \ScanLink132[13] , \ScanLink132[12] , \ScanLink132[11] , 
        \ScanLink132[10] , \ScanLink132[9] , \ScanLink132[8] , 
        \ScanLink132[7] , \ScanLink132[6] , \ScanLink132[5] , \ScanLink132[4] , 
        \ScanLink132[3] , \ScanLink132[2] , \ScanLink132[1] , \ScanLink132[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_5[31] , 
        \wRegOut_7_5[30] , \wRegOut_7_5[29] , \wRegOut_7_5[28] , 
        \wRegOut_7_5[27] , \wRegOut_7_5[26] , \wRegOut_7_5[25] , 
        \wRegOut_7_5[24] , \wRegOut_7_5[23] , \wRegOut_7_5[22] , 
        \wRegOut_7_5[21] , \wRegOut_7_5[20] , \wRegOut_7_5[19] , 
        \wRegOut_7_5[18] , \wRegOut_7_5[17] , \wRegOut_7_5[16] , 
        \wRegOut_7_5[15] , \wRegOut_7_5[14] , \wRegOut_7_5[13] , 
        \wRegOut_7_5[12] , \wRegOut_7_5[11] , \wRegOut_7_5[10] , 
        \wRegOut_7_5[9] , \wRegOut_7_5[8] , \wRegOut_7_5[7] , \wRegOut_7_5[6] , 
        \wRegOut_7_5[5] , \wRegOut_7_5[4] , \wRegOut_7_5[3] , \wRegOut_7_5[2] , 
        \wRegOut_7_5[1] , \wRegOut_7_5[0] }), .Enable1(\wRegEnTop_7_5[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_5[31] , \wRegInTop_7_5[30] , 
        \wRegInTop_7_5[29] , \wRegInTop_7_5[28] , \wRegInTop_7_5[27] , 
        \wRegInTop_7_5[26] , \wRegInTop_7_5[25] , \wRegInTop_7_5[24] , 
        \wRegInTop_7_5[23] , \wRegInTop_7_5[22] , \wRegInTop_7_5[21] , 
        \wRegInTop_7_5[20] , \wRegInTop_7_5[19] , \wRegInTop_7_5[18] , 
        \wRegInTop_7_5[17] , \wRegInTop_7_5[16] , \wRegInTop_7_5[15] , 
        \wRegInTop_7_5[14] , \wRegInTop_7_5[13] , \wRegInTop_7_5[12] , 
        \wRegInTop_7_5[11] , \wRegInTop_7_5[10] , \wRegInTop_7_5[9] , 
        \wRegInTop_7_5[8] , \wRegInTop_7_5[7] , \wRegInTop_7_5[6] , 
        \wRegInTop_7_5[5] , \wRegInTop_7_5[4] , \wRegInTop_7_5[3] , 
        \wRegInTop_7_5[2] , \wRegInTop_7_5[1] , \wRegInTop_7_5[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_43 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink171[31] , \ScanLink171[30] , \ScanLink171[29] , 
        \ScanLink171[28] , \ScanLink171[27] , \ScanLink171[26] , 
        \ScanLink171[25] , \ScanLink171[24] , \ScanLink171[23] , 
        \ScanLink171[22] , \ScanLink171[21] , \ScanLink171[20] , 
        \ScanLink171[19] , \ScanLink171[18] , \ScanLink171[17] , 
        \ScanLink171[16] , \ScanLink171[15] , \ScanLink171[14] , 
        \ScanLink171[13] , \ScanLink171[12] , \ScanLink171[11] , 
        \ScanLink171[10] , \ScanLink171[9] , \ScanLink171[8] , 
        \ScanLink171[7] , \ScanLink171[6] , \ScanLink171[5] , \ScanLink171[4] , 
        \ScanLink171[3] , \ScanLink171[2] , \ScanLink171[1] , \ScanLink171[0] 
        }), .ScanOut({\ScanLink170[31] , \ScanLink170[30] , \ScanLink170[29] , 
        \ScanLink170[28] , \ScanLink170[27] , \ScanLink170[26] , 
        \ScanLink170[25] , \ScanLink170[24] , \ScanLink170[23] , 
        \ScanLink170[22] , \ScanLink170[21] , \ScanLink170[20] , 
        \ScanLink170[19] , \ScanLink170[18] , \ScanLink170[17] , 
        \ScanLink170[16] , \ScanLink170[15] , \ScanLink170[14] , 
        \ScanLink170[13] , \ScanLink170[12] , \ScanLink170[11] , 
        \ScanLink170[10] , \ScanLink170[9] , \ScanLink170[8] , 
        \ScanLink170[7] , \ScanLink170[6] , \ScanLink170[5] , \ScanLink170[4] , 
        \ScanLink170[3] , \ScanLink170[2] , \ScanLink170[1] , \ScanLink170[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_43[31] , 
        \wRegOut_7_43[30] , \wRegOut_7_43[29] , \wRegOut_7_43[28] , 
        \wRegOut_7_43[27] , \wRegOut_7_43[26] , \wRegOut_7_43[25] , 
        \wRegOut_7_43[24] , \wRegOut_7_43[23] , \wRegOut_7_43[22] , 
        \wRegOut_7_43[21] , \wRegOut_7_43[20] , \wRegOut_7_43[19] , 
        \wRegOut_7_43[18] , \wRegOut_7_43[17] , \wRegOut_7_43[16] , 
        \wRegOut_7_43[15] , \wRegOut_7_43[14] , \wRegOut_7_43[13] , 
        \wRegOut_7_43[12] , \wRegOut_7_43[11] , \wRegOut_7_43[10] , 
        \wRegOut_7_43[9] , \wRegOut_7_43[8] , \wRegOut_7_43[7] , 
        \wRegOut_7_43[6] , \wRegOut_7_43[5] , \wRegOut_7_43[4] , 
        \wRegOut_7_43[3] , \wRegOut_7_43[2] , \wRegOut_7_43[1] , 
        \wRegOut_7_43[0] }), .Enable1(\wRegEnTop_7_43[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_43[31] , \wRegInTop_7_43[30] , \wRegInTop_7_43[29] , 
        \wRegInTop_7_43[28] , \wRegInTop_7_43[27] , \wRegInTop_7_43[26] , 
        \wRegInTop_7_43[25] , \wRegInTop_7_43[24] , \wRegInTop_7_43[23] , 
        \wRegInTop_7_43[22] , \wRegInTop_7_43[21] , \wRegInTop_7_43[20] , 
        \wRegInTop_7_43[19] , \wRegInTop_7_43[18] , \wRegInTop_7_43[17] , 
        \wRegInTop_7_43[16] , \wRegInTop_7_43[15] , \wRegInTop_7_43[14] , 
        \wRegInTop_7_43[13] , \wRegInTop_7_43[12] , \wRegInTop_7_43[11] , 
        \wRegInTop_7_43[10] , \wRegInTop_7_43[9] , \wRegInTop_7_43[8] , 
        \wRegInTop_7_43[7] , \wRegInTop_7_43[6] , \wRegInTop_7_43[5] , 
        \wRegInTop_7_43[4] , \wRegInTop_7_43[3] , \wRegInTop_7_43[2] , 
        \wRegInTop_7_43[1] , \wRegInTop_7_43[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink11[31] , \ScanLink11[30] , \ScanLink11[29] , 
        \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , \ScanLink11[25] , 
        \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , \ScanLink11[21] , 
        \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , \ScanLink11[17] , 
        \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , \ScanLink11[13] , 
        \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , \ScanLink11[9] , 
        \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , \ScanLink11[5] , 
        \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , \ScanLink11[1] , 
        \ScanLink11[0] }), .ScanOut({\ScanLink10[31] , \ScanLink10[30] , 
        \ScanLink10[29] , \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , 
        \ScanLink10[25] , \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , 
        \ScanLink10[21] , \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , 
        \ScanLink10[17] , \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , 
        \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , 
        \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , 
        \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , 
        \ScanLink10[1] , \ScanLink10[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_3[31] , \wRegOut_3_3[30] , \wRegOut_3_3[29] , 
        \wRegOut_3_3[28] , \wRegOut_3_3[27] , \wRegOut_3_3[26] , 
        \wRegOut_3_3[25] , \wRegOut_3_3[24] , \wRegOut_3_3[23] , 
        \wRegOut_3_3[22] , \wRegOut_3_3[21] , \wRegOut_3_3[20] , 
        \wRegOut_3_3[19] , \wRegOut_3_3[18] , \wRegOut_3_3[17] , 
        \wRegOut_3_3[16] , \wRegOut_3_3[15] , \wRegOut_3_3[14] , 
        \wRegOut_3_3[13] , \wRegOut_3_3[12] , \wRegOut_3_3[11] , 
        \wRegOut_3_3[10] , \wRegOut_3_3[9] , \wRegOut_3_3[8] , 
        \wRegOut_3_3[7] , \wRegOut_3_3[6] , \wRegOut_3_3[5] , \wRegOut_3_3[4] , 
        \wRegOut_3_3[3] , \wRegOut_3_3[2] , \wRegOut_3_3[1] , \wRegOut_3_3[0] 
        }), .Enable1(\wRegEnTop_3_3[0] ), .Enable2(\wRegEnBot_3_3[0] ), .In1({
        \wRegInTop_3_3[31] , \wRegInTop_3_3[30] , \wRegInTop_3_3[29] , 
        \wRegInTop_3_3[28] , \wRegInTop_3_3[27] , \wRegInTop_3_3[26] , 
        \wRegInTop_3_3[25] , \wRegInTop_3_3[24] , \wRegInTop_3_3[23] , 
        \wRegInTop_3_3[22] , \wRegInTop_3_3[21] , \wRegInTop_3_3[20] , 
        \wRegInTop_3_3[19] , \wRegInTop_3_3[18] , \wRegInTop_3_3[17] , 
        \wRegInTop_3_3[16] , \wRegInTop_3_3[15] , \wRegInTop_3_3[14] , 
        \wRegInTop_3_3[13] , \wRegInTop_3_3[12] , \wRegInTop_3_3[11] , 
        \wRegInTop_3_3[10] , \wRegInTop_3_3[9] , \wRegInTop_3_3[8] , 
        \wRegInTop_3_3[7] , \wRegInTop_3_3[6] , \wRegInTop_3_3[5] , 
        \wRegInTop_3_3[4] , \wRegInTop_3_3[3] , \wRegInTop_3_3[2] , 
        \wRegInTop_3_3[1] , \wRegInTop_3_3[0] }), .In2({\wRegInBot_3_3[31] , 
        \wRegInBot_3_3[30] , \wRegInBot_3_3[29] , \wRegInBot_3_3[28] , 
        \wRegInBot_3_3[27] , \wRegInBot_3_3[26] , \wRegInBot_3_3[25] , 
        \wRegInBot_3_3[24] , \wRegInBot_3_3[23] , \wRegInBot_3_3[22] , 
        \wRegInBot_3_3[21] , \wRegInBot_3_3[20] , \wRegInBot_3_3[19] , 
        \wRegInBot_3_3[18] , \wRegInBot_3_3[17] , \wRegInBot_3_3[16] , 
        \wRegInBot_3_3[15] , \wRegInBot_3_3[14] , \wRegInBot_3_3[13] , 
        \wRegInBot_3_3[12] , \wRegInBot_3_3[11] , \wRegInBot_3_3[10] , 
        \wRegInBot_3_3[9] , \wRegInBot_3_3[8] , \wRegInBot_3_3[7] , 
        \wRegInBot_3_3[6] , \wRegInBot_3_3[5] , \wRegInBot_3_3[4] , 
        \wRegInBot_3_3[3] , \wRegInBot_3_3[2] , \wRegInBot_3_3[1] , 
        \wRegInBot_3_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink41[31] , \ScanLink41[30] , \ScanLink41[29] , 
        \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , \ScanLink41[25] , 
        \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , \ScanLink41[21] , 
        \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , \ScanLink41[17] , 
        \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , \ScanLink41[13] , 
        \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , \ScanLink41[9] , 
        \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , \ScanLink41[5] , 
        \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , \ScanLink41[1] , 
        \ScanLink41[0] }), .ScanOut({\ScanLink40[31] , \ScanLink40[30] , 
        \ScanLink40[29] , \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , 
        \ScanLink40[25] , \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , 
        \ScanLink40[21] , \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , 
        \ScanLink40[17] , \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , 
        \ScanLink40[13] , \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , 
        \ScanLink40[9] , \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , 
        \ScanLink40[5] , \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , 
        \ScanLink40[1] , \ScanLink40[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_9[31] , \wRegOut_5_9[30] , \wRegOut_5_9[29] , 
        \wRegOut_5_9[28] , \wRegOut_5_9[27] , \wRegOut_5_9[26] , 
        \wRegOut_5_9[25] , \wRegOut_5_9[24] , \wRegOut_5_9[23] , 
        \wRegOut_5_9[22] , \wRegOut_5_9[21] , \wRegOut_5_9[20] , 
        \wRegOut_5_9[19] , \wRegOut_5_9[18] , \wRegOut_5_9[17] , 
        \wRegOut_5_9[16] , \wRegOut_5_9[15] , \wRegOut_5_9[14] , 
        \wRegOut_5_9[13] , \wRegOut_5_9[12] , \wRegOut_5_9[11] , 
        \wRegOut_5_9[10] , \wRegOut_5_9[9] , \wRegOut_5_9[8] , 
        \wRegOut_5_9[7] , \wRegOut_5_9[6] , \wRegOut_5_9[5] , \wRegOut_5_9[4] , 
        \wRegOut_5_9[3] , \wRegOut_5_9[2] , \wRegOut_5_9[1] , \wRegOut_5_9[0] 
        }), .Enable1(\wRegEnTop_5_9[0] ), .Enable2(\wRegEnBot_5_9[0] ), .In1({
        \wRegInTop_5_9[31] , \wRegInTop_5_9[30] , \wRegInTop_5_9[29] , 
        \wRegInTop_5_9[28] , \wRegInTop_5_9[27] , \wRegInTop_5_9[26] , 
        \wRegInTop_5_9[25] , \wRegInTop_5_9[24] , \wRegInTop_5_9[23] , 
        \wRegInTop_5_9[22] , \wRegInTop_5_9[21] , \wRegInTop_5_9[20] , 
        \wRegInTop_5_9[19] , \wRegInTop_5_9[18] , \wRegInTop_5_9[17] , 
        \wRegInTop_5_9[16] , \wRegInTop_5_9[15] , \wRegInTop_5_9[14] , 
        \wRegInTop_5_9[13] , \wRegInTop_5_9[12] , \wRegInTop_5_9[11] , 
        \wRegInTop_5_9[10] , \wRegInTop_5_9[9] , \wRegInTop_5_9[8] , 
        \wRegInTop_5_9[7] , \wRegInTop_5_9[6] , \wRegInTop_5_9[5] , 
        \wRegInTop_5_9[4] , \wRegInTop_5_9[3] , \wRegInTop_5_9[2] , 
        \wRegInTop_5_9[1] , \wRegInTop_5_9[0] }), .In2({\wRegInBot_5_9[31] , 
        \wRegInBot_5_9[30] , \wRegInBot_5_9[29] , \wRegInBot_5_9[28] , 
        \wRegInBot_5_9[27] , \wRegInBot_5_9[26] , \wRegInBot_5_9[25] , 
        \wRegInBot_5_9[24] , \wRegInBot_5_9[23] , \wRegInBot_5_9[22] , 
        \wRegInBot_5_9[21] , \wRegInBot_5_9[20] , \wRegInBot_5_9[19] , 
        \wRegInBot_5_9[18] , \wRegInBot_5_9[17] , \wRegInBot_5_9[16] , 
        \wRegInBot_5_9[15] , \wRegInBot_5_9[14] , \wRegInBot_5_9[13] , 
        \wRegInBot_5_9[12] , \wRegInBot_5_9[11] , \wRegInBot_5_9[10] , 
        \wRegInBot_5_9[9] , \wRegInBot_5_9[8] , \wRegInBot_5_9[7] , 
        \wRegInBot_5_9[6] , \wRegInBot_5_9[5] , \wRegInBot_5_9[4] , 
        \wRegInBot_5_9[3] , \wRegInBot_5_9[2] , \wRegInBot_5_9[1] , 
        \wRegInBot_5_9[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_20 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink52[31] , \ScanLink52[30] , \ScanLink52[29] , 
        \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , \ScanLink52[25] , 
        \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , \ScanLink52[21] , 
        \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , \ScanLink52[17] , 
        \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , \ScanLink52[13] , 
        \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , \ScanLink52[9] , 
        \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , \ScanLink52[5] , 
        \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , \ScanLink52[1] , 
        \ScanLink52[0] }), .ScanOut({\ScanLink51[31] , \ScanLink51[30] , 
        \ScanLink51[29] , \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , 
        \ScanLink51[25] , \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , 
        \ScanLink51[21] , \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , 
        \ScanLink51[17] , \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , 
        \ScanLink51[13] , \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , 
        \ScanLink51[9] , \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , 
        \ScanLink51[5] , \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , 
        \ScanLink51[1] , \ScanLink51[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_20[31] , \wRegOut_5_20[30] , 
        \wRegOut_5_20[29] , \wRegOut_5_20[28] , \wRegOut_5_20[27] , 
        \wRegOut_5_20[26] , \wRegOut_5_20[25] , \wRegOut_5_20[24] , 
        \wRegOut_5_20[23] , \wRegOut_5_20[22] , \wRegOut_5_20[21] , 
        \wRegOut_5_20[20] , \wRegOut_5_20[19] , \wRegOut_5_20[18] , 
        \wRegOut_5_20[17] , \wRegOut_5_20[16] , \wRegOut_5_20[15] , 
        \wRegOut_5_20[14] , \wRegOut_5_20[13] , \wRegOut_5_20[12] , 
        \wRegOut_5_20[11] , \wRegOut_5_20[10] , \wRegOut_5_20[9] , 
        \wRegOut_5_20[8] , \wRegOut_5_20[7] , \wRegOut_5_20[6] , 
        \wRegOut_5_20[5] , \wRegOut_5_20[4] , \wRegOut_5_20[3] , 
        \wRegOut_5_20[2] , \wRegOut_5_20[1] , \wRegOut_5_20[0] }), .Enable1(
        \wRegEnTop_5_20[0] ), .Enable2(\wRegEnBot_5_20[0] ), .In1({
        \wRegInTop_5_20[31] , \wRegInTop_5_20[30] , \wRegInTop_5_20[29] , 
        \wRegInTop_5_20[28] , \wRegInTop_5_20[27] , \wRegInTop_5_20[26] , 
        \wRegInTop_5_20[25] , \wRegInTop_5_20[24] , \wRegInTop_5_20[23] , 
        \wRegInTop_5_20[22] , \wRegInTop_5_20[21] , \wRegInTop_5_20[20] , 
        \wRegInTop_5_20[19] , \wRegInTop_5_20[18] , \wRegInTop_5_20[17] , 
        \wRegInTop_5_20[16] , \wRegInTop_5_20[15] , \wRegInTop_5_20[14] , 
        \wRegInTop_5_20[13] , \wRegInTop_5_20[12] , \wRegInTop_5_20[11] , 
        \wRegInTop_5_20[10] , \wRegInTop_5_20[9] , \wRegInTop_5_20[8] , 
        \wRegInTop_5_20[7] , \wRegInTop_5_20[6] , \wRegInTop_5_20[5] , 
        \wRegInTop_5_20[4] , \wRegInTop_5_20[3] , \wRegInTop_5_20[2] , 
        \wRegInTop_5_20[1] , \wRegInTop_5_20[0] }), .In2({\wRegInBot_5_20[31] , 
        \wRegInBot_5_20[30] , \wRegInBot_5_20[29] , \wRegInBot_5_20[28] , 
        \wRegInBot_5_20[27] , \wRegInBot_5_20[26] , \wRegInBot_5_20[25] , 
        \wRegInBot_5_20[24] , \wRegInBot_5_20[23] , \wRegInBot_5_20[22] , 
        \wRegInBot_5_20[21] , \wRegInBot_5_20[20] , \wRegInBot_5_20[19] , 
        \wRegInBot_5_20[18] , \wRegInBot_5_20[17] , \wRegInBot_5_20[16] , 
        \wRegInBot_5_20[15] , \wRegInBot_5_20[14] , \wRegInBot_5_20[13] , 
        \wRegInBot_5_20[12] , \wRegInBot_5_20[11] , \wRegInBot_5_20[10] , 
        \wRegInBot_5_20[9] , \wRegInBot_5_20[8] , \wRegInBot_5_20[7] , 
        \wRegInBot_5_20[6] , \wRegInBot_5_20[5] , \wRegInBot_5_20[4] , 
        \wRegInBot_5_20[3] , \wRegInBot_5_20[2] , \wRegInBot_5_20[1] , 
        \wRegInBot_5_20[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink74[31] , \ScanLink74[30] , \ScanLink74[29] , 
        \ScanLink74[28] , \ScanLink74[27] , \ScanLink74[26] , \ScanLink74[25] , 
        \ScanLink74[24] , \ScanLink74[23] , \ScanLink74[22] , \ScanLink74[21] , 
        \ScanLink74[20] , \ScanLink74[19] , \ScanLink74[18] , \ScanLink74[17] , 
        \ScanLink74[16] , \ScanLink74[15] , \ScanLink74[14] , \ScanLink74[13] , 
        \ScanLink74[12] , \ScanLink74[11] , \ScanLink74[10] , \ScanLink74[9] , 
        \ScanLink74[8] , \ScanLink74[7] , \ScanLink74[6] , \ScanLink74[5] , 
        \ScanLink74[4] , \ScanLink74[3] , \ScanLink74[2] , \ScanLink74[1] , 
        \ScanLink74[0] }), .ScanOut({\ScanLink73[31] , \ScanLink73[30] , 
        \ScanLink73[29] , \ScanLink73[28] , \ScanLink73[27] , \ScanLink73[26] , 
        \ScanLink73[25] , \ScanLink73[24] , \ScanLink73[23] , \ScanLink73[22] , 
        \ScanLink73[21] , \ScanLink73[20] , \ScanLink73[19] , \ScanLink73[18] , 
        \ScanLink73[17] , \ScanLink73[16] , \ScanLink73[15] , \ScanLink73[14] , 
        \ScanLink73[13] , \ScanLink73[12] , \ScanLink73[11] , \ScanLink73[10] , 
        \ScanLink73[9] , \ScanLink73[8] , \ScanLink73[7] , \ScanLink73[6] , 
        \ScanLink73[5] , \ScanLink73[4] , \ScanLink73[3] , \ScanLink73[2] , 
        \ScanLink73[1] , \ScanLink73[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_10[31] , \wRegOut_6_10[30] , 
        \wRegOut_6_10[29] , \wRegOut_6_10[28] , \wRegOut_6_10[27] , 
        \wRegOut_6_10[26] , \wRegOut_6_10[25] , \wRegOut_6_10[24] , 
        \wRegOut_6_10[23] , \wRegOut_6_10[22] , \wRegOut_6_10[21] , 
        \wRegOut_6_10[20] , \wRegOut_6_10[19] , \wRegOut_6_10[18] , 
        \wRegOut_6_10[17] , \wRegOut_6_10[16] , \wRegOut_6_10[15] , 
        \wRegOut_6_10[14] , \wRegOut_6_10[13] , \wRegOut_6_10[12] , 
        \wRegOut_6_10[11] , \wRegOut_6_10[10] , \wRegOut_6_10[9] , 
        \wRegOut_6_10[8] , \wRegOut_6_10[7] , \wRegOut_6_10[6] , 
        \wRegOut_6_10[5] , \wRegOut_6_10[4] , \wRegOut_6_10[3] , 
        \wRegOut_6_10[2] , \wRegOut_6_10[1] , \wRegOut_6_10[0] }), .Enable1(
        \wRegEnTop_6_10[0] ), .Enable2(\wRegEnBot_6_10[0] ), .In1({
        \wRegInTop_6_10[31] , \wRegInTop_6_10[30] , \wRegInTop_6_10[29] , 
        \wRegInTop_6_10[28] , \wRegInTop_6_10[27] , \wRegInTop_6_10[26] , 
        \wRegInTop_6_10[25] , \wRegInTop_6_10[24] , \wRegInTop_6_10[23] , 
        \wRegInTop_6_10[22] , \wRegInTop_6_10[21] , \wRegInTop_6_10[20] , 
        \wRegInTop_6_10[19] , \wRegInTop_6_10[18] , \wRegInTop_6_10[17] , 
        \wRegInTop_6_10[16] , \wRegInTop_6_10[15] , \wRegInTop_6_10[14] , 
        \wRegInTop_6_10[13] , \wRegInTop_6_10[12] , \wRegInTop_6_10[11] , 
        \wRegInTop_6_10[10] , \wRegInTop_6_10[9] , \wRegInTop_6_10[8] , 
        \wRegInTop_6_10[7] , \wRegInTop_6_10[6] , \wRegInTop_6_10[5] , 
        \wRegInTop_6_10[4] , \wRegInTop_6_10[3] , \wRegInTop_6_10[2] , 
        \wRegInTop_6_10[1] , \wRegInTop_6_10[0] }), .In2({\wRegInBot_6_10[31] , 
        \wRegInBot_6_10[30] , \wRegInBot_6_10[29] , \wRegInBot_6_10[28] , 
        \wRegInBot_6_10[27] , \wRegInBot_6_10[26] , \wRegInBot_6_10[25] , 
        \wRegInBot_6_10[24] , \wRegInBot_6_10[23] , \wRegInBot_6_10[22] , 
        \wRegInBot_6_10[21] , \wRegInBot_6_10[20] , \wRegInBot_6_10[19] , 
        \wRegInBot_6_10[18] , \wRegInBot_6_10[17] , \wRegInBot_6_10[16] , 
        \wRegInBot_6_10[15] , \wRegInBot_6_10[14] , \wRegInBot_6_10[13] , 
        \wRegInBot_6_10[12] , \wRegInBot_6_10[11] , \wRegInBot_6_10[10] , 
        \wRegInBot_6_10[9] , \wRegInBot_6_10[8] , \wRegInBot_6_10[7] , 
        \wRegInBot_6_10[6] , \wRegInBot_6_10[5] , \wRegInBot_6_10[4] , 
        \wRegInBot_6_10[3] , \wRegInBot_6_10[2] , \wRegInBot_6_10[1] , 
        \wRegInBot_6_10[0] }) );
    BHeap_Node_WIDTH32 BHN_6_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_38[0] ), .P_In({\wRegOut_6_38[31] , 
        \wRegOut_6_38[30] , \wRegOut_6_38[29] , \wRegOut_6_38[28] , 
        \wRegOut_6_38[27] , \wRegOut_6_38[26] , \wRegOut_6_38[25] , 
        \wRegOut_6_38[24] , \wRegOut_6_38[23] , \wRegOut_6_38[22] , 
        \wRegOut_6_38[21] , \wRegOut_6_38[20] , \wRegOut_6_38[19] , 
        \wRegOut_6_38[18] , \wRegOut_6_38[17] , \wRegOut_6_38[16] , 
        \wRegOut_6_38[15] , \wRegOut_6_38[14] , \wRegOut_6_38[13] , 
        \wRegOut_6_38[12] , \wRegOut_6_38[11] , \wRegOut_6_38[10] , 
        \wRegOut_6_38[9] , \wRegOut_6_38[8] , \wRegOut_6_38[7] , 
        \wRegOut_6_38[6] , \wRegOut_6_38[5] , \wRegOut_6_38[4] , 
        \wRegOut_6_38[3] , \wRegOut_6_38[2] , \wRegOut_6_38[1] , 
        \wRegOut_6_38[0] }), .P_Out({\wRegInBot_6_38[31] , 
        \wRegInBot_6_38[30] , \wRegInBot_6_38[29] , \wRegInBot_6_38[28] , 
        \wRegInBot_6_38[27] , \wRegInBot_6_38[26] , \wRegInBot_6_38[25] , 
        \wRegInBot_6_38[24] , \wRegInBot_6_38[23] , \wRegInBot_6_38[22] , 
        \wRegInBot_6_38[21] , \wRegInBot_6_38[20] , \wRegInBot_6_38[19] , 
        \wRegInBot_6_38[18] , \wRegInBot_6_38[17] , \wRegInBot_6_38[16] , 
        \wRegInBot_6_38[15] , \wRegInBot_6_38[14] , \wRegInBot_6_38[13] , 
        \wRegInBot_6_38[12] , \wRegInBot_6_38[11] , \wRegInBot_6_38[10] , 
        \wRegInBot_6_38[9] , \wRegInBot_6_38[8] , \wRegInBot_6_38[7] , 
        \wRegInBot_6_38[6] , \wRegInBot_6_38[5] , \wRegInBot_6_38[4] , 
        \wRegInBot_6_38[3] , \wRegInBot_6_38[2] , \wRegInBot_6_38[1] , 
        \wRegInBot_6_38[0] }), .L_WR(\wRegEnTop_7_76[0] ), .L_In({
        \wRegOut_7_76[31] , \wRegOut_7_76[30] , \wRegOut_7_76[29] , 
        \wRegOut_7_76[28] , \wRegOut_7_76[27] , \wRegOut_7_76[26] , 
        \wRegOut_7_76[25] , \wRegOut_7_76[24] , \wRegOut_7_76[23] , 
        \wRegOut_7_76[22] , \wRegOut_7_76[21] , \wRegOut_7_76[20] , 
        \wRegOut_7_76[19] , \wRegOut_7_76[18] , \wRegOut_7_76[17] , 
        \wRegOut_7_76[16] , \wRegOut_7_76[15] , \wRegOut_7_76[14] , 
        \wRegOut_7_76[13] , \wRegOut_7_76[12] , \wRegOut_7_76[11] , 
        \wRegOut_7_76[10] , \wRegOut_7_76[9] , \wRegOut_7_76[8] , 
        \wRegOut_7_76[7] , \wRegOut_7_76[6] , \wRegOut_7_76[5] , 
        \wRegOut_7_76[4] , \wRegOut_7_76[3] , \wRegOut_7_76[2] , 
        \wRegOut_7_76[1] , \wRegOut_7_76[0] }), .L_Out({\wRegInTop_7_76[31] , 
        \wRegInTop_7_76[30] , \wRegInTop_7_76[29] , \wRegInTop_7_76[28] , 
        \wRegInTop_7_76[27] , \wRegInTop_7_76[26] , \wRegInTop_7_76[25] , 
        \wRegInTop_7_76[24] , \wRegInTop_7_76[23] , \wRegInTop_7_76[22] , 
        \wRegInTop_7_76[21] , \wRegInTop_7_76[20] , \wRegInTop_7_76[19] , 
        \wRegInTop_7_76[18] , \wRegInTop_7_76[17] , \wRegInTop_7_76[16] , 
        \wRegInTop_7_76[15] , \wRegInTop_7_76[14] , \wRegInTop_7_76[13] , 
        \wRegInTop_7_76[12] , \wRegInTop_7_76[11] , \wRegInTop_7_76[10] , 
        \wRegInTop_7_76[9] , \wRegInTop_7_76[8] , \wRegInTop_7_76[7] , 
        \wRegInTop_7_76[6] , \wRegInTop_7_76[5] , \wRegInTop_7_76[4] , 
        \wRegInTop_7_76[3] , \wRegInTop_7_76[2] , \wRegInTop_7_76[1] , 
        \wRegInTop_7_76[0] }), .R_WR(\wRegEnTop_7_77[0] ), .R_In({
        \wRegOut_7_77[31] , \wRegOut_7_77[30] , \wRegOut_7_77[29] , 
        \wRegOut_7_77[28] , \wRegOut_7_77[27] , \wRegOut_7_77[26] , 
        \wRegOut_7_77[25] , \wRegOut_7_77[24] , \wRegOut_7_77[23] , 
        \wRegOut_7_77[22] , \wRegOut_7_77[21] , \wRegOut_7_77[20] , 
        \wRegOut_7_77[19] , \wRegOut_7_77[18] , \wRegOut_7_77[17] , 
        \wRegOut_7_77[16] , \wRegOut_7_77[15] , \wRegOut_7_77[14] , 
        \wRegOut_7_77[13] , \wRegOut_7_77[12] , \wRegOut_7_77[11] , 
        \wRegOut_7_77[10] , \wRegOut_7_77[9] , \wRegOut_7_77[8] , 
        \wRegOut_7_77[7] , \wRegOut_7_77[6] , \wRegOut_7_77[5] , 
        \wRegOut_7_77[4] , \wRegOut_7_77[3] , \wRegOut_7_77[2] , 
        \wRegOut_7_77[1] , \wRegOut_7_77[0] }), .R_Out({\wRegInTop_7_77[31] , 
        \wRegInTop_7_77[30] , \wRegInTop_7_77[29] , \wRegInTop_7_77[28] , 
        \wRegInTop_7_77[27] , \wRegInTop_7_77[26] , \wRegInTop_7_77[25] , 
        \wRegInTop_7_77[24] , \wRegInTop_7_77[23] , \wRegInTop_7_77[22] , 
        \wRegInTop_7_77[21] , \wRegInTop_7_77[20] , \wRegInTop_7_77[19] , 
        \wRegInTop_7_77[18] , \wRegInTop_7_77[17] , \wRegInTop_7_77[16] , 
        \wRegInTop_7_77[15] , \wRegInTop_7_77[14] , \wRegInTop_7_77[13] , 
        \wRegInTop_7_77[12] , \wRegInTop_7_77[11] , \wRegInTop_7_77[10] , 
        \wRegInTop_7_77[9] , \wRegInTop_7_77[8] , \wRegInTop_7_77[7] , 
        \wRegInTop_7_77[6] , \wRegInTop_7_77[5] , \wRegInTop_7_77[4] , 
        \wRegInTop_7_77[3] , \wRegInTop_7_77[2] , \wRegInTop_7_77[1] , 
        \wRegInTop_7_77[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_64 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink192[31] , \ScanLink192[30] , \ScanLink192[29] , 
        \ScanLink192[28] , \ScanLink192[27] , \ScanLink192[26] , 
        \ScanLink192[25] , \ScanLink192[24] , \ScanLink192[23] , 
        \ScanLink192[22] , \ScanLink192[21] , \ScanLink192[20] , 
        \ScanLink192[19] , \ScanLink192[18] , \ScanLink192[17] , 
        \ScanLink192[16] , \ScanLink192[15] , \ScanLink192[14] , 
        \ScanLink192[13] , \ScanLink192[12] , \ScanLink192[11] , 
        \ScanLink192[10] , \ScanLink192[9] , \ScanLink192[8] , 
        \ScanLink192[7] , \ScanLink192[6] , \ScanLink192[5] , \ScanLink192[4] , 
        \ScanLink192[3] , \ScanLink192[2] , \ScanLink192[1] , \ScanLink192[0] 
        }), .ScanOut({\ScanLink191[31] , \ScanLink191[30] , \ScanLink191[29] , 
        \ScanLink191[28] , \ScanLink191[27] , \ScanLink191[26] , 
        \ScanLink191[25] , \ScanLink191[24] , \ScanLink191[23] , 
        \ScanLink191[22] , \ScanLink191[21] , \ScanLink191[20] , 
        \ScanLink191[19] , \ScanLink191[18] , \ScanLink191[17] , 
        \ScanLink191[16] , \ScanLink191[15] , \ScanLink191[14] , 
        \ScanLink191[13] , \ScanLink191[12] , \ScanLink191[11] , 
        \ScanLink191[10] , \ScanLink191[9] , \ScanLink191[8] , 
        \ScanLink191[7] , \ScanLink191[6] , \ScanLink191[5] , \ScanLink191[4] , 
        \ScanLink191[3] , \ScanLink191[2] , \ScanLink191[1] , \ScanLink191[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_64[31] , 
        \wRegOut_7_64[30] , \wRegOut_7_64[29] , \wRegOut_7_64[28] , 
        \wRegOut_7_64[27] , \wRegOut_7_64[26] , \wRegOut_7_64[25] , 
        \wRegOut_7_64[24] , \wRegOut_7_64[23] , \wRegOut_7_64[22] , 
        \wRegOut_7_64[21] , \wRegOut_7_64[20] , \wRegOut_7_64[19] , 
        \wRegOut_7_64[18] , \wRegOut_7_64[17] , \wRegOut_7_64[16] , 
        \wRegOut_7_64[15] , \wRegOut_7_64[14] , \wRegOut_7_64[13] , 
        \wRegOut_7_64[12] , \wRegOut_7_64[11] , \wRegOut_7_64[10] , 
        \wRegOut_7_64[9] , \wRegOut_7_64[8] , \wRegOut_7_64[7] , 
        \wRegOut_7_64[6] , \wRegOut_7_64[5] , \wRegOut_7_64[4] , 
        \wRegOut_7_64[3] , \wRegOut_7_64[2] , \wRegOut_7_64[1] , 
        \wRegOut_7_64[0] }), .Enable1(\wRegEnTop_7_64[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_64[31] , \wRegInTop_7_64[30] , \wRegInTop_7_64[29] , 
        \wRegInTop_7_64[28] , \wRegInTop_7_64[27] , \wRegInTop_7_64[26] , 
        \wRegInTop_7_64[25] , \wRegInTop_7_64[24] , \wRegInTop_7_64[23] , 
        \wRegInTop_7_64[22] , \wRegInTop_7_64[21] , \wRegInTop_7_64[20] , 
        \wRegInTop_7_64[19] , \wRegInTop_7_64[18] , \wRegInTop_7_64[17] , 
        \wRegInTop_7_64[16] , \wRegInTop_7_64[15] , \wRegInTop_7_64[14] , 
        \wRegInTop_7_64[13] , \wRegInTop_7_64[12] , \wRegInTop_7_64[11] , 
        \wRegInTop_7_64[10] , \wRegInTop_7_64[9] , \wRegInTop_7_64[8] , 
        \wRegInTop_7_64[7] , \wRegInTop_7_64[6] , \wRegInTop_7_64[5] , 
        \wRegInTop_7_64[4] , \wRegInTop_7_64[3] , \wRegInTop_7_64[2] , 
        \wRegInTop_7_64[1] , \wRegInTop_7_64[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_42 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink106[31] , \ScanLink106[30] , \ScanLink106[29] , 
        \ScanLink106[28] , \ScanLink106[27] , \ScanLink106[26] , 
        \ScanLink106[25] , \ScanLink106[24] , \ScanLink106[23] , 
        \ScanLink106[22] , \ScanLink106[21] , \ScanLink106[20] , 
        \ScanLink106[19] , \ScanLink106[18] , \ScanLink106[17] , 
        \ScanLink106[16] , \ScanLink106[15] , \ScanLink106[14] , 
        \ScanLink106[13] , \ScanLink106[12] , \ScanLink106[11] , 
        \ScanLink106[10] , \ScanLink106[9] , \ScanLink106[8] , 
        \ScanLink106[7] , \ScanLink106[6] , \ScanLink106[5] , \ScanLink106[4] , 
        \ScanLink106[3] , \ScanLink106[2] , \ScanLink106[1] , \ScanLink106[0] 
        }), .ScanOut({\ScanLink105[31] , \ScanLink105[30] , \ScanLink105[29] , 
        \ScanLink105[28] , \ScanLink105[27] , \ScanLink105[26] , 
        \ScanLink105[25] , \ScanLink105[24] , \ScanLink105[23] , 
        \ScanLink105[22] , \ScanLink105[21] , \ScanLink105[20] , 
        \ScanLink105[19] , \ScanLink105[18] , \ScanLink105[17] , 
        \ScanLink105[16] , \ScanLink105[15] , \ScanLink105[14] , 
        \ScanLink105[13] , \ScanLink105[12] , \ScanLink105[11] , 
        \ScanLink105[10] , \ScanLink105[9] , \ScanLink105[8] , 
        \ScanLink105[7] , \ScanLink105[6] , \ScanLink105[5] , \ScanLink105[4] , 
        \ScanLink105[3] , \ScanLink105[2] , \ScanLink105[1] , \ScanLink105[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_42[31] , 
        \wRegOut_6_42[30] , \wRegOut_6_42[29] , \wRegOut_6_42[28] , 
        \wRegOut_6_42[27] , \wRegOut_6_42[26] , \wRegOut_6_42[25] , 
        \wRegOut_6_42[24] , \wRegOut_6_42[23] , \wRegOut_6_42[22] , 
        \wRegOut_6_42[21] , \wRegOut_6_42[20] , \wRegOut_6_42[19] , 
        \wRegOut_6_42[18] , \wRegOut_6_42[17] , \wRegOut_6_42[16] , 
        \wRegOut_6_42[15] , \wRegOut_6_42[14] , \wRegOut_6_42[13] , 
        \wRegOut_6_42[12] , \wRegOut_6_42[11] , \wRegOut_6_42[10] , 
        \wRegOut_6_42[9] , \wRegOut_6_42[8] , \wRegOut_6_42[7] , 
        \wRegOut_6_42[6] , \wRegOut_6_42[5] , \wRegOut_6_42[4] , 
        \wRegOut_6_42[3] , \wRegOut_6_42[2] , \wRegOut_6_42[1] , 
        \wRegOut_6_42[0] }), .Enable1(\wRegEnTop_6_42[0] ), .Enable2(
        \wRegEnBot_6_42[0] ), .In1({\wRegInTop_6_42[31] , \wRegInTop_6_42[30] , 
        \wRegInTop_6_42[29] , \wRegInTop_6_42[28] , \wRegInTop_6_42[27] , 
        \wRegInTop_6_42[26] , \wRegInTop_6_42[25] , \wRegInTop_6_42[24] , 
        \wRegInTop_6_42[23] , \wRegInTop_6_42[22] , \wRegInTop_6_42[21] , 
        \wRegInTop_6_42[20] , \wRegInTop_6_42[19] , \wRegInTop_6_42[18] , 
        \wRegInTop_6_42[17] , \wRegInTop_6_42[16] , \wRegInTop_6_42[15] , 
        \wRegInTop_6_42[14] , \wRegInTop_6_42[13] , \wRegInTop_6_42[12] , 
        \wRegInTop_6_42[11] , \wRegInTop_6_42[10] , \wRegInTop_6_42[9] , 
        \wRegInTop_6_42[8] , \wRegInTop_6_42[7] , \wRegInTop_6_42[6] , 
        \wRegInTop_6_42[5] , \wRegInTop_6_42[4] , \wRegInTop_6_42[3] , 
        \wRegInTop_6_42[2] , \wRegInTop_6_42[1] , \wRegInTop_6_42[0] }), .In2(
        {\wRegInBot_6_42[31] , \wRegInBot_6_42[30] , \wRegInBot_6_42[29] , 
        \wRegInBot_6_42[28] , \wRegInBot_6_42[27] , \wRegInBot_6_42[26] , 
        \wRegInBot_6_42[25] , \wRegInBot_6_42[24] , \wRegInBot_6_42[23] , 
        \wRegInBot_6_42[22] , \wRegInBot_6_42[21] , \wRegInBot_6_42[20] , 
        \wRegInBot_6_42[19] , \wRegInBot_6_42[18] , \wRegInBot_6_42[17] , 
        \wRegInBot_6_42[16] , \wRegInBot_6_42[15] , \wRegInBot_6_42[14] , 
        \wRegInBot_6_42[13] , \wRegInBot_6_42[12] , \wRegInBot_6_42[11] , 
        \wRegInBot_6_42[10] , \wRegInBot_6_42[9] , \wRegInBot_6_42[8] , 
        \wRegInBot_6_42[7] , \wRegInBot_6_42[6] , \wRegInBot_6_42[5] , 
        \wRegInBot_6_42[4] , \wRegInBot_6_42[3] , \wRegInBot_6_42[2] , 
        \wRegInBot_6_42[1] , \wRegInBot_6_42[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_59 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink123[31] , \ScanLink123[30] , \ScanLink123[29] , 
        \ScanLink123[28] , \ScanLink123[27] , \ScanLink123[26] , 
        \ScanLink123[25] , \ScanLink123[24] , \ScanLink123[23] , 
        \ScanLink123[22] , \ScanLink123[21] , \ScanLink123[20] , 
        \ScanLink123[19] , \ScanLink123[18] , \ScanLink123[17] , 
        \ScanLink123[16] , \ScanLink123[15] , \ScanLink123[14] , 
        \ScanLink123[13] , \ScanLink123[12] , \ScanLink123[11] , 
        \ScanLink123[10] , \ScanLink123[9] , \ScanLink123[8] , 
        \ScanLink123[7] , \ScanLink123[6] , \ScanLink123[5] , \ScanLink123[4] , 
        \ScanLink123[3] , \ScanLink123[2] , \ScanLink123[1] , \ScanLink123[0] 
        }), .ScanOut({\ScanLink122[31] , \ScanLink122[30] , \ScanLink122[29] , 
        \ScanLink122[28] , \ScanLink122[27] , \ScanLink122[26] , 
        \ScanLink122[25] , \ScanLink122[24] , \ScanLink122[23] , 
        \ScanLink122[22] , \ScanLink122[21] , \ScanLink122[20] , 
        \ScanLink122[19] , \ScanLink122[18] , \ScanLink122[17] , 
        \ScanLink122[16] , \ScanLink122[15] , \ScanLink122[14] , 
        \ScanLink122[13] , \ScanLink122[12] , \ScanLink122[11] , 
        \ScanLink122[10] , \ScanLink122[9] , \ScanLink122[8] , 
        \ScanLink122[7] , \ScanLink122[6] , \ScanLink122[5] , \ScanLink122[4] , 
        \ScanLink122[3] , \ScanLink122[2] , \ScanLink122[1] , \ScanLink122[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_59[31] , 
        \wRegOut_6_59[30] , \wRegOut_6_59[29] , \wRegOut_6_59[28] , 
        \wRegOut_6_59[27] , \wRegOut_6_59[26] , \wRegOut_6_59[25] , 
        \wRegOut_6_59[24] , \wRegOut_6_59[23] , \wRegOut_6_59[22] , 
        \wRegOut_6_59[21] , \wRegOut_6_59[20] , \wRegOut_6_59[19] , 
        \wRegOut_6_59[18] , \wRegOut_6_59[17] , \wRegOut_6_59[16] , 
        \wRegOut_6_59[15] , \wRegOut_6_59[14] , \wRegOut_6_59[13] , 
        \wRegOut_6_59[12] , \wRegOut_6_59[11] , \wRegOut_6_59[10] , 
        \wRegOut_6_59[9] , \wRegOut_6_59[8] , \wRegOut_6_59[7] , 
        \wRegOut_6_59[6] , \wRegOut_6_59[5] , \wRegOut_6_59[4] , 
        \wRegOut_6_59[3] , \wRegOut_6_59[2] , \wRegOut_6_59[1] , 
        \wRegOut_6_59[0] }), .Enable1(\wRegEnTop_6_59[0] ), .Enable2(
        \wRegEnBot_6_59[0] ), .In1({\wRegInTop_6_59[31] , \wRegInTop_6_59[30] , 
        \wRegInTop_6_59[29] , \wRegInTop_6_59[28] , \wRegInTop_6_59[27] , 
        \wRegInTop_6_59[26] , \wRegInTop_6_59[25] , \wRegInTop_6_59[24] , 
        \wRegInTop_6_59[23] , \wRegInTop_6_59[22] , \wRegInTop_6_59[21] , 
        \wRegInTop_6_59[20] , \wRegInTop_6_59[19] , \wRegInTop_6_59[18] , 
        \wRegInTop_6_59[17] , \wRegInTop_6_59[16] , \wRegInTop_6_59[15] , 
        \wRegInTop_6_59[14] , \wRegInTop_6_59[13] , \wRegInTop_6_59[12] , 
        \wRegInTop_6_59[11] , \wRegInTop_6_59[10] , \wRegInTop_6_59[9] , 
        \wRegInTop_6_59[8] , \wRegInTop_6_59[7] , \wRegInTop_6_59[6] , 
        \wRegInTop_6_59[5] , \wRegInTop_6_59[4] , \wRegInTop_6_59[3] , 
        \wRegInTop_6_59[2] , \wRegInTop_6_59[1] , \wRegInTop_6_59[0] }), .In2(
        {\wRegInBot_6_59[31] , \wRegInBot_6_59[30] , \wRegInBot_6_59[29] , 
        \wRegInBot_6_59[28] , \wRegInBot_6_59[27] , \wRegInBot_6_59[26] , 
        \wRegInBot_6_59[25] , \wRegInBot_6_59[24] , \wRegInBot_6_59[23] , 
        \wRegInBot_6_59[22] , \wRegInBot_6_59[21] , \wRegInBot_6_59[20] , 
        \wRegInBot_6_59[19] , \wRegInBot_6_59[18] , \wRegInBot_6_59[17] , 
        \wRegInBot_6_59[16] , \wRegInBot_6_59[15] , \wRegInBot_6_59[14] , 
        \wRegInBot_6_59[13] , \wRegInBot_6_59[12] , \wRegInBot_6_59[11] , 
        \wRegInBot_6_59[10] , \wRegInBot_6_59[9] , \wRegInBot_6_59[8] , 
        \wRegInBot_6_59[7] , \wRegInBot_6_59[6] , \wRegInBot_6_59[5] , 
        \wRegInBot_6_59[4] , \wRegInBot_6_59[3] , \wRegInBot_6_59[2] , 
        \wRegInBot_6_59[1] , \wRegInBot_6_59[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_81 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink209[31] , \ScanLink209[30] , \ScanLink209[29] , 
        \ScanLink209[28] , \ScanLink209[27] , \ScanLink209[26] , 
        \ScanLink209[25] , \ScanLink209[24] , \ScanLink209[23] , 
        \ScanLink209[22] , \ScanLink209[21] , \ScanLink209[20] , 
        \ScanLink209[19] , \ScanLink209[18] , \ScanLink209[17] , 
        \ScanLink209[16] , \ScanLink209[15] , \ScanLink209[14] , 
        \ScanLink209[13] , \ScanLink209[12] , \ScanLink209[11] , 
        \ScanLink209[10] , \ScanLink209[9] , \ScanLink209[8] , 
        \ScanLink209[7] , \ScanLink209[6] , \ScanLink209[5] , \ScanLink209[4] , 
        \ScanLink209[3] , \ScanLink209[2] , \ScanLink209[1] , \ScanLink209[0] 
        }), .ScanOut({\ScanLink208[31] , \ScanLink208[30] , \ScanLink208[29] , 
        \ScanLink208[28] , \ScanLink208[27] , \ScanLink208[26] , 
        \ScanLink208[25] , \ScanLink208[24] , \ScanLink208[23] , 
        \ScanLink208[22] , \ScanLink208[21] , \ScanLink208[20] , 
        \ScanLink208[19] , \ScanLink208[18] , \ScanLink208[17] , 
        \ScanLink208[16] , \ScanLink208[15] , \ScanLink208[14] , 
        \ScanLink208[13] , \ScanLink208[12] , \ScanLink208[11] , 
        \ScanLink208[10] , \ScanLink208[9] , \ScanLink208[8] , 
        \ScanLink208[7] , \ScanLink208[6] , \ScanLink208[5] , \ScanLink208[4] , 
        \ScanLink208[3] , \ScanLink208[2] , \ScanLink208[1] , \ScanLink208[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_81[31] , 
        \wRegOut_7_81[30] , \wRegOut_7_81[29] , \wRegOut_7_81[28] , 
        \wRegOut_7_81[27] , \wRegOut_7_81[26] , \wRegOut_7_81[25] , 
        \wRegOut_7_81[24] , \wRegOut_7_81[23] , \wRegOut_7_81[22] , 
        \wRegOut_7_81[21] , \wRegOut_7_81[20] , \wRegOut_7_81[19] , 
        \wRegOut_7_81[18] , \wRegOut_7_81[17] , \wRegOut_7_81[16] , 
        \wRegOut_7_81[15] , \wRegOut_7_81[14] , \wRegOut_7_81[13] , 
        \wRegOut_7_81[12] , \wRegOut_7_81[11] , \wRegOut_7_81[10] , 
        \wRegOut_7_81[9] , \wRegOut_7_81[8] , \wRegOut_7_81[7] , 
        \wRegOut_7_81[6] , \wRegOut_7_81[5] , \wRegOut_7_81[4] , 
        \wRegOut_7_81[3] , \wRegOut_7_81[2] , \wRegOut_7_81[1] , 
        \wRegOut_7_81[0] }), .Enable1(\wRegEnTop_7_81[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_81[31] , \wRegInTop_7_81[30] , \wRegInTop_7_81[29] , 
        \wRegInTop_7_81[28] , \wRegInTop_7_81[27] , \wRegInTop_7_81[26] , 
        \wRegInTop_7_81[25] , \wRegInTop_7_81[24] , \wRegInTop_7_81[23] , 
        \wRegInTop_7_81[22] , \wRegInTop_7_81[21] , \wRegInTop_7_81[20] , 
        \wRegInTop_7_81[19] , \wRegInTop_7_81[18] , \wRegInTop_7_81[17] , 
        \wRegInTop_7_81[16] , \wRegInTop_7_81[15] , \wRegInTop_7_81[14] , 
        \wRegInTop_7_81[13] , \wRegInTop_7_81[12] , \wRegInTop_7_81[11] , 
        \wRegInTop_7_81[10] , \wRegInTop_7_81[9] , \wRegInTop_7_81[8] , 
        \wRegInTop_7_81[7] , \wRegInTop_7_81[6] , \wRegInTop_7_81[5] , 
        \wRegInTop_7_81[4] , \wRegInTop_7_81[3] , \wRegInTop_7_81[2] , 
        \wRegInTop_7_81[1] , \wRegInTop_7_81[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_1[0] ), .P_In({\wRegOut_3_1[31] , 
        \wRegOut_3_1[30] , \wRegOut_3_1[29] , \wRegOut_3_1[28] , 
        \wRegOut_3_1[27] , \wRegOut_3_1[26] , \wRegOut_3_1[25] , 
        \wRegOut_3_1[24] , \wRegOut_3_1[23] , \wRegOut_3_1[22] , 
        \wRegOut_3_1[21] , \wRegOut_3_1[20] , \wRegOut_3_1[19] , 
        \wRegOut_3_1[18] , \wRegOut_3_1[17] , \wRegOut_3_1[16] , 
        \wRegOut_3_1[15] , \wRegOut_3_1[14] , \wRegOut_3_1[13] , 
        \wRegOut_3_1[12] , \wRegOut_3_1[11] , \wRegOut_3_1[10] , 
        \wRegOut_3_1[9] , \wRegOut_3_1[8] , \wRegOut_3_1[7] , \wRegOut_3_1[6] , 
        \wRegOut_3_1[5] , \wRegOut_3_1[4] , \wRegOut_3_1[3] , \wRegOut_3_1[2] , 
        \wRegOut_3_1[1] , \wRegOut_3_1[0] }), .P_Out({\wRegInBot_3_1[31] , 
        \wRegInBot_3_1[30] , \wRegInBot_3_1[29] , \wRegInBot_3_1[28] , 
        \wRegInBot_3_1[27] , \wRegInBot_3_1[26] , \wRegInBot_3_1[25] , 
        \wRegInBot_3_1[24] , \wRegInBot_3_1[23] , \wRegInBot_3_1[22] , 
        \wRegInBot_3_1[21] , \wRegInBot_3_1[20] , \wRegInBot_3_1[19] , 
        \wRegInBot_3_1[18] , \wRegInBot_3_1[17] , \wRegInBot_3_1[16] , 
        \wRegInBot_3_1[15] , \wRegInBot_3_1[14] , \wRegInBot_3_1[13] , 
        \wRegInBot_3_1[12] , \wRegInBot_3_1[11] , \wRegInBot_3_1[10] , 
        \wRegInBot_3_1[9] , \wRegInBot_3_1[8] , \wRegInBot_3_1[7] , 
        \wRegInBot_3_1[6] , \wRegInBot_3_1[5] , \wRegInBot_3_1[4] , 
        \wRegInBot_3_1[3] , \wRegInBot_3_1[2] , \wRegInBot_3_1[1] , 
        \wRegInBot_3_1[0] }), .L_WR(\wRegEnTop_4_2[0] ), .L_In({
        \wRegOut_4_2[31] , \wRegOut_4_2[30] , \wRegOut_4_2[29] , 
        \wRegOut_4_2[28] , \wRegOut_4_2[27] , \wRegOut_4_2[26] , 
        \wRegOut_4_2[25] , \wRegOut_4_2[24] , \wRegOut_4_2[23] , 
        \wRegOut_4_2[22] , \wRegOut_4_2[21] , \wRegOut_4_2[20] , 
        \wRegOut_4_2[19] , \wRegOut_4_2[18] , \wRegOut_4_2[17] , 
        \wRegOut_4_2[16] , \wRegOut_4_2[15] , \wRegOut_4_2[14] , 
        \wRegOut_4_2[13] , \wRegOut_4_2[12] , \wRegOut_4_2[11] , 
        \wRegOut_4_2[10] , \wRegOut_4_2[9] , \wRegOut_4_2[8] , 
        \wRegOut_4_2[7] , \wRegOut_4_2[6] , \wRegOut_4_2[5] , \wRegOut_4_2[4] , 
        \wRegOut_4_2[3] , \wRegOut_4_2[2] , \wRegOut_4_2[1] , \wRegOut_4_2[0] 
        }), .L_Out({\wRegInTop_4_2[31] , \wRegInTop_4_2[30] , 
        \wRegInTop_4_2[29] , \wRegInTop_4_2[28] , \wRegInTop_4_2[27] , 
        \wRegInTop_4_2[26] , \wRegInTop_4_2[25] , \wRegInTop_4_2[24] , 
        \wRegInTop_4_2[23] , \wRegInTop_4_2[22] , \wRegInTop_4_2[21] , 
        \wRegInTop_4_2[20] , \wRegInTop_4_2[19] , \wRegInTop_4_2[18] , 
        \wRegInTop_4_2[17] , \wRegInTop_4_2[16] , \wRegInTop_4_2[15] , 
        \wRegInTop_4_2[14] , \wRegInTop_4_2[13] , \wRegInTop_4_2[12] , 
        \wRegInTop_4_2[11] , \wRegInTop_4_2[10] , \wRegInTop_4_2[9] , 
        \wRegInTop_4_2[8] , \wRegInTop_4_2[7] , \wRegInTop_4_2[6] , 
        \wRegInTop_4_2[5] , \wRegInTop_4_2[4] , \wRegInTop_4_2[3] , 
        \wRegInTop_4_2[2] , \wRegInTop_4_2[1] , \wRegInTop_4_2[0] }), .R_WR(
        \wRegEnTop_4_3[0] ), .R_In({\wRegOut_4_3[31] , \wRegOut_4_3[30] , 
        \wRegOut_4_3[29] , \wRegOut_4_3[28] , \wRegOut_4_3[27] , 
        \wRegOut_4_3[26] , \wRegOut_4_3[25] , \wRegOut_4_3[24] , 
        \wRegOut_4_3[23] , \wRegOut_4_3[22] , \wRegOut_4_3[21] , 
        \wRegOut_4_3[20] , \wRegOut_4_3[19] , \wRegOut_4_3[18] , 
        \wRegOut_4_3[17] , \wRegOut_4_3[16] , \wRegOut_4_3[15] , 
        \wRegOut_4_3[14] , \wRegOut_4_3[13] , \wRegOut_4_3[12] , 
        \wRegOut_4_3[11] , \wRegOut_4_3[10] , \wRegOut_4_3[9] , 
        \wRegOut_4_3[8] , \wRegOut_4_3[7] , \wRegOut_4_3[6] , \wRegOut_4_3[5] , 
        \wRegOut_4_3[4] , \wRegOut_4_3[3] , \wRegOut_4_3[2] , \wRegOut_4_3[1] , 
        \wRegOut_4_3[0] }), .R_Out({\wRegInTop_4_3[31] , \wRegInTop_4_3[30] , 
        \wRegInTop_4_3[29] , \wRegInTop_4_3[28] , \wRegInTop_4_3[27] , 
        \wRegInTop_4_3[26] , \wRegInTop_4_3[25] , \wRegInTop_4_3[24] , 
        \wRegInTop_4_3[23] , \wRegInTop_4_3[22] , \wRegInTop_4_3[21] , 
        \wRegInTop_4_3[20] , \wRegInTop_4_3[19] , \wRegInTop_4_3[18] , 
        \wRegInTop_4_3[17] , \wRegInTop_4_3[16] , \wRegInTop_4_3[15] , 
        \wRegInTop_4_3[14] , \wRegInTop_4_3[13] , \wRegInTop_4_3[12] , 
        \wRegInTop_4_3[11] , \wRegInTop_4_3[10] , \wRegInTop_4_3[9] , 
        \wRegInTop_4_3[8] , \wRegInTop_4_3[7] , \wRegInTop_4_3[6] , 
        \wRegInTop_4_3[5] , \wRegInTop_4_3[4] , \wRegInTop_4_3[3] , 
        \wRegInTop_4_3[2] , \wRegInTop_4_3[1] , \wRegInTop_4_3[0] }) );
    BHeap_Node_WIDTH32 BHN_4_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_12[0] ), .P_In({\wRegOut_4_12[31] , 
        \wRegOut_4_12[30] , \wRegOut_4_12[29] , \wRegOut_4_12[28] , 
        \wRegOut_4_12[27] , \wRegOut_4_12[26] , \wRegOut_4_12[25] , 
        \wRegOut_4_12[24] , \wRegOut_4_12[23] , \wRegOut_4_12[22] , 
        \wRegOut_4_12[21] , \wRegOut_4_12[20] , \wRegOut_4_12[19] , 
        \wRegOut_4_12[18] , \wRegOut_4_12[17] , \wRegOut_4_12[16] , 
        \wRegOut_4_12[15] , \wRegOut_4_12[14] , \wRegOut_4_12[13] , 
        \wRegOut_4_12[12] , \wRegOut_4_12[11] , \wRegOut_4_12[10] , 
        \wRegOut_4_12[9] , \wRegOut_4_12[8] , \wRegOut_4_12[7] , 
        \wRegOut_4_12[6] , \wRegOut_4_12[5] , \wRegOut_4_12[4] , 
        \wRegOut_4_12[3] , \wRegOut_4_12[2] , \wRegOut_4_12[1] , 
        \wRegOut_4_12[0] }), .P_Out({\wRegInBot_4_12[31] , 
        \wRegInBot_4_12[30] , \wRegInBot_4_12[29] , \wRegInBot_4_12[28] , 
        \wRegInBot_4_12[27] , \wRegInBot_4_12[26] , \wRegInBot_4_12[25] , 
        \wRegInBot_4_12[24] , \wRegInBot_4_12[23] , \wRegInBot_4_12[22] , 
        \wRegInBot_4_12[21] , \wRegInBot_4_12[20] , \wRegInBot_4_12[19] , 
        \wRegInBot_4_12[18] , \wRegInBot_4_12[17] , \wRegInBot_4_12[16] , 
        \wRegInBot_4_12[15] , \wRegInBot_4_12[14] , \wRegInBot_4_12[13] , 
        \wRegInBot_4_12[12] , \wRegInBot_4_12[11] , \wRegInBot_4_12[10] , 
        \wRegInBot_4_12[9] , \wRegInBot_4_12[8] , \wRegInBot_4_12[7] , 
        \wRegInBot_4_12[6] , \wRegInBot_4_12[5] , \wRegInBot_4_12[4] , 
        \wRegInBot_4_12[3] , \wRegInBot_4_12[2] , \wRegInBot_4_12[1] , 
        \wRegInBot_4_12[0] }), .L_WR(\wRegEnTop_5_24[0] ), .L_In({
        \wRegOut_5_24[31] , \wRegOut_5_24[30] , \wRegOut_5_24[29] , 
        \wRegOut_5_24[28] , \wRegOut_5_24[27] , \wRegOut_5_24[26] , 
        \wRegOut_5_24[25] , \wRegOut_5_24[24] , \wRegOut_5_24[23] , 
        \wRegOut_5_24[22] , \wRegOut_5_24[21] , \wRegOut_5_24[20] , 
        \wRegOut_5_24[19] , \wRegOut_5_24[18] , \wRegOut_5_24[17] , 
        \wRegOut_5_24[16] , \wRegOut_5_24[15] , \wRegOut_5_24[14] , 
        \wRegOut_5_24[13] , \wRegOut_5_24[12] , \wRegOut_5_24[11] , 
        \wRegOut_5_24[10] , \wRegOut_5_24[9] , \wRegOut_5_24[8] , 
        \wRegOut_5_24[7] , \wRegOut_5_24[6] , \wRegOut_5_24[5] , 
        \wRegOut_5_24[4] , \wRegOut_5_24[3] , \wRegOut_5_24[2] , 
        \wRegOut_5_24[1] , \wRegOut_5_24[0] }), .L_Out({\wRegInTop_5_24[31] , 
        \wRegInTop_5_24[30] , \wRegInTop_5_24[29] , \wRegInTop_5_24[28] , 
        \wRegInTop_5_24[27] , \wRegInTop_5_24[26] , \wRegInTop_5_24[25] , 
        \wRegInTop_5_24[24] , \wRegInTop_5_24[23] , \wRegInTop_5_24[22] , 
        \wRegInTop_5_24[21] , \wRegInTop_5_24[20] , \wRegInTop_5_24[19] , 
        \wRegInTop_5_24[18] , \wRegInTop_5_24[17] , \wRegInTop_5_24[16] , 
        \wRegInTop_5_24[15] , \wRegInTop_5_24[14] , \wRegInTop_5_24[13] , 
        \wRegInTop_5_24[12] , \wRegInTop_5_24[11] , \wRegInTop_5_24[10] , 
        \wRegInTop_5_24[9] , \wRegInTop_5_24[8] , \wRegInTop_5_24[7] , 
        \wRegInTop_5_24[6] , \wRegInTop_5_24[5] , \wRegInTop_5_24[4] , 
        \wRegInTop_5_24[3] , \wRegInTop_5_24[2] , \wRegInTop_5_24[1] , 
        \wRegInTop_5_24[0] }), .R_WR(\wRegEnTop_5_25[0] ), .R_In({
        \wRegOut_5_25[31] , \wRegOut_5_25[30] , \wRegOut_5_25[29] , 
        \wRegOut_5_25[28] , \wRegOut_5_25[27] , \wRegOut_5_25[26] , 
        \wRegOut_5_25[25] , \wRegOut_5_25[24] , \wRegOut_5_25[23] , 
        \wRegOut_5_25[22] , \wRegOut_5_25[21] , \wRegOut_5_25[20] , 
        \wRegOut_5_25[19] , \wRegOut_5_25[18] , \wRegOut_5_25[17] , 
        \wRegOut_5_25[16] , \wRegOut_5_25[15] , \wRegOut_5_25[14] , 
        \wRegOut_5_25[13] , \wRegOut_5_25[12] , \wRegOut_5_25[11] , 
        \wRegOut_5_25[10] , \wRegOut_5_25[9] , \wRegOut_5_25[8] , 
        \wRegOut_5_25[7] , \wRegOut_5_25[6] , \wRegOut_5_25[5] , 
        \wRegOut_5_25[4] , \wRegOut_5_25[3] , \wRegOut_5_25[2] , 
        \wRegOut_5_25[1] , \wRegOut_5_25[0] }), .R_Out({\wRegInTop_5_25[31] , 
        \wRegInTop_5_25[30] , \wRegInTop_5_25[29] , \wRegInTop_5_25[28] , 
        \wRegInTop_5_25[27] , \wRegInTop_5_25[26] , \wRegInTop_5_25[25] , 
        \wRegInTop_5_25[24] , \wRegInTop_5_25[23] , \wRegInTop_5_25[22] , 
        \wRegInTop_5_25[21] , \wRegInTop_5_25[20] , \wRegInTop_5_25[19] , 
        \wRegInTop_5_25[18] , \wRegInTop_5_25[17] , \wRegInTop_5_25[16] , 
        \wRegInTop_5_25[15] , \wRegInTop_5_25[14] , \wRegInTop_5_25[13] , 
        \wRegInTop_5_25[12] , \wRegInTop_5_25[11] , \wRegInTop_5_25[10] , 
        \wRegInTop_5_25[9] , \wRegInTop_5_25[8] , \wRegInTop_5_25[7] , 
        \wRegInTop_5_25[6] , \wRegInTop_5_25[5] , \wRegInTop_5_25[4] , 
        \wRegInTop_5_25[3] , \wRegInTop_5_25[2] , \wRegInTop_5_25[1] , 
        \wRegInTop_5_25[0] }) );
    BHeap_Node_WIDTH32 BHN_6_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_7[0] ), .P_In({\wRegOut_6_7[31] , 
        \wRegOut_6_7[30] , \wRegOut_6_7[29] , \wRegOut_6_7[28] , 
        \wRegOut_6_7[27] , \wRegOut_6_7[26] , \wRegOut_6_7[25] , 
        \wRegOut_6_7[24] , \wRegOut_6_7[23] , \wRegOut_6_7[22] , 
        \wRegOut_6_7[21] , \wRegOut_6_7[20] , \wRegOut_6_7[19] , 
        \wRegOut_6_7[18] , \wRegOut_6_7[17] , \wRegOut_6_7[16] , 
        \wRegOut_6_7[15] , \wRegOut_6_7[14] , \wRegOut_6_7[13] , 
        \wRegOut_6_7[12] , \wRegOut_6_7[11] , \wRegOut_6_7[10] , 
        \wRegOut_6_7[9] , \wRegOut_6_7[8] , \wRegOut_6_7[7] , \wRegOut_6_7[6] , 
        \wRegOut_6_7[5] , \wRegOut_6_7[4] , \wRegOut_6_7[3] , \wRegOut_6_7[2] , 
        \wRegOut_6_7[1] , \wRegOut_6_7[0] }), .P_Out({\wRegInBot_6_7[31] , 
        \wRegInBot_6_7[30] , \wRegInBot_6_7[29] , \wRegInBot_6_7[28] , 
        \wRegInBot_6_7[27] , \wRegInBot_6_7[26] , \wRegInBot_6_7[25] , 
        \wRegInBot_6_7[24] , \wRegInBot_6_7[23] , \wRegInBot_6_7[22] , 
        \wRegInBot_6_7[21] , \wRegInBot_6_7[20] , \wRegInBot_6_7[19] , 
        \wRegInBot_6_7[18] , \wRegInBot_6_7[17] , \wRegInBot_6_7[16] , 
        \wRegInBot_6_7[15] , \wRegInBot_6_7[14] , \wRegInBot_6_7[13] , 
        \wRegInBot_6_7[12] , \wRegInBot_6_7[11] , \wRegInBot_6_7[10] , 
        \wRegInBot_6_7[9] , \wRegInBot_6_7[8] , \wRegInBot_6_7[7] , 
        \wRegInBot_6_7[6] , \wRegInBot_6_7[5] , \wRegInBot_6_7[4] , 
        \wRegInBot_6_7[3] , \wRegInBot_6_7[2] , \wRegInBot_6_7[1] , 
        \wRegInBot_6_7[0] }), .L_WR(\wRegEnTop_7_14[0] ), .L_In({
        \wRegOut_7_14[31] , \wRegOut_7_14[30] , \wRegOut_7_14[29] , 
        \wRegOut_7_14[28] , \wRegOut_7_14[27] , \wRegOut_7_14[26] , 
        \wRegOut_7_14[25] , \wRegOut_7_14[24] , \wRegOut_7_14[23] , 
        \wRegOut_7_14[22] , \wRegOut_7_14[21] , \wRegOut_7_14[20] , 
        \wRegOut_7_14[19] , \wRegOut_7_14[18] , \wRegOut_7_14[17] , 
        \wRegOut_7_14[16] , \wRegOut_7_14[15] , \wRegOut_7_14[14] , 
        \wRegOut_7_14[13] , \wRegOut_7_14[12] , \wRegOut_7_14[11] , 
        \wRegOut_7_14[10] , \wRegOut_7_14[9] , \wRegOut_7_14[8] , 
        \wRegOut_7_14[7] , \wRegOut_7_14[6] , \wRegOut_7_14[5] , 
        \wRegOut_7_14[4] , \wRegOut_7_14[3] , \wRegOut_7_14[2] , 
        \wRegOut_7_14[1] , \wRegOut_7_14[0] }), .L_Out({\wRegInTop_7_14[31] , 
        \wRegInTop_7_14[30] , \wRegInTop_7_14[29] , \wRegInTop_7_14[28] , 
        \wRegInTop_7_14[27] , \wRegInTop_7_14[26] , \wRegInTop_7_14[25] , 
        \wRegInTop_7_14[24] , \wRegInTop_7_14[23] , \wRegInTop_7_14[22] , 
        \wRegInTop_7_14[21] , \wRegInTop_7_14[20] , \wRegInTop_7_14[19] , 
        \wRegInTop_7_14[18] , \wRegInTop_7_14[17] , \wRegInTop_7_14[16] , 
        \wRegInTop_7_14[15] , \wRegInTop_7_14[14] , \wRegInTop_7_14[13] , 
        \wRegInTop_7_14[12] , \wRegInTop_7_14[11] , \wRegInTop_7_14[10] , 
        \wRegInTop_7_14[9] , \wRegInTop_7_14[8] , \wRegInTop_7_14[7] , 
        \wRegInTop_7_14[6] , \wRegInTop_7_14[5] , \wRegInTop_7_14[4] , 
        \wRegInTop_7_14[3] , \wRegInTop_7_14[2] , \wRegInTop_7_14[1] , 
        \wRegInTop_7_14[0] }), .R_WR(\wRegEnTop_7_15[0] ), .R_In({
        \wRegOut_7_15[31] , \wRegOut_7_15[30] , \wRegOut_7_15[29] , 
        \wRegOut_7_15[28] , \wRegOut_7_15[27] , \wRegOut_7_15[26] , 
        \wRegOut_7_15[25] , \wRegOut_7_15[24] , \wRegOut_7_15[23] , 
        \wRegOut_7_15[22] , \wRegOut_7_15[21] , \wRegOut_7_15[20] , 
        \wRegOut_7_15[19] , \wRegOut_7_15[18] , \wRegOut_7_15[17] , 
        \wRegOut_7_15[16] , \wRegOut_7_15[15] , \wRegOut_7_15[14] , 
        \wRegOut_7_15[13] , \wRegOut_7_15[12] , \wRegOut_7_15[11] , 
        \wRegOut_7_15[10] , \wRegOut_7_15[9] , \wRegOut_7_15[8] , 
        \wRegOut_7_15[7] , \wRegOut_7_15[6] , \wRegOut_7_15[5] , 
        \wRegOut_7_15[4] , \wRegOut_7_15[3] , \wRegOut_7_15[2] , 
        \wRegOut_7_15[1] , \wRegOut_7_15[0] }), .R_Out({\wRegInTop_7_15[31] , 
        \wRegInTop_7_15[30] , \wRegInTop_7_15[29] , \wRegInTop_7_15[28] , 
        \wRegInTop_7_15[27] , \wRegInTop_7_15[26] , \wRegInTop_7_15[25] , 
        \wRegInTop_7_15[24] , \wRegInTop_7_15[23] , \wRegInTop_7_15[22] , 
        \wRegInTop_7_15[21] , \wRegInTop_7_15[20] , \wRegInTop_7_15[19] , 
        \wRegInTop_7_15[18] , \wRegInTop_7_15[17] , \wRegInTop_7_15[16] , 
        \wRegInTop_7_15[15] , \wRegInTop_7_15[14] , \wRegInTop_7_15[13] , 
        \wRegInTop_7_15[12] , \wRegInTop_7_15[11] , \wRegInTop_7_15[10] , 
        \wRegInTop_7_15[9] , \wRegInTop_7_15[8] , \wRegInTop_7_15[7] , 
        \wRegInTop_7_15[6] , \wRegInTop_7_15[5] , \wRegInTop_7_15[4] , 
        \wRegInTop_7_15[3] , \wRegInTop_7_15[2] , \wRegInTop_7_15[1] , 
        \wRegInTop_7_15[0] }) );
    BHeap_Node_WIDTH32 BHN_6_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_56[0] ), .P_In({\wRegOut_6_56[31] , 
        \wRegOut_6_56[30] , \wRegOut_6_56[29] , \wRegOut_6_56[28] , 
        \wRegOut_6_56[27] , \wRegOut_6_56[26] , \wRegOut_6_56[25] , 
        \wRegOut_6_56[24] , \wRegOut_6_56[23] , \wRegOut_6_56[22] , 
        \wRegOut_6_56[21] , \wRegOut_6_56[20] , \wRegOut_6_56[19] , 
        \wRegOut_6_56[18] , \wRegOut_6_56[17] , \wRegOut_6_56[16] , 
        \wRegOut_6_56[15] , \wRegOut_6_56[14] , \wRegOut_6_56[13] , 
        \wRegOut_6_56[12] , \wRegOut_6_56[11] , \wRegOut_6_56[10] , 
        \wRegOut_6_56[9] , \wRegOut_6_56[8] , \wRegOut_6_56[7] , 
        \wRegOut_6_56[6] , \wRegOut_6_56[5] , \wRegOut_6_56[4] , 
        \wRegOut_6_56[3] , \wRegOut_6_56[2] , \wRegOut_6_56[1] , 
        \wRegOut_6_56[0] }), .P_Out({\wRegInBot_6_56[31] , 
        \wRegInBot_6_56[30] , \wRegInBot_6_56[29] , \wRegInBot_6_56[28] , 
        \wRegInBot_6_56[27] , \wRegInBot_6_56[26] , \wRegInBot_6_56[25] , 
        \wRegInBot_6_56[24] , \wRegInBot_6_56[23] , \wRegInBot_6_56[22] , 
        \wRegInBot_6_56[21] , \wRegInBot_6_56[20] , \wRegInBot_6_56[19] , 
        \wRegInBot_6_56[18] , \wRegInBot_6_56[17] , \wRegInBot_6_56[16] , 
        \wRegInBot_6_56[15] , \wRegInBot_6_56[14] , \wRegInBot_6_56[13] , 
        \wRegInBot_6_56[12] , \wRegInBot_6_56[11] , \wRegInBot_6_56[10] , 
        \wRegInBot_6_56[9] , \wRegInBot_6_56[8] , \wRegInBot_6_56[7] , 
        \wRegInBot_6_56[6] , \wRegInBot_6_56[5] , \wRegInBot_6_56[4] , 
        \wRegInBot_6_56[3] , \wRegInBot_6_56[2] , \wRegInBot_6_56[1] , 
        \wRegInBot_6_56[0] }), .L_WR(\wRegEnTop_7_112[0] ), .L_In({
        \wRegOut_7_112[31] , \wRegOut_7_112[30] , \wRegOut_7_112[29] , 
        \wRegOut_7_112[28] , \wRegOut_7_112[27] , \wRegOut_7_112[26] , 
        \wRegOut_7_112[25] , \wRegOut_7_112[24] , \wRegOut_7_112[23] , 
        \wRegOut_7_112[22] , \wRegOut_7_112[21] , \wRegOut_7_112[20] , 
        \wRegOut_7_112[19] , \wRegOut_7_112[18] , \wRegOut_7_112[17] , 
        \wRegOut_7_112[16] , \wRegOut_7_112[15] , \wRegOut_7_112[14] , 
        \wRegOut_7_112[13] , \wRegOut_7_112[12] , \wRegOut_7_112[11] , 
        \wRegOut_7_112[10] , \wRegOut_7_112[9] , \wRegOut_7_112[8] , 
        \wRegOut_7_112[7] , \wRegOut_7_112[6] , \wRegOut_7_112[5] , 
        \wRegOut_7_112[4] , \wRegOut_7_112[3] , \wRegOut_7_112[2] , 
        \wRegOut_7_112[1] , \wRegOut_7_112[0] }), .L_Out({
        \wRegInTop_7_112[31] , \wRegInTop_7_112[30] , \wRegInTop_7_112[29] , 
        \wRegInTop_7_112[28] , \wRegInTop_7_112[27] , \wRegInTop_7_112[26] , 
        \wRegInTop_7_112[25] , \wRegInTop_7_112[24] , \wRegInTop_7_112[23] , 
        \wRegInTop_7_112[22] , \wRegInTop_7_112[21] , \wRegInTop_7_112[20] , 
        \wRegInTop_7_112[19] , \wRegInTop_7_112[18] , \wRegInTop_7_112[17] , 
        \wRegInTop_7_112[16] , \wRegInTop_7_112[15] , \wRegInTop_7_112[14] , 
        \wRegInTop_7_112[13] , \wRegInTop_7_112[12] , \wRegInTop_7_112[11] , 
        \wRegInTop_7_112[10] , \wRegInTop_7_112[9] , \wRegInTop_7_112[8] , 
        \wRegInTop_7_112[7] , \wRegInTop_7_112[6] , \wRegInTop_7_112[5] , 
        \wRegInTop_7_112[4] , \wRegInTop_7_112[3] , \wRegInTop_7_112[2] , 
        \wRegInTop_7_112[1] , \wRegInTop_7_112[0] }), .R_WR(
        \wRegEnTop_7_113[0] ), .R_In({\wRegOut_7_113[31] , \wRegOut_7_113[30] , 
        \wRegOut_7_113[29] , \wRegOut_7_113[28] , \wRegOut_7_113[27] , 
        \wRegOut_7_113[26] , \wRegOut_7_113[25] , \wRegOut_7_113[24] , 
        \wRegOut_7_113[23] , \wRegOut_7_113[22] , \wRegOut_7_113[21] , 
        \wRegOut_7_113[20] , \wRegOut_7_113[19] , \wRegOut_7_113[18] , 
        \wRegOut_7_113[17] , \wRegOut_7_113[16] , \wRegOut_7_113[15] , 
        \wRegOut_7_113[14] , \wRegOut_7_113[13] , \wRegOut_7_113[12] , 
        \wRegOut_7_113[11] , \wRegOut_7_113[10] , \wRegOut_7_113[9] , 
        \wRegOut_7_113[8] , \wRegOut_7_113[7] , \wRegOut_7_113[6] , 
        \wRegOut_7_113[5] , \wRegOut_7_113[4] , \wRegOut_7_113[3] , 
        \wRegOut_7_113[2] , \wRegOut_7_113[1] , \wRegOut_7_113[0] }), .R_Out({
        \wRegInTop_7_113[31] , \wRegInTop_7_113[30] , \wRegInTop_7_113[29] , 
        \wRegInTop_7_113[28] , \wRegInTop_7_113[27] , \wRegInTop_7_113[26] , 
        \wRegInTop_7_113[25] , \wRegInTop_7_113[24] , \wRegInTop_7_113[23] , 
        \wRegInTop_7_113[22] , \wRegInTop_7_113[21] , \wRegInTop_7_113[20] , 
        \wRegInTop_7_113[19] , \wRegInTop_7_113[18] , \wRegInTop_7_113[17] , 
        \wRegInTop_7_113[16] , \wRegInTop_7_113[15] , \wRegInTop_7_113[14] , 
        \wRegInTop_7_113[13] , \wRegInTop_7_113[12] , \wRegInTop_7_113[11] , 
        \wRegInTop_7_113[10] , \wRegInTop_7_113[9] , \wRegInTop_7_113[8] , 
        \wRegInTop_7_113[7] , \wRegInTop_7_113[6] , \wRegInTop_7_113[5] , 
        \wRegInTop_7_113[4] , \wRegInTop_7_113[3] , \wRegInTop_7_113[2] , 
        \wRegInTop_7_113[1] , \wRegInTop_7_113[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_36 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink164[31] , \ScanLink164[30] , \ScanLink164[29] , 
        \ScanLink164[28] , \ScanLink164[27] , \ScanLink164[26] , 
        \ScanLink164[25] , \ScanLink164[24] , \ScanLink164[23] , 
        \ScanLink164[22] , \ScanLink164[21] , \ScanLink164[20] , 
        \ScanLink164[19] , \ScanLink164[18] , \ScanLink164[17] , 
        \ScanLink164[16] , \ScanLink164[15] , \ScanLink164[14] , 
        \ScanLink164[13] , \ScanLink164[12] , \ScanLink164[11] , 
        \ScanLink164[10] , \ScanLink164[9] , \ScanLink164[8] , 
        \ScanLink164[7] , \ScanLink164[6] , \ScanLink164[5] , \ScanLink164[4] , 
        \ScanLink164[3] , \ScanLink164[2] , \ScanLink164[1] , \ScanLink164[0] 
        }), .ScanOut({\ScanLink163[31] , \ScanLink163[30] , \ScanLink163[29] , 
        \ScanLink163[28] , \ScanLink163[27] , \ScanLink163[26] , 
        \ScanLink163[25] , \ScanLink163[24] , \ScanLink163[23] , 
        \ScanLink163[22] , \ScanLink163[21] , \ScanLink163[20] , 
        \ScanLink163[19] , \ScanLink163[18] , \ScanLink163[17] , 
        \ScanLink163[16] , \ScanLink163[15] , \ScanLink163[14] , 
        \ScanLink163[13] , \ScanLink163[12] , \ScanLink163[11] , 
        \ScanLink163[10] , \ScanLink163[9] , \ScanLink163[8] , 
        \ScanLink163[7] , \ScanLink163[6] , \ScanLink163[5] , \ScanLink163[4] , 
        \ScanLink163[3] , \ScanLink163[2] , \ScanLink163[1] , \ScanLink163[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_36[31] , 
        \wRegOut_7_36[30] , \wRegOut_7_36[29] , \wRegOut_7_36[28] , 
        \wRegOut_7_36[27] , \wRegOut_7_36[26] , \wRegOut_7_36[25] , 
        \wRegOut_7_36[24] , \wRegOut_7_36[23] , \wRegOut_7_36[22] , 
        \wRegOut_7_36[21] , \wRegOut_7_36[20] , \wRegOut_7_36[19] , 
        \wRegOut_7_36[18] , \wRegOut_7_36[17] , \wRegOut_7_36[16] , 
        \wRegOut_7_36[15] , \wRegOut_7_36[14] , \wRegOut_7_36[13] , 
        \wRegOut_7_36[12] , \wRegOut_7_36[11] , \wRegOut_7_36[10] , 
        \wRegOut_7_36[9] , \wRegOut_7_36[8] , \wRegOut_7_36[7] , 
        \wRegOut_7_36[6] , \wRegOut_7_36[5] , \wRegOut_7_36[4] , 
        \wRegOut_7_36[3] , \wRegOut_7_36[2] , \wRegOut_7_36[1] , 
        \wRegOut_7_36[0] }), .Enable1(\wRegEnTop_7_36[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_36[31] , \wRegInTop_7_36[30] , \wRegInTop_7_36[29] , 
        \wRegInTop_7_36[28] , \wRegInTop_7_36[27] , \wRegInTop_7_36[26] , 
        \wRegInTop_7_36[25] , \wRegInTop_7_36[24] , \wRegInTop_7_36[23] , 
        \wRegInTop_7_36[22] , \wRegInTop_7_36[21] , \wRegInTop_7_36[20] , 
        \wRegInTop_7_36[19] , \wRegInTop_7_36[18] , \wRegInTop_7_36[17] , 
        \wRegInTop_7_36[16] , \wRegInTop_7_36[15] , \wRegInTop_7_36[14] , 
        \wRegInTop_7_36[13] , \wRegInTop_7_36[12] , \wRegInTop_7_36[11] , 
        \wRegInTop_7_36[10] , \wRegInTop_7_36[9] , \wRegInTop_7_36[8] , 
        \wRegInTop_7_36[7] , \wRegInTop_7_36[6] , \wRegInTop_7_36[5] , 
        \wRegInTop_7_36[4] , \wRegInTop_7_36[3] , \wRegInTop_7_36[2] , 
        \wRegInTop_7_36[1] , \wRegInTop_7_36[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink139[31] , \ScanLink139[30] , \ScanLink139[29] , 
        \ScanLink139[28] , \ScanLink139[27] , \ScanLink139[26] , 
        \ScanLink139[25] , \ScanLink139[24] , \ScanLink139[23] , 
        \ScanLink139[22] , \ScanLink139[21] , \ScanLink139[20] , 
        \ScanLink139[19] , \ScanLink139[18] , \ScanLink139[17] , 
        \ScanLink139[16] , \ScanLink139[15] , \ScanLink139[14] , 
        \ScanLink139[13] , \ScanLink139[12] , \ScanLink139[11] , 
        \ScanLink139[10] , \ScanLink139[9] , \ScanLink139[8] , 
        \ScanLink139[7] , \ScanLink139[6] , \ScanLink139[5] , \ScanLink139[4] , 
        \ScanLink139[3] , \ScanLink139[2] , \ScanLink139[1] , \ScanLink139[0] 
        }), .ScanOut({\ScanLink138[31] , \ScanLink138[30] , \ScanLink138[29] , 
        \ScanLink138[28] , \ScanLink138[27] , \ScanLink138[26] , 
        \ScanLink138[25] , \ScanLink138[24] , \ScanLink138[23] , 
        \ScanLink138[22] , \ScanLink138[21] , \ScanLink138[20] , 
        \ScanLink138[19] , \ScanLink138[18] , \ScanLink138[17] , 
        \ScanLink138[16] , \ScanLink138[15] , \ScanLink138[14] , 
        \ScanLink138[13] , \ScanLink138[12] , \ScanLink138[11] , 
        \ScanLink138[10] , \ScanLink138[9] , \ScanLink138[8] , 
        \ScanLink138[7] , \ScanLink138[6] , \ScanLink138[5] , \ScanLink138[4] , 
        \ScanLink138[3] , \ScanLink138[2] , \ScanLink138[1] , \ScanLink138[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_11[31] , 
        \wRegOut_7_11[30] , \wRegOut_7_11[29] , \wRegOut_7_11[28] , 
        \wRegOut_7_11[27] , \wRegOut_7_11[26] , \wRegOut_7_11[25] , 
        \wRegOut_7_11[24] , \wRegOut_7_11[23] , \wRegOut_7_11[22] , 
        \wRegOut_7_11[21] , \wRegOut_7_11[20] , \wRegOut_7_11[19] , 
        \wRegOut_7_11[18] , \wRegOut_7_11[17] , \wRegOut_7_11[16] , 
        \wRegOut_7_11[15] , \wRegOut_7_11[14] , \wRegOut_7_11[13] , 
        \wRegOut_7_11[12] , \wRegOut_7_11[11] , \wRegOut_7_11[10] , 
        \wRegOut_7_11[9] , \wRegOut_7_11[8] , \wRegOut_7_11[7] , 
        \wRegOut_7_11[6] , \wRegOut_7_11[5] , \wRegOut_7_11[4] , 
        \wRegOut_7_11[3] , \wRegOut_7_11[2] , \wRegOut_7_11[1] , 
        \wRegOut_7_11[0] }), .Enable1(\wRegEnTop_7_11[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_11[31] , \wRegInTop_7_11[30] , \wRegInTop_7_11[29] , 
        \wRegInTop_7_11[28] , \wRegInTop_7_11[27] , \wRegInTop_7_11[26] , 
        \wRegInTop_7_11[25] , \wRegInTop_7_11[24] , \wRegInTop_7_11[23] , 
        \wRegInTop_7_11[22] , \wRegInTop_7_11[21] , \wRegInTop_7_11[20] , 
        \wRegInTop_7_11[19] , \wRegInTop_7_11[18] , \wRegInTop_7_11[17] , 
        \wRegInTop_7_11[16] , \wRegInTop_7_11[15] , \wRegInTop_7_11[14] , 
        \wRegInTop_7_11[13] , \wRegInTop_7_11[12] , \wRegInTop_7_11[11] , 
        \wRegInTop_7_11[10] , \wRegInTop_7_11[9] , \wRegInTop_7_11[8] , 
        \wRegInTop_7_11[7] , \wRegInTop_7_11[6] , \wRegInTop_7_11[5] , 
        \wRegInTop_7_11[4] , \wRegInTop_7_11[3] , \wRegInTop_7_11[2] , 
        \wRegInTop_7_11[1] , \wRegInTop_7_11[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_122 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink250[31] , \ScanLink250[30] , \ScanLink250[29] , 
        \ScanLink250[28] , \ScanLink250[27] , \ScanLink250[26] , 
        \ScanLink250[25] , \ScanLink250[24] , \ScanLink250[23] , 
        \ScanLink250[22] , \ScanLink250[21] , \ScanLink250[20] , 
        \ScanLink250[19] , \ScanLink250[18] , \ScanLink250[17] , 
        \ScanLink250[16] , \ScanLink250[15] , \ScanLink250[14] , 
        \ScanLink250[13] , \ScanLink250[12] , \ScanLink250[11] , 
        \ScanLink250[10] , \ScanLink250[9] , \ScanLink250[8] , 
        \ScanLink250[7] , \ScanLink250[6] , \ScanLink250[5] , \ScanLink250[4] , 
        \ScanLink250[3] , \ScanLink250[2] , \ScanLink250[1] , \ScanLink250[0] 
        }), .ScanOut({\ScanLink249[31] , \ScanLink249[30] , \ScanLink249[29] , 
        \ScanLink249[28] , \ScanLink249[27] , \ScanLink249[26] , 
        \ScanLink249[25] , \ScanLink249[24] , \ScanLink249[23] , 
        \ScanLink249[22] , \ScanLink249[21] , \ScanLink249[20] , 
        \ScanLink249[19] , \ScanLink249[18] , \ScanLink249[17] , 
        \ScanLink249[16] , \ScanLink249[15] , \ScanLink249[14] , 
        \ScanLink249[13] , \ScanLink249[12] , \ScanLink249[11] , 
        \ScanLink249[10] , \ScanLink249[9] , \ScanLink249[8] , 
        \ScanLink249[7] , \ScanLink249[6] , \ScanLink249[5] , \ScanLink249[4] , 
        \ScanLink249[3] , \ScanLink249[2] , \ScanLink249[1] , \ScanLink249[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_122[31] , 
        \wRegOut_7_122[30] , \wRegOut_7_122[29] , \wRegOut_7_122[28] , 
        \wRegOut_7_122[27] , \wRegOut_7_122[26] , \wRegOut_7_122[25] , 
        \wRegOut_7_122[24] , \wRegOut_7_122[23] , \wRegOut_7_122[22] , 
        \wRegOut_7_122[21] , \wRegOut_7_122[20] , \wRegOut_7_122[19] , 
        \wRegOut_7_122[18] , \wRegOut_7_122[17] , \wRegOut_7_122[16] , 
        \wRegOut_7_122[15] , \wRegOut_7_122[14] , \wRegOut_7_122[13] , 
        \wRegOut_7_122[12] , \wRegOut_7_122[11] , \wRegOut_7_122[10] , 
        \wRegOut_7_122[9] , \wRegOut_7_122[8] , \wRegOut_7_122[7] , 
        \wRegOut_7_122[6] , \wRegOut_7_122[5] , \wRegOut_7_122[4] , 
        \wRegOut_7_122[3] , \wRegOut_7_122[2] , \wRegOut_7_122[1] , 
        \wRegOut_7_122[0] }), .Enable1(\wRegEnTop_7_122[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_122[31] , \wRegInTop_7_122[30] , 
        \wRegInTop_7_122[29] , \wRegInTop_7_122[28] , \wRegInTop_7_122[27] , 
        \wRegInTop_7_122[26] , \wRegInTop_7_122[25] , \wRegInTop_7_122[24] , 
        \wRegInTop_7_122[23] , \wRegInTop_7_122[22] , \wRegInTop_7_122[21] , 
        \wRegInTop_7_122[20] , \wRegInTop_7_122[19] , \wRegInTop_7_122[18] , 
        \wRegInTop_7_122[17] , \wRegInTop_7_122[16] , \wRegInTop_7_122[15] , 
        \wRegInTop_7_122[14] , \wRegInTop_7_122[13] , \wRegInTop_7_122[12] , 
        \wRegInTop_7_122[11] , \wRegInTop_7_122[10] , \wRegInTop_7_122[9] , 
        \wRegInTop_7_122[8] , \wRegInTop_7_122[7] , \wRegInTop_7_122[6] , 
        \wRegInTop_7_122[5] , \wRegInTop_7_122[4] , \wRegInTop_7_122[3] , 
        \wRegInTop_7_122[2] , \wRegInTop_7_122[1] , \wRegInTop_7_122[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_105 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink233[31] , \ScanLink233[30] , \ScanLink233[29] , 
        \ScanLink233[28] , \ScanLink233[27] , \ScanLink233[26] , 
        \ScanLink233[25] , \ScanLink233[24] , \ScanLink233[23] , 
        \ScanLink233[22] , \ScanLink233[21] , \ScanLink233[20] , 
        \ScanLink233[19] , \ScanLink233[18] , \ScanLink233[17] , 
        \ScanLink233[16] , \ScanLink233[15] , \ScanLink233[14] , 
        \ScanLink233[13] , \ScanLink233[12] , \ScanLink233[11] , 
        \ScanLink233[10] , \ScanLink233[9] , \ScanLink233[8] , 
        \ScanLink233[7] , \ScanLink233[6] , \ScanLink233[5] , \ScanLink233[4] , 
        \ScanLink233[3] , \ScanLink233[2] , \ScanLink233[1] , \ScanLink233[0] 
        }), .ScanOut({\ScanLink232[31] , \ScanLink232[30] , \ScanLink232[29] , 
        \ScanLink232[28] , \ScanLink232[27] , \ScanLink232[26] , 
        \ScanLink232[25] , \ScanLink232[24] , \ScanLink232[23] , 
        \ScanLink232[22] , \ScanLink232[21] , \ScanLink232[20] , 
        \ScanLink232[19] , \ScanLink232[18] , \ScanLink232[17] , 
        \ScanLink232[16] , \ScanLink232[15] , \ScanLink232[14] , 
        \ScanLink232[13] , \ScanLink232[12] , \ScanLink232[11] , 
        \ScanLink232[10] , \ScanLink232[9] , \ScanLink232[8] , 
        \ScanLink232[7] , \ScanLink232[6] , \ScanLink232[5] , \ScanLink232[4] , 
        \ScanLink232[3] , \ScanLink232[2] , \ScanLink232[1] , \ScanLink232[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_105[31] , 
        \wRegOut_7_105[30] , \wRegOut_7_105[29] , \wRegOut_7_105[28] , 
        \wRegOut_7_105[27] , \wRegOut_7_105[26] , \wRegOut_7_105[25] , 
        \wRegOut_7_105[24] , \wRegOut_7_105[23] , \wRegOut_7_105[22] , 
        \wRegOut_7_105[21] , \wRegOut_7_105[20] , \wRegOut_7_105[19] , 
        \wRegOut_7_105[18] , \wRegOut_7_105[17] , \wRegOut_7_105[16] , 
        \wRegOut_7_105[15] , \wRegOut_7_105[14] , \wRegOut_7_105[13] , 
        \wRegOut_7_105[12] , \wRegOut_7_105[11] , \wRegOut_7_105[10] , 
        \wRegOut_7_105[9] , \wRegOut_7_105[8] , \wRegOut_7_105[7] , 
        \wRegOut_7_105[6] , \wRegOut_7_105[5] , \wRegOut_7_105[4] , 
        \wRegOut_7_105[3] , \wRegOut_7_105[2] , \wRegOut_7_105[1] , 
        \wRegOut_7_105[0] }), .Enable1(\wRegEnTop_7_105[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_105[31] , \wRegInTop_7_105[30] , 
        \wRegInTop_7_105[29] , \wRegInTop_7_105[28] , \wRegInTop_7_105[27] , 
        \wRegInTop_7_105[26] , \wRegInTop_7_105[25] , \wRegInTop_7_105[24] , 
        \wRegInTop_7_105[23] , \wRegInTop_7_105[22] , \wRegInTop_7_105[21] , 
        \wRegInTop_7_105[20] , \wRegInTop_7_105[19] , \wRegInTop_7_105[18] , 
        \wRegInTop_7_105[17] , \wRegInTop_7_105[16] , \wRegInTop_7_105[15] , 
        \wRegInTop_7_105[14] , \wRegInTop_7_105[13] , \wRegInTop_7_105[12] , 
        \wRegInTop_7_105[11] , \wRegInTop_7_105[10] , \wRegInTop_7_105[9] , 
        \wRegInTop_7_105[8] , \wRegInTop_7_105[7] , \wRegInTop_7_105[6] , 
        \wRegInTop_7_105[5] , \wRegInTop_7_105[4] , \wRegInTop_7_105[3] , 
        \wRegInTop_7_105[2] , \wRegInTop_7_105[1] , \wRegInTop_7_105[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_CtrlReg_WIDTH32 BHCR_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_6[0] ), 
        .Out(\wCtrlOut_5[0] ), .Enable(\wEnable_5[0] ) );
    BHeap_Node_WIDTH32 BHN_2_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_2[0] ), .P_WR(\wRegEnBot_2_1[0] ), .P_In({\wRegOut_2_1[31] , 
        \wRegOut_2_1[30] , \wRegOut_2_1[29] , \wRegOut_2_1[28] , 
        \wRegOut_2_1[27] , \wRegOut_2_1[26] , \wRegOut_2_1[25] , 
        \wRegOut_2_1[24] , \wRegOut_2_1[23] , \wRegOut_2_1[22] , 
        \wRegOut_2_1[21] , \wRegOut_2_1[20] , \wRegOut_2_1[19] , 
        \wRegOut_2_1[18] , \wRegOut_2_1[17] , \wRegOut_2_1[16] , 
        \wRegOut_2_1[15] , \wRegOut_2_1[14] , \wRegOut_2_1[13] , 
        \wRegOut_2_1[12] , \wRegOut_2_1[11] , \wRegOut_2_1[10] , 
        \wRegOut_2_1[9] , \wRegOut_2_1[8] , \wRegOut_2_1[7] , \wRegOut_2_1[6] , 
        \wRegOut_2_1[5] , \wRegOut_2_1[4] , \wRegOut_2_1[3] , \wRegOut_2_1[2] , 
        \wRegOut_2_1[1] , \wRegOut_2_1[0] }), .P_Out({\wRegInBot_2_1[31] , 
        \wRegInBot_2_1[30] , \wRegInBot_2_1[29] , \wRegInBot_2_1[28] , 
        \wRegInBot_2_1[27] , \wRegInBot_2_1[26] , \wRegInBot_2_1[25] , 
        \wRegInBot_2_1[24] , \wRegInBot_2_1[23] , \wRegInBot_2_1[22] , 
        \wRegInBot_2_1[21] , \wRegInBot_2_1[20] , \wRegInBot_2_1[19] , 
        \wRegInBot_2_1[18] , \wRegInBot_2_1[17] , \wRegInBot_2_1[16] , 
        \wRegInBot_2_1[15] , \wRegInBot_2_1[14] , \wRegInBot_2_1[13] , 
        \wRegInBot_2_1[12] , \wRegInBot_2_1[11] , \wRegInBot_2_1[10] , 
        \wRegInBot_2_1[9] , \wRegInBot_2_1[8] , \wRegInBot_2_1[7] , 
        \wRegInBot_2_1[6] , \wRegInBot_2_1[5] , \wRegInBot_2_1[4] , 
        \wRegInBot_2_1[3] , \wRegInBot_2_1[2] , \wRegInBot_2_1[1] , 
        \wRegInBot_2_1[0] }), .L_WR(\wRegEnTop_3_2[0] ), .L_In({
        \wRegOut_3_2[31] , \wRegOut_3_2[30] , \wRegOut_3_2[29] , 
        \wRegOut_3_2[28] , \wRegOut_3_2[27] , \wRegOut_3_2[26] , 
        \wRegOut_3_2[25] , \wRegOut_3_2[24] , \wRegOut_3_2[23] , 
        \wRegOut_3_2[22] , \wRegOut_3_2[21] , \wRegOut_3_2[20] , 
        \wRegOut_3_2[19] , \wRegOut_3_2[18] , \wRegOut_3_2[17] , 
        \wRegOut_3_2[16] , \wRegOut_3_2[15] , \wRegOut_3_2[14] , 
        \wRegOut_3_2[13] , \wRegOut_3_2[12] , \wRegOut_3_2[11] , 
        \wRegOut_3_2[10] , \wRegOut_3_2[9] , \wRegOut_3_2[8] , 
        \wRegOut_3_2[7] , \wRegOut_3_2[6] , \wRegOut_3_2[5] , \wRegOut_3_2[4] , 
        \wRegOut_3_2[3] , \wRegOut_3_2[2] , \wRegOut_3_2[1] , \wRegOut_3_2[0] 
        }), .L_Out({\wRegInTop_3_2[31] , \wRegInTop_3_2[30] , 
        \wRegInTop_3_2[29] , \wRegInTop_3_2[28] , \wRegInTop_3_2[27] , 
        \wRegInTop_3_2[26] , \wRegInTop_3_2[25] , \wRegInTop_3_2[24] , 
        \wRegInTop_3_2[23] , \wRegInTop_3_2[22] , \wRegInTop_3_2[21] , 
        \wRegInTop_3_2[20] , \wRegInTop_3_2[19] , \wRegInTop_3_2[18] , 
        \wRegInTop_3_2[17] , \wRegInTop_3_2[16] , \wRegInTop_3_2[15] , 
        \wRegInTop_3_2[14] , \wRegInTop_3_2[13] , \wRegInTop_3_2[12] , 
        \wRegInTop_3_2[11] , \wRegInTop_3_2[10] , \wRegInTop_3_2[9] , 
        \wRegInTop_3_2[8] , \wRegInTop_3_2[7] , \wRegInTop_3_2[6] , 
        \wRegInTop_3_2[5] , \wRegInTop_3_2[4] , \wRegInTop_3_2[3] , 
        \wRegInTop_3_2[2] , \wRegInTop_3_2[1] , \wRegInTop_3_2[0] }), .R_WR(
        \wRegEnTop_3_3[0] ), .R_In({\wRegOut_3_3[31] , \wRegOut_3_3[30] , 
        \wRegOut_3_3[29] , \wRegOut_3_3[28] , \wRegOut_3_3[27] , 
        \wRegOut_3_3[26] , \wRegOut_3_3[25] , \wRegOut_3_3[24] , 
        \wRegOut_3_3[23] , \wRegOut_3_3[22] , \wRegOut_3_3[21] , 
        \wRegOut_3_3[20] , \wRegOut_3_3[19] , \wRegOut_3_3[18] , 
        \wRegOut_3_3[17] , \wRegOut_3_3[16] , \wRegOut_3_3[15] , 
        \wRegOut_3_3[14] , \wRegOut_3_3[13] , \wRegOut_3_3[12] , 
        \wRegOut_3_3[11] , \wRegOut_3_3[10] , \wRegOut_3_3[9] , 
        \wRegOut_3_3[8] , \wRegOut_3_3[7] , \wRegOut_3_3[6] , \wRegOut_3_3[5] , 
        \wRegOut_3_3[4] , \wRegOut_3_3[3] , \wRegOut_3_3[2] , \wRegOut_3_3[1] , 
        \wRegOut_3_3[0] }), .R_Out({\wRegInTop_3_3[31] , \wRegInTop_3_3[30] , 
        \wRegInTop_3_3[29] , \wRegInTop_3_3[28] , \wRegInTop_3_3[27] , 
        \wRegInTop_3_3[26] , \wRegInTop_3_3[25] , \wRegInTop_3_3[24] , 
        \wRegInTop_3_3[23] , \wRegInTop_3_3[22] , \wRegInTop_3_3[21] , 
        \wRegInTop_3_3[20] , \wRegInTop_3_3[19] , \wRegInTop_3_3[18] , 
        \wRegInTop_3_3[17] , \wRegInTop_3_3[16] , \wRegInTop_3_3[15] , 
        \wRegInTop_3_3[14] , \wRegInTop_3_3[13] , \wRegInTop_3_3[12] , 
        \wRegInTop_3_3[11] , \wRegInTop_3_3[10] , \wRegInTop_3_3[9] , 
        \wRegInTop_3_3[8] , \wRegInTop_3_3[7] , \wRegInTop_3_3[6] , 
        \wRegInTop_3_3[5] , \wRegInTop_3_3[4] , \wRegInTop_3_3[3] , 
        \wRegInTop_3_3[2] , \wRegInTop_3_3[1] , \wRegInTop_3_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink12[31] , \ScanLink12[30] , \ScanLink12[29] , 
        \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , \ScanLink12[25] , 
        \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , \ScanLink12[21] , 
        \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , \ScanLink12[17] , 
        \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , \ScanLink12[13] , 
        \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , \ScanLink12[9] , 
        \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , \ScanLink12[5] , 
        \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , \ScanLink12[1] , 
        \ScanLink12[0] }), .ScanOut({\ScanLink11[31] , \ScanLink11[30] , 
        \ScanLink11[29] , \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , 
        \ScanLink11[25] , \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , 
        \ScanLink11[21] , \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , 
        \ScanLink11[17] , \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , 
        \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , 
        \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , 
        \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , 
        \ScanLink11[1] , \ScanLink11[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_4[31] , \wRegOut_3_4[30] , \wRegOut_3_4[29] , 
        \wRegOut_3_4[28] , \wRegOut_3_4[27] , \wRegOut_3_4[26] , 
        \wRegOut_3_4[25] , \wRegOut_3_4[24] , \wRegOut_3_4[23] , 
        \wRegOut_3_4[22] , \wRegOut_3_4[21] , \wRegOut_3_4[20] , 
        \wRegOut_3_4[19] , \wRegOut_3_4[18] , \wRegOut_3_4[17] , 
        \wRegOut_3_4[16] , \wRegOut_3_4[15] , \wRegOut_3_4[14] , 
        \wRegOut_3_4[13] , \wRegOut_3_4[12] , \wRegOut_3_4[11] , 
        \wRegOut_3_4[10] , \wRegOut_3_4[9] , \wRegOut_3_4[8] , 
        \wRegOut_3_4[7] , \wRegOut_3_4[6] , \wRegOut_3_4[5] , \wRegOut_3_4[4] , 
        \wRegOut_3_4[3] , \wRegOut_3_4[2] , \wRegOut_3_4[1] , \wRegOut_3_4[0] 
        }), .Enable1(\wRegEnTop_3_4[0] ), .Enable2(\wRegEnBot_3_4[0] ), .In1({
        \wRegInTop_3_4[31] , \wRegInTop_3_4[30] , \wRegInTop_3_4[29] , 
        \wRegInTop_3_4[28] , \wRegInTop_3_4[27] , \wRegInTop_3_4[26] , 
        \wRegInTop_3_4[25] , \wRegInTop_3_4[24] , \wRegInTop_3_4[23] , 
        \wRegInTop_3_4[22] , \wRegInTop_3_4[21] , \wRegInTop_3_4[20] , 
        \wRegInTop_3_4[19] , \wRegInTop_3_4[18] , \wRegInTop_3_4[17] , 
        \wRegInTop_3_4[16] , \wRegInTop_3_4[15] , \wRegInTop_3_4[14] , 
        \wRegInTop_3_4[13] , \wRegInTop_3_4[12] , \wRegInTop_3_4[11] , 
        \wRegInTop_3_4[10] , \wRegInTop_3_4[9] , \wRegInTop_3_4[8] , 
        \wRegInTop_3_4[7] , \wRegInTop_3_4[6] , \wRegInTop_3_4[5] , 
        \wRegInTop_3_4[4] , \wRegInTop_3_4[3] , \wRegInTop_3_4[2] , 
        \wRegInTop_3_4[1] , \wRegInTop_3_4[0] }), .In2({\wRegInBot_3_4[31] , 
        \wRegInBot_3_4[30] , \wRegInBot_3_4[29] , \wRegInBot_3_4[28] , 
        \wRegInBot_3_4[27] , \wRegInBot_3_4[26] , \wRegInBot_3_4[25] , 
        \wRegInBot_3_4[24] , \wRegInBot_3_4[23] , \wRegInBot_3_4[22] , 
        \wRegInBot_3_4[21] , \wRegInBot_3_4[20] , \wRegInBot_3_4[19] , 
        \wRegInBot_3_4[18] , \wRegInBot_3_4[17] , \wRegInBot_3_4[16] , 
        \wRegInBot_3_4[15] , \wRegInBot_3_4[14] , \wRegInBot_3_4[13] , 
        \wRegInBot_3_4[12] , \wRegInBot_3_4[11] , \wRegInBot_3_4[10] , 
        \wRegInBot_3_4[9] , \wRegInBot_3_4[8] , \wRegInBot_3_4[7] , 
        \wRegInBot_3_4[6] , \wRegInBot_3_4[5] , \wRegInBot_3_4[4] , 
        \wRegInBot_3_4[3] , \wRegInBot_3_4[2] , \wRegInBot_3_4[1] , 
        \wRegInBot_3_4[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink25[31] , \ScanLink25[30] , \ScanLink25[29] , 
        \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , \ScanLink25[25] , 
        \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , \ScanLink25[21] , 
        \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , \ScanLink25[17] , 
        \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , \ScanLink25[13] , 
        \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , \ScanLink25[9] , 
        \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , \ScanLink25[5] , 
        \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , \ScanLink25[1] , 
        \ScanLink25[0] }), .ScanOut({\ScanLink24[31] , \ScanLink24[30] , 
        \ScanLink24[29] , \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , 
        \ScanLink24[25] , \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , 
        \ScanLink24[21] , \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , 
        \ScanLink24[17] , \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , 
        \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , 
        \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , 
        \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , 
        \ScanLink24[1] , \ScanLink24[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_9[31] , \wRegOut_4_9[30] , \wRegOut_4_9[29] , 
        \wRegOut_4_9[28] , \wRegOut_4_9[27] , \wRegOut_4_9[26] , 
        \wRegOut_4_9[25] , \wRegOut_4_9[24] , \wRegOut_4_9[23] , 
        \wRegOut_4_9[22] , \wRegOut_4_9[21] , \wRegOut_4_9[20] , 
        \wRegOut_4_9[19] , \wRegOut_4_9[18] , \wRegOut_4_9[17] , 
        \wRegOut_4_9[16] , \wRegOut_4_9[15] , \wRegOut_4_9[14] , 
        \wRegOut_4_9[13] , \wRegOut_4_9[12] , \wRegOut_4_9[11] , 
        \wRegOut_4_9[10] , \wRegOut_4_9[9] , \wRegOut_4_9[8] , 
        \wRegOut_4_9[7] , \wRegOut_4_9[6] , \wRegOut_4_9[5] , \wRegOut_4_9[4] , 
        \wRegOut_4_9[3] , \wRegOut_4_9[2] , \wRegOut_4_9[1] , \wRegOut_4_9[0] 
        }), .Enable1(\wRegEnTop_4_9[0] ), .Enable2(\wRegEnBot_4_9[0] ), .In1({
        \wRegInTop_4_9[31] , \wRegInTop_4_9[30] , \wRegInTop_4_9[29] , 
        \wRegInTop_4_9[28] , \wRegInTop_4_9[27] , \wRegInTop_4_9[26] , 
        \wRegInTop_4_9[25] , \wRegInTop_4_9[24] , \wRegInTop_4_9[23] , 
        \wRegInTop_4_9[22] , \wRegInTop_4_9[21] , \wRegInTop_4_9[20] , 
        \wRegInTop_4_9[19] , \wRegInTop_4_9[18] , \wRegInTop_4_9[17] , 
        \wRegInTop_4_9[16] , \wRegInTop_4_9[15] , \wRegInTop_4_9[14] , 
        \wRegInTop_4_9[13] , \wRegInTop_4_9[12] , \wRegInTop_4_9[11] , 
        \wRegInTop_4_9[10] , \wRegInTop_4_9[9] , \wRegInTop_4_9[8] , 
        \wRegInTop_4_9[7] , \wRegInTop_4_9[6] , \wRegInTop_4_9[5] , 
        \wRegInTop_4_9[4] , \wRegInTop_4_9[3] , \wRegInTop_4_9[2] , 
        \wRegInTop_4_9[1] , \wRegInTop_4_9[0] }), .In2({\wRegInBot_4_9[31] , 
        \wRegInBot_4_9[30] , \wRegInBot_4_9[29] , \wRegInBot_4_9[28] , 
        \wRegInBot_4_9[27] , \wRegInBot_4_9[26] , \wRegInBot_4_9[25] , 
        \wRegInBot_4_9[24] , \wRegInBot_4_9[23] , \wRegInBot_4_9[22] , 
        \wRegInBot_4_9[21] , \wRegInBot_4_9[20] , \wRegInBot_4_9[19] , 
        \wRegInBot_4_9[18] , \wRegInBot_4_9[17] , \wRegInBot_4_9[16] , 
        \wRegInBot_4_9[15] , \wRegInBot_4_9[14] , \wRegInBot_4_9[13] , 
        \wRegInBot_4_9[12] , \wRegInBot_4_9[11] , \wRegInBot_4_9[10] , 
        \wRegInBot_4_9[9] , \wRegInBot_4_9[8] , \wRegInBot_4_9[7] , 
        \wRegInBot_4_9[6] , \wRegInBot_4_9[5] , \wRegInBot_4_9[4] , 
        \wRegInBot_4_9[3] , \wRegInBot_4_9[2] , \wRegInBot_4_9[1] , 
        \wRegInBot_4_9[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink69[31] , \ScanLink69[30] , \ScanLink69[29] , 
        \ScanLink69[28] , \ScanLink69[27] , \ScanLink69[26] , \ScanLink69[25] , 
        \ScanLink69[24] , \ScanLink69[23] , \ScanLink69[22] , \ScanLink69[21] , 
        \ScanLink69[20] , \ScanLink69[19] , \ScanLink69[18] , \ScanLink69[17] , 
        \ScanLink69[16] , \ScanLink69[15] , \ScanLink69[14] , \ScanLink69[13] , 
        \ScanLink69[12] , \ScanLink69[11] , \ScanLink69[10] , \ScanLink69[9] , 
        \ScanLink69[8] , \ScanLink69[7] , \ScanLink69[6] , \ScanLink69[5] , 
        \ScanLink69[4] , \ScanLink69[3] , \ScanLink69[2] , \ScanLink69[1] , 
        \ScanLink69[0] }), .ScanOut({\ScanLink68[31] , \ScanLink68[30] , 
        \ScanLink68[29] , \ScanLink68[28] , \ScanLink68[27] , \ScanLink68[26] , 
        \ScanLink68[25] , \ScanLink68[24] , \ScanLink68[23] , \ScanLink68[22] , 
        \ScanLink68[21] , \ScanLink68[20] , \ScanLink68[19] , \ScanLink68[18] , 
        \ScanLink68[17] , \ScanLink68[16] , \ScanLink68[15] , \ScanLink68[14] , 
        \ScanLink68[13] , \ScanLink68[12] , \ScanLink68[11] , \ScanLink68[10] , 
        \ScanLink68[9] , \ScanLink68[8] , \ScanLink68[7] , \ScanLink68[6] , 
        \ScanLink68[5] , \ScanLink68[4] , \ScanLink68[3] , \ScanLink68[2] , 
        \ScanLink68[1] , \ScanLink68[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_5[31] , \wRegOut_6_5[30] , \wRegOut_6_5[29] , 
        \wRegOut_6_5[28] , \wRegOut_6_5[27] , \wRegOut_6_5[26] , 
        \wRegOut_6_5[25] , \wRegOut_6_5[24] , \wRegOut_6_5[23] , 
        \wRegOut_6_5[22] , \wRegOut_6_5[21] , \wRegOut_6_5[20] , 
        \wRegOut_6_5[19] , \wRegOut_6_5[18] , \wRegOut_6_5[17] , 
        \wRegOut_6_5[16] , \wRegOut_6_5[15] , \wRegOut_6_5[14] , 
        \wRegOut_6_5[13] , \wRegOut_6_5[12] , \wRegOut_6_5[11] , 
        \wRegOut_6_5[10] , \wRegOut_6_5[9] , \wRegOut_6_5[8] , 
        \wRegOut_6_5[7] , \wRegOut_6_5[6] , \wRegOut_6_5[5] , \wRegOut_6_5[4] , 
        \wRegOut_6_5[3] , \wRegOut_6_5[2] , \wRegOut_6_5[1] , \wRegOut_6_5[0] 
        }), .Enable1(\wRegEnTop_6_5[0] ), .Enable2(\wRegEnBot_6_5[0] ), .In1({
        \wRegInTop_6_5[31] , \wRegInTop_6_5[30] , \wRegInTop_6_5[29] , 
        \wRegInTop_6_5[28] , \wRegInTop_6_5[27] , \wRegInTop_6_5[26] , 
        \wRegInTop_6_5[25] , \wRegInTop_6_5[24] , \wRegInTop_6_5[23] , 
        \wRegInTop_6_5[22] , \wRegInTop_6_5[21] , \wRegInTop_6_5[20] , 
        \wRegInTop_6_5[19] , \wRegInTop_6_5[18] , \wRegInTop_6_5[17] , 
        \wRegInTop_6_5[16] , \wRegInTop_6_5[15] , \wRegInTop_6_5[14] , 
        \wRegInTop_6_5[13] , \wRegInTop_6_5[12] , \wRegInTop_6_5[11] , 
        \wRegInTop_6_5[10] , \wRegInTop_6_5[9] , \wRegInTop_6_5[8] , 
        \wRegInTop_6_5[7] , \wRegInTop_6_5[6] , \wRegInTop_6_5[5] , 
        \wRegInTop_6_5[4] , \wRegInTop_6_5[3] , \wRegInTop_6_5[2] , 
        \wRegInTop_6_5[1] , \wRegInTop_6_5[0] }), .In2({\wRegInBot_6_5[31] , 
        \wRegInBot_6_5[30] , \wRegInBot_6_5[29] , \wRegInBot_6_5[28] , 
        \wRegInBot_6_5[27] , \wRegInBot_6_5[26] , \wRegInBot_6_5[25] , 
        \wRegInBot_6_5[24] , \wRegInBot_6_5[23] , \wRegInBot_6_5[22] , 
        \wRegInBot_6_5[21] , \wRegInBot_6_5[20] , \wRegInBot_6_5[19] , 
        \wRegInBot_6_5[18] , \wRegInBot_6_5[17] , \wRegInBot_6_5[16] , 
        \wRegInBot_6_5[15] , \wRegInBot_6_5[14] , \wRegInBot_6_5[13] , 
        \wRegInBot_6_5[12] , \wRegInBot_6_5[11] , \wRegInBot_6_5[10] , 
        \wRegInBot_6_5[9] , \wRegInBot_6_5[8] , \wRegInBot_6_5[7] , 
        \wRegInBot_6_5[6] , \wRegInBot_6_5[5] , \wRegInBot_6_5[4] , 
        \wRegInBot_6_5[3] , \wRegInBot_6_5[2] , \wRegInBot_6_5[1] , 
        \wRegInBot_6_5[0] }) );
    BHeap_Node_WIDTH32 BHN_5_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_13[0] ), .P_In({\wRegOut_5_13[31] , 
        \wRegOut_5_13[30] , \wRegOut_5_13[29] , \wRegOut_5_13[28] , 
        \wRegOut_5_13[27] , \wRegOut_5_13[26] , \wRegOut_5_13[25] , 
        \wRegOut_5_13[24] , \wRegOut_5_13[23] , \wRegOut_5_13[22] , 
        \wRegOut_5_13[21] , \wRegOut_5_13[20] , \wRegOut_5_13[19] , 
        \wRegOut_5_13[18] , \wRegOut_5_13[17] , \wRegOut_5_13[16] , 
        \wRegOut_5_13[15] , \wRegOut_5_13[14] , \wRegOut_5_13[13] , 
        \wRegOut_5_13[12] , \wRegOut_5_13[11] , \wRegOut_5_13[10] , 
        \wRegOut_5_13[9] , \wRegOut_5_13[8] , \wRegOut_5_13[7] , 
        \wRegOut_5_13[6] , \wRegOut_5_13[5] , \wRegOut_5_13[4] , 
        \wRegOut_5_13[3] , \wRegOut_5_13[2] , \wRegOut_5_13[1] , 
        \wRegOut_5_13[0] }), .P_Out({\wRegInBot_5_13[31] , 
        \wRegInBot_5_13[30] , \wRegInBot_5_13[29] , \wRegInBot_5_13[28] , 
        \wRegInBot_5_13[27] , \wRegInBot_5_13[26] , \wRegInBot_5_13[25] , 
        \wRegInBot_5_13[24] , \wRegInBot_5_13[23] , \wRegInBot_5_13[22] , 
        \wRegInBot_5_13[21] , \wRegInBot_5_13[20] , \wRegInBot_5_13[19] , 
        \wRegInBot_5_13[18] , \wRegInBot_5_13[17] , \wRegInBot_5_13[16] , 
        \wRegInBot_5_13[15] , \wRegInBot_5_13[14] , \wRegInBot_5_13[13] , 
        \wRegInBot_5_13[12] , \wRegInBot_5_13[11] , \wRegInBot_5_13[10] , 
        \wRegInBot_5_13[9] , \wRegInBot_5_13[8] , \wRegInBot_5_13[7] , 
        \wRegInBot_5_13[6] , \wRegInBot_5_13[5] , \wRegInBot_5_13[4] , 
        \wRegInBot_5_13[3] , \wRegInBot_5_13[2] , \wRegInBot_5_13[1] , 
        \wRegInBot_5_13[0] }), .L_WR(\wRegEnTop_6_26[0] ), .L_In({
        \wRegOut_6_26[31] , \wRegOut_6_26[30] , \wRegOut_6_26[29] , 
        \wRegOut_6_26[28] , \wRegOut_6_26[27] , \wRegOut_6_26[26] , 
        \wRegOut_6_26[25] , \wRegOut_6_26[24] , \wRegOut_6_26[23] , 
        \wRegOut_6_26[22] , \wRegOut_6_26[21] , \wRegOut_6_26[20] , 
        \wRegOut_6_26[19] , \wRegOut_6_26[18] , \wRegOut_6_26[17] , 
        \wRegOut_6_26[16] , \wRegOut_6_26[15] , \wRegOut_6_26[14] , 
        \wRegOut_6_26[13] , \wRegOut_6_26[12] , \wRegOut_6_26[11] , 
        \wRegOut_6_26[10] , \wRegOut_6_26[9] , \wRegOut_6_26[8] , 
        \wRegOut_6_26[7] , \wRegOut_6_26[6] , \wRegOut_6_26[5] , 
        \wRegOut_6_26[4] , \wRegOut_6_26[3] , \wRegOut_6_26[2] , 
        \wRegOut_6_26[1] , \wRegOut_6_26[0] }), .L_Out({\wRegInTop_6_26[31] , 
        \wRegInTop_6_26[30] , \wRegInTop_6_26[29] , \wRegInTop_6_26[28] , 
        \wRegInTop_6_26[27] , \wRegInTop_6_26[26] , \wRegInTop_6_26[25] , 
        \wRegInTop_6_26[24] , \wRegInTop_6_26[23] , \wRegInTop_6_26[22] , 
        \wRegInTop_6_26[21] , \wRegInTop_6_26[20] , \wRegInTop_6_26[19] , 
        \wRegInTop_6_26[18] , \wRegInTop_6_26[17] , \wRegInTop_6_26[16] , 
        \wRegInTop_6_26[15] , \wRegInTop_6_26[14] , \wRegInTop_6_26[13] , 
        \wRegInTop_6_26[12] , \wRegInTop_6_26[11] , \wRegInTop_6_26[10] , 
        \wRegInTop_6_26[9] , \wRegInTop_6_26[8] , \wRegInTop_6_26[7] , 
        \wRegInTop_6_26[6] , \wRegInTop_6_26[5] , \wRegInTop_6_26[4] , 
        \wRegInTop_6_26[3] , \wRegInTop_6_26[2] , \wRegInTop_6_26[1] , 
        \wRegInTop_6_26[0] }), .R_WR(\wRegEnTop_6_27[0] ), .R_In({
        \wRegOut_6_27[31] , \wRegOut_6_27[30] , \wRegOut_6_27[29] , 
        \wRegOut_6_27[28] , \wRegOut_6_27[27] , \wRegOut_6_27[26] , 
        \wRegOut_6_27[25] , \wRegOut_6_27[24] , \wRegOut_6_27[23] , 
        \wRegOut_6_27[22] , \wRegOut_6_27[21] , \wRegOut_6_27[20] , 
        \wRegOut_6_27[19] , \wRegOut_6_27[18] , \wRegOut_6_27[17] , 
        \wRegOut_6_27[16] , \wRegOut_6_27[15] , \wRegOut_6_27[14] , 
        \wRegOut_6_27[13] , \wRegOut_6_27[12] , \wRegOut_6_27[11] , 
        \wRegOut_6_27[10] , \wRegOut_6_27[9] , \wRegOut_6_27[8] , 
        \wRegOut_6_27[7] , \wRegOut_6_27[6] , \wRegOut_6_27[5] , 
        \wRegOut_6_27[4] , \wRegOut_6_27[3] , \wRegOut_6_27[2] , 
        \wRegOut_6_27[1] , \wRegOut_6_27[0] }), .R_Out({\wRegInTop_6_27[31] , 
        \wRegInTop_6_27[30] , \wRegInTop_6_27[29] , \wRegInTop_6_27[28] , 
        \wRegInTop_6_27[27] , \wRegInTop_6_27[26] , \wRegInTop_6_27[25] , 
        \wRegInTop_6_27[24] , \wRegInTop_6_27[23] , \wRegInTop_6_27[22] , 
        \wRegInTop_6_27[21] , \wRegInTop_6_27[20] , \wRegInTop_6_27[19] , 
        \wRegInTop_6_27[18] , \wRegInTop_6_27[17] , \wRegInTop_6_27[16] , 
        \wRegInTop_6_27[15] , \wRegInTop_6_27[14] , \wRegInTop_6_27[13] , 
        \wRegInTop_6_27[12] , \wRegInTop_6_27[11] , \wRegInTop_6_27[10] , 
        \wRegInTop_6_27[9] , \wRegInTop_6_27[8] , \wRegInTop_6_27[7] , 
        \wRegInTop_6_27[6] , \wRegInTop_6_27[5] , \wRegInTop_6_27[4] , 
        \wRegInTop_6_27[3] , \wRegInTop_6_27[2] , \wRegInTop_6_27[1] , 
        \wRegInTop_6_27[0] }) );
    BHeap_Node_WIDTH32 BHN_6_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_23[0] ), .P_In({\wRegOut_6_23[31] , 
        \wRegOut_6_23[30] , \wRegOut_6_23[29] , \wRegOut_6_23[28] , 
        \wRegOut_6_23[27] , \wRegOut_6_23[26] , \wRegOut_6_23[25] , 
        \wRegOut_6_23[24] , \wRegOut_6_23[23] , \wRegOut_6_23[22] , 
        \wRegOut_6_23[21] , \wRegOut_6_23[20] , \wRegOut_6_23[19] , 
        \wRegOut_6_23[18] , \wRegOut_6_23[17] , \wRegOut_6_23[16] , 
        \wRegOut_6_23[15] , \wRegOut_6_23[14] , \wRegOut_6_23[13] , 
        \wRegOut_6_23[12] , \wRegOut_6_23[11] , \wRegOut_6_23[10] , 
        \wRegOut_6_23[9] , \wRegOut_6_23[8] , \wRegOut_6_23[7] , 
        \wRegOut_6_23[6] , \wRegOut_6_23[5] , \wRegOut_6_23[4] , 
        \wRegOut_6_23[3] , \wRegOut_6_23[2] , \wRegOut_6_23[1] , 
        \wRegOut_6_23[0] }), .P_Out({\wRegInBot_6_23[31] , 
        \wRegInBot_6_23[30] , \wRegInBot_6_23[29] , \wRegInBot_6_23[28] , 
        \wRegInBot_6_23[27] , \wRegInBot_6_23[26] , \wRegInBot_6_23[25] , 
        \wRegInBot_6_23[24] , \wRegInBot_6_23[23] , \wRegInBot_6_23[22] , 
        \wRegInBot_6_23[21] , \wRegInBot_6_23[20] , \wRegInBot_6_23[19] , 
        \wRegInBot_6_23[18] , \wRegInBot_6_23[17] , \wRegInBot_6_23[16] , 
        \wRegInBot_6_23[15] , \wRegInBot_6_23[14] , \wRegInBot_6_23[13] , 
        \wRegInBot_6_23[12] , \wRegInBot_6_23[11] , \wRegInBot_6_23[10] , 
        \wRegInBot_6_23[9] , \wRegInBot_6_23[8] , \wRegInBot_6_23[7] , 
        \wRegInBot_6_23[6] , \wRegInBot_6_23[5] , \wRegInBot_6_23[4] , 
        \wRegInBot_6_23[3] , \wRegInBot_6_23[2] , \wRegInBot_6_23[1] , 
        \wRegInBot_6_23[0] }), .L_WR(\wRegEnTop_7_46[0] ), .L_In({
        \wRegOut_7_46[31] , \wRegOut_7_46[30] , \wRegOut_7_46[29] , 
        \wRegOut_7_46[28] , \wRegOut_7_46[27] , \wRegOut_7_46[26] , 
        \wRegOut_7_46[25] , \wRegOut_7_46[24] , \wRegOut_7_46[23] , 
        \wRegOut_7_46[22] , \wRegOut_7_46[21] , \wRegOut_7_46[20] , 
        \wRegOut_7_46[19] , \wRegOut_7_46[18] , \wRegOut_7_46[17] , 
        \wRegOut_7_46[16] , \wRegOut_7_46[15] , \wRegOut_7_46[14] , 
        \wRegOut_7_46[13] , \wRegOut_7_46[12] , \wRegOut_7_46[11] , 
        \wRegOut_7_46[10] , \wRegOut_7_46[9] , \wRegOut_7_46[8] , 
        \wRegOut_7_46[7] , \wRegOut_7_46[6] , \wRegOut_7_46[5] , 
        \wRegOut_7_46[4] , \wRegOut_7_46[3] , \wRegOut_7_46[2] , 
        \wRegOut_7_46[1] , \wRegOut_7_46[0] }), .L_Out({\wRegInTop_7_46[31] , 
        \wRegInTop_7_46[30] , \wRegInTop_7_46[29] , \wRegInTop_7_46[28] , 
        \wRegInTop_7_46[27] , \wRegInTop_7_46[26] , \wRegInTop_7_46[25] , 
        \wRegInTop_7_46[24] , \wRegInTop_7_46[23] , \wRegInTop_7_46[22] , 
        \wRegInTop_7_46[21] , \wRegInTop_7_46[20] , \wRegInTop_7_46[19] , 
        \wRegInTop_7_46[18] , \wRegInTop_7_46[17] , \wRegInTop_7_46[16] , 
        \wRegInTop_7_46[15] , \wRegInTop_7_46[14] , \wRegInTop_7_46[13] , 
        \wRegInTop_7_46[12] , \wRegInTop_7_46[11] , \wRegInTop_7_46[10] , 
        \wRegInTop_7_46[9] , \wRegInTop_7_46[8] , \wRegInTop_7_46[7] , 
        \wRegInTop_7_46[6] , \wRegInTop_7_46[5] , \wRegInTop_7_46[4] , 
        \wRegInTop_7_46[3] , \wRegInTop_7_46[2] , \wRegInTop_7_46[1] , 
        \wRegInTop_7_46[0] }), .R_WR(\wRegEnTop_7_47[0] ), .R_In({
        \wRegOut_7_47[31] , \wRegOut_7_47[30] , \wRegOut_7_47[29] , 
        \wRegOut_7_47[28] , \wRegOut_7_47[27] , \wRegOut_7_47[26] , 
        \wRegOut_7_47[25] , \wRegOut_7_47[24] , \wRegOut_7_47[23] , 
        \wRegOut_7_47[22] , \wRegOut_7_47[21] , \wRegOut_7_47[20] , 
        \wRegOut_7_47[19] , \wRegOut_7_47[18] , \wRegOut_7_47[17] , 
        \wRegOut_7_47[16] , \wRegOut_7_47[15] , \wRegOut_7_47[14] , 
        \wRegOut_7_47[13] , \wRegOut_7_47[12] , \wRegOut_7_47[11] , 
        \wRegOut_7_47[10] , \wRegOut_7_47[9] , \wRegOut_7_47[8] , 
        \wRegOut_7_47[7] , \wRegOut_7_47[6] , \wRegOut_7_47[5] , 
        \wRegOut_7_47[4] , \wRegOut_7_47[3] , \wRegOut_7_47[2] , 
        \wRegOut_7_47[1] , \wRegOut_7_47[0] }), .R_Out({\wRegInTop_7_47[31] , 
        \wRegInTop_7_47[30] , \wRegInTop_7_47[29] , \wRegInTop_7_47[28] , 
        \wRegInTop_7_47[27] , \wRegInTop_7_47[26] , \wRegInTop_7_47[25] , 
        \wRegInTop_7_47[24] , \wRegInTop_7_47[23] , \wRegInTop_7_47[22] , 
        \wRegInTop_7_47[21] , \wRegInTop_7_47[20] , \wRegInTop_7_47[19] , 
        \wRegInTop_7_47[18] , \wRegInTop_7_47[17] , \wRegInTop_7_47[16] , 
        \wRegInTop_7_47[15] , \wRegInTop_7_47[14] , \wRegInTop_7_47[13] , 
        \wRegInTop_7_47[12] , \wRegInTop_7_47[11] , \wRegInTop_7_47[10] , 
        \wRegInTop_7_47[9] , \wRegInTop_7_47[8] , \wRegInTop_7_47[7] , 
        \wRegInTop_7_47[6] , \wRegInTop_7_47[5] , \wRegInTop_7_47[4] , 
        \wRegInTop_7_47[3] , \wRegInTop_7_47[2] , \wRegInTop_7_47[1] , 
        \wRegInTop_7_47[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink66[31] , \ScanLink66[30] , \ScanLink66[29] , 
        \ScanLink66[28] , \ScanLink66[27] , \ScanLink66[26] , \ScanLink66[25] , 
        \ScanLink66[24] , \ScanLink66[23] , \ScanLink66[22] , \ScanLink66[21] , 
        \ScanLink66[20] , \ScanLink66[19] , \ScanLink66[18] , \ScanLink66[17] , 
        \ScanLink66[16] , \ScanLink66[15] , \ScanLink66[14] , \ScanLink66[13] , 
        \ScanLink66[12] , \ScanLink66[11] , \ScanLink66[10] , \ScanLink66[9] , 
        \ScanLink66[8] , \ScanLink66[7] , \ScanLink66[6] , \ScanLink66[5] , 
        \ScanLink66[4] , \ScanLink66[3] , \ScanLink66[2] , \ScanLink66[1] , 
        \ScanLink66[0] }), .ScanOut({\ScanLink65[31] , \ScanLink65[30] , 
        \ScanLink65[29] , \ScanLink65[28] , \ScanLink65[27] , \ScanLink65[26] , 
        \ScanLink65[25] , \ScanLink65[24] , \ScanLink65[23] , \ScanLink65[22] , 
        \ScanLink65[21] , \ScanLink65[20] , \ScanLink65[19] , \ScanLink65[18] , 
        \ScanLink65[17] , \ScanLink65[16] , \ScanLink65[15] , \ScanLink65[14] , 
        \ScanLink65[13] , \ScanLink65[12] , \ScanLink65[11] , \ScanLink65[10] , 
        \ScanLink65[9] , \ScanLink65[8] , \ScanLink65[7] , \ScanLink65[6] , 
        \ScanLink65[5] , \ScanLink65[4] , \ScanLink65[3] , \ScanLink65[2] , 
        \ScanLink65[1] , \ScanLink65[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_2[31] , \wRegOut_6_2[30] , \wRegOut_6_2[29] , 
        \wRegOut_6_2[28] , \wRegOut_6_2[27] , \wRegOut_6_2[26] , 
        \wRegOut_6_2[25] , \wRegOut_6_2[24] , \wRegOut_6_2[23] , 
        \wRegOut_6_2[22] , \wRegOut_6_2[21] , \wRegOut_6_2[20] , 
        \wRegOut_6_2[19] , \wRegOut_6_2[18] , \wRegOut_6_2[17] , 
        \wRegOut_6_2[16] , \wRegOut_6_2[15] , \wRegOut_6_2[14] , 
        \wRegOut_6_2[13] , \wRegOut_6_2[12] , \wRegOut_6_2[11] , 
        \wRegOut_6_2[10] , \wRegOut_6_2[9] , \wRegOut_6_2[8] , 
        \wRegOut_6_2[7] , \wRegOut_6_2[6] , \wRegOut_6_2[5] , \wRegOut_6_2[4] , 
        \wRegOut_6_2[3] , \wRegOut_6_2[2] , \wRegOut_6_2[1] , \wRegOut_6_2[0] 
        }), .Enable1(\wRegEnTop_6_2[0] ), .Enable2(\wRegEnBot_6_2[0] ), .In1({
        \wRegInTop_6_2[31] , \wRegInTop_6_2[30] , \wRegInTop_6_2[29] , 
        \wRegInTop_6_2[28] , \wRegInTop_6_2[27] , \wRegInTop_6_2[26] , 
        \wRegInTop_6_2[25] , \wRegInTop_6_2[24] , \wRegInTop_6_2[23] , 
        \wRegInTop_6_2[22] , \wRegInTop_6_2[21] , \wRegInTop_6_2[20] , 
        \wRegInTop_6_2[19] , \wRegInTop_6_2[18] , \wRegInTop_6_2[17] , 
        \wRegInTop_6_2[16] , \wRegInTop_6_2[15] , \wRegInTop_6_2[14] , 
        \wRegInTop_6_2[13] , \wRegInTop_6_2[12] , \wRegInTop_6_2[11] , 
        \wRegInTop_6_2[10] , \wRegInTop_6_2[9] , \wRegInTop_6_2[8] , 
        \wRegInTop_6_2[7] , \wRegInTop_6_2[6] , \wRegInTop_6_2[5] , 
        \wRegInTop_6_2[4] , \wRegInTop_6_2[3] , \wRegInTop_6_2[2] , 
        \wRegInTop_6_2[1] , \wRegInTop_6_2[0] }), .In2({\wRegInBot_6_2[31] , 
        \wRegInBot_6_2[30] , \wRegInBot_6_2[29] , \wRegInBot_6_2[28] , 
        \wRegInBot_6_2[27] , \wRegInBot_6_2[26] , \wRegInBot_6_2[25] , 
        \wRegInBot_6_2[24] , \wRegInBot_6_2[23] , \wRegInBot_6_2[22] , 
        \wRegInBot_6_2[21] , \wRegInBot_6_2[20] , \wRegInBot_6_2[19] , 
        \wRegInBot_6_2[18] , \wRegInBot_6_2[17] , \wRegInBot_6_2[16] , 
        \wRegInBot_6_2[15] , \wRegInBot_6_2[14] , \wRegInBot_6_2[13] , 
        \wRegInBot_6_2[12] , \wRegInBot_6_2[11] , \wRegInBot_6_2[10] , 
        \wRegInBot_6_2[9] , \wRegInBot_6_2[8] , \wRegInBot_6_2[7] , 
        \wRegInBot_6_2[6] , \wRegInBot_6_2[5] , \wRegInBot_6_2[4] , 
        \wRegInBot_6_2[3] , \wRegInBot_6_2[2] , \wRegInBot_6_2[1] , 
        \wRegInBot_6_2[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_58 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink186[31] , \ScanLink186[30] , \ScanLink186[29] , 
        \ScanLink186[28] , \ScanLink186[27] , \ScanLink186[26] , 
        \ScanLink186[25] , \ScanLink186[24] , \ScanLink186[23] , 
        \ScanLink186[22] , \ScanLink186[21] , \ScanLink186[20] , 
        \ScanLink186[19] , \ScanLink186[18] , \ScanLink186[17] , 
        \ScanLink186[16] , \ScanLink186[15] , \ScanLink186[14] , 
        \ScanLink186[13] , \ScanLink186[12] , \ScanLink186[11] , 
        \ScanLink186[10] , \ScanLink186[9] , \ScanLink186[8] , 
        \ScanLink186[7] , \ScanLink186[6] , \ScanLink186[5] , \ScanLink186[4] , 
        \ScanLink186[3] , \ScanLink186[2] , \ScanLink186[1] , \ScanLink186[0] 
        }), .ScanOut({\ScanLink185[31] , \ScanLink185[30] , \ScanLink185[29] , 
        \ScanLink185[28] , \ScanLink185[27] , \ScanLink185[26] , 
        \ScanLink185[25] , \ScanLink185[24] , \ScanLink185[23] , 
        \ScanLink185[22] , \ScanLink185[21] , \ScanLink185[20] , 
        \ScanLink185[19] , \ScanLink185[18] , \ScanLink185[17] , 
        \ScanLink185[16] , \ScanLink185[15] , \ScanLink185[14] , 
        \ScanLink185[13] , \ScanLink185[12] , \ScanLink185[11] , 
        \ScanLink185[10] , \ScanLink185[9] , \ScanLink185[8] , 
        \ScanLink185[7] , \ScanLink185[6] , \ScanLink185[5] , \ScanLink185[4] , 
        \ScanLink185[3] , \ScanLink185[2] , \ScanLink185[1] , \ScanLink185[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_58[31] , 
        \wRegOut_7_58[30] , \wRegOut_7_58[29] , \wRegOut_7_58[28] , 
        \wRegOut_7_58[27] , \wRegOut_7_58[26] , \wRegOut_7_58[25] , 
        \wRegOut_7_58[24] , \wRegOut_7_58[23] , \wRegOut_7_58[22] , 
        \wRegOut_7_58[21] , \wRegOut_7_58[20] , \wRegOut_7_58[19] , 
        \wRegOut_7_58[18] , \wRegOut_7_58[17] , \wRegOut_7_58[16] , 
        \wRegOut_7_58[15] , \wRegOut_7_58[14] , \wRegOut_7_58[13] , 
        \wRegOut_7_58[12] , \wRegOut_7_58[11] , \wRegOut_7_58[10] , 
        \wRegOut_7_58[9] , \wRegOut_7_58[8] , \wRegOut_7_58[7] , 
        \wRegOut_7_58[6] , \wRegOut_7_58[5] , \wRegOut_7_58[4] , 
        \wRegOut_7_58[3] , \wRegOut_7_58[2] , \wRegOut_7_58[1] , 
        \wRegOut_7_58[0] }), .Enable1(\wRegEnTop_7_58[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_58[31] , \wRegInTop_7_58[30] , \wRegInTop_7_58[29] , 
        \wRegInTop_7_58[28] , \wRegInTop_7_58[27] , \wRegInTop_7_58[26] , 
        \wRegInTop_7_58[25] , \wRegInTop_7_58[24] , \wRegInTop_7_58[23] , 
        \wRegInTop_7_58[22] , \wRegInTop_7_58[21] , \wRegInTop_7_58[20] , 
        \wRegInTop_7_58[19] , \wRegInTop_7_58[18] , \wRegInTop_7_58[17] , 
        \wRegInTop_7_58[16] , \wRegInTop_7_58[15] , \wRegInTop_7_58[14] , 
        \wRegInTop_7_58[13] , \wRegInTop_7_58[12] , \wRegInTop_7_58[11] , 
        \wRegInTop_7_58[10] , \wRegInTop_7_58[9] , \wRegInTop_7_58[8] , 
        \wRegInTop_7_58[7] , \wRegInTop_7_58[6] , \wRegInTop_7_58[5] , 
        \wRegInTop_7_58[4] , \wRegInTop_7_58[3] , \wRegInTop_7_58[2] , 
        \wRegInTop_7_58[1] , \wRegInTop_7_58[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink23[31] , \ScanLink23[30] , \ScanLink23[29] , 
        \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , \ScanLink23[25] , 
        \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , \ScanLink23[21] , 
        \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , \ScanLink23[17] , 
        \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , \ScanLink23[13] , 
        \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , \ScanLink23[9] , 
        \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , \ScanLink23[5] , 
        \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , \ScanLink23[1] , 
        \ScanLink23[0] }), .ScanOut({\ScanLink22[31] , \ScanLink22[30] , 
        \ScanLink22[29] , \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , 
        \ScanLink22[25] , \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , 
        \ScanLink22[21] , \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , 
        \ScanLink22[17] , \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , 
        \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , 
        \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , 
        \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , 
        \ScanLink22[1] , \ScanLink22[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_7[31] , \wRegOut_4_7[30] , \wRegOut_4_7[29] , 
        \wRegOut_4_7[28] , \wRegOut_4_7[27] , \wRegOut_4_7[26] , 
        \wRegOut_4_7[25] , \wRegOut_4_7[24] , \wRegOut_4_7[23] , 
        \wRegOut_4_7[22] , \wRegOut_4_7[21] , \wRegOut_4_7[20] , 
        \wRegOut_4_7[19] , \wRegOut_4_7[18] , \wRegOut_4_7[17] , 
        \wRegOut_4_7[16] , \wRegOut_4_7[15] , \wRegOut_4_7[14] , 
        \wRegOut_4_7[13] , \wRegOut_4_7[12] , \wRegOut_4_7[11] , 
        \wRegOut_4_7[10] , \wRegOut_4_7[9] , \wRegOut_4_7[8] , 
        \wRegOut_4_7[7] , \wRegOut_4_7[6] , \wRegOut_4_7[5] , \wRegOut_4_7[4] , 
        \wRegOut_4_7[3] , \wRegOut_4_7[2] , \wRegOut_4_7[1] , \wRegOut_4_7[0] 
        }), .Enable1(\wRegEnTop_4_7[0] ), .Enable2(\wRegEnBot_4_7[0] ), .In1({
        \wRegInTop_4_7[31] , \wRegInTop_4_7[30] , \wRegInTop_4_7[29] , 
        \wRegInTop_4_7[28] , \wRegInTop_4_7[27] , \wRegInTop_4_7[26] , 
        \wRegInTop_4_7[25] , \wRegInTop_4_7[24] , \wRegInTop_4_7[23] , 
        \wRegInTop_4_7[22] , \wRegInTop_4_7[21] , \wRegInTop_4_7[20] , 
        \wRegInTop_4_7[19] , \wRegInTop_4_7[18] , \wRegInTop_4_7[17] , 
        \wRegInTop_4_7[16] , \wRegInTop_4_7[15] , \wRegInTop_4_7[14] , 
        \wRegInTop_4_7[13] , \wRegInTop_4_7[12] , \wRegInTop_4_7[11] , 
        \wRegInTop_4_7[10] , \wRegInTop_4_7[9] , \wRegInTop_4_7[8] , 
        \wRegInTop_4_7[7] , \wRegInTop_4_7[6] , \wRegInTop_4_7[5] , 
        \wRegInTop_4_7[4] , \wRegInTop_4_7[3] , \wRegInTop_4_7[2] , 
        \wRegInTop_4_7[1] , \wRegInTop_4_7[0] }), .In2({\wRegInBot_4_7[31] , 
        \wRegInBot_4_7[30] , \wRegInBot_4_7[29] , \wRegInBot_4_7[28] , 
        \wRegInBot_4_7[27] , \wRegInBot_4_7[26] , \wRegInBot_4_7[25] , 
        \wRegInBot_4_7[24] , \wRegInBot_4_7[23] , \wRegInBot_4_7[22] , 
        \wRegInBot_4_7[21] , \wRegInBot_4_7[20] , \wRegInBot_4_7[19] , 
        \wRegInBot_4_7[18] , \wRegInBot_4_7[17] , \wRegInBot_4_7[16] , 
        \wRegInBot_4_7[15] , \wRegInBot_4_7[14] , \wRegInBot_4_7[13] , 
        \wRegInBot_4_7[12] , \wRegInBot_4_7[11] , \wRegInBot_4_7[10] , 
        \wRegInBot_4_7[9] , \wRegInBot_4_7[8] , \wRegInBot_4_7[7] , 
        \wRegInBot_4_7[6] , \wRegInBot_4_7[5] , \wRegInBot_4_7[4] , 
        \wRegInBot_4_7[3] , \wRegInBot_4_7[2] , \wRegInBot_4_7[1] , 
        \wRegInBot_4_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_27 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink59[31] , \ScanLink59[30] , \ScanLink59[29] , 
        \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , \ScanLink59[25] , 
        \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , \ScanLink59[21] , 
        \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , \ScanLink59[17] , 
        \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , \ScanLink59[13] , 
        \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , \ScanLink59[9] , 
        \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , \ScanLink59[5] , 
        \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , \ScanLink59[1] , 
        \ScanLink59[0] }), .ScanOut({\ScanLink58[31] , \ScanLink58[30] , 
        \ScanLink58[29] , \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , 
        \ScanLink58[25] , \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , 
        \ScanLink58[21] , \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , 
        \ScanLink58[17] , \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , 
        \ScanLink58[13] , \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , 
        \ScanLink58[9] , \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , 
        \ScanLink58[5] , \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , 
        \ScanLink58[1] , \ScanLink58[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_27[31] , \wRegOut_5_27[30] , 
        \wRegOut_5_27[29] , \wRegOut_5_27[28] , \wRegOut_5_27[27] , 
        \wRegOut_5_27[26] , \wRegOut_5_27[25] , \wRegOut_5_27[24] , 
        \wRegOut_5_27[23] , \wRegOut_5_27[22] , \wRegOut_5_27[21] , 
        \wRegOut_5_27[20] , \wRegOut_5_27[19] , \wRegOut_5_27[18] , 
        \wRegOut_5_27[17] , \wRegOut_5_27[16] , \wRegOut_5_27[15] , 
        \wRegOut_5_27[14] , \wRegOut_5_27[13] , \wRegOut_5_27[12] , 
        \wRegOut_5_27[11] , \wRegOut_5_27[10] , \wRegOut_5_27[9] , 
        \wRegOut_5_27[8] , \wRegOut_5_27[7] , \wRegOut_5_27[6] , 
        \wRegOut_5_27[5] , \wRegOut_5_27[4] , \wRegOut_5_27[3] , 
        \wRegOut_5_27[2] , \wRegOut_5_27[1] , \wRegOut_5_27[0] }), .Enable1(
        \wRegEnTop_5_27[0] ), .Enable2(\wRegEnBot_5_27[0] ), .In1({
        \wRegInTop_5_27[31] , \wRegInTop_5_27[30] , \wRegInTop_5_27[29] , 
        \wRegInTop_5_27[28] , \wRegInTop_5_27[27] , \wRegInTop_5_27[26] , 
        \wRegInTop_5_27[25] , \wRegInTop_5_27[24] , \wRegInTop_5_27[23] , 
        \wRegInTop_5_27[22] , \wRegInTop_5_27[21] , \wRegInTop_5_27[20] , 
        \wRegInTop_5_27[19] , \wRegInTop_5_27[18] , \wRegInTop_5_27[17] , 
        \wRegInTop_5_27[16] , \wRegInTop_5_27[15] , \wRegInTop_5_27[14] , 
        \wRegInTop_5_27[13] , \wRegInTop_5_27[12] , \wRegInTop_5_27[11] , 
        \wRegInTop_5_27[10] , \wRegInTop_5_27[9] , \wRegInTop_5_27[8] , 
        \wRegInTop_5_27[7] , \wRegInTop_5_27[6] , \wRegInTop_5_27[5] , 
        \wRegInTop_5_27[4] , \wRegInTop_5_27[3] , \wRegInTop_5_27[2] , 
        \wRegInTop_5_27[1] , \wRegInTop_5_27[0] }), .In2({\wRegInBot_5_27[31] , 
        \wRegInBot_5_27[30] , \wRegInBot_5_27[29] , \wRegInBot_5_27[28] , 
        \wRegInBot_5_27[27] , \wRegInBot_5_27[26] , \wRegInBot_5_27[25] , 
        \wRegInBot_5_27[24] , \wRegInBot_5_27[23] , \wRegInBot_5_27[22] , 
        \wRegInBot_5_27[21] , \wRegInBot_5_27[20] , \wRegInBot_5_27[19] , 
        \wRegInBot_5_27[18] , \wRegInBot_5_27[17] , \wRegInBot_5_27[16] , 
        \wRegInBot_5_27[15] , \wRegInBot_5_27[14] , \wRegInBot_5_27[13] , 
        \wRegInBot_5_27[12] , \wRegInBot_5_27[11] , \wRegInBot_5_27[10] , 
        \wRegInBot_5_27[9] , \wRegInBot_5_27[8] , \wRegInBot_5_27[7] , 
        \wRegInBot_5_27[6] , \wRegInBot_5_27[5] , \wRegInBot_5_27[4] , 
        \wRegInBot_5_27[3] , \wRegInBot_5_27[2] , \wRegInBot_5_27[1] , 
        \wRegInBot_5_27[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_45 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink109[31] , \ScanLink109[30] , \ScanLink109[29] , 
        \ScanLink109[28] , \ScanLink109[27] , \ScanLink109[26] , 
        \ScanLink109[25] , \ScanLink109[24] , \ScanLink109[23] , 
        \ScanLink109[22] , \ScanLink109[21] , \ScanLink109[20] , 
        \ScanLink109[19] , \ScanLink109[18] , \ScanLink109[17] , 
        \ScanLink109[16] , \ScanLink109[15] , \ScanLink109[14] , 
        \ScanLink109[13] , \ScanLink109[12] , \ScanLink109[11] , 
        \ScanLink109[10] , \ScanLink109[9] , \ScanLink109[8] , 
        \ScanLink109[7] , \ScanLink109[6] , \ScanLink109[5] , \ScanLink109[4] , 
        \ScanLink109[3] , \ScanLink109[2] , \ScanLink109[1] , \ScanLink109[0] 
        }), .ScanOut({\ScanLink108[31] , \ScanLink108[30] , \ScanLink108[29] , 
        \ScanLink108[28] , \ScanLink108[27] , \ScanLink108[26] , 
        \ScanLink108[25] , \ScanLink108[24] , \ScanLink108[23] , 
        \ScanLink108[22] , \ScanLink108[21] , \ScanLink108[20] , 
        \ScanLink108[19] , \ScanLink108[18] , \ScanLink108[17] , 
        \ScanLink108[16] , \ScanLink108[15] , \ScanLink108[14] , 
        \ScanLink108[13] , \ScanLink108[12] , \ScanLink108[11] , 
        \ScanLink108[10] , \ScanLink108[9] , \ScanLink108[8] , 
        \ScanLink108[7] , \ScanLink108[6] , \ScanLink108[5] , \ScanLink108[4] , 
        \ScanLink108[3] , \ScanLink108[2] , \ScanLink108[1] , \ScanLink108[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_45[31] , 
        \wRegOut_6_45[30] , \wRegOut_6_45[29] , \wRegOut_6_45[28] , 
        \wRegOut_6_45[27] , \wRegOut_6_45[26] , \wRegOut_6_45[25] , 
        \wRegOut_6_45[24] , \wRegOut_6_45[23] , \wRegOut_6_45[22] , 
        \wRegOut_6_45[21] , \wRegOut_6_45[20] , \wRegOut_6_45[19] , 
        \wRegOut_6_45[18] , \wRegOut_6_45[17] , \wRegOut_6_45[16] , 
        \wRegOut_6_45[15] , \wRegOut_6_45[14] , \wRegOut_6_45[13] , 
        \wRegOut_6_45[12] , \wRegOut_6_45[11] , \wRegOut_6_45[10] , 
        \wRegOut_6_45[9] , \wRegOut_6_45[8] , \wRegOut_6_45[7] , 
        \wRegOut_6_45[6] , \wRegOut_6_45[5] , \wRegOut_6_45[4] , 
        \wRegOut_6_45[3] , \wRegOut_6_45[2] , \wRegOut_6_45[1] , 
        \wRegOut_6_45[0] }), .Enable1(\wRegEnTop_6_45[0] ), .Enable2(
        \wRegEnBot_6_45[0] ), .In1({\wRegInTop_6_45[31] , \wRegInTop_6_45[30] , 
        \wRegInTop_6_45[29] , \wRegInTop_6_45[28] , \wRegInTop_6_45[27] , 
        \wRegInTop_6_45[26] , \wRegInTop_6_45[25] , \wRegInTop_6_45[24] , 
        \wRegInTop_6_45[23] , \wRegInTop_6_45[22] , \wRegInTop_6_45[21] , 
        \wRegInTop_6_45[20] , \wRegInTop_6_45[19] , \wRegInTop_6_45[18] , 
        \wRegInTop_6_45[17] , \wRegInTop_6_45[16] , \wRegInTop_6_45[15] , 
        \wRegInTop_6_45[14] , \wRegInTop_6_45[13] , \wRegInTop_6_45[12] , 
        \wRegInTop_6_45[11] , \wRegInTop_6_45[10] , \wRegInTop_6_45[9] , 
        \wRegInTop_6_45[8] , \wRegInTop_6_45[7] , \wRegInTop_6_45[6] , 
        \wRegInTop_6_45[5] , \wRegInTop_6_45[4] , \wRegInTop_6_45[3] , 
        \wRegInTop_6_45[2] , \wRegInTop_6_45[1] , \wRegInTop_6_45[0] }), .In2(
        {\wRegInBot_6_45[31] , \wRegInBot_6_45[30] , \wRegInBot_6_45[29] , 
        \wRegInBot_6_45[28] , \wRegInBot_6_45[27] , \wRegInBot_6_45[26] , 
        \wRegInBot_6_45[25] , \wRegInBot_6_45[24] , \wRegInBot_6_45[23] , 
        \wRegInBot_6_45[22] , \wRegInBot_6_45[21] , \wRegInBot_6_45[20] , 
        \wRegInBot_6_45[19] , \wRegInBot_6_45[18] , \wRegInBot_6_45[17] , 
        \wRegInBot_6_45[16] , \wRegInBot_6_45[15] , \wRegInBot_6_45[14] , 
        \wRegInBot_6_45[13] , \wRegInBot_6_45[12] , \wRegInBot_6_45[11] , 
        \wRegInBot_6_45[10] , \wRegInBot_6_45[9] , \wRegInBot_6_45[8] , 
        \wRegInBot_6_45[7] , \wRegInBot_6_45[6] , \wRegInBot_6_45[5] , 
        \wRegInBot_6_45[4] , \wRegInBot_6_45[3] , \wRegInBot_6_45[2] , 
        \wRegInBot_6_45[1] , \wRegInBot_6_45[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_62 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink126[31] , \ScanLink126[30] , \ScanLink126[29] , 
        \ScanLink126[28] , \ScanLink126[27] , \ScanLink126[26] , 
        \ScanLink126[25] , \ScanLink126[24] , \ScanLink126[23] , 
        \ScanLink126[22] , \ScanLink126[21] , \ScanLink126[20] , 
        \ScanLink126[19] , \ScanLink126[18] , \ScanLink126[17] , 
        \ScanLink126[16] , \ScanLink126[15] , \ScanLink126[14] , 
        \ScanLink126[13] , \ScanLink126[12] , \ScanLink126[11] , 
        \ScanLink126[10] , \ScanLink126[9] , \ScanLink126[8] , 
        \ScanLink126[7] , \ScanLink126[6] , \ScanLink126[5] , \ScanLink126[4] , 
        \ScanLink126[3] , \ScanLink126[2] , \ScanLink126[1] , \ScanLink126[0] 
        }), .ScanOut({\ScanLink125[31] , \ScanLink125[30] , \ScanLink125[29] , 
        \ScanLink125[28] , \ScanLink125[27] , \ScanLink125[26] , 
        \ScanLink125[25] , \ScanLink125[24] , \ScanLink125[23] , 
        \ScanLink125[22] , \ScanLink125[21] , \ScanLink125[20] , 
        \ScanLink125[19] , \ScanLink125[18] , \ScanLink125[17] , 
        \ScanLink125[16] , \ScanLink125[15] , \ScanLink125[14] , 
        \ScanLink125[13] , \ScanLink125[12] , \ScanLink125[11] , 
        \ScanLink125[10] , \ScanLink125[9] , \ScanLink125[8] , 
        \ScanLink125[7] , \ScanLink125[6] , \ScanLink125[5] , \ScanLink125[4] , 
        \ScanLink125[3] , \ScanLink125[2] , \ScanLink125[1] , \ScanLink125[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_62[31] , 
        \wRegOut_6_62[30] , \wRegOut_6_62[29] , \wRegOut_6_62[28] , 
        \wRegOut_6_62[27] , \wRegOut_6_62[26] , \wRegOut_6_62[25] , 
        \wRegOut_6_62[24] , \wRegOut_6_62[23] , \wRegOut_6_62[22] , 
        \wRegOut_6_62[21] , \wRegOut_6_62[20] , \wRegOut_6_62[19] , 
        \wRegOut_6_62[18] , \wRegOut_6_62[17] , \wRegOut_6_62[16] , 
        \wRegOut_6_62[15] , \wRegOut_6_62[14] , \wRegOut_6_62[13] , 
        \wRegOut_6_62[12] , \wRegOut_6_62[11] , \wRegOut_6_62[10] , 
        \wRegOut_6_62[9] , \wRegOut_6_62[8] , \wRegOut_6_62[7] , 
        \wRegOut_6_62[6] , \wRegOut_6_62[5] , \wRegOut_6_62[4] , 
        \wRegOut_6_62[3] , \wRegOut_6_62[2] , \wRegOut_6_62[1] , 
        \wRegOut_6_62[0] }), .Enable1(\wRegEnTop_6_62[0] ), .Enable2(
        \wRegEnBot_6_62[0] ), .In1({\wRegInTop_6_62[31] , \wRegInTop_6_62[30] , 
        \wRegInTop_6_62[29] , \wRegInTop_6_62[28] , \wRegInTop_6_62[27] , 
        \wRegInTop_6_62[26] , \wRegInTop_6_62[25] , \wRegInTop_6_62[24] , 
        \wRegInTop_6_62[23] , \wRegInTop_6_62[22] , \wRegInTop_6_62[21] , 
        \wRegInTop_6_62[20] , \wRegInTop_6_62[19] , \wRegInTop_6_62[18] , 
        \wRegInTop_6_62[17] , \wRegInTop_6_62[16] , \wRegInTop_6_62[15] , 
        \wRegInTop_6_62[14] , \wRegInTop_6_62[13] , \wRegInTop_6_62[12] , 
        \wRegInTop_6_62[11] , \wRegInTop_6_62[10] , \wRegInTop_6_62[9] , 
        \wRegInTop_6_62[8] , \wRegInTop_6_62[7] , \wRegInTop_6_62[6] , 
        \wRegInTop_6_62[5] , \wRegInTop_6_62[4] , \wRegInTop_6_62[3] , 
        \wRegInTop_6_62[2] , \wRegInTop_6_62[1] , \wRegInTop_6_62[0] }), .In2(
        {\wRegInBot_6_62[31] , \wRegInBot_6_62[30] , \wRegInBot_6_62[29] , 
        \wRegInBot_6_62[28] , \wRegInBot_6_62[27] , \wRegInBot_6_62[26] , 
        \wRegInBot_6_62[25] , \wRegInBot_6_62[24] , \wRegInBot_6_62[23] , 
        \wRegInBot_6_62[22] , \wRegInBot_6_62[21] , \wRegInBot_6_62[20] , 
        \wRegInBot_6_62[19] , \wRegInBot_6_62[18] , \wRegInBot_6_62[17] , 
        \wRegInBot_6_62[16] , \wRegInBot_6_62[15] , \wRegInBot_6_62[14] , 
        \wRegInBot_6_62[13] , \wRegInBot_6_62[12] , \wRegInBot_6_62[11] , 
        \wRegInBot_6_62[10] , \wRegInBot_6_62[9] , \wRegInBot_6_62[8] , 
        \wRegInBot_6_62[7] , \wRegInBot_6_62[6] , \wRegInBot_6_62[5] , 
        \wRegInBot_6_62[4] , \wRegInBot_6_62[3] , \wRegInBot_6_62[2] , 
        \wRegInBot_6_62[1] , \wRegInBot_6_62[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_78 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink206[31] , \ScanLink206[30] , \ScanLink206[29] , 
        \ScanLink206[28] , \ScanLink206[27] , \ScanLink206[26] , 
        \ScanLink206[25] , \ScanLink206[24] , \ScanLink206[23] , 
        \ScanLink206[22] , \ScanLink206[21] , \ScanLink206[20] , 
        \ScanLink206[19] , \ScanLink206[18] , \ScanLink206[17] , 
        \ScanLink206[16] , \ScanLink206[15] , \ScanLink206[14] , 
        \ScanLink206[13] , \ScanLink206[12] , \ScanLink206[11] , 
        \ScanLink206[10] , \ScanLink206[9] , \ScanLink206[8] , 
        \ScanLink206[7] , \ScanLink206[6] , \ScanLink206[5] , \ScanLink206[4] , 
        \ScanLink206[3] , \ScanLink206[2] , \ScanLink206[1] , \ScanLink206[0] 
        }), .ScanOut({\ScanLink205[31] , \ScanLink205[30] , \ScanLink205[29] , 
        \ScanLink205[28] , \ScanLink205[27] , \ScanLink205[26] , 
        \ScanLink205[25] , \ScanLink205[24] , \ScanLink205[23] , 
        \ScanLink205[22] , \ScanLink205[21] , \ScanLink205[20] , 
        \ScanLink205[19] , \ScanLink205[18] , \ScanLink205[17] , 
        \ScanLink205[16] , \ScanLink205[15] , \ScanLink205[14] , 
        \ScanLink205[13] , \ScanLink205[12] , \ScanLink205[11] , 
        \ScanLink205[10] , \ScanLink205[9] , \ScanLink205[8] , 
        \ScanLink205[7] , \ScanLink205[6] , \ScanLink205[5] , \ScanLink205[4] , 
        \ScanLink205[3] , \ScanLink205[2] , \ScanLink205[1] , \ScanLink205[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_78[31] , 
        \wRegOut_7_78[30] , \wRegOut_7_78[29] , \wRegOut_7_78[28] , 
        \wRegOut_7_78[27] , \wRegOut_7_78[26] , \wRegOut_7_78[25] , 
        \wRegOut_7_78[24] , \wRegOut_7_78[23] , \wRegOut_7_78[22] , 
        \wRegOut_7_78[21] , \wRegOut_7_78[20] , \wRegOut_7_78[19] , 
        \wRegOut_7_78[18] , \wRegOut_7_78[17] , \wRegOut_7_78[16] , 
        \wRegOut_7_78[15] , \wRegOut_7_78[14] , \wRegOut_7_78[13] , 
        \wRegOut_7_78[12] , \wRegOut_7_78[11] , \wRegOut_7_78[10] , 
        \wRegOut_7_78[9] , \wRegOut_7_78[8] , \wRegOut_7_78[7] , 
        \wRegOut_7_78[6] , \wRegOut_7_78[5] , \wRegOut_7_78[4] , 
        \wRegOut_7_78[3] , \wRegOut_7_78[2] , \wRegOut_7_78[1] , 
        \wRegOut_7_78[0] }), .Enable1(\wRegEnTop_7_78[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_78[31] , \wRegInTop_7_78[30] , \wRegInTop_7_78[29] , 
        \wRegInTop_7_78[28] , \wRegInTop_7_78[27] , \wRegInTop_7_78[26] , 
        \wRegInTop_7_78[25] , \wRegInTop_7_78[24] , \wRegInTop_7_78[23] , 
        \wRegInTop_7_78[22] , \wRegInTop_7_78[21] , \wRegInTop_7_78[20] , 
        \wRegInTop_7_78[19] , \wRegInTop_7_78[18] , \wRegInTop_7_78[17] , 
        \wRegInTop_7_78[16] , \wRegInTop_7_78[15] , \wRegInTop_7_78[14] , 
        \wRegInTop_7_78[13] , \wRegInTop_7_78[12] , \wRegInTop_7_78[11] , 
        \wRegInTop_7_78[10] , \wRegInTop_7_78[9] , \wRegInTop_7_78[8] , 
        \wRegInTop_7_78[7] , \wRegInTop_7_78[6] , \wRegInTop_7_78[5] , 
        \wRegInTop_7_78[4] , \wRegInTop_7_78[3] , \wRegInTop_7_78[2] , 
        \wRegInTop_7_78[1] , \wRegInTop_7_78[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_14[0] ), .P_In({\wRegOut_5_14[31] , 
        \wRegOut_5_14[30] , \wRegOut_5_14[29] , \wRegOut_5_14[28] , 
        \wRegOut_5_14[27] , \wRegOut_5_14[26] , \wRegOut_5_14[25] , 
        \wRegOut_5_14[24] , \wRegOut_5_14[23] , \wRegOut_5_14[22] , 
        \wRegOut_5_14[21] , \wRegOut_5_14[20] , \wRegOut_5_14[19] , 
        \wRegOut_5_14[18] , \wRegOut_5_14[17] , \wRegOut_5_14[16] , 
        \wRegOut_5_14[15] , \wRegOut_5_14[14] , \wRegOut_5_14[13] , 
        \wRegOut_5_14[12] , \wRegOut_5_14[11] , \wRegOut_5_14[10] , 
        \wRegOut_5_14[9] , \wRegOut_5_14[8] , \wRegOut_5_14[7] , 
        \wRegOut_5_14[6] , \wRegOut_5_14[5] , \wRegOut_5_14[4] , 
        \wRegOut_5_14[3] , \wRegOut_5_14[2] , \wRegOut_5_14[1] , 
        \wRegOut_5_14[0] }), .P_Out({\wRegInBot_5_14[31] , 
        \wRegInBot_5_14[30] , \wRegInBot_5_14[29] , \wRegInBot_5_14[28] , 
        \wRegInBot_5_14[27] , \wRegInBot_5_14[26] , \wRegInBot_5_14[25] , 
        \wRegInBot_5_14[24] , \wRegInBot_5_14[23] , \wRegInBot_5_14[22] , 
        \wRegInBot_5_14[21] , \wRegInBot_5_14[20] , \wRegInBot_5_14[19] , 
        \wRegInBot_5_14[18] , \wRegInBot_5_14[17] , \wRegInBot_5_14[16] , 
        \wRegInBot_5_14[15] , \wRegInBot_5_14[14] , \wRegInBot_5_14[13] , 
        \wRegInBot_5_14[12] , \wRegInBot_5_14[11] , \wRegInBot_5_14[10] , 
        \wRegInBot_5_14[9] , \wRegInBot_5_14[8] , \wRegInBot_5_14[7] , 
        \wRegInBot_5_14[6] , \wRegInBot_5_14[5] , \wRegInBot_5_14[4] , 
        \wRegInBot_5_14[3] , \wRegInBot_5_14[2] , \wRegInBot_5_14[1] , 
        \wRegInBot_5_14[0] }), .L_WR(\wRegEnTop_6_28[0] ), .L_In({
        \wRegOut_6_28[31] , \wRegOut_6_28[30] , \wRegOut_6_28[29] , 
        \wRegOut_6_28[28] , \wRegOut_6_28[27] , \wRegOut_6_28[26] , 
        \wRegOut_6_28[25] , \wRegOut_6_28[24] , \wRegOut_6_28[23] , 
        \wRegOut_6_28[22] , \wRegOut_6_28[21] , \wRegOut_6_28[20] , 
        \wRegOut_6_28[19] , \wRegOut_6_28[18] , \wRegOut_6_28[17] , 
        \wRegOut_6_28[16] , \wRegOut_6_28[15] , \wRegOut_6_28[14] , 
        \wRegOut_6_28[13] , \wRegOut_6_28[12] , \wRegOut_6_28[11] , 
        \wRegOut_6_28[10] , \wRegOut_6_28[9] , \wRegOut_6_28[8] , 
        \wRegOut_6_28[7] , \wRegOut_6_28[6] , \wRegOut_6_28[5] , 
        \wRegOut_6_28[4] , \wRegOut_6_28[3] , \wRegOut_6_28[2] , 
        \wRegOut_6_28[1] , \wRegOut_6_28[0] }), .L_Out({\wRegInTop_6_28[31] , 
        \wRegInTop_6_28[30] , \wRegInTop_6_28[29] , \wRegInTop_6_28[28] , 
        \wRegInTop_6_28[27] , \wRegInTop_6_28[26] , \wRegInTop_6_28[25] , 
        \wRegInTop_6_28[24] , \wRegInTop_6_28[23] , \wRegInTop_6_28[22] , 
        \wRegInTop_6_28[21] , \wRegInTop_6_28[20] , \wRegInTop_6_28[19] , 
        \wRegInTop_6_28[18] , \wRegInTop_6_28[17] , \wRegInTop_6_28[16] , 
        \wRegInTop_6_28[15] , \wRegInTop_6_28[14] , \wRegInTop_6_28[13] , 
        \wRegInTop_6_28[12] , \wRegInTop_6_28[11] , \wRegInTop_6_28[10] , 
        \wRegInTop_6_28[9] , \wRegInTop_6_28[8] , \wRegInTop_6_28[7] , 
        \wRegInTop_6_28[6] , \wRegInTop_6_28[5] , \wRegInTop_6_28[4] , 
        \wRegInTop_6_28[3] , \wRegInTop_6_28[2] , \wRegInTop_6_28[1] , 
        \wRegInTop_6_28[0] }), .R_WR(\wRegEnTop_6_29[0] ), .R_In({
        \wRegOut_6_29[31] , \wRegOut_6_29[30] , \wRegOut_6_29[29] , 
        \wRegOut_6_29[28] , \wRegOut_6_29[27] , \wRegOut_6_29[26] , 
        \wRegOut_6_29[25] , \wRegOut_6_29[24] , \wRegOut_6_29[23] , 
        \wRegOut_6_29[22] , \wRegOut_6_29[21] , \wRegOut_6_29[20] , 
        \wRegOut_6_29[19] , \wRegOut_6_29[18] , \wRegOut_6_29[17] , 
        \wRegOut_6_29[16] , \wRegOut_6_29[15] , \wRegOut_6_29[14] , 
        \wRegOut_6_29[13] , \wRegOut_6_29[12] , \wRegOut_6_29[11] , 
        \wRegOut_6_29[10] , \wRegOut_6_29[9] , \wRegOut_6_29[8] , 
        \wRegOut_6_29[7] , \wRegOut_6_29[6] , \wRegOut_6_29[5] , 
        \wRegOut_6_29[4] , \wRegOut_6_29[3] , \wRegOut_6_29[2] , 
        \wRegOut_6_29[1] , \wRegOut_6_29[0] }), .R_Out({\wRegInTop_6_29[31] , 
        \wRegInTop_6_29[30] , \wRegInTop_6_29[29] , \wRegInTop_6_29[28] , 
        \wRegInTop_6_29[27] , \wRegInTop_6_29[26] , \wRegInTop_6_29[25] , 
        \wRegInTop_6_29[24] , \wRegInTop_6_29[23] , \wRegInTop_6_29[22] , 
        \wRegInTop_6_29[21] , \wRegInTop_6_29[20] , \wRegInTop_6_29[19] , 
        \wRegInTop_6_29[18] , \wRegInTop_6_29[17] , \wRegInTop_6_29[16] , 
        \wRegInTop_6_29[15] , \wRegInTop_6_29[14] , \wRegInTop_6_29[13] , 
        \wRegInTop_6_29[12] , \wRegInTop_6_29[11] , \wRegInTop_6_29[10] , 
        \wRegInTop_6_29[9] , \wRegInTop_6_29[8] , \wRegInTop_6_29[7] , 
        \wRegInTop_6_29[6] , \wRegInTop_6_29[5] , \wRegInTop_6_29[4] , 
        \wRegInTop_6_29[3] , \wRegInTop_6_29[2] , \wRegInTop_6_29[1] , 
        \wRegInTop_6_29[0] }) );
    BHeap_Node_WIDTH32 BHN_6_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_24[0] ), .P_In({\wRegOut_6_24[31] , 
        \wRegOut_6_24[30] , \wRegOut_6_24[29] , \wRegOut_6_24[28] , 
        \wRegOut_6_24[27] , \wRegOut_6_24[26] , \wRegOut_6_24[25] , 
        \wRegOut_6_24[24] , \wRegOut_6_24[23] , \wRegOut_6_24[22] , 
        \wRegOut_6_24[21] , \wRegOut_6_24[20] , \wRegOut_6_24[19] , 
        \wRegOut_6_24[18] , \wRegOut_6_24[17] , \wRegOut_6_24[16] , 
        \wRegOut_6_24[15] , \wRegOut_6_24[14] , \wRegOut_6_24[13] , 
        \wRegOut_6_24[12] , \wRegOut_6_24[11] , \wRegOut_6_24[10] , 
        \wRegOut_6_24[9] , \wRegOut_6_24[8] , \wRegOut_6_24[7] , 
        \wRegOut_6_24[6] , \wRegOut_6_24[5] , \wRegOut_6_24[4] , 
        \wRegOut_6_24[3] , \wRegOut_6_24[2] , \wRegOut_6_24[1] , 
        \wRegOut_6_24[0] }), .P_Out({\wRegInBot_6_24[31] , 
        \wRegInBot_6_24[30] , \wRegInBot_6_24[29] , \wRegInBot_6_24[28] , 
        \wRegInBot_6_24[27] , \wRegInBot_6_24[26] , \wRegInBot_6_24[25] , 
        \wRegInBot_6_24[24] , \wRegInBot_6_24[23] , \wRegInBot_6_24[22] , 
        \wRegInBot_6_24[21] , \wRegInBot_6_24[20] , \wRegInBot_6_24[19] , 
        \wRegInBot_6_24[18] , \wRegInBot_6_24[17] , \wRegInBot_6_24[16] , 
        \wRegInBot_6_24[15] , \wRegInBot_6_24[14] , \wRegInBot_6_24[13] , 
        \wRegInBot_6_24[12] , \wRegInBot_6_24[11] , \wRegInBot_6_24[10] , 
        \wRegInBot_6_24[9] , \wRegInBot_6_24[8] , \wRegInBot_6_24[7] , 
        \wRegInBot_6_24[6] , \wRegInBot_6_24[5] , \wRegInBot_6_24[4] , 
        \wRegInBot_6_24[3] , \wRegInBot_6_24[2] , \wRegInBot_6_24[1] , 
        \wRegInBot_6_24[0] }), .L_WR(\wRegEnTop_7_48[0] ), .L_In({
        \wRegOut_7_48[31] , \wRegOut_7_48[30] , \wRegOut_7_48[29] , 
        \wRegOut_7_48[28] , \wRegOut_7_48[27] , \wRegOut_7_48[26] , 
        \wRegOut_7_48[25] , \wRegOut_7_48[24] , \wRegOut_7_48[23] , 
        \wRegOut_7_48[22] , \wRegOut_7_48[21] , \wRegOut_7_48[20] , 
        \wRegOut_7_48[19] , \wRegOut_7_48[18] , \wRegOut_7_48[17] , 
        \wRegOut_7_48[16] , \wRegOut_7_48[15] , \wRegOut_7_48[14] , 
        \wRegOut_7_48[13] , \wRegOut_7_48[12] , \wRegOut_7_48[11] , 
        \wRegOut_7_48[10] , \wRegOut_7_48[9] , \wRegOut_7_48[8] , 
        \wRegOut_7_48[7] , \wRegOut_7_48[6] , \wRegOut_7_48[5] , 
        \wRegOut_7_48[4] , \wRegOut_7_48[3] , \wRegOut_7_48[2] , 
        \wRegOut_7_48[1] , \wRegOut_7_48[0] }), .L_Out({\wRegInTop_7_48[31] , 
        \wRegInTop_7_48[30] , \wRegInTop_7_48[29] , \wRegInTop_7_48[28] , 
        \wRegInTop_7_48[27] , \wRegInTop_7_48[26] , \wRegInTop_7_48[25] , 
        \wRegInTop_7_48[24] , \wRegInTop_7_48[23] , \wRegInTop_7_48[22] , 
        \wRegInTop_7_48[21] , \wRegInTop_7_48[20] , \wRegInTop_7_48[19] , 
        \wRegInTop_7_48[18] , \wRegInTop_7_48[17] , \wRegInTop_7_48[16] , 
        \wRegInTop_7_48[15] , \wRegInTop_7_48[14] , \wRegInTop_7_48[13] , 
        \wRegInTop_7_48[12] , \wRegInTop_7_48[11] , \wRegInTop_7_48[10] , 
        \wRegInTop_7_48[9] , \wRegInTop_7_48[8] , \wRegInTop_7_48[7] , 
        \wRegInTop_7_48[6] , \wRegInTop_7_48[5] , \wRegInTop_7_48[4] , 
        \wRegInTop_7_48[3] , \wRegInTop_7_48[2] , \wRegInTop_7_48[1] , 
        \wRegInTop_7_48[0] }), .R_WR(\wRegEnTop_7_49[0] ), .R_In({
        \wRegOut_7_49[31] , \wRegOut_7_49[30] , \wRegOut_7_49[29] , 
        \wRegOut_7_49[28] , \wRegOut_7_49[27] , \wRegOut_7_49[26] , 
        \wRegOut_7_49[25] , \wRegOut_7_49[24] , \wRegOut_7_49[23] , 
        \wRegOut_7_49[22] , \wRegOut_7_49[21] , \wRegOut_7_49[20] , 
        \wRegOut_7_49[19] , \wRegOut_7_49[18] , \wRegOut_7_49[17] , 
        \wRegOut_7_49[16] , \wRegOut_7_49[15] , \wRegOut_7_49[14] , 
        \wRegOut_7_49[13] , \wRegOut_7_49[12] , \wRegOut_7_49[11] , 
        \wRegOut_7_49[10] , \wRegOut_7_49[9] , \wRegOut_7_49[8] , 
        \wRegOut_7_49[7] , \wRegOut_7_49[6] , \wRegOut_7_49[5] , 
        \wRegOut_7_49[4] , \wRegOut_7_49[3] , \wRegOut_7_49[2] , 
        \wRegOut_7_49[1] , \wRegOut_7_49[0] }), .R_Out({\wRegInTop_7_49[31] , 
        \wRegInTop_7_49[30] , \wRegInTop_7_49[29] , \wRegInTop_7_49[28] , 
        \wRegInTop_7_49[27] , \wRegInTop_7_49[26] , \wRegInTop_7_49[25] , 
        \wRegInTop_7_49[24] , \wRegInTop_7_49[23] , \wRegInTop_7_49[22] , 
        \wRegInTop_7_49[21] , \wRegInTop_7_49[20] , \wRegInTop_7_49[19] , 
        \wRegInTop_7_49[18] , \wRegInTop_7_49[17] , \wRegInTop_7_49[16] , 
        \wRegInTop_7_49[15] , \wRegInTop_7_49[14] , \wRegInTop_7_49[13] , 
        \wRegInTop_7_49[12] , \wRegInTop_7_49[11] , \wRegInTop_7_49[10] , 
        \wRegInTop_7_49[9] , \wRegInTop_7_49[8] , \wRegInTop_7_49[7] , 
        \wRegInTop_7_49[6] , \wRegInTop_7_49[5] , \wRegInTop_7_49[4] , 
        \wRegInTop_7_49[3] , \wRegInTop_7_49[2] , \wRegInTop_7_49[1] , 
        \wRegInTop_7_49[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_102 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink230[31] , \ScanLink230[30] , \ScanLink230[29] , 
        \ScanLink230[28] , \ScanLink230[27] , \ScanLink230[26] , 
        \ScanLink230[25] , \ScanLink230[24] , \ScanLink230[23] , 
        \ScanLink230[22] , \ScanLink230[21] , \ScanLink230[20] , 
        \ScanLink230[19] , \ScanLink230[18] , \ScanLink230[17] , 
        \ScanLink230[16] , \ScanLink230[15] , \ScanLink230[14] , 
        \ScanLink230[13] , \ScanLink230[12] , \ScanLink230[11] , 
        \ScanLink230[10] , \ScanLink230[9] , \ScanLink230[8] , 
        \ScanLink230[7] , \ScanLink230[6] , \ScanLink230[5] , \ScanLink230[4] , 
        \ScanLink230[3] , \ScanLink230[2] , \ScanLink230[1] , \ScanLink230[0] 
        }), .ScanOut({\ScanLink229[31] , \ScanLink229[30] , \ScanLink229[29] , 
        \ScanLink229[28] , \ScanLink229[27] , \ScanLink229[26] , 
        \ScanLink229[25] , \ScanLink229[24] , \ScanLink229[23] , 
        \ScanLink229[22] , \ScanLink229[21] , \ScanLink229[20] , 
        \ScanLink229[19] , \ScanLink229[18] , \ScanLink229[17] , 
        \ScanLink229[16] , \ScanLink229[15] , \ScanLink229[14] , 
        \ScanLink229[13] , \ScanLink229[12] , \ScanLink229[11] , 
        \ScanLink229[10] , \ScanLink229[9] , \ScanLink229[8] , 
        \ScanLink229[7] , \ScanLink229[6] , \ScanLink229[5] , \ScanLink229[4] , 
        \ScanLink229[3] , \ScanLink229[2] , \ScanLink229[1] , \ScanLink229[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_102[31] , 
        \wRegOut_7_102[30] , \wRegOut_7_102[29] , \wRegOut_7_102[28] , 
        \wRegOut_7_102[27] , \wRegOut_7_102[26] , \wRegOut_7_102[25] , 
        \wRegOut_7_102[24] , \wRegOut_7_102[23] , \wRegOut_7_102[22] , 
        \wRegOut_7_102[21] , \wRegOut_7_102[20] , \wRegOut_7_102[19] , 
        \wRegOut_7_102[18] , \wRegOut_7_102[17] , \wRegOut_7_102[16] , 
        \wRegOut_7_102[15] , \wRegOut_7_102[14] , \wRegOut_7_102[13] , 
        \wRegOut_7_102[12] , \wRegOut_7_102[11] , \wRegOut_7_102[10] , 
        \wRegOut_7_102[9] , \wRegOut_7_102[8] , \wRegOut_7_102[7] , 
        \wRegOut_7_102[6] , \wRegOut_7_102[5] , \wRegOut_7_102[4] , 
        \wRegOut_7_102[3] , \wRegOut_7_102[2] , \wRegOut_7_102[1] , 
        \wRegOut_7_102[0] }), .Enable1(\wRegEnTop_7_102[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_102[31] , \wRegInTop_7_102[30] , 
        \wRegInTop_7_102[29] , \wRegInTop_7_102[28] , \wRegInTop_7_102[27] , 
        \wRegInTop_7_102[26] , \wRegInTop_7_102[25] , \wRegInTop_7_102[24] , 
        \wRegInTop_7_102[23] , \wRegInTop_7_102[22] , \wRegInTop_7_102[21] , 
        \wRegInTop_7_102[20] , \wRegInTop_7_102[19] , \wRegInTop_7_102[18] , 
        \wRegInTop_7_102[17] , \wRegInTop_7_102[16] , \wRegInTop_7_102[15] , 
        \wRegInTop_7_102[14] , \wRegInTop_7_102[13] , \wRegInTop_7_102[12] , 
        \wRegInTop_7_102[11] , \wRegInTop_7_102[10] , \wRegInTop_7_102[9] , 
        \wRegInTop_7_102[8] , \wRegInTop_7_102[7] , \wRegInTop_7_102[6] , 
        \wRegInTop_7_102[5] , \wRegInTop_7_102[4] , \wRegInTop_7_102[3] , 
        \wRegInTop_7_102[2] , \wRegInTop_7_102[1] , \wRegInTop_7_102[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_16 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink144[31] , \ScanLink144[30] , \ScanLink144[29] , 
        \ScanLink144[28] , \ScanLink144[27] , \ScanLink144[26] , 
        \ScanLink144[25] , \ScanLink144[24] , \ScanLink144[23] , 
        \ScanLink144[22] , \ScanLink144[21] , \ScanLink144[20] , 
        \ScanLink144[19] , \ScanLink144[18] , \ScanLink144[17] , 
        \ScanLink144[16] , \ScanLink144[15] , \ScanLink144[14] , 
        \ScanLink144[13] , \ScanLink144[12] , \ScanLink144[11] , 
        \ScanLink144[10] , \ScanLink144[9] , \ScanLink144[8] , 
        \ScanLink144[7] , \ScanLink144[6] , \ScanLink144[5] , \ScanLink144[4] , 
        \ScanLink144[3] , \ScanLink144[2] , \ScanLink144[1] , \ScanLink144[0] 
        }), .ScanOut({\ScanLink143[31] , \ScanLink143[30] , \ScanLink143[29] , 
        \ScanLink143[28] , \ScanLink143[27] , \ScanLink143[26] , 
        \ScanLink143[25] , \ScanLink143[24] , \ScanLink143[23] , 
        \ScanLink143[22] , \ScanLink143[21] , \ScanLink143[20] , 
        \ScanLink143[19] , \ScanLink143[18] , \ScanLink143[17] , 
        \ScanLink143[16] , \ScanLink143[15] , \ScanLink143[14] , 
        \ScanLink143[13] , \ScanLink143[12] , \ScanLink143[11] , 
        \ScanLink143[10] , \ScanLink143[9] , \ScanLink143[8] , 
        \ScanLink143[7] , \ScanLink143[6] , \ScanLink143[5] , \ScanLink143[4] , 
        \ScanLink143[3] , \ScanLink143[2] , \ScanLink143[1] , \ScanLink143[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_16[31] , 
        \wRegOut_7_16[30] , \wRegOut_7_16[29] , \wRegOut_7_16[28] , 
        \wRegOut_7_16[27] , \wRegOut_7_16[26] , \wRegOut_7_16[25] , 
        \wRegOut_7_16[24] , \wRegOut_7_16[23] , \wRegOut_7_16[22] , 
        \wRegOut_7_16[21] , \wRegOut_7_16[20] , \wRegOut_7_16[19] , 
        \wRegOut_7_16[18] , \wRegOut_7_16[17] , \wRegOut_7_16[16] , 
        \wRegOut_7_16[15] , \wRegOut_7_16[14] , \wRegOut_7_16[13] , 
        \wRegOut_7_16[12] , \wRegOut_7_16[11] , \wRegOut_7_16[10] , 
        \wRegOut_7_16[9] , \wRegOut_7_16[8] , \wRegOut_7_16[7] , 
        \wRegOut_7_16[6] , \wRegOut_7_16[5] , \wRegOut_7_16[4] , 
        \wRegOut_7_16[3] , \wRegOut_7_16[2] , \wRegOut_7_16[1] , 
        \wRegOut_7_16[0] }), .Enable1(\wRegEnTop_7_16[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_16[31] , \wRegInTop_7_16[30] , \wRegInTop_7_16[29] , 
        \wRegInTop_7_16[28] , \wRegInTop_7_16[27] , \wRegInTop_7_16[26] , 
        \wRegInTop_7_16[25] , \wRegInTop_7_16[24] , \wRegInTop_7_16[23] , 
        \wRegInTop_7_16[22] , \wRegInTop_7_16[21] , \wRegInTop_7_16[20] , 
        \wRegInTop_7_16[19] , \wRegInTop_7_16[18] , \wRegInTop_7_16[17] , 
        \wRegInTop_7_16[16] , \wRegInTop_7_16[15] , \wRegInTop_7_16[14] , 
        \wRegInTop_7_16[13] , \wRegInTop_7_16[12] , \wRegInTop_7_16[11] , 
        \wRegInTop_7_16[10] , \wRegInTop_7_16[9] , \wRegInTop_7_16[8] , 
        \wRegInTop_7_16[7] , \wRegInTop_7_16[6] , \wRegInTop_7_16[5] , 
        \wRegInTop_7_16[4] , \wRegInTop_7_16[3] , \wRegInTop_7_16[2] , 
        \wRegInTop_7_16[1] , \wRegInTop_7_16[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_CtrlReg_WIDTH32 BHCR_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_3[0] ), 
        .Out(\wCtrlOut_2[0] ), .Enable(\wEnable_2[0] ) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_31 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink159[31] , \ScanLink159[30] , \ScanLink159[29] , 
        \ScanLink159[28] , \ScanLink159[27] , \ScanLink159[26] , 
        \ScanLink159[25] , \ScanLink159[24] , \ScanLink159[23] , 
        \ScanLink159[22] , \ScanLink159[21] , \ScanLink159[20] , 
        \ScanLink159[19] , \ScanLink159[18] , \ScanLink159[17] , 
        \ScanLink159[16] , \ScanLink159[15] , \ScanLink159[14] , 
        \ScanLink159[13] , \ScanLink159[12] , \ScanLink159[11] , 
        \ScanLink159[10] , \ScanLink159[9] , \ScanLink159[8] , 
        \ScanLink159[7] , \ScanLink159[6] , \ScanLink159[5] , \ScanLink159[4] , 
        \ScanLink159[3] , \ScanLink159[2] , \ScanLink159[1] , \ScanLink159[0] 
        }), .ScanOut({\ScanLink158[31] , \ScanLink158[30] , \ScanLink158[29] , 
        \ScanLink158[28] , \ScanLink158[27] , \ScanLink158[26] , 
        \ScanLink158[25] , \ScanLink158[24] , \ScanLink158[23] , 
        \ScanLink158[22] , \ScanLink158[21] , \ScanLink158[20] , 
        \ScanLink158[19] , \ScanLink158[18] , \ScanLink158[17] , 
        \ScanLink158[16] , \ScanLink158[15] , \ScanLink158[14] , 
        \ScanLink158[13] , \ScanLink158[12] , \ScanLink158[11] , 
        \ScanLink158[10] , \ScanLink158[9] , \ScanLink158[8] , 
        \ScanLink158[7] , \ScanLink158[6] , \ScanLink158[5] , \ScanLink158[4] , 
        \ScanLink158[3] , \ScanLink158[2] , \ScanLink158[1] , \ScanLink158[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_31[31] , 
        \wRegOut_7_31[30] , \wRegOut_7_31[29] , \wRegOut_7_31[28] , 
        \wRegOut_7_31[27] , \wRegOut_7_31[26] , \wRegOut_7_31[25] , 
        \wRegOut_7_31[24] , \wRegOut_7_31[23] , \wRegOut_7_31[22] , 
        \wRegOut_7_31[21] , \wRegOut_7_31[20] , \wRegOut_7_31[19] , 
        \wRegOut_7_31[18] , \wRegOut_7_31[17] , \wRegOut_7_31[16] , 
        \wRegOut_7_31[15] , \wRegOut_7_31[14] , \wRegOut_7_31[13] , 
        \wRegOut_7_31[12] , \wRegOut_7_31[11] , \wRegOut_7_31[10] , 
        \wRegOut_7_31[9] , \wRegOut_7_31[8] , \wRegOut_7_31[7] , 
        \wRegOut_7_31[6] , \wRegOut_7_31[5] , \wRegOut_7_31[4] , 
        \wRegOut_7_31[3] , \wRegOut_7_31[2] , \wRegOut_7_31[1] , 
        \wRegOut_7_31[0] }), .Enable1(\wRegEnTop_7_31[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_31[31] , \wRegInTop_7_31[30] , \wRegInTop_7_31[29] , 
        \wRegInTop_7_31[28] , \wRegInTop_7_31[27] , \wRegInTop_7_31[26] , 
        \wRegInTop_7_31[25] , \wRegInTop_7_31[24] , \wRegInTop_7_31[23] , 
        \wRegInTop_7_31[22] , \wRegInTop_7_31[21] , \wRegInTop_7_31[20] , 
        \wRegInTop_7_31[19] , \wRegInTop_7_31[18] , \wRegInTop_7_31[17] , 
        \wRegInTop_7_31[16] , \wRegInTop_7_31[15] , \wRegInTop_7_31[14] , 
        \wRegInTop_7_31[13] , \wRegInTop_7_31[12] , \wRegInTop_7_31[11] , 
        \wRegInTop_7_31[10] , \wRegInTop_7_31[9] , \wRegInTop_7_31[8] , 
        \wRegInTop_7_31[7] , \wRegInTop_7_31[6] , \wRegInTop_7_31[5] , 
        \wRegInTop_7_31[4] , \wRegInTop_7_31[3] , \wRegInTop_7_31[2] , 
        \wRegInTop_7_31[1] , \wRegInTop_7_31[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_125 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink253[31] , \ScanLink253[30] , \ScanLink253[29] , 
        \ScanLink253[28] , \ScanLink253[27] , \ScanLink253[26] , 
        \ScanLink253[25] , \ScanLink253[24] , \ScanLink253[23] , 
        \ScanLink253[22] , \ScanLink253[21] , \ScanLink253[20] , 
        \ScanLink253[19] , \ScanLink253[18] , \ScanLink253[17] , 
        \ScanLink253[16] , \ScanLink253[15] , \ScanLink253[14] , 
        \ScanLink253[13] , \ScanLink253[12] , \ScanLink253[11] , 
        \ScanLink253[10] , \ScanLink253[9] , \ScanLink253[8] , 
        \ScanLink253[7] , \ScanLink253[6] , \ScanLink253[5] , \ScanLink253[4] , 
        \ScanLink253[3] , \ScanLink253[2] , \ScanLink253[1] , \ScanLink253[0] 
        }), .ScanOut({\ScanLink252[31] , \ScanLink252[30] , \ScanLink252[29] , 
        \ScanLink252[28] , \ScanLink252[27] , \ScanLink252[26] , 
        \ScanLink252[25] , \ScanLink252[24] , \ScanLink252[23] , 
        \ScanLink252[22] , \ScanLink252[21] , \ScanLink252[20] , 
        \ScanLink252[19] , \ScanLink252[18] , \ScanLink252[17] , 
        \ScanLink252[16] , \ScanLink252[15] , \ScanLink252[14] , 
        \ScanLink252[13] , \ScanLink252[12] , \ScanLink252[11] , 
        \ScanLink252[10] , \ScanLink252[9] , \ScanLink252[8] , 
        \ScanLink252[7] , \ScanLink252[6] , \ScanLink252[5] , \ScanLink252[4] , 
        \ScanLink252[3] , \ScanLink252[2] , \ScanLink252[1] , \ScanLink252[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_125[31] , 
        \wRegOut_7_125[30] , \wRegOut_7_125[29] , \wRegOut_7_125[28] , 
        \wRegOut_7_125[27] , \wRegOut_7_125[26] , \wRegOut_7_125[25] , 
        \wRegOut_7_125[24] , \wRegOut_7_125[23] , \wRegOut_7_125[22] , 
        \wRegOut_7_125[21] , \wRegOut_7_125[20] , \wRegOut_7_125[19] , 
        \wRegOut_7_125[18] , \wRegOut_7_125[17] , \wRegOut_7_125[16] , 
        \wRegOut_7_125[15] , \wRegOut_7_125[14] , \wRegOut_7_125[13] , 
        \wRegOut_7_125[12] , \wRegOut_7_125[11] , \wRegOut_7_125[10] , 
        \wRegOut_7_125[9] , \wRegOut_7_125[8] , \wRegOut_7_125[7] , 
        \wRegOut_7_125[6] , \wRegOut_7_125[5] , \wRegOut_7_125[4] , 
        \wRegOut_7_125[3] , \wRegOut_7_125[2] , \wRegOut_7_125[1] , 
        \wRegOut_7_125[0] }), .Enable1(\wRegEnTop_7_125[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_125[31] , \wRegInTop_7_125[30] , 
        \wRegInTop_7_125[29] , \wRegInTop_7_125[28] , \wRegInTop_7_125[27] , 
        \wRegInTop_7_125[26] , \wRegInTop_7_125[25] , \wRegInTop_7_125[24] , 
        \wRegInTop_7_125[23] , \wRegInTop_7_125[22] , \wRegInTop_7_125[21] , 
        \wRegInTop_7_125[20] , \wRegInTop_7_125[19] , \wRegInTop_7_125[18] , 
        \wRegInTop_7_125[17] , \wRegInTop_7_125[16] , \wRegInTop_7_125[15] , 
        \wRegInTop_7_125[14] , \wRegInTop_7_125[13] , \wRegInTop_7_125[12] , 
        \wRegInTop_7_125[11] , \wRegInTop_7_125[10] , \wRegInTop_7_125[9] , 
        \wRegInTop_7_125[8] , \wRegInTop_7_125[7] , \wRegInTop_7_125[6] , 
        \wRegInTop_7_125[5] , \wRegInTop_7_125[4] , \wRegInTop_7_125[3] , 
        \wRegInTop_7_125[2] , \wRegInTop_7_125[1] , \wRegInTop_7_125[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_63 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink191[31] , \ScanLink191[30] , \ScanLink191[29] , 
        \ScanLink191[28] , \ScanLink191[27] , \ScanLink191[26] , 
        \ScanLink191[25] , \ScanLink191[24] , \ScanLink191[23] , 
        \ScanLink191[22] , \ScanLink191[21] , \ScanLink191[20] , 
        \ScanLink191[19] , \ScanLink191[18] , \ScanLink191[17] , 
        \ScanLink191[16] , \ScanLink191[15] , \ScanLink191[14] , 
        \ScanLink191[13] , \ScanLink191[12] , \ScanLink191[11] , 
        \ScanLink191[10] , \ScanLink191[9] , \ScanLink191[8] , 
        \ScanLink191[7] , \ScanLink191[6] , \ScanLink191[5] , \ScanLink191[4] , 
        \ScanLink191[3] , \ScanLink191[2] , \ScanLink191[1] , \ScanLink191[0] 
        }), .ScanOut({\ScanLink190[31] , \ScanLink190[30] , \ScanLink190[29] , 
        \ScanLink190[28] , \ScanLink190[27] , \ScanLink190[26] , 
        \ScanLink190[25] , \ScanLink190[24] , \ScanLink190[23] , 
        \ScanLink190[22] , \ScanLink190[21] , \ScanLink190[20] , 
        \ScanLink190[19] , \ScanLink190[18] , \ScanLink190[17] , 
        \ScanLink190[16] , \ScanLink190[15] , \ScanLink190[14] , 
        \ScanLink190[13] , \ScanLink190[12] , \ScanLink190[11] , 
        \ScanLink190[10] , \ScanLink190[9] , \ScanLink190[8] , 
        \ScanLink190[7] , \ScanLink190[6] , \ScanLink190[5] , \ScanLink190[4] , 
        \ScanLink190[3] , \ScanLink190[2] , \ScanLink190[1] , \ScanLink190[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_63[31] , 
        \wRegOut_7_63[30] , \wRegOut_7_63[29] , \wRegOut_7_63[28] , 
        \wRegOut_7_63[27] , \wRegOut_7_63[26] , \wRegOut_7_63[25] , 
        \wRegOut_7_63[24] , \wRegOut_7_63[23] , \wRegOut_7_63[22] , 
        \wRegOut_7_63[21] , \wRegOut_7_63[20] , \wRegOut_7_63[19] , 
        \wRegOut_7_63[18] , \wRegOut_7_63[17] , \wRegOut_7_63[16] , 
        \wRegOut_7_63[15] , \wRegOut_7_63[14] , \wRegOut_7_63[13] , 
        \wRegOut_7_63[12] , \wRegOut_7_63[11] , \wRegOut_7_63[10] , 
        \wRegOut_7_63[9] , \wRegOut_7_63[8] , \wRegOut_7_63[7] , 
        \wRegOut_7_63[6] , \wRegOut_7_63[5] , \wRegOut_7_63[4] , 
        \wRegOut_7_63[3] , \wRegOut_7_63[2] , \wRegOut_7_63[1] , 
        \wRegOut_7_63[0] }), .Enable1(\wRegEnTop_7_63[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_63[31] , \wRegInTop_7_63[30] , \wRegInTop_7_63[29] , 
        \wRegInTop_7_63[28] , \wRegInTop_7_63[27] , \wRegInTop_7_63[26] , 
        \wRegInTop_7_63[25] , \wRegInTop_7_63[24] , \wRegInTop_7_63[23] , 
        \wRegInTop_7_63[22] , \wRegInTop_7_63[21] , \wRegInTop_7_63[20] , 
        \wRegInTop_7_63[19] , \wRegInTop_7_63[18] , \wRegInTop_7_63[17] , 
        \wRegInTop_7_63[16] , \wRegInTop_7_63[15] , \wRegInTop_7_63[14] , 
        \wRegInTop_7_63[13] , \wRegInTop_7_63[12] , \wRegInTop_7_63[11] , 
        \wRegInTop_7_63[10] , \wRegInTop_7_63[9] , \wRegInTop_7_63[8] , 
        \wRegInTop_7_63[7] , \wRegInTop_7_63[6] , \wRegInTop_7_63[5] , 
        \wRegInTop_7_63[4] , \wRegInTop_7_63[3] , \wRegInTop_7_63[2] , 
        \wRegInTop_7_63[1] , \wRegInTop_7_63[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_86 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink214[31] , \ScanLink214[30] , \ScanLink214[29] , 
        \ScanLink214[28] , \ScanLink214[27] , \ScanLink214[26] , 
        \ScanLink214[25] , \ScanLink214[24] , \ScanLink214[23] , 
        \ScanLink214[22] , \ScanLink214[21] , \ScanLink214[20] , 
        \ScanLink214[19] , \ScanLink214[18] , \ScanLink214[17] , 
        \ScanLink214[16] , \ScanLink214[15] , \ScanLink214[14] , 
        \ScanLink214[13] , \ScanLink214[12] , \ScanLink214[11] , 
        \ScanLink214[10] , \ScanLink214[9] , \ScanLink214[8] , 
        \ScanLink214[7] , \ScanLink214[6] , \ScanLink214[5] , \ScanLink214[4] , 
        \ScanLink214[3] , \ScanLink214[2] , \ScanLink214[1] , \ScanLink214[0] 
        }), .ScanOut({\ScanLink213[31] , \ScanLink213[30] , \ScanLink213[29] , 
        \ScanLink213[28] , \ScanLink213[27] , \ScanLink213[26] , 
        \ScanLink213[25] , \ScanLink213[24] , \ScanLink213[23] , 
        \ScanLink213[22] , \ScanLink213[21] , \ScanLink213[20] , 
        \ScanLink213[19] , \ScanLink213[18] , \ScanLink213[17] , 
        \ScanLink213[16] , \ScanLink213[15] , \ScanLink213[14] , 
        \ScanLink213[13] , \ScanLink213[12] , \ScanLink213[11] , 
        \ScanLink213[10] , \ScanLink213[9] , \ScanLink213[8] , 
        \ScanLink213[7] , \ScanLink213[6] , \ScanLink213[5] , \ScanLink213[4] , 
        \ScanLink213[3] , \ScanLink213[2] , \ScanLink213[1] , \ScanLink213[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_86[31] , 
        \wRegOut_7_86[30] , \wRegOut_7_86[29] , \wRegOut_7_86[28] , 
        \wRegOut_7_86[27] , \wRegOut_7_86[26] , \wRegOut_7_86[25] , 
        \wRegOut_7_86[24] , \wRegOut_7_86[23] , \wRegOut_7_86[22] , 
        \wRegOut_7_86[21] , \wRegOut_7_86[20] , \wRegOut_7_86[19] , 
        \wRegOut_7_86[18] , \wRegOut_7_86[17] , \wRegOut_7_86[16] , 
        \wRegOut_7_86[15] , \wRegOut_7_86[14] , \wRegOut_7_86[13] , 
        \wRegOut_7_86[12] , \wRegOut_7_86[11] , \wRegOut_7_86[10] , 
        \wRegOut_7_86[9] , \wRegOut_7_86[8] , \wRegOut_7_86[7] , 
        \wRegOut_7_86[6] , \wRegOut_7_86[5] , \wRegOut_7_86[4] , 
        \wRegOut_7_86[3] , \wRegOut_7_86[2] , \wRegOut_7_86[1] , 
        \wRegOut_7_86[0] }), .Enable1(\wRegEnTop_7_86[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_86[31] , \wRegInTop_7_86[30] , \wRegInTop_7_86[29] , 
        \wRegInTop_7_86[28] , \wRegInTop_7_86[27] , \wRegInTop_7_86[26] , 
        \wRegInTop_7_86[25] , \wRegInTop_7_86[24] , \wRegInTop_7_86[23] , 
        \wRegInTop_7_86[22] , \wRegInTop_7_86[21] , \wRegInTop_7_86[20] , 
        \wRegInTop_7_86[19] , \wRegInTop_7_86[18] , \wRegInTop_7_86[17] , 
        \wRegInTop_7_86[16] , \wRegInTop_7_86[15] , \wRegInTop_7_86[14] , 
        \wRegInTop_7_86[13] , \wRegInTop_7_86[12] , \wRegInTop_7_86[11] , 
        \wRegInTop_7_86[10] , \wRegInTop_7_86[9] , \wRegInTop_7_86[8] , 
        \wRegInTop_7_86[7] , \wRegInTop_7_86[6] , \wRegInTop_7_86[5] , 
        \wRegInTop_7_86[4] , \wRegInTop_7_86[3] , \wRegInTop_7_86[2] , 
        \wRegInTop_7_86[1] , \wRegInTop_7_86[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_0[0] ), .P_In({\wRegOut_6_0[31] , 
        \wRegOut_6_0[30] , \wRegOut_6_0[29] , \wRegOut_6_0[28] , 
        \wRegOut_6_0[27] , \wRegOut_6_0[26] , \wRegOut_6_0[25] , 
        \wRegOut_6_0[24] , \wRegOut_6_0[23] , \wRegOut_6_0[22] , 
        \wRegOut_6_0[21] , \wRegOut_6_0[20] , \wRegOut_6_0[19] , 
        \wRegOut_6_0[18] , \wRegOut_6_0[17] , \wRegOut_6_0[16] , 
        \wRegOut_6_0[15] , \wRegOut_6_0[14] , \wRegOut_6_0[13] , 
        \wRegOut_6_0[12] , \wRegOut_6_0[11] , \wRegOut_6_0[10] , 
        \wRegOut_6_0[9] , \wRegOut_6_0[8] , \wRegOut_6_0[7] , \wRegOut_6_0[6] , 
        \wRegOut_6_0[5] , \wRegOut_6_0[4] , \wRegOut_6_0[3] , \wRegOut_6_0[2] , 
        \wRegOut_6_0[1] , \wRegOut_6_0[0] }), .P_Out({\wRegInBot_6_0[31] , 
        \wRegInBot_6_0[30] , \wRegInBot_6_0[29] , \wRegInBot_6_0[28] , 
        \wRegInBot_6_0[27] , \wRegInBot_6_0[26] , \wRegInBot_6_0[25] , 
        \wRegInBot_6_0[24] , \wRegInBot_6_0[23] , \wRegInBot_6_0[22] , 
        \wRegInBot_6_0[21] , \wRegInBot_6_0[20] , \wRegInBot_6_0[19] , 
        \wRegInBot_6_0[18] , \wRegInBot_6_0[17] , \wRegInBot_6_0[16] , 
        \wRegInBot_6_0[15] , \wRegInBot_6_0[14] , \wRegInBot_6_0[13] , 
        \wRegInBot_6_0[12] , \wRegInBot_6_0[11] , \wRegInBot_6_0[10] , 
        \wRegInBot_6_0[9] , \wRegInBot_6_0[8] , \wRegInBot_6_0[7] , 
        \wRegInBot_6_0[6] , \wRegInBot_6_0[5] , \wRegInBot_6_0[4] , 
        \wRegInBot_6_0[3] , \wRegInBot_6_0[2] , \wRegInBot_6_0[1] , 
        \wRegInBot_6_0[0] }), .L_WR(\wRegEnTop_7_0[0] ), .L_In({
        \wRegOut_7_0[31] , \wRegOut_7_0[30] , \wRegOut_7_0[29] , 
        \wRegOut_7_0[28] , \wRegOut_7_0[27] , \wRegOut_7_0[26] , 
        \wRegOut_7_0[25] , \wRegOut_7_0[24] , \wRegOut_7_0[23] , 
        \wRegOut_7_0[22] , \wRegOut_7_0[21] , \wRegOut_7_0[20] , 
        \wRegOut_7_0[19] , \wRegOut_7_0[18] , \wRegOut_7_0[17] , 
        \wRegOut_7_0[16] , \wRegOut_7_0[15] , \wRegOut_7_0[14] , 
        \wRegOut_7_0[13] , \wRegOut_7_0[12] , \wRegOut_7_0[11] , 
        \wRegOut_7_0[10] , \wRegOut_7_0[9] , \wRegOut_7_0[8] , 
        \wRegOut_7_0[7] , \wRegOut_7_0[6] , \wRegOut_7_0[5] , \wRegOut_7_0[4] , 
        \wRegOut_7_0[3] , \wRegOut_7_0[2] , \wRegOut_7_0[1] , \wRegOut_7_0[0] 
        }), .L_Out({\wRegInTop_7_0[31] , \wRegInTop_7_0[30] , 
        \wRegInTop_7_0[29] , \wRegInTop_7_0[28] , \wRegInTop_7_0[27] , 
        \wRegInTop_7_0[26] , \wRegInTop_7_0[25] , \wRegInTop_7_0[24] , 
        \wRegInTop_7_0[23] , \wRegInTop_7_0[22] , \wRegInTop_7_0[21] , 
        \wRegInTop_7_0[20] , \wRegInTop_7_0[19] , \wRegInTop_7_0[18] , 
        \wRegInTop_7_0[17] , \wRegInTop_7_0[16] , \wRegInTop_7_0[15] , 
        \wRegInTop_7_0[14] , \wRegInTop_7_0[13] , \wRegInTop_7_0[12] , 
        \wRegInTop_7_0[11] , \wRegInTop_7_0[10] , \wRegInTop_7_0[9] , 
        \wRegInTop_7_0[8] , \wRegInTop_7_0[7] , \wRegInTop_7_0[6] , 
        \wRegInTop_7_0[5] , \wRegInTop_7_0[4] , \wRegInTop_7_0[3] , 
        \wRegInTop_7_0[2] , \wRegInTop_7_0[1] , \wRegInTop_7_0[0] }), .R_WR(
        \wRegEnTop_7_1[0] ), .R_In({\wRegOut_7_1[31] , \wRegOut_7_1[30] , 
        \wRegOut_7_1[29] , \wRegOut_7_1[28] , \wRegOut_7_1[27] , 
        \wRegOut_7_1[26] , \wRegOut_7_1[25] , \wRegOut_7_1[24] , 
        \wRegOut_7_1[23] , \wRegOut_7_1[22] , \wRegOut_7_1[21] , 
        \wRegOut_7_1[20] , \wRegOut_7_1[19] , \wRegOut_7_1[18] , 
        \wRegOut_7_1[17] , \wRegOut_7_1[16] , \wRegOut_7_1[15] , 
        \wRegOut_7_1[14] , \wRegOut_7_1[13] , \wRegOut_7_1[12] , 
        \wRegOut_7_1[11] , \wRegOut_7_1[10] , \wRegOut_7_1[9] , 
        \wRegOut_7_1[8] , \wRegOut_7_1[7] , \wRegOut_7_1[6] , \wRegOut_7_1[5] , 
        \wRegOut_7_1[4] , \wRegOut_7_1[3] , \wRegOut_7_1[2] , \wRegOut_7_1[1] , 
        \wRegOut_7_1[0] }), .R_Out({\wRegInTop_7_1[31] , \wRegInTop_7_1[30] , 
        \wRegInTop_7_1[29] , \wRegInTop_7_1[28] , \wRegInTop_7_1[27] , 
        \wRegInTop_7_1[26] , \wRegInTop_7_1[25] , \wRegInTop_7_1[24] , 
        \wRegInTop_7_1[23] , \wRegInTop_7_1[22] , \wRegInTop_7_1[21] , 
        \wRegInTop_7_1[20] , \wRegInTop_7_1[19] , \wRegInTop_7_1[18] , 
        \wRegInTop_7_1[17] , \wRegInTop_7_1[16] , \wRegInTop_7_1[15] , 
        \wRegInTop_7_1[14] , \wRegInTop_7_1[13] , \wRegInTop_7_1[12] , 
        \wRegInTop_7_1[11] , \wRegInTop_7_1[10] , \wRegInTop_7_1[9] , 
        \wRegInTop_7_1[8] , \wRegInTop_7_1[7] , \wRegInTop_7_1[6] , 
        \wRegInTop_7_1[5] , \wRegInTop_7_1[4] , \wRegInTop_7_1[3] , 
        \wRegInTop_7_1[2] , \wRegInTop_7_1[1] , \wRegInTop_7_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_119 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink247[31] , \ScanLink247[30] , \ScanLink247[29] , 
        \ScanLink247[28] , \ScanLink247[27] , \ScanLink247[26] , 
        \ScanLink247[25] , \ScanLink247[24] , \ScanLink247[23] , 
        \ScanLink247[22] , \ScanLink247[21] , \ScanLink247[20] , 
        \ScanLink247[19] , \ScanLink247[18] , \ScanLink247[17] , 
        \ScanLink247[16] , \ScanLink247[15] , \ScanLink247[14] , 
        \ScanLink247[13] , \ScanLink247[12] , \ScanLink247[11] , 
        \ScanLink247[10] , \ScanLink247[9] , \ScanLink247[8] , 
        \ScanLink247[7] , \ScanLink247[6] , \ScanLink247[5] , \ScanLink247[4] , 
        \ScanLink247[3] , \ScanLink247[2] , \ScanLink247[1] , \ScanLink247[0] 
        }), .ScanOut({\ScanLink246[31] , \ScanLink246[30] , \ScanLink246[29] , 
        \ScanLink246[28] , \ScanLink246[27] , \ScanLink246[26] , 
        \ScanLink246[25] , \ScanLink246[24] , \ScanLink246[23] , 
        \ScanLink246[22] , \ScanLink246[21] , \ScanLink246[20] , 
        \ScanLink246[19] , \ScanLink246[18] , \ScanLink246[17] , 
        \ScanLink246[16] , \ScanLink246[15] , \ScanLink246[14] , 
        \ScanLink246[13] , \ScanLink246[12] , \ScanLink246[11] , 
        \ScanLink246[10] , \ScanLink246[9] , \ScanLink246[8] , 
        \ScanLink246[7] , \ScanLink246[6] , \ScanLink246[5] , \ScanLink246[4] , 
        \ScanLink246[3] , \ScanLink246[2] , \ScanLink246[1] , \ScanLink246[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_119[31] , 
        \wRegOut_7_119[30] , \wRegOut_7_119[29] , \wRegOut_7_119[28] , 
        \wRegOut_7_119[27] , \wRegOut_7_119[26] , \wRegOut_7_119[25] , 
        \wRegOut_7_119[24] , \wRegOut_7_119[23] , \wRegOut_7_119[22] , 
        \wRegOut_7_119[21] , \wRegOut_7_119[20] , \wRegOut_7_119[19] , 
        \wRegOut_7_119[18] , \wRegOut_7_119[17] , \wRegOut_7_119[16] , 
        \wRegOut_7_119[15] , \wRegOut_7_119[14] , \wRegOut_7_119[13] , 
        \wRegOut_7_119[12] , \wRegOut_7_119[11] , \wRegOut_7_119[10] , 
        \wRegOut_7_119[9] , \wRegOut_7_119[8] , \wRegOut_7_119[7] , 
        \wRegOut_7_119[6] , \wRegOut_7_119[5] , \wRegOut_7_119[4] , 
        \wRegOut_7_119[3] , \wRegOut_7_119[2] , \wRegOut_7_119[1] , 
        \wRegOut_7_119[0] }), .Enable1(\wRegEnTop_7_119[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_119[31] , \wRegInTop_7_119[30] , 
        \wRegInTop_7_119[29] , \wRegInTop_7_119[28] , \wRegInTop_7_119[27] , 
        \wRegInTop_7_119[26] , \wRegInTop_7_119[25] , \wRegInTop_7_119[24] , 
        \wRegInTop_7_119[23] , \wRegInTop_7_119[22] , \wRegInTop_7_119[21] , 
        \wRegInTop_7_119[20] , \wRegInTop_7_119[19] , \wRegInTop_7_119[18] , 
        \wRegInTop_7_119[17] , \wRegInTop_7_119[16] , \wRegInTop_7_119[15] , 
        \wRegInTop_7_119[14] , \wRegInTop_7_119[13] , \wRegInTop_7_119[12] , 
        \wRegInTop_7_119[11] , \wRegInTop_7_119[10] , \wRegInTop_7_119[9] , 
        \wRegInTop_7_119[8] , \wRegInTop_7_119[7] , \wRegInTop_7_119[6] , 
        \wRegInTop_7_119[5] , \wRegInTop_7_119[4] , \wRegInTop_7_119[3] , 
        \wRegInTop_7_119[2] , \wRegInTop_7_119[1] , \wRegInTop_7_119[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_6[0] ), .P_In({\wRegOut_3_6[31] , 
        \wRegOut_3_6[30] , \wRegOut_3_6[29] , \wRegOut_3_6[28] , 
        \wRegOut_3_6[27] , \wRegOut_3_6[26] , \wRegOut_3_6[25] , 
        \wRegOut_3_6[24] , \wRegOut_3_6[23] , \wRegOut_3_6[22] , 
        \wRegOut_3_6[21] , \wRegOut_3_6[20] , \wRegOut_3_6[19] , 
        \wRegOut_3_6[18] , \wRegOut_3_6[17] , \wRegOut_3_6[16] , 
        \wRegOut_3_6[15] , \wRegOut_3_6[14] , \wRegOut_3_6[13] , 
        \wRegOut_3_6[12] , \wRegOut_3_6[11] , \wRegOut_3_6[10] , 
        \wRegOut_3_6[9] , \wRegOut_3_6[8] , \wRegOut_3_6[7] , \wRegOut_3_6[6] , 
        \wRegOut_3_6[5] , \wRegOut_3_6[4] , \wRegOut_3_6[3] , \wRegOut_3_6[2] , 
        \wRegOut_3_6[1] , \wRegOut_3_6[0] }), .P_Out({\wRegInBot_3_6[31] , 
        \wRegInBot_3_6[30] , \wRegInBot_3_6[29] , \wRegInBot_3_6[28] , 
        \wRegInBot_3_6[27] , \wRegInBot_3_6[26] , \wRegInBot_3_6[25] , 
        \wRegInBot_3_6[24] , \wRegInBot_3_6[23] , \wRegInBot_3_6[22] , 
        \wRegInBot_3_6[21] , \wRegInBot_3_6[20] , \wRegInBot_3_6[19] , 
        \wRegInBot_3_6[18] , \wRegInBot_3_6[17] , \wRegInBot_3_6[16] , 
        \wRegInBot_3_6[15] , \wRegInBot_3_6[14] , \wRegInBot_3_6[13] , 
        \wRegInBot_3_6[12] , \wRegInBot_3_6[11] , \wRegInBot_3_6[10] , 
        \wRegInBot_3_6[9] , \wRegInBot_3_6[8] , \wRegInBot_3_6[7] , 
        \wRegInBot_3_6[6] , \wRegInBot_3_6[5] , \wRegInBot_3_6[4] , 
        \wRegInBot_3_6[3] , \wRegInBot_3_6[2] , \wRegInBot_3_6[1] , 
        \wRegInBot_3_6[0] }), .L_WR(\wRegEnTop_4_12[0] ), .L_In({
        \wRegOut_4_12[31] , \wRegOut_4_12[30] , \wRegOut_4_12[29] , 
        \wRegOut_4_12[28] , \wRegOut_4_12[27] , \wRegOut_4_12[26] , 
        \wRegOut_4_12[25] , \wRegOut_4_12[24] , \wRegOut_4_12[23] , 
        \wRegOut_4_12[22] , \wRegOut_4_12[21] , \wRegOut_4_12[20] , 
        \wRegOut_4_12[19] , \wRegOut_4_12[18] , \wRegOut_4_12[17] , 
        \wRegOut_4_12[16] , \wRegOut_4_12[15] , \wRegOut_4_12[14] , 
        \wRegOut_4_12[13] , \wRegOut_4_12[12] , \wRegOut_4_12[11] , 
        \wRegOut_4_12[10] , \wRegOut_4_12[9] , \wRegOut_4_12[8] , 
        \wRegOut_4_12[7] , \wRegOut_4_12[6] , \wRegOut_4_12[5] , 
        \wRegOut_4_12[4] , \wRegOut_4_12[3] , \wRegOut_4_12[2] , 
        \wRegOut_4_12[1] , \wRegOut_4_12[0] }), .L_Out({\wRegInTop_4_12[31] , 
        \wRegInTop_4_12[30] , \wRegInTop_4_12[29] , \wRegInTop_4_12[28] , 
        \wRegInTop_4_12[27] , \wRegInTop_4_12[26] , \wRegInTop_4_12[25] , 
        \wRegInTop_4_12[24] , \wRegInTop_4_12[23] , \wRegInTop_4_12[22] , 
        \wRegInTop_4_12[21] , \wRegInTop_4_12[20] , \wRegInTop_4_12[19] , 
        \wRegInTop_4_12[18] , \wRegInTop_4_12[17] , \wRegInTop_4_12[16] , 
        \wRegInTop_4_12[15] , \wRegInTop_4_12[14] , \wRegInTop_4_12[13] , 
        \wRegInTop_4_12[12] , \wRegInTop_4_12[11] , \wRegInTop_4_12[10] , 
        \wRegInTop_4_12[9] , \wRegInTop_4_12[8] , \wRegInTop_4_12[7] , 
        \wRegInTop_4_12[6] , \wRegInTop_4_12[5] , \wRegInTop_4_12[4] , 
        \wRegInTop_4_12[3] , \wRegInTop_4_12[2] , \wRegInTop_4_12[1] , 
        \wRegInTop_4_12[0] }), .R_WR(\wRegEnTop_4_13[0] ), .R_In({
        \wRegOut_4_13[31] , \wRegOut_4_13[30] , \wRegOut_4_13[29] , 
        \wRegOut_4_13[28] , \wRegOut_4_13[27] , \wRegOut_4_13[26] , 
        \wRegOut_4_13[25] , \wRegOut_4_13[24] , \wRegOut_4_13[23] , 
        \wRegOut_4_13[22] , \wRegOut_4_13[21] , \wRegOut_4_13[20] , 
        \wRegOut_4_13[19] , \wRegOut_4_13[18] , \wRegOut_4_13[17] , 
        \wRegOut_4_13[16] , \wRegOut_4_13[15] , \wRegOut_4_13[14] , 
        \wRegOut_4_13[13] , \wRegOut_4_13[12] , \wRegOut_4_13[11] , 
        \wRegOut_4_13[10] , \wRegOut_4_13[9] , \wRegOut_4_13[8] , 
        \wRegOut_4_13[7] , \wRegOut_4_13[6] , \wRegOut_4_13[5] , 
        \wRegOut_4_13[4] , \wRegOut_4_13[3] , \wRegOut_4_13[2] , 
        \wRegOut_4_13[1] , \wRegOut_4_13[0] }), .R_Out({\wRegInTop_4_13[31] , 
        \wRegInTop_4_13[30] , \wRegInTop_4_13[29] , \wRegInTop_4_13[28] , 
        \wRegInTop_4_13[27] , \wRegInTop_4_13[26] , \wRegInTop_4_13[25] , 
        \wRegInTop_4_13[24] , \wRegInTop_4_13[23] , \wRegInTop_4_13[22] , 
        \wRegInTop_4_13[21] , \wRegInTop_4_13[20] , \wRegInTop_4_13[19] , 
        \wRegInTop_4_13[18] , \wRegInTop_4_13[17] , \wRegInTop_4_13[16] , 
        \wRegInTop_4_13[15] , \wRegInTop_4_13[14] , \wRegInTop_4_13[13] , 
        \wRegInTop_4_13[12] , \wRegInTop_4_13[11] , \wRegInTop_4_13[10] , 
        \wRegInTop_4_13[9] , \wRegInTop_4_13[8] , \wRegInTop_4_13[7] , 
        \wRegInTop_4_13[6] , \wRegInTop_4_13[5] , \wRegInTop_4_13[4] , 
        \wRegInTop_4_13[3] , \wRegInTop_4_13[2] , \wRegInTop_4_13[1] , 
        \wRegInTop_4_13[0] }) );
    BHeap_Node_WIDTH32 BHN_4_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_15[0] ), .P_In({\wRegOut_4_15[31] , 
        \wRegOut_4_15[30] , \wRegOut_4_15[29] , \wRegOut_4_15[28] , 
        \wRegOut_4_15[27] , \wRegOut_4_15[26] , \wRegOut_4_15[25] , 
        \wRegOut_4_15[24] , \wRegOut_4_15[23] , \wRegOut_4_15[22] , 
        \wRegOut_4_15[21] , \wRegOut_4_15[20] , \wRegOut_4_15[19] , 
        \wRegOut_4_15[18] , \wRegOut_4_15[17] , \wRegOut_4_15[16] , 
        \wRegOut_4_15[15] , \wRegOut_4_15[14] , \wRegOut_4_15[13] , 
        \wRegOut_4_15[12] , \wRegOut_4_15[11] , \wRegOut_4_15[10] , 
        \wRegOut_4_15[9] , \wRegOut_4_15[8] , \wRegOut_4_15[7] , 
        \wRegOut_4_15[6] , \wRegOut_4_15[5] , \wRegOut_4_15[4] , 
        \wRegOut_4_15[3] , \wRegOut_4_15[2] , \wRegOut_4_15[1] , 
        \wRegOut_4_15[0] }), .P_Out({\wRegInBot_4_15[31] , 
        \wRegInBot_4_15[30] , \wRegInBot_4_15[29] , \wRegInBot_4_15[28] , 
        \wRegInBot_4_15[27] , \wRegInBot_4_15[26] , \wRegInBot_4_15[25] , 
        \wRegInBot_4_15[24] , \wRegInBot_4_15[23] , \wRegInBot_4_15[22] , 
        \wRegInBot_4_15[21] , \wRegInBot_4_15[20] , \wRegInBot_4_15[19] , 
        \wRegInBot_4_15[18] , \wRegInBot_4_15[17] , \wRegInBot_4_15[16] , 
        \wRegInBot_4_15[15] , \wRegInBot_4_15[14] , \wRegInBot_4_15[13] , 
        \wRegInBot_4_15[12] , \wRegInBot_4_15[11] , \wRegInBot_4_15[10] , 
        \wRegInBot_4_15[9] , \wRegInBot_4_15[8] , \wRegInBot_4_15[7] , 
        \wRegInBot_4_15[6] , \wRegInBot_4_15[5] , \wRegInBot_4_15[4] , 
        \wRegInBot_4_15[3] , \wRegInBot_4_15[2] , \wRegInBot_4_15[1] , 
        \wRegInBot_4_15[0] }), .L_WR(\wRegEnTop_5_30[0] ), .L_In({
        \wRegOut_5_30[31] , \wRegOut_5_30[30] , \wRegOut_5_30[29] , 
        \wRegOut_5_30[28] , \wRegOut_5_30[27] , \wRegOut_5_30[26] , 
        \wRegOut_5_30[25] , \wRegOut_5_30[24] , \wRegOut_5_30[23] , 
        \wRegOut_5_30[22] , \wRegOut_5_30[21] , \wRegOut_5_30[20] , 
        \wRegOut_5_30[19] , \wRegOut_5_30[18] , \wRegOut_5_30[17] , 
        \wRegOut_5_30[16] , \wRegOut_5_30[15] , \wRegOut_5_30[14] , 
        \wRegOut_5_30[13] , \wRegOut_5_30[12] , \wRegOut_5_30[11] , 
        \wRegOut_5_30[10] , \wRegOut_5_30[9] , \wRegOut_5_30[8] , 
        \wRegOut_5_30[7] , \wRegOut_5_30[6] , \wRegOut_5_30[5] , 
        \wRegOut_5_30[4] , \wRegOut_5_30[3] , \wRegOut_5_30[2] , 
        \wRegOut_5_30[1] , \wRegOut_5_30[0] }), .L_Out({\wRegInTop_5_30[31] , 
        \wRegInTop_5_30[30] , \wRegInTop_5_30[29] , \wRegInTop_5_30[28] , 
        \wRegInTop_5_30[27] , \wRegInTop_5_30[26] , \wRegInTop_5_30[25] , 
        \wRegInTop_5_30[24] , \wRegInTop_5_30[23] , \wRegInTop_5_30[22] , 
        \wRegInTop_5_30[21] , \wRegInTop_5_30[20] , \wRegInTop_5_30[19] , 
        \wRegInTop_5_30[18] , \wRegInTop_5_30[17] , \wRegInTop_5_30[16] , 
        \wRegInTop_5_30[15] , \wRegInTop_5_30[14] , \wRegInTop_5_30[13] , 
        \wRegInTop_5_30[12] , \wRegInTop_5_30[11] , \wRegInTop_5_30[10] , 
        \wRegInTop_5_30[9] , \wRegInTop_5_30[8] , \wRegInTop_5_30[7] , 
        \wRegInTop_5_30[6] , \wRegInTop_5_30[5] , \wRegInTop_5_30[4] , 
        \wRegInTop_5_30[3] , \wRegInTop_5_30[2] , \wRegInTop_5_30[1] , 
        \wRegInTop_5_30[0] }), .R_WR(\wRegEnTop_5_31[0] ), .R_In({
        \wRegOut_5_31[31] , \wRegOut_5_31[30] , \wRegOut_5_31[29] , 
        \wRegOut_5_31[28] , \wRegOut_5_31[27] , \wRegOut_5_31[26] , 
        \wRegOut_5_31[25] , \wRegOut_5_31[24] , \wRegOut_5_31[23] , 
        \wRegOut_5_31[22] , \wRegOut_5_31[21] , \wRegOut_5_31[20] , 
        \wRegOut_5_31[19] , \wRegOut_5_31[18] , \wRegOut_5_31[17] , 
        \wRegOut_5_31[16] , \wRegOut_5_31[15] , \wRegOut_5_31[14] , 
        \wRegOut_5_31[13] , \wRegOut_5_31[12] , \wRegOut_5_31[11] , 
        \wRegOut_5_31[10] , \wRegOut_5_31[9] , \wRegOut_5_31[8] , 
        \wRegOut_5_31[7] , \wRegOut_5_31[6] , \wRegOut_5_31[5] , 
        \wRegOut_5_31[4] , \wRegOut_5_31[3] , \wRegOut_5_31[2] , 
        \wRegOut_5_31[1] , \wRegOut_5_31[0] }), .R_Out({\wRegInTop_5_31[31] , 
        \wRegInTop_5_31[30] , \wRegInTop_5_31[29] , \wRegInTop_5_31[28] , 
        \wRegInTop_5_31[27] , \wRegInTop_5_31[26] , \wRegInTop_5_31[25] , 
        \wRegInTop_5_31[24] , \wRegInTop_5_31[23] , \wRegInTop_5_31[22] , 
        \wRegInTop_5_31[21] , \wRegInTop_5_31[20] , \wRegInTop_5_31[19] , 
        \wRegInTop_5_31[18] , \wRegInTop_5_31[17] , \wRegInTop_5_31[16] , 
        \wRegInTop_5_31[15] , \wRegInTop_5_31[14] , \wRegInTop_5_31[13] , 
        \wRegInTop_5_31[12] , \wRegInTop_5_31[11] , \wRegInTop_5_31[10] , 
        \wRegInTop_5_31[9] , \wRegInTop_5_31[8] , \wRegInTop_5_31[7] , 
        \wRegInTop_5_31[6] , \wRegInTop_5_31[5] , \wRegInTop_5_31[4] , 
        \wRegInTop_5_31[3] , \wRegInTop_5_31[2] , \wRegInTop_5_31[1] , 
        \wRegInTop_5_31[0] }) );
    BHeap_Node_WIDTH32 BHN_6_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_51[0] ), .P_In({\wRegOut_6_51[31] , 
        \wRegOut_6_51[30] , \wRegOut_6_51[29] , \wRegOut_6_51[28] , 
        \wRegOut_6_51[27] , \wRegOut_6_51[26] , \wRegOut_6_51[25] , 
        \wRegOut_6_51[24] , \wRegOut_6_51[23] , \wRegOut_6_51[22] , 
        \wRegOut_6_51[21] , \wRegOut_6_51[20] , \wRegOut_6_51[19] , 
        \wRegOut_6_51[18] , \wRegOut_6_51[17] , \wRegOut_6_51[16] , 
        \wRegOut_6_51[15] , \wRegOut_6_51[14] , \wRegOut_6_51[13] , 
        \wRegOut_6_51[12] , \wRegOut_6_51[11] , \wRegOut_6_51[10] , 
        \wRegOut_6_51[9] , \wRegOut_6_51[8] , \wRegOut_6_51[7] , 
        \wRegOut_6_51[6] , \wRegOut_6_51[5] , \wRegOut_6_51[4] , 
        \wRegOut_6_51[3] , \wRegOut_6_51[2] , \wRegOut_6_51[1] , 
        \wRegOut_6_51[0] }), .P_Out({\wRegInBot_6_51[31] , 
        \wRegInBot_6_51[30] , \wRegInBot_6_51[29] , \wRegInBot_6_51[28] , 
        \wRegInBot_6_51[27] , \wRegInBot_6_51[26] , \wRegInBot_6_51[25] , 
        \wRegInBot_6_51[24] , \wRegInBot_6_51[23] , \wRegInBot_6_51[22] , 
        \wRegInBot_6_51[21] , \wRegInBot_6_51[20] , \wRegInBot_6_51[19] , 
        \wRegInBot_6_51[18] , \wRegInBot_6_51[17] , \wRegInBot_6_51[16] , 
        \wRegInBot_6_51[15] , \wRegInBot_6_51[14] , \wRegInBot_6_51[13] , 
        \wRegInBot_6_51[12] , \wRegInBot_6_51[11] , \wRegInBot_6_51[10] , 
        \wRegInBot_6_51[9] , \wRegInBot_6_51[8] , \wRegInBot_6_51[7] , 
        \wRegInBot_6_51[6] , \wRegInBot_6_51[5] , \wRegInBot_6_51[4] , 
        \wRegInBot_6_51[3] , \wRegInBot_6_51[2] , \wRegInBot_6_51[1] , 
        \wRegInBot_6_51[0] }), .L_WR(\wRegEnTop_7_102[0] ), .L_In({
        \wRegOut_7_102[31] , \wRegOut_7_102[30] , \wRegOut_7_102[29] , 
        \wRegOut_7_102[28] , \wRegOut_7_102[27] , \wRegOut_7_102[26] , 
        \wRegOut_7_102[25] , \wRegOut_7_102[24] , \wRegOut_7_102[23] , 
        \wRegOut_7_102[22] , \wRegOut_7_102[21] , \wRegOut_7_102[20] , 
        \wRegOut_7_102[19] , \wRegOut_7_102[18] , \wRegOut_7_102[17] , 
        \wRegOut_7_102[16] , \wRegOut_7_102[15] , \wRegOut_7_102[14] , 
        \wRegOut_7_102[13] , \wRegOut_7_102[12] , \wRegOut_7_102[11] , 
        \wRegOut_7_102[10] , \wRegOut_7_102[9] , \wRegOut_7_102[8] , 
        \wRegOut_7_102[7] , \wRegOut_7_102[6] , \wRegOut_7_102[5] , 
        \wRegOut_7_102[4] , \wRegOut_7_102[3] , \wRegOut_7_102[2] , 
        \wRegOut_7_102[1] , \wRegOut_7_102[0] }), .L_Out({
        \wRegInTop_7_102[31] , \wRegInTop_7_102[30] , \wRegInTop_7_102[29] , 
        \wRegInTop_7_102[28] , \wRegInTop_7_102[27] , \wRegInTop_7_102[26] , 
        \wRegInTop_7_102[25] , \wRegInTop_7_102[24] , \wRegInTop_7_102[23] , 
        \wRegInTop_7_102[22] , \wRegInTop_7_102[21] , \wRegInTop_7_102[20] , 
        \wRegInTop_7_102[19] , \wRegInTop_7_102[18] , \wRegInTop_7_102[17] , 
        \wRegInTop_7_102[16] , \wRegInTop_7_102[15] , \wRegInTop_7_102[14] , 
        \wRegInTop_7_102[13] , \wRegInTop_7_102[12] , \wRegInTop_7_102[11] , 
        \wRegInTop_7_102[10] , \wRegInTop_7_102[9] , \wRegInTop_7_102[8] , 
        \wRegInTop_7_102[7] , \wRegInTop_7_102[6] , \wRegInTop_7_102[5] , 
        \wRegInTop_7_102[4] , \wRegInTop_7_102[3] , \wRegInTop_7_102[2] , 
        \wRegInTop_7_102[1] , \wRegInTop_7_102[0] }), .R_WR(
        \wRegEnTop_7_103[0] ), .R_In({\wRegOut_7_103[31] , \wRegOut_7_103[30] , 
        \wRegOut_7_103[29] , \wRegOut_7_103[28] , \wRegOut_7_103[27] , 
        \wRegOut_7_103[26] , \wRegOut_7_103[25] , \wRegOut_7_103[24] , 
        \wRegOut_7_103[23] , \wRegOut_7_103[22] , \wRegOut_7_103[21] , 
        \wRegOut_7_103[20] , \wRegOut_7_103[19] , \wRegOut_7_103[18] , 
        \wRegOut_7_103[17] , \wRegOut_7_103[16] , \wRegOut_7_103[15] , 
        \wRegOut_7_103[14] , \wRegOut_7_103[13] , \wRegOut_7_103[12] , 
        \wRegOut_7_103[11] , \wRegOut_7_103[10] , \wRegOut_7_103[9] , 
        \wRegOut_7_103[8] , \wRegOut_7_103[7] , \wRegOut_7_103[6] , 
        \wRegOut_7_103[5] , \wRegOut_7_103[4] , \wRegOut_7_103[3] , 
        \wRegOut_7_103[2] , \wRegOut_7_103[1] , \wRegOut_7_103[0] }), .R_Out({
        \wRegInTop_7_103[31] , \wRegInTop_7_103[30] , \wRegInTop_7_103[29] , 
        \wRegInTop_7_103[28] , \wRegInTop_7_103[27] , \wRegInTop_7_103[26] , 
        \wRegInTop_7_103[25] , \wRegInTop_7_103[24] , \wRegInTop_7_103[23] , 
        \wRegInTop_7_103[22] , \wRegInTop_7_103[21] , \wRegInTop_7_103[20] , 
        \wRegInTop_7_103[19] , \wRegInTop_7_103[18] , \wRegInTop_7_103[17] , 
        \wRegInTop_7_103[16] , \wRegInTop_7_103[15] , \wRegInTop_7_103[14] , 
        \wRegInTop_7_103[13] , \wRegInTop_7_103[12] , \wRegInTop_7_103[11] , 
        \wRegInTop_7_103[10] , \wRegInTop_7_103[9] , \wRegInTop_7_103[8] , 
        \wRegInTop_7_103[7] , \wRegInTop_7_103[6] , \wRegInTop_7_103[5] , 
        \wRegInTop_7_103[4] , \wRegInTop_7_103[3] , \wRegInTop_7_103[2] , 
        \wRegInTop_7_103[1] , \wRegInTop_7_103[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_17 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink81[31] , \ScanLink81[30] , \ScanLink81[29] , 
        \ScanLink81[28] , \ScanLink81[27] , \ScanLink81[26] , \ScanLink81[25] , 
        \ScanLink81[24] , \ScanLink81[23] , \ScanLink81[22] , \ScanLink81[21] , 
        \ScanLink81[20] , \ScanLink81[19] , \ScanLink81[18] , \ScanLink81[17] , 
        \ScanLink81[16] , \ScanLink81[15] , \ScanLink81[14] , \ScanLink81[13] , 
        \ScanLink81[12] , \ScanLink81[11] , \ScanLink81[10] , \ScanLink81[9] , 
        \ScanLink81[8] , \ScanLink81[7] , \ScanLink81[6] , \ScanLink81[5] , 
        \ScanLink81[4] , \ScanLink81[3] , \ScanLink81[2] , \ScanLink81[1] , 
        \ScanLink81[0] }), .ScanOut({\ScanLink80[31] , \ScanLink80[30] , 
        \ScanLink80[29] , \ScanLink80[28] , \ScanLink80[27] , \ScanLink80[26] , 
        \ScanLink80[25] , \ScanLink80[24] , \ScanLink80[23] , \ScanLink80[22] , 
        \ScanLink80[21] , \ScanLink80[20] , \ScanLink80[19] , \ScanLink80[18] , 
        \ScanLink80[17] , \ScanLink80[16] , \ScanLink80[15] , \ScanLink80[14] , 
        \ScanLink80[13] , \ScanLink80[12] , \ScanLink80[11] , \ScanLink80[10] , 
        \ScanLink80[9] , \ScanLink80[8] , \ScanLink80[7] , \ScanLink80[6] , 
        \ScanLink80[5] , \ScanLink80[4] , \ScanLink80[3] , \ScanLink80[2] , 
        \ScanLink80[1] , \ScanLink80[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_17[31] , \wRegOut_6_17[30] , 
        \wRegOut_6_17[29] , \wRegOut_6_17[28] , \wRegOut_6_17[27] , 
        \wRegOut_6_17[26] , \wRegOut_6_17[25] , \wRegOut_6_17[24] , 
        \wRegOut_6_17[23] , \wRegOut_6_17[22] , \wRegOut_6_17[21] , 
        \wRegOut_6_17[20] , \wRegOut_6_17[19] , \wRegOut_6_17[18] , 
        \wRegOut_6_17[17] , \wRegOut_6_17[16] , \wRegOut_6_17[15] , 
        \wRegOut_6_17[14] , \wRegOut_6_17[13] , \wRegOut_6_17[12] , 
        \wRegOut_6_17[11] , \wRegOut_6_17[10] , \wRegOut_6_17[9] , 
        \wRegOut_6_17[8] , \wRegOut_6_17[7] , \wRegOut_6_17[6] , 
        \wRegOut_6_17[5] , \wRegOut_6_17[4] , \wRegOut_6_17[3] , 
        \wRegOut_6_17[2] , \wRegOut_6_17[1] , \wRegOut_6_17[0] }), .Enable1(
        \wRegEnTop_6_17[0] ), .Enable2(\wRegEnBot_6_17[0] ), .In1({
        \wRegInTop_6_17[31] , \wRegInTop_6_17[30] , \wRegInTop_6_17[29] , 
        \wRegInTop_6_17[28] , \wRegInTop_6_17[27] , \wRegInTop_6_17[26] , 
        \wRegInTop_6_17[25] , \wRegInTop_6_17[24] , \wRegInTop_6_17[23] , 
        \wRegInTop_6_17[22] , \wRegInTop_6_17[21] , \wRegInTop_6_17[20] , 
        \wRegInTop_6_17[19] , \wRegInTop_6_17[18] , \wRegInTop_6_17[17] , 
        \wRegInTop_6_17[16] , \wRegInTop_6_17[15] , \wRegInTop_6_17[14] , 
        \wRegInTop_6_17[13] , \wRegInTop_6_17[12] , \wRegInTop_6_17[11] , 
        \wRegInTop_6_17[10] , \wRegInTop_6_17[9] , \wRegInTop_6_17[8] , 
        \wRegInTop_6_17[7] , \wRegInTop_6_17[6] , \wRegInTop_6_17[5] , 
        \wRegInTop_6_17[4] , \wRegInTop_6_17[3] , \wRegInTop_6_17[2] , 
        \wRegInTop_6_17[1] , \wRegInTop_6_17[0] }), .In2({\wRegInBot_6_17[31] , 
        \wRegInBot_6_17[30] , \wRegInBot_6_17[29] , \wRegInBot_6_17[28] , 
        \wRegInBot_6_17[27] , \wRegInBot_6_17[26] , \wRegInBot_6_17[25] , 
        \wRegInBot_6_17[24] , \wRegInBot_6_17[23] , \wRegInBot_6_17[22] , 
        \wRegInBot_6_17[21] , \wRegInBot_6_17[20] , \wRegInBot_6_17[19] , 
        \wRegInBot_6_17[18] , \wRegInBot_6_17[17] , \wRegInBot_6_17[16] , 
        \wRegInBot_6_17[15] , \wRegInBot_6_17[14] , \wRegInBot_6_17[13] , 
        \wRegInBot_6_17[12] , \wRegInBot_6_17[11] , \wRegInBot_6_17[10] , 
        \wRegInBot_6_17[9] , \wRegInBot_6_17[8] , \wRegInBot_6_17[7] , 
        \wRegInBot_6_17[6] , \wRegInBot_6_17[5] , \wRegInBot_6_17[4] , 
        \wRegInBot_6_17[3] , \wRegInBot_6_17[2] , \wRegInBot_6_17[1] , 
        \wRegInBot_6_17[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_30 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink94[31] , \ScanLink94[30] , \ScanLink94[29] , 
        \ScanLink94[28] , \ScanLink94[27] , \ScanLink94[26] , \ScanLink94[25] , 
        \ScanLink94[24] , \ScanLink94[23] , \ScanLink94[22] , \ScanLink94[21] , 
        \ScanLink94[20] , \ScanLink94[19] , \ScanLink94[18] , \ScanLink94[17] , 
        \ScanLink94[16] , \ScanLink94[15] , \ScanLink94[14] , \ScanLink94[13] , 
        \ScanLink94[12] , \ScanLink94[11] , \ScanLink94[10] , \ScanLink94[9] , 
        \ScanLink94[8] , \ScanLink94[7] , \ScanLink94[6] , \ScanLink94[5] , 
        \ScanLink94[4] , \ScanLink94[3] , \ScanLink94[2] , \ScanLink94[1] , 
        \ScanLink94[0] }), .ScanOut({\ScanLink93[31] , \ScanLink93[30] , 
        \ScanLink93[29] , \ScanLink93[28] , \ScanLink93[27] , \ScanLink93[26] , 
        \ScanLink93[25] , \ScanLink93[24] , \ScanLink93[23] , \ScanLink93[22] , 
        \ScanLink93[21] , \ScanLink93[20] , \ScanLink93[19] , \ScanLink93[18] , 
        \ScanLink93[17] , \ScanLink93[16] , \ScanLink93[15] , \ScanLink93[14] , 
        \ScanLink93[13] , \ScanLink93[12] , \ScanLink93[11] , \ScanLink93[10] , 
        \ScanLink93[9] , \ScanLink93[8] , \ScanLink93[7] , \ScanLink93[6] , 
        \ScanLink93[5] , \ScanLink93[4] , \ScanLink93[3] , \ScanLink93[2] , 
        \ScanLink93[1] , \ScanLink93[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_30[31] , \wRegOut_6_30[30] , 
        \wRegOut_6_30[29] , \wRegOut_6_30[28] , \wRegOut_6_30[27] , 
        \wRegOut_6_30[26] , \wRegOut_6_30[25] , \wRegOut_6_30[24] , 
        \wRegOut_6_30[23] , \wRegOut_6_30[22] , \wRegOut_6_30[21] , 
        \wRegOut_6_30[20] , \wRegOut_6_30[19] , \wRegOut_6_30[18] , 
        \wRegOut_6_30[17] , \wRegOut_6_30[16] , \wRegOut_6_30[15] , 
        \wRegOut_6_30[14] , \wRegOut_6_30[13] , \wRegOut_6_30[12] , 
        \wRegOut_6_30[11] , \wRegOut_6_30[10] , \wRegOut_6_30[9] , 
        \wRegOut_6_30[8] , \wRegOut_6_30[7] , \wRegOut_6_30[6] , 
        \wRegOut_6_30[5] , \wRegOut_6_30[4] , \wRegOut_6_30[3] , 
        \wRegOut_6_30[2] , \wRegOut_6_30[1] , \wRegOut_6_30[0] }), .Enable1(
        \wRegEnTop_6_30[0] ), .Enable2(\wRegEnBot_6_30[0] ), .In1({
        \wRegInTop_6_30[31] , \wRegInTop_6_30[30] , \wRegInTop_6_30[29] , 
        \wRegInTop_6_30[28] , \wRegInTop_6_30[27] , \wRegInTop_6_30[26] , 
        \wRegInTop_6_30[25] , \wRegInTop_6_30[24] , \wRegInTop_6_30[23] , 
        \wRegInTop_6_30[22] , \wRegInTop_6_30[21] , \wRegInTop_6_30[20] , 
        \wRegInTop_6_30[19] , \wRegInTop_6_30[18] , \wRegInTop_6_30[17] , 
        \wRegInTop_6_30[16] , \wRegInTop_6_30[15] , \wRegInTop_6_30[14] , 
        \wRegInTop_6_30[13] , \wRegInTop_6_30[12] , \wRegInTop_6_30[11] , 
        \wRegInTop_6_30[10] , \wRegInTop_6_30[9] , \wRegInTop_6_30[8] , 
        \wRegInTop_6_30[7] , \wRegInTop_6_30[6] , \wRegInTop_6_30[5] , 
        \wRegInTop_6_30[4] , \wRegInTop_6_30[3] , \wRegInTop_6_30[2] , 
        \wRegInTop_6_30[1] , \wRegInTop_6_30[0] }), .In2({\wRegInBot_6_30[31] , 
        \wRegInBot_6_30[30] , \wRegInBot_6_30[29] , \wRegInBot_6_30[28] , 
        \wRegInBot_6_30[27] , \wRegInBot_6_30[26] , \wRegInBot_6_30[25] , 
        \wRegInBot_6_30[24] , \wRegInBot_6_30[23] , \wRegInBot_6_30[22] , 
        \wRegInBot_6_30[21] , \wRegInBot_6_30[20] , \wRegInBot_6_30[19] , 
        \wRegInBot_6_30[18] , \wRegInBot_6_30[17] , \wRegInBot_6_30[16] , 
        \wRegInBot_6_30[15] , \wRegInBot_6_30[14] , \wRegInBot_6_30[13] , 
        \wRegInBot_6_30[12] , \wRegInBot_6_30[11] , \wRegInBot_6_30[10] , 
        \wRegInBot_6_30[9] , \wRegInBot_6_30[8] , \wRegInBot_6_30[7] , 
        \wRegInBot_6_30[6] , \wRegInBot_6_30[5] , \wRegInBot_6_30[4] , 
        \wRegInBot_6_30[3] , \wRegInBot_6_30[2] , \wRegInBot_6_30[1] , 
        \wRegInBot_6_30[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink130[31] , \ScanLink130[30] , \ScanLink130[29] , 
        \ScanLink130[28] , \ScanLink130[27] , \ScanLink130[26] , 
        \ScanLink130[25] , \ScanLink130[24] , \ScanLink130[23] , 
        \ScanLink130[22] , \ScanLink130[21] , \ScanLink130[20] , 
        \ScanLink130[19] , \ScanLink130[18] , \ScanLink130[17] , 
        \ScanLink130[16] , \ScanLink130[15] , \ScanLink130[14] , 
        \ScanLink130[13] , \ScanLink130[12] , \ScanLink130[11] , 
        \ScanLink130[10] , \ScanLink130[9] , \ScanLink130[8] , 
        \ScanLink130[7] , \ScanLink130[6] , \ScanLink130[5] , \ScanLink130[4] , 
        \ScanLink130[3] , \ScanLink130[2] , \ScanLink130[1] , \ScanLink130[0] 
        }), .ScanOut({\ScanLink129[31] , \ScanLink129[30] , \ScanLink129[29] , 
        \ScanLink129[28] , \ScanLink129[27] , \ScanLink129[26] , 
        \ScanLink129[25] , \ScanLink129[24] , \ScanLink129[23] , 
        \ScanLink129[22] , \ScanLink129[21] , \ScanLink129[20] , 
        \ScanLink129[19] , \ScanLink129[18] , \ScanLink129[17] , 
        \ScanLink129[16] , \ScanLink129[15] , \ScanLink129[14] , 
        \ScanLink129[13] , \ScanLink129[12] , \ScanLink129[11] , 
        \ScanLink129[10] , \ScanLink129[9] , \ScanLink129[8] , 
        \ScanLink129[7] , \ScanLink129[6] , \ScanLink129[5] , \ScanLink129[4] , 
        \ScanLink129[3] , \ScanLink129[2] , \ScanLink129[1] , \ScanLink129[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_2[31] , 
        \wRegOut_7_2[30] , \wRegOut_7_2[29] , \wRegOut_7_2[28] , 
        \wRegOut_7_2[27] , \wRegOut_7_2[26] , \wRegOut_7_2[25] , 
        \wRegOut_7_2[24] , \wRegOut_7_2[23] , \wRegOut_7_2[22] , 
        \wRegOut_7_2[21] , \wRegOut_7_2[20] , \wRegOut_7_2[19] , 
        \wRegOut_7_2[18] , \wRegOut_7_2[17] , \wRegOut_7_2[16] , 
        \wRegOut_7_2[15] , \wRegOut_7_2[14] , \wRegOut_7_2[13] , 
        \wRegOut_7_2[12] , \wRegOut_7_2[11] , \wRegOut_7_2[10] , 
        \wRegOut_7_2[9] , \wRegOut_7_2[8] , \wRegOut_7_2[7] , \wRegOut_7_2[6] , 
        \wRegOut_7_2[5] , \wRegOut_7_2[4] , \wRegOut_7_2[3] , \wRegOut_7_2[2] , 
        \wRegOut_7_2[1] , \wRegOut_7_2[0] }), .Enable1(\wRegEnTop_7_2[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_2[31] , \wRegInTop_7_2[30] , 
        \wRegInTop_7_2[29] , \wRegInTop_7_2[28] , \wRegInTop_7_2[27] , 
        \wRegInTop_7_2[26] , \wRegInTop_7_2[25] , \wRegInTop_7_2[24] , 
        \wRegInTop_7_2[23] , \wRegInTop_7_2[22] , \wRegInTop_7_2[21] , 
        \wRegInTop_7_2[20] , \wRegInTop_7_2[19] , \wRegInTop_7_2[18] , 
        \wRegInTop_7_2[17] , \wRegInTop_7_2[16] , \wRegInTop_7_2[15] , 
        \wRegInTop_7_2[14] , \wRegInTop_7_2[13] , \wRegInTop_7_2[12] , 
        \wRegInTop_7_2[11] , \wRegInTop_7_2[10] , \wRegInTop_7_2[9] , 
        \wRegInTop_7_2[8] , \wRegInTop_7_2[7] , \wRegInTop_7_2[6] , 
        \wRegInTop_7_2[5] , \wRegInTop_7_2[4] , \wRegInTop_7_2[3] , 
        \wRegInTop_7_2[2] , \wRegInTop_7_2[1] , \wRegInTop_7_2[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_44 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink172[31] , \ScanLink172[30] , \ScanLink172[29] , 
        \ScanLink172[28] , \ScanLink172[27] , \ScanLink172[26] , 
        \ScanLink172[25] , \ScanLink172[24] , \ScanLink172[23] , 
        \ScanLink172[22] , \ScanLink172[21] , \ScanLink172[20] , 
        \ScanLink172[19] , \ScanLink172[18] , \ScanLink172[17] , 
        \ScanLink172[16] , \ScanLink172[15] , \ScanLink172[14] , 
        \ScanLink172[13] , \ScanLink172[12] , \ScanLink172[11] , 
        \ScanLink172[10] , \ScanLink172[9] , \ScanLink172[8] , 
        \ScanLink172[7] , \ScanLink172[6] , \ScanLink172[5] , \ScanLink172[4] , 
        \ScanLink172[3] , \ScanLink172[2] , \ScanLink172[1] , \ScanLink172[0] 
        }), .ScanOut({\ScanLink171[31] , \ScanLink171[30] , \ScanLink171[29] , 
        \ScanLink171[28] , \ScanLink171[27] , \ScanLink171[26] , 
        \ScanLink171[25] , \ScanLink171[24] , \ScanLink171[23] , 
        \ScanLink171[22] , \ScanLink171[21] , \ScanLink171[20] , 
        \ScanLink171[19] , \ScanLink171[18] , \ScanLink171[17] , 
        \ScanLink171[16] , \ScanLink171[15] , \ScanLink171[14] , 
        \ScanLink171[13] , \ScanLink171[12] , \ScanLink171[11] , 
        \ScanLink171[10] , \ScanLink171[9] , \ScanLink171[8] , 
        \ScanLink171[7] , \ScanLink171[6] , \ScanLink171[5] , \ScanLink171[4] , 
        \ScanLink171[3] , \ScanLink171[2] , \ScanLink171[1] , \ScanLink171[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_44[31] , 
        \wRegOut_7_44[30] , \wRegOut_7_44[29] , \wRegOut_7_44[28] , 
        \wRegOut_7_44[27] , \wRegOut_7_44[26] , \wRegOut_7_44[25] , 
        \wRegOut_7_44[24] , \wRegOut_7_44[23] , \wRegOut_7_44[22] , 
        \wRegOut_7_44[21] , \wRegOut_7_44[20] , \wRegOut_7_44[19] , 
        \wRegOut_7_44[18] , \wRegOut_7_44[17] , \wRegOut_7_44[16] , 
        \wRegOut_7_44[15] , \wRegOut_7_44[14] , \wRegOut_7_44[13] , 
        \wRegOut_7_44[12] , \wRegOut_7_44[11] , \wRegOut_7_44[10] , 
        \wRegOut_7_44[9] , \wRegOut_7_44[8] , \wRegOut_7_44[7] , 
        \wRegOut_7_44[6] , \wRegOut_7_44[5] , \wRegOut_7_44[4] , 
        \wRegOut_7_44[3] , \wRegOut_7_44[2] , \wRegOut_7_44[1] , 
        \wRegOut_7_44[0] }), .Enable1(\wRegEnTop_7_44[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_44[31] , \wRegInTop_7_44[30] , \wRegInTop_7_44[29] , 
        \wRegInTop_7_44[28] , \wRegInTop_7_44[27] , \wRegInTop_7_44[26] , 
        \wRegInTop_7_44[25] , \wRegInTop_7_44[24] , \wRegInTop_7_44[23] , 
        \wRegInTop_7_44[22] , \wRegInTop_7_44[21] , \wRegInTop_7_44[20] , 
        \wRegInTop_7_44[19] , \wRegInTop_7_44[18] , \wRegInTop_7_44[17] , 
        \wRegInTop_7_44[16] , \wRegInTop_7_44[15] , \wRegInTop_7_44[14] , 
        \wRegInTop_7_44[13] , \wRegInTop_7_44[12] , \wRegInTop_7_44[11] , 
        \wRegInTop_7_44[10] , \wRegInTop_7_44[9] , \wRegInTop_7_44[8] , 
        \wRegInTop_7_44[7] , \wRegInTop_7_44[6] , \wRegInTop_7_44[5] , 
        \wRegInTop_7_44[4] , \wRegInTop_7_44[3] , \wRegInTop_7_44[2] , 
        \wRegInTop_7_44[1] , \wRegInTop_7_44[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_18[0] ), .P_In({\wRegOut_6_18[31] , 
        \wRegOut_6_18[30] , \wRegOut_6_18[29] , \wRegOut_6_18[28] , 
        \wRegOut_6_18[27] , \wRegOut_6_18[26] , \wRegOut_6_18[25] , 
        \wRegOut_6_18[24] , \wRegOut_6_18[23] , \wRegOut_6_18[22] , 
        \wRegOut_6_18[21] , \wRegOut_6_18[20] , \wRegOut_6_18[19] , 
        \wRegOut_6_18[18] , \wRegOut_6_18[17] , \wRegOut_6_18[16] , 
        \wRegOut_6_18[15] , \wRegOut_6_18[14] , \wRegOut_6_18[13] , 
        \wRegOut_6_18[12] , \wRegOut_6_18[11] , \wRegOut_6_18[10] , 
        \wRegOut_6_18[9] , \wRegOut_6_18[8] , \wRegOut_6_18[7] , 
        \wRegOut_6_18[6] , \wRegOut_6_18[5] , \wRegOut_6_18[4] , 
        \wRegOut_6_18[3] , \wRegOut_6_18[2] , \wRegOut_6_18[1] , 
        \wRegOut_6_18[0] }), .P_Out({\wRegInBot_6_18[31] , 
        \wRegInBot_6_18[30] , \wRegInBot_6_18[29] , \wRegInBot_6_18[28] , 
        \wRegInBot_6_18[27] , \wRegInBot_6_18[26] , \wRegInBot_6_18[25] , 
        \wRegInBot_6_18[24] , \wRegInBot_6_18[23] , \wRegInBot_6_18[22] , 
        \wRegInBot_6_18[21] , \wRegInBot_6_18[20] , \wRegInBot_6_18[19] , 
        \wRegInBot_6_18[18] , \wRegInBot_6_18[17] , \wRegInBot_6_18[16] , 
        \wRegInBot_6_18[15] , \wRegInBot_6_18[14] , \wRegInBot_6_18[13] , 
        \wRegInBot_6_18[12] , \wRegInBot_6_18[11] , \wRegInBot_6_18[10] , 
        \wRegInBot_6_18[9] , \wRegInBot_6_18[8] , \wRegInBot_6_18[7] , 
        \wRegInBot_6_18[6] , \wRegInBot_6_18[5] , \wRegInBot_6_18[4] , 
        \wRegInBot_6_18[3] , \wRegInBot_6_18[2] , \wRegInBot_6_18[1] , 
        \wRegInBot_6_18[0] }), .L_WR(\wRegEnTop_7_36[0] ), .L_In({
        \wRegOut_7_36[31] , \wRegOut_7_36[30] , \wRegOut_7_36[29] , 
        \wRegOut_7_36[28] , \wRegOut_7_36[27] , \wRegOut_7_36[26] , 
        \wRegOut_7_36[25] , \wRegOut_7_36[24] , \wRegOut_7_36[23] , 
        \wRegOut_7_36[22] , \wRegOut_7_36[21] , \wRegOut_7_36[20] , 
        \wRegOut_7_36[19] , \wRegOut_7_36[18] , \wRegOut_7_36[17] , 
        \wRegOut_7_36[16] , \wRegOut_7_36[15] , \wRegOut_7_36[14] , 
        \wRegOut_7_36[13] , \wRegOut_7_36[12] , \wRegOut_7_36[11] , 
        \wRegOut_7_36[10] , \wRegOut_7_36[9] , \wRegOut_7_36[8] , 
        \wRegOut_7_36[7] , \wRegOut_7_36[6] , \wRegOut_7_36[5] , 
        \wRegOut_7_36[4] , \wRegOut_7_36[3] , \wRegOut_7_36[2] , 
        \wRegOut_7_36[1] , \wRegOut_7_36[0] }), .L_Out({\wRegInTop_7_36[31] , 
        \wRegInTop_7_36[30] , \wRegInTop_7_36[29] , \wRegInTop_7_36[28] , 
        \wRegInTop_7_36[27] , \wRegInTop_7_36[26] , \wRegInTop_7_36[25] , 
        \wRegInTop_7_36[24] , \wRegInTop_7_36[23] , \wRegInTop_7_36[22] , 
        \wRegInTop_7_36[21] , \wRegInTop_7_36[20] , \wRegInTop_7_36[19] , 
        \wRegInTop_7_36[18] , \wRegInTop_7_36[17] , \wRegInTop_7_36[16] , 
        \wRegInTop_7_36[15] , \wRegInTop_7_36[14] , \wRegInTop_7_36[13] , 
        \wRegInTop_7_36[12] , \wRegInTop_7_36[11] , \wRegInTop_7_36[10] , 
        \wRegInTop_7_36[9] , \wRegInTop_7_36[8] , \wRegInTop_7_36[7] , 
        \wRegInTop_7_36[6] , \wRegInTop_7_36[5] , \wRegInTop_7_36[4] , 
        \wRegInTop_7_36[3] , \wRegInTop_7_36[2] , \wRegInTop_7_36[1] , 
        \wRegInTop_7_36[0] }), .R_WR(\wRegEnTop_7_37[0] ), .R_In({
        \wRegOut_7_37[31] , \wRegOut_7_37[30] , \wRegOut_7_37[29] , 
        \wRegOut_7_37[28] , \wRegOut_7_37[27] , \wRegOut_7_37[26] , 
        \wRegOut_7_37[25] , \wRegOut_7_37[24] , \wRegOut_7_37[23] , 
        \wRegOut_7_37[22] , \wRegOut_7_37[21] , \wRegOut_7_37[20] , 
        \wRegOut_7_37[19] , \wRegOut_7_37[18] , \wRegOut_7_37[17] , 
        \wRegOut_7_37[16] , \wRegOut_7_37[15] , \wRegOut_7_37[14] , 
        \wRegOut_7_37[13] , \wRegOut_7_37[12] , \wRegOut_7_37[11] , 
        \wRegOut_7_37[10] , \wRegOut_7_37[9] , \wRegOut_7_37[8] , 
        \wRegOut_7_37[7] , \wRegOut_7_37[6] , \wRegOut_7_37[5] , 
        \wRegOut_7_37[4] , \wRegOut_7_37[3] , \wRegOut_7_37[2] , 
        \wRegOut_7_37[1] , \wRegOut_7_37[0] }), .R_Out({\wRegInTop_7_37[31] , 
        \wRegInTop_7_37[30] , \wRegInTop_7_37[29] , \wRegInTop_7_37[28] , 
        \wRegInTop_7_37[27] , \wRegInTop_7_37[26] , \wRegInTop_7_37[25] , 
        \wRegInTop_7_37[24] , \wRegInTop_7_37[23] , \wRegInTop_7_37[22] , 
        \wRegInTop_7_37[21] , \wRegInTop_7_37[20] , \wRegInTop_7_37[19] , 
        \wRegInTop_7_37[18] , \wRegInTop_7_37[17] , \wRegInTop_7_37[16] , 
        \wRegInTop_7_37[15] , \wRegInTop_7_37[14] , \wRegInTop_7_37[13] , 
        \wRegInTop_7_37[12] , \wRegInTop_7_37[11] , \wRegInTop_7_37[10] , 
        \wRegInTop_7_37[9] , \wRegInTop_7_37[8] , \wRegInTop_7_37[7] , 
        \wRegInTop_7_37[6] , \wRegInTop_7_37[5] , \wRegInTop_7_37[4] , 
        \wRegInTop_7_37[3] , \wRegInTop_7_37[2] , \wRegInTop_7_37[1] , 
        \wRegInTop_7_37[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_71 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink199[31] , \ScanLink199[30] , \ScanLink199[29] , 
        \ScanLink199[28] , \ScanLink199[27] , \ScanLink199[26] , 
        \ScanLink199[25] , \ScanLink199[24] , \ScanLink199[23] , 
        \ScanLink199[22] , \ScanLink199[21] , \ScanLink199[20] , 
        \ScanLink199[19] , \ScanLink199[18] , \ScanLink199[17] , 
        \ScanLink199[16] , \ScanLink199[15] , \ScanLink199[14] , 
        \ScanLink199[13] , \ScanLink199[12] , \ScanLink199[11] , 
        \ScanLink199[10] , \ScanLink199[9] , \ScanLink199[8] , 
        \ScanLink199[7] , \ScanLink199[6] , \ScanLink199[5] , \ScanLink199[4] , 
        \ScanLink199[3] , \ScanLink199[2] , \ScanLink199[1] , \ScanLink199[0] 
        }), .ScanOut({\ScanLink198[31] , \ScanLink198[30] , \ScanLink198[29] , 
        \ScanLink198[28] , \ScanLink198[27] , \ScanLink198[26] , 
        \ScanLink198[25] , \ScanLink198[24] , \ScanLink198[23] , 
        \ScanLink198[22] , \ScanLink198[21] , \ScanLink198[20] , 
        \ScanLink198[19] , \ScanLink198[18] , \ScanLink198[17] , 
        \ScanLink198[16] , \ScanLink198[15] , \ScanLink198[14] , 
        \ScanLink198[13] , \ScanLink198[12] , \ScanLink198[11] , 
        \ScanLink198[10] , \ScanLink198[9] , \ScanLink198[8] , 
        \ScanLink198[7] , \ScanLink198[6] , \ScanLink198[5] , \ScanLink198[4] , 
        \ScanLink198[3] , \ScanLink198[2] , \ScanLink198[1] , \ScanLink198[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_71[31] , 
        \wRegOut_7_71[30] , \wRegOut_7_71[29] , \wRegOut_7_71[28] , 
        \wRegOut_7_71[27] , \wRegOut_7_71[26] , \wRegOut_7_71[25] , 
        \wRegOut_7_71[24] , \wRegOut_7_71[23] , \wRegOut_7_71[22] , 
        \wRegOut_7_71[21] , \wRegOut_7_71[20] , \wRegOut_7_71[19] , 
        \wRegOut_7_71[18] , \wRegOut_7_71[17] , \wRegOut_7_71[16] , 
        \wRegOut_7_71[15] , \wRegOut_7_71[14] , \wRegOut_7_71[13] , 
        \wRegOut_7_71[12] , \wRegOut_7_71[11] , \wRegOut_7_71[10] , 
        \wRegOut_7_71[9] , \wRegOut_7_71[8] , \wRegOut_7_71[7] , 
        \wRegOut_7_71[6] , \wRegOut_7_71[5] , \wRegOut_7_71[4] , 
        \wRegOut_7_71[3] , \wRegOut_7_71[2] , \wRegOut_7_71[1] , 
        \wRegOut_7_71[0] }), .Enable1(\wRegEnTop_7_71[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_71[31] , \wRegInTop_7_71[30] , \wRegInTop_7_71[29] , 
        \wRegInTop_7_71[28] , \wRegInTop_7_71[27] , \wRegInTop_7_71[26] , 
        \wRegInTop_7_71[25] , \wRegInTop_7_71[24] , \wRegInTop_7_71[23] , 
        \wRegInTop_7_71[22] , \wRegInTop_7_71[21] , \wRegInTop_7_71[20] , 
        \wRegInTop_7_71[19] , \wRegInTop_7_71[18] , \wRegInTop_7_71[17] , 
        \wRegInTop_7_71[16] , \wRegInTop_7_71[15] , \wRegInTop_7_71[14] , 
        \wRegInTop_7_71[13] , \wRegInTop_7_71[12] , \wRegInTop_7_71[11] , 
        \wRegInTop_7_71[10] , \wRegInTop_7_71[9] , \wRegInTop_7_71[8] , 
        \wRegInTop_7_71[7] , \wRegInTop_7_71[6] , \wRegInTop_7_71[5] , 
        \wRegInTop_7_71[4] , \wRegInTop_7_71[3] , \wRegInTop_7_71[2] , 
        \wRegInTop_7_71[1] , \wRegInTop_7_71[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_28[0] ), .P_In({\wRegOut_5_28[31] , 
        \wRegOut_5_28[30] , \wRegOut_5_28[29] , \wRegOut_5_28[28] , 
        \wRegOut_5_28[27] , \wRegOut_5_28[26] , \wRegOut_5_28[25] , 
        \wRegOut_5_28[24] , \wRegOut_5_28[23] , \wRegOut_5_28[22] , 
        \wRegOut_5_28[21] , \wRegOut_5_28[20] , \wRegOut_5_28[19] , 
        \wRegOut_5_28[18] , \wRegOut_5_28[17] , \wRegOut_5_28[16] , 
        \wRegOut_5_28[15] , \wRegOut_5_28[14] , \wRegOut_5_28[13] , 
        \wRegOut_5_28[12] , \wRegOut_5_28[11] , \wRegOut_5_28[10] , 
        \wRegOut_5_28[9] , \wRegOut_5_28[8] , \wRegOut_5_28[7] , 
        \wRegOut_5_28[6] , \wRegOut_5_28[5] , \wRegOut_5_28[4] , 
        \wRegOut_5_28[3] , \wRegOut_5_28[2] , \wRegOut_5_28[1] , 
        \wRegOut_5_28[0] }), .P_Out({\wRegInBot_5_28[31] , 
        \wRegInBot_5_28[30] , \wRegInBot_5_28[29] , \wRegInBot_5_28[28] , 
        \wRegInBot_5_28[27] , \wRegInBot_5_28[26] , \wRegInBot_5_28[25] , 
        \wRegInBot_5_28[24] , \wRegInBot_5_28[23] , \wRegInBot_5_28[22] , 
        \wRegInBot_5_28[21] , \wRegInBot_5_28[20] , \wRegInBot_5_28[19] , 
        \wRegInBot_5_28[18] , \wRegInBot_5_28[17] , \wRegInBot_5_28[16] , 
        \wRegInBot_5_28[15] , \wRegInBot_5_28[14] , \wRegInBot_5_28[13] , 
        \wRegInBot_5_28[12] , \wRegInBot_5_28[11] , \wRegInBot_5_28[10] , 
        \wRegInBot_5_28[9] , \wRegInBot_5_28[8] , \wRegInBot_5_28[7] , 
        \wRegInBot_5_28[6] , \wRegInBot_5_28[5] , \wRegInBot_5_28[4] , 
        \wRegInBot_5_28[3] , \wRegInBot_5_28[2] , \wRegInBot_5_28[1] , 
        \wRegInBot_5_28[0] }), .L_WR(\wRegEnTop_6_56[0] ), .L_In({
        \wRegOut_6_56[31] , \wRegOut_6_56[30] , \wRegOut_6_56[29] , 
        \wRegOut_6_56[28] , \wRegOut_6_56[27] , \wRegOut_6_56[26] , 
        \wRegOut_6_56[25] , \wRegOut_6_56[24] , \wRegOut_6_56[23] , 
        \wRegOut_6_56[22] , \wRegOut_6_56[21] , \wRegOut_6_56[20] , 
        \wRegOut_6_56[19] , \wRegOut_6_56[18] , \wRegOut_6_56[17] , 
        \wRegOut_6_56[16] , \wRegOut_6_56[15] , \wRegOut_6_56[14] , 
        \wRegOut_6_56[13] , \wRegOut_6_56[12] , \wRegOut_6_56[11] , 
        \wRegOut_6_56[10] , \wRegOut_6_56[9] , \wRegOut_6_56[8] , 
        \wRegOut_6_56[7] , \wRegOut_6_56[6] , \wRegOut_6_56[5] , 
        \wRegOut_6_56[4] , \wRegOut_6_56[3] , \wRegOut_6_56[2] , 
        \wRegOut_6_56[1] , \wRegOut_6_56[0] }), .L_Out({\wRegInTop_6_56[31] , 
        \wRegInTop_6_56[30] , \wRegInTop_6_56[29] , \wRegInTop_6_56[28] , 
        \wRegInTop_6_56[27] , \wRegInTop_6_56[26] , \wRegInTop_6_56[25] , 
        \wRegInTop_6_56[24] , \wRegInTop_6_56[23] , \wRegInTop_6_56[22] , 
        \wRegInTop_6_56[21] , \wRegInTop_6_56[20] , \wRegInTop_6_56[19] , 
        \wRegInTop_6_56[18] , \wRegInTop_6_56[17] , \wRegInTop_6_56[16] , 
        \wRegInTop_6_56[15] , \wRegInTop_6_56[14] , \wRegInTop_6_56[13] , 
        \wRegInTop_6_56[12] , \wRegInTop_6_56[11] , \wRegInTop_6_56[10] , 
        \wRegInTop_6_56[9] , \wRegInTop_6_56[8] , \wRegInTop_6_56[7] , 
        \wRegInTop_6_56[6] , \wRegInTop_6_56[5] , \wRegInTop_6_56[4] , 
        \wRegInTop_6_56[3] , \wRegInTop_6_56[2] , \wRegInTop_6_56[1] , 
        \wRegInTop_6_56[0] }), .R_WR(\wRegEnTop_6_57[0] ), .R_In({
        \wRegOut_6_57[31] , \wRegOut_6_57[30] , \wRegOut_6_57[29] , 
        \wRegOut_6_57[28] , \wRegOut_6_57[27] , \wRegOut_6_57[26] , 
        \wRegOut_6_57[25] , \wRegOut_6_57[24] , \wRegOut_6_57[23] , 
        \wRegOut_6_57[22] , \wRegOut_6_57[21] , \wRegOut_6_57[20] , 
        \wRegOut_6_57[19] , \wRegOut_6_57[18] , \wRegOut_6_57[17] , 
        \wRegOut_6_57[16] , \wRegOut_6_57[15] , \wRegOut_6_57[14] , 
        \wRegOut_6_57[13] , \wRegOut_6_57[12] , \wRegOut_6_57[11] , 
        \wRegOut_6_57[10] , \wRegOut_6_57[9] , \wRegOut_6_57[8] , 
        \wRegOut_6_57[7] , \wRegOut_6_57[6] , \wRegOut_6_57[5] , 
        \wRegOut_6_57[4] , \wRegOut_6_57[3] , \wRegOut_6_57[2] , 
        \wRegOut_6_57[1] , \wRegOut_6_57[0] }), .R_Out({\wRegInTop_6_57[31] , 
        \wRegInTop_6_57[30] , \wRegInTop_6_57[29] , \wRegInTop_6_57[28] , 
        \wRegInTop_6_57[27] , \wRegInTop_6_57[26] , \wRegInTop_6_57[25] , 
        \wRegInTop_6_57[24] , \wRegInTop_6_57[23] , \wRegInTop_6_57[22] , 
        \wRegInTop_6_57[21] , \wRegInTop_6_57[20] , \wRegInTop_6_57[19] , 
        \wRegInTop_6_57[18] , \wRegInTop_6_57[17] , \wRegInTop_6_57[16] , 
        \wRegInTop_6_57[15] , \wRegInTop_6_57[14] , \wRegInTop_6_57[13] , 
        \wRegInTop_6_57[12] , \wRegInTop_6_57[11] , \wRegInTop_6_57[10] , 
        \wRegInTop_6_57[9] , \wRegInTop_6_57[8] , \wRegInTop_6_57[7] , 
        \wRegInTop_6_57[6] , \wRegInTop_6_57[5] , \wRegInTop_6_57[4] , 
        \wRegInTop_6_57[3] , \wRegInTop_6_57[2] , \wRegInTop_6_57[1] , 
        \wRegInTop_6_57[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink44[31] , \ScanLink44[30] , \ScanLink44[29] , 
        \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , \ScanLink44[25] , 
        \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , \ScanLink44[21] , 
        \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , \ScanLink44[17] , 
        \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , \ScanLink44[13] , 
        \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , \ScanLink44[9] , 
        \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , \ScanLink44[5] , 
        \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , \ScanLink44[1] , 
        \ScanLink44[0] }), .ScanOut({\ScanLink43[31] , \ScanLink43[30] , 
        \ScanLink43[29] , \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , 
        \ScanLink43[25] , \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , 
        \ScanLink43[21] , \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , 
        \ScanLink43[17] , \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , 
        \ScanLink43[13] , \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , 
        \ScanLink43[9] , \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , 
        \ScanLink43[5] , \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , 
        \ScanLink43[1] , \ScanLink43[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_12[31] , \wRegOut_5_12[30] , 
        \wRegOut_5_12[29] , \wRegOut_5_12[28] , \wRegOut_5_12[27] , 
        \wRegOut_5_12[26] , \wRegOut_5_12[25] , \wRegOut_5_12[24] , 
        \wRegOut_5_12[23] , \wRegOut_5_12[22] , \wRegOut_5_12[21] , 
        \wRegOut_5_12[20] , \wRegOut_5_12[19] , \wRegOut_5_12[18] , 
        \wRegOut_5_12[17] , \wRegOut_5_12[16] , \wRegOut_5_12[15] , 
        \wRegOut_5_12[14] , \wRegOut_5_12[13] , \wRegOut_5_12[12] , 
        \wRegOut_5_12[11] , \wRegOut_5_12[10] , \wRegOut_5_12[9] , 
        \wRegOut_5_12[8] , \wRegOut_5_12[7] , \wRegOut_5_12[6] , 
        \wRegOut_5_12[5] , \wRegOut_5_12[4] , \wRegOut_5_12[3] , 
        \wRegOut_5_12[2] , \wRegOut_5_12[1] , \wRegOut_5_12[0] }), .Enable1(
        \wRegEnTop_5_12[0] ), .Enable2(\wRegEnBot_5_12[0] ), .In1({
        \wRegInTop_5_12[31] , \wRegInTop_5_12[30] , \wRegInTop_5_12[29] , 
        \wRegInTop_5_12[28] , \wRegInTop_5_12[27] , \wRegInTop_5_12[26] , 
        \wRegInTop_5_12[25] , \wRegInTop_5_12[24] , \wRegInTop_5_12[23] , 
        \wRegInTop_5_12[22] , \wRegInTop_5_12[21] , \wRegInTop_5_12[20] , 
        \wRegInTop_5_12[19] , \wRegInTop_5_12[18] , \wRegInTop_5_12[17] , 
        \wRegInTop_5_12[16] , \wRegInTop_5_12[15] , \wRegInTop_5_12[14] , 
        \wRegInTop_5_12[13] , \wRegInTop_5_12[12] , \wRegInTop_5_12[11] , 
        \wRegInTop_5_12[10] , \wRegInTop_5_12[9] , \wRegInTop_5_12[8] , 
        \wRegInTop_5_12[7] , \wRegInTop_5_12[6] , \wRegInTop_5_12[5] , 
        \wRegInTop_5_12[4] , \wRegInTop_5_12[3] , \wRegInTop_5_12[2] , 
        \wRegInTop_5_12[1] , \wRegInTop_5_12[0] }), .In2({\wRegInBot_5_12[31] , 
        \wRegInBot_5_12[30] , \wRegInBot_5_12[29] , \wRegInBot_5_12[28] , 
        \wRegInBot_5_12[27] , \wRegInBot_5_12[26] , \wRegInBot_5_12[25] , 
        \wRegInBot_5_12[24] , \wRegInBot_5_12[23] , \wRegInBot_5_12[22] , 
        \wRegInBot_5_12[21] , \wRegInBot_5_12[20] , \wRegInBot_5_12[19] , 
        \wRegInBot_5_12[18] , \wRegInBot_5_12[17] , \wRegInBot_5_12[16] , 
        \wRegInBot_5_12[15] , \wRegInBot_5_12[14] , \wRegInBot_5_12[13] , 
        \wRegInBot_5_12[12] , \wRegInBot_5_12[11] , \wRegInBot_5_12[10] , 
        \wRegInBot_5_12[9] , \wRegInBot_5_12[8] , \wRegInBot_5_12[7] , 
        \wRegInBot_5_12[6] , \wRegInBot_5_12[5] , \wRegInBot_5_12[4] , 
        \wRegInBot_5_12[3] , \wRegInBot_5_12[2] , \wRegInBot_5_12[1] , 
        \wRegInBot_5_12[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_2_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink4[31] , \ScanLink4[30] , \ScanLink4[29] , 
        \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , \ScanLink4[25] , 
        \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , \ScanLink4[21] , 
        \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , \ScanLink4[17] , 
        \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , \ScanLink4[13] , 
        \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , \ScanLink4[9] , 
        \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , \ScanLink4[5] , 
        \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , \ScanLink4[1] , 
        \ScanLink4[0] }), .ScanOut({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_2_0[31] , \wRegOut_2_0[30] , \wRegOut_2_0[29] , 
        \wRegOut_2_0[28] , \wRegOut_2_0[27] , \wRegOut_2_0[26] , 
        \wRegOut_2_0[25] , \wRegOut_2_0[24] , \wRegOut_2_0[23] , 
        \wRegOut_2_0[22] , \wRegOut_2_0[21] , \wRegOut_2_0[20] , 
        \wRegOut_2_0[19] , \wRegOut_2_0[18] , \wRegOut_2_0[17] , 
        \wRegOut_2_0[16] , \wRegOut_2_0[15] , \wRegOut_2_0[14] , 
        \wRegOut_2_0[13] , \wRegOut_2_0[12] , \wRegOut_2_0[11] , 
        \wRegOut_2_0[10] , \wRegOut_2_0[9] , \wRegOut_2_0[8] , 
        \wRegOut_2_0[7] , \wRegOut_2_0[6] , \wRegOut_2_0[5] , \wRegOut_2_0[4] , 
        \wRegOut_2_0[3] , \wRegOut_2_0[2] , \wRegOut_2_0[1] , \wRegOut_2_0[0] 
        }), .Enable1(\wRegEnTop_2_0[0] ), .Enable2(\wRegEnBot_2_0[0] ), .In1({
        \wRegInTop_2_0[31] , \wRegInTop_2_0[30] , \wRegInTop_2_0[29] , 
        \wRegInTop_2_0[28] , \wRegInTop_2_0[27] , \wRegInTop_2_0[26] , 
        \wRegInTop_2_0[25] , \wRegInTop_2_0[24] , \wRegInTop_2_0[23] , 
        \wRegInTop_2_0[22] , \wRegInTop_2_0[21] , \wRegInTop_2_0[20] , 
        \wRegInTop_2_0[19] , \wRegInTop_2_0[18] , \wRegInTop_2_0[17] , 
        \wRegInTop_2_0[16] , \wRegInTop_2_0[15] , \wRegInTop_2_0[14] , 
        \wRegInTop_2_0[13] , \wRegInTop_2_0[12] , \wRegInTop_2_0[11] , 
        \wRegInTop_2_0[10] , \wRegInTop_2_0[9] , \wRegInTop_2_0[8] , 
        \wRegInTop_2_0[7] , \wRegInTop_2_0[6] , \wRegInTop_2_0[5] , 
        \wRegInTop_2_0[4] , \wRegInTop_2_0[3] , \wRegInTop_2_0[2] , 
        \wRegInTop_2_0[1] , \wRegInTop_2_0[0] }), .In2({\wRegInBot_2_0[31] , 
        \wRegInBot_2_0[30] , \wRegInBot_2_0[29] , \wRegInBot_2_0[28] , 
        \wRegInBot_2_0[27] , \wRegInBot_2_0[26] , \wRegInBot_2_0[25] , 
        \wRegInBot_2_0[24] , \wRegInBot_2_0[23] , \wRegInBot_2_0[22] , 
        \wRegInBot_2_0[21] , \wRegInBot_2_0[20] , \wRegInBot_2_0[19] , 
        \wRegInBot_2_0[18] , \wRegInBot_2_0[17] , \wRegInBot_2_0[16] , 
        \wRegInBot_2_0[15] , \wRegInBot_2_0[14] , \wRegInBot_2_0[13] , 
        \wRegInBot_2_0[12] , \wRegInBot_2_0[11] , \wRegInBot_2_0[10] , 
        \wRegInBot_2_0[9] , \wRegInBot_2_0[8] , \wRegInBot_2_0[7] , 
        \wRegInBot_2_0[6] , \wRegInBot_2_0[5] , \wRegInBot_2_0[4] , 
        \wRegInBot_2_0[3] , \wRegInBot_2_0[2] , \wRegInBot_2_0[1] , 
        \wRegInBot_2_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_2_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink5[31] , \ScanLink5[30] , \ScanLink5[29] , 
        \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , \ScanLink5[25] , 
        \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , \ScanLink5[21] , 
        \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , \ScanLink5[17] , 
        \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , \ScanLink5[13] , 
        \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , \ScanLink5[9] , 
        \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , \ScanLink5[5] , 
        \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , \ScanLink5[1] , 
        \ScanLink5[0] }), .ScanOut({\ScanLink4[31] , \ScanLink4[30] , 
        \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , 
        \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , 
        \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , 
        \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , 
        \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , 
        \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_2_1[31] , \wRegOut_2_1[30] , \wRegOut_2_1[29] , 
        \wRegOut_2_1[28] , \wRegOut_2_1[27] , \wRegOut_2_1[26] , 
        \wRegOut_2_1[25] , \wRegOut_2_1[24] , \wRegOut_2_1[23] , 
        \wRegOut_2_1[22] , \wRegOut_2_1[21] , \wRegOut_2_1[20] , 
        \wRegOut_2_1[19] , \wRegOut_2_1[18] , \wRegOut_2_1[17] , 
        \wRegOut_2_1[16] , \wRegOut_2_1[15] , \wRegOut_2_1[14] , 
        \wRegOut_2_1[13] , \wRegOut_2_1[12] , \wRegOut_2_1[11] , 
        \wRegOut_2_1[10] , \wRegOut_2_1[9] , \wRegOut_2_1[8] , 
        \wRegOut_2_1[7] , \wRegOut_2_1[6] , \wRegOut_2_1[5] , \wRegOut_2_1[4] , 
        \wRegOut_2_1[3] , \wRegOut_2_1[2] , \wRegOut_2_1[1] , \wRegOut_2_1[0] 
        }), .Enable1(\wRegEnTop_2_1[0] ), .Enable2(\wRegEnBot_2_1[0] ), .In1({
        \wRegInTop_2_1[31] , \wRegInTop_2_1[30] , \wRegInTop_2_1[29] , 
        \wRegInTop_2_1[28] , \wRegInTop_2_1[27] , \wRegInTop_2_1[26] , 
        \wRegInTop_2_1[25] , \wRegInTop_2_1[24] , \wRegInTop_2_1[23] , 
        \wRegInTop_2_1[22] , \wRegInTop_2_1[21] , \wRegInTop_2_1[20] , 
        \wRegInTop_2_1[19] , \wRegInTop_2_1[18] , \wRegInTop_2_1[17] , 
        \wRegInTop_2_1[16] , \wRegInTop_2_1[15] , \wRegInTop_2_1[14] , 
        \wRegInTop_2_1[13] , \wRegInTop_2_1[12] , \wRegInTop_2_1[11] , 
        \wRegInTop_2_1[10] , \wRegInTop_2_1[9] , \wRegInTop_2_1[8] , 
        \wRegInTop_2_1[7] , \wRegInTop_2_1[6] , \wRegInTop_2_1[5] , 
        \wRegInTop_2_1[4] , \wRegInTop_2_1[3] , \wRegInTop_2_1[2] , 
        \wRegInTop_2_1[1] , \wRegInTop_2_1[0] }), .In2({\wRegInBot_2_1[31] , 
        \wRegInBot_2_1[30] , \wRegInBot_2_1[29] , \wRegInBot_2_1[28] , 
        \wRegInBot_2_1[27] , \wRegInBot_2_1[26] , \wRegInBot_2_1[25] , 
        \wRegInBot_2_1[24] , \wRegInBot_2_1[23] , \wRegInBot_2_1[22] , 
        \wRegInBot_2_1[21] , \wRegInBot_2_1[20] , \wRegInBot_2_1[19] , 
        \wRegInBot_2_1[18] , \wRegInBot_2_1[17] , \wRegInBot_2_1[16] , 
        \wRegInBot_2_1[15] , \wRegInBot_2_1[14] , \wRegInBot_2_1[13] , 
        \wRegInBot_2_1[12] , \wRegInBot_2_1[11] , \wRegInBot_2_1[10] , 
        \wRegInBot_2_1[9] , \wRegInBot_2_1[8] , \wRegInBot_2_1[7] , 
        \wRegInBot_2_1[6] , \wRegInBot_2_1[5] , \wRegInBot_2_1[4] , 
        \wRegInBot_2_1[3] , \wRegInBot_2_1[2] , \wRegInBot_2_1[1] , 
        \wRegInBot_2_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink9[31] , \ScanLink9[30] , \ScanLink9[29] , 
        \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , \ScanLink9[25] , 
        \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , \ScanLink9[21] , 
        \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , \ScanLink9[17] , 
        \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , \ScanLink9[13] , 
        \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , \ScanLink9[9] , 
        \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , \ScanLink9[5] , 
        \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , \ScanLink9[1] , 
        \ScanLink9[0] }), .ScanOut({\ScanLink8[31] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , 
        \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , 
        \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , 
        \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , 
        \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , 
        \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_1[31] , \wRegOut_3_1[30] , \wRegOut_3_1[29] , 
        \wRegOut_3_1[28] , \wRegOut_3_1[27] , \wRegOut_3_1[26] , 
        \wRegOut_3_1[25] , \wRegOut_3_1[24] , \wRegOut_3_1[23] , 
        \wRegOut_3_1[22] , \wRegOut_3_1[21] , \wRegOut_3_1[20] , 
        \wRegOut_3_1[19] , \wRegOut_3_1[18] , \wRegOut_3_1[17] , 
        \wRegOut_3_1[16] , \wRegOut_3_1[15] , \wRegOut_3_1[14] , 
        \wRegOut_3_1[13] , \wRegOut_3_1[12] , \wRegOut_3_1[11] , 
        \wRegOut_3_1[10] , \wRegOut_3_1[9] , \wRegOut_3_1[8] , 
        \wRegOut_3_1[7] , \wRegOut_3_1[6] , \wRegOut_3_1[5] , \wRegOut_3_1[4] , 
        \wRegOut_3_1[3] , \wRegOut_3_1[2] , \wRegOut_3_1[1] , \wRegOut_3_1[0] 
        }), .Enable1(\wRegEnTop_3_1[0] ), .Enable2(\wRegEnBot_3_1[0] ), .In1({
        \wRegInTop_3_1[31] , \wRegInTop_3_1[30] , \wRegInTop_3_1[29] , 
        \wRegInTop_3_1[28] , \wRegInTop_3_1[27] , \wRegInTop_3_1[26] , 
        \wRegInTop_3_1[25] , \wRegInTop_3_1[24] , \wRegInTop_3_1[23] , 
        \wRegInTop_3_1[22] , \wRegInTop_3_1[21] , \wRegInTop_3_1[20] , 
        \wRegInTop_3_1[19] , \wRegInTop_3_1[18] , \wRegInTop_3_1[17] , 
        \wRegInTop_3_1[16] , \wRegInTop_3_1[15] , \wRegInTop_3_1[14] , 
        \wRegInTop_3_1[13] , \wRegInTop_3_1[12] , \wRegInTop_3_1[11] , 
        \wRegInTop_3_1[10] , \wRegInTop_3_1[9] , \wRegInTop_3_1[8] , 
        \wRegInTop_3_1[7] , \wRegInTop_3_1[6] , \wRegInTop_3_1[5] , 
        \wRegInTop_3_1[4] , \wRegInTop_3_1[3] , \wRegInTop_3_1[2] , 
        \wRegInTop_3_1[1] , \wRegInTop_3_1[0] }), .In2({\wRegInBot_3_1[31] , 
        \wRegInBot_3_1[30] , \wRegInBot_3_1[29] , \wRegInBot_3_1[28] , 
        \wRegInBot_3_1[27] , \wRegInBot_3_1[26] , \wRegInBot_3_1[25] , 
        \wRegInBot_3_1[24] , \wRegInBot_3_1[23] , \wRegInBot_3_1[22] , 
        \wRegInBot_3_1[21] , \wRegInBot_3_1[20] , \wRegInBot_3_1[19] , 
        \wRegInBot_3_1[18] , \wRegInBot_3_1[17] , \wRegInBot_3_1[16] , 
        \wRegInBot_3_1[15] , \wRegInBot_3_1[14] , \wRegInBot_3_1[13] , 
        \wRegInBot_3_1[12] , \wRegInBot_3_1[11] , \wRegInBot_3_1[10] , 
        \wRegInBot_3_1[9] , \wRegInBot_3_1[8] , \wRegInBot_3_1[7] , 
        \wRegInBot_3_1[6] , \wRegInBot_3_1[5] , \wRegInBot_3_1[4] , 
        \wRegInBot_3_1[3] , \wRegInBot_3_1[2] , \wRegInBot_3_1[1] , 
        \wRegInBot_3_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink14[31] , \ScanLink14[30] , \ScanLink14[29] , 
        \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , \ScanLink14[25] , 
        \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , \ScanLink14[21] , 
        \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , \ScanLink14[17] , 
        \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , \ScanLink14[13] , 
        \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , \ScanLink14[9] , 
        \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , \ScanLink14[5] , 
        \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , \ScanLink14[1] , 
        \ScanLink14[0] }), .ScanOut({\ScanLink13[31] , \ScanLink13[30] , 
        \ScanLink13[29] , \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , 
        \ScanLink13[25] , \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , 
        \ScanLink13[21] , \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , 
        \ScanLink13[17] , \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , 
        \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , 
        \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , 
        \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , 
        \ScanLink13[1] , \ScanLink13[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_6[31] , \wRegOut_3_6[30] , \wRegOut_3_6[29] , 
        \wRegOut_3_6[28] , \wRegOut_3_6[27] , \wRegOut_3_6[26] , 
        \wRegOut_3_6[25] , \wRegOut_3_6[24] , \wRegOut_3_6[23] , 
        \wRegOut_3_6[22] , \wRegOut_3_6[21] , \wRegOut_3_6[20] , 
        \wRegOut_3_6[19] , \wRegOut_3_6[18] , \wRegOut_3_6[17] , 
        \wRegOut_3_6[16] , \wRegOut_3_6[15] , \wRegOut_3_6[14] , 
        \wRegOut_3_6[13] , \wRegOut_3_6[12] , \wRegOut_3_6[11] , 
        \wRegOut_3_6[10] , \wRegOut_3_6[9] , \wRegOut_3_6[8] , 
        \wRegOut_3_6[7] , \wRegOut_3_6[6] , \wRegOut_3_6[5] , \wRegOut_3_6[4] , 
        \wRegOut_3_6[3] , \wRegOut_3_6[2] , \wRegOut_3_6[1] , \wRegOut_3_6[0] 
        }), .Enable1(\wRegEnTop_3_6[0] ), .Enable2(\wRegEnBot_3_6[0] ), .In1({
        \wRegInTop_3_6[31] , \wRegInTop_3_6[30] , \wRegInTop_3_6[29] , 
        \wRegInTop_3_6[28] , \wRegInTop_3_6[27] , \wRegInTop_3_6[26] , 
        \wRegInTop_3_6[25] , \wRegInTop_3_6[24] , \wRegInTop_3_6[23] , 
        \wRegInTop_3_6[22] , \wRegInTop_3_6[21] , \wRegInTop_3_6[20] , 
        \wRegInTop_3_6[19] , \wRegInTop_3_6[18] , \wRegInTop_3_6[17] , 
        \wRegInTop_3_6[16] , \wRegInTop_3_6[15] , \wRegInTop_3_6[14] , 
        \wRegInTop_3_6[13] , \wRegInTop_3_6[12] , \wRegInTop_3_6[11] , 
        \wRegInTop_3_6[10] , \wRegInTop_3_6[9] , \wRegInTop_3_6[8] , 
        \wRegInTop_3_6[7] , \wRegInTop_3_6[6] , \wRegInTop_3_6[5] , 
        \wRegInTop_3_6[4] , \wRegInTop_3_6[3] , \wRegInTop_3_6[2] , 
        \wRegInTop_3_6[1] , \wRegInTop_3_6[0] }), .In2({\wRegInBot_3_6[31] , 
        \wRegInBot_3_6[30] , \wRegInBot_3_6[29] , \wRegInBot_3_6[28] , 
        \wRegInBot_3_6[27] , \wRegInBot_3_6[26] , \wRegInBot_3_6[25] , 
        \wRegInBot_3_6[24] , \wRegInBot_3_6[23] , \wRegInBot_3_6[22] , 
        \wRegInBot_3_6[21] , \wRegInBot_3_6[20] , \wRegInBot_3_6[19] , 
        \wRegInBot_3_6[18] , \wRegInBot_3_6[17] , \wRegInBot_3_6[16] , 
        \wRegInBot_3_6[15] , \wRegInBot_3_6[14] , \wRegInBot_3_6[13] , 
        \wRegInBot_3_6[12] , \wRegInBot_3_6[11] , \wRegInBot_3_6[10] , 
        \wRegInBot_3_6[9] , \wRegInBot_3_6[8] , \wRegInBot_3_6[7] , 
        \wRegInBot_3_6[6] , \wRegInBot_3_6[5] , \wRegInBot_3_6[4] , 
        \wRegInBot_3_6[3] , \wRegInBot_3_6[2] , \wRegInBot_3_6[1] , 
        \wRegInBot_3_6[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink29[31] , \ScanLink29[30] , \ScanLink29[29] , 
        \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , \ScanLink29[25] , 
        \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , \ScanLink29[21] , 
        \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , \ScanLink29[17] , 
        \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , \ScanLink29[13] , 
        \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , \ScanLink29[9] , 
        \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , \ScanLink29[5] , 
        \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , \ScanLink29[1] , 
        \ScanLink29[0] }), .ScanOut({\ScanLink28[31] , \ScanLink28[30] , 
        \ScanLink28[29] , \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , 
        \ScanLink28[25] , \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , 
        \ScanLink28[21] , \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , 
        \ScanLink28[17] , \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , 
        \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , 
        \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , 
        \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , 
        \ScanLink28[1] , \ScanLink28[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_13[31] , \wRegOut_4_13[30] , 
        \wRegOut_4_13[29] , \wRegOut_4_13[28] , \wRegOut_4_13[27] , 
        \wRegOut_4_13[26] , \wRegOut_4_13[25] , \wRegOut_4_13[24] , 
        \wRegOut_4_13[23] , \wRegOut_4_13[22] , \wRegOut_4_13[21] , 
        \wRegOut_4_13[20] , \wRegOut_4_13[19] , \wRegOut_4_13[18] , 
        \wRegOut_4_13[17] , \wRegOut_4_13[16] , \wRegOut_4_13[15] , 
        \wRegOut_4_13[14] , \wRegOut_4_13[13] , \wRegOut_4_13[12] , 
        \wRegOut_4_13[11] , \wRegOut_4_13[10] , \wRegOut_4_13[9] , 
        \wRegOut_4_13[8] , \wRegOut_4_13[7] , \wRegOut_4_13[6] , 
        \wRegOut_4_13[5] , \wRegOut_4_13[4] , \wRegOut_4_13[3] , 
        \wRegOut_4_13[2] , \wRegOut_4_13[1] , \wRegOut_4_13[0] }), .Enable1(
        \wRegEnTop_4_13[0] ), .Enable2(\wRegEnBot_4_13[0] ), .In1({
        \wRegInTop_4_13[31] , \wRegInTop_4_13[30] , \wRegInTop_4_13[29] , 
        \wRegInTop_4_13[28] , \wRegInTop_4_13[27] , \wRegInTop_4_13[26] , 
        \wRegInTop_4_13[25] , \wRegInTop_4_13[24] , \wRegInTop_4_13[23] , 
        \wRegInTop_4_13[22] , \wRegInTop_4_13[21] , \wRegInTop_4_13[20] , 
        \wRegInTop_4_13[19] , \wRegInTop_4_13[18] , \wRegInTop_4_13[17] , 
        \wRegInTop_4_13[16] , \wRegInTop_4_13[15] , \wRegInTop_4_13[14] , 
        \wRegInTop_4_13[13] , \wRegInTop_4_13[12] , \wRegInTop_4_13[11] , 
        \wRegInTop_4_13[10] , \wRegInTop_4_13[9] , \wRegInTop_4_13[8] , 
        \wRegInTop_4_13[7] , \wRegInTop_4_13[6] , \wRegInTop_4_13[5] , 
        \wRegInTop_4_13[4] , \wRegInTop_4_13[3] , \wRegInTop_4_13[2] , 
        \wRegInTop_4_13[1] , \wRegInTop_4_13[0] }), .In2({\wRegInBot_4_13[31] , 
        \wRegInBot_4_13[30] , \wRegInBot_4_13[29] , \wRegInBot_4_13[28] , 
        \wRegInBot_4_13[27] , \wRegInBot_4_13[26] , \wRegInBot_4_13[25] , 
        \wRegInBot_4_13[24] , \wRegInBot_4_13[23] , \wRegInBot_4_13[22] , 
        \wRegInBot_4_13[21] , \wRegInBot_4_13[20] , \wRegInBot_4_13[19] , 
        \wRegInBot_4_13[18] , \wRegInBot_4_13[17] , \wRegInBot_4_13[16] , 
        \wRegInBot_4_13[15] , \wRegInBot_4_13[14] , \wRegInBot_4_13[13] , 
        \wRegInBot_4_13[12] , \wRegInBot_4_13[11] , \wRegInBot_4_13[10] , 
        \wRegInBot_4_13[9] , \wRegInBot_4_13[8] , \wRegInBot_4_13[7] , 
        \wRegInBot_4_13[6] , \wRegInBot_4_13[5] , \wRegInBot_4_13[4] , 
        \wRegInBot_4_13[3] , \wRegInBot_4_13[2] , \wRegInBot_4_13[1] , 
        \wRegInBot_4_13[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_22 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink86[31] , \ScanLink86[30] , \ScanLink86[29] , 
        \ScanLink86[28] , \ScanLink86[27] , \ScanLink86[26] , \ScanLink86[25] , 
        \ScanLink86[24] , \ScanLink86[23] , \ScanLink86[22] , \ScanLink86[21] , 
        \ScanLink86[20] , \ScanLink86[19] , \ScanLink86[18] , \ScanLink86[17] , 
        \ScanLink86[16] , \ScanLink86[15] , \ScanLink86[14] , \ScanLink86[13] , 
        \ScanLink86[12] , \ScanLink86[11] , \ScanLink86[10] , \ScanLink86[9] , 
        \ScanLink86[8] , \ScanLink86[7] , \ScanLink86[6] , \ScanLink86[5] , 
        \ScanLink86[4] , \ScanLink86[3] , \ScanLink86[2] , \ScanLink86[1] , 
        \ScanLink86[0] }), .ScanOut({\ScanLink85[31] , \ScanLink85[30] , 
        \ScanLink85[29] , \ScanLink85[28] , \ScanLink85[27] , \ScanLink85[26] , 
        \ScanLink85[25] , \ScanLink85[24] , \ScanLink85[23] , \ScanLink85[22] , 
        \ScanLink85[21] , \ScanLink85[20] , \ScanLink85[19] , \ScanLink85[18] , 
        \ScanLink85[17] , \ScanLink85[16] , \ScanLink85[15] , \ScanLink85[14] , 
        \ScanLink85[13] , \ScanLink85[12] , \ScanLink85[11] , \ScanLink85[10] , 
        \ScanLink85[9] , \ScanLink85[8] , \ScanLink85[7] , \ScanLink85[6] , 
        \ScanLink85[5] , \ScanLink85[4] , \ScanLink85[3] , \ScanLink85[2] , 
        \ScanLink85[1] , \ScanLink85[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_22[31] , \wRegOut_6_22[30] , 
        \wRegOut_6_22[29] , \wRegOut_6_22[28] , \wRegOut_6_22[27] , 
        \wRegOut_6_22[26] , \wRegOut_6_22[25] , \wRegOut_6_22[24] , 
        \wRegOut_6_22[23] , \wRegOut_6_22[22] , \wRegOut_6_22[21] , 
        \wRegOut_6_22[20] , \wRegOut_6_22[19] , \wRegOut_6_22[18] , 
        \wRegOut_6_22[17] , \wRegOut_6_22[16] , \wRegOut_6_22[15] , 
        \wRegOut_6_22[14] , \wRegOut_6_22[13] , \wRegOut_6_22[12] , 
        \wRegOut_6_22[11] , \wRegOut_6_22[10] , \wRegOut_6_22[9] , 
        \wRegOut_6_22[8] , \wRegOut_6_22[7] , \wRegOut_6_22[6] , 
        \wRegOut_6_22[5] , \wRegOut_6_22[4] , \wRegOut_6_22[3] , 
        \wRegOut_6_22[2] , \wRegOut_6_22[1] , \wRegOut_6_22[0] }), .Enable1(
        \wRegEnTop_6_22[0] ), .Enable2(\wRegEnBot_6_22[0] ), .In1({
        \wRegInTop_6_22[31] , \wRegInTop_6_22[30] , \wRegInTop_6_22[29] , 
        \wRegInTop_6_22[28] , \wRegInTop_6_22[27] , \wRegInTop_6_22[26] , 
        \wRegInTop_6_22[25] , \wRegInTop_6_22[24] , \wRegInTop_6_22[23] , 
        \wRegInTop_6_22[22] , \wRegInTop_6_22[21] , \wRegInTop_6_22[20] , 
        \wRegInTop_6_22[19] , \wRegInTop_6_22[18] , \wRegInTop_6_22[17] , 
        \wRegInTop_6_22[16] , \wRegInTop_6_22[15] , \wRegInTop_6_22[14] , 
        \wRegInTop_6_22[13] , \wRegInTop_6_22[12] , \wRegInTop_6_22[11] , 
        \wRegInTop_6_22[10] , \wRegInTop_6_22[9] , \wRegInTop_6_22[8] , 
        \wRegInTop_6_22[7] , \wRegInTop_6_22[6] , \wRegInTop_6_22[5] , 
        \wRegInTop_6_22[4] , \wRegInTop_6_22[3] , \wRegInTop_6_22[2] , 
        \wRegInTop_6_22[1] , \wRegInTop_6_22[0] }), .In2({\wRegInBot_6_22[31] , 
        \wRegInBot_6_22[30] , \wRegInBot_6_22[29] , \wRegInBot_6_22[28] , 
        \wRegInBot_6_22[27] , \wRegInBot_6_22[26] , \wRegInBot_6_22[25] , 
        \wRegInBot_6_22[24] , \wRegInBot_6_22[23] , \wRegInBot_6_22[22] , 
        \wRegInBot_6_22[21] , \wRegInBot_6_22[20] , \wRegInBot_6_22[19] , 
        \wRegInBot_6_22[18] , \wRegInBot_6_22[17] , \wRegInBot_6_22[16] , 
        \wRegInBot_6_22[15] , \wRegInBot_6_22[14] , \wRegInBot_6_22[13] , 
        \wRegInBot_6_22[12] , \wRegInBot_6_22[11] , \wRegInBot_6_22[10] , 
        \wRegInBot_6_22[9] , \wRegInBot_6_22[8] , \wRegInBot_6_22[7] , 
        \wRegInBot_6_22[6] , \wRegInBot_6_22[5] , \wRegInBot_6_22[4] , 
        \wRegInBot_6_22[3] , \wRegInBot_6_22[2] , \wRegInBot_6_22[1] , 
        \wRegInBot_6_22[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_56 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink184[31] , \ScanLink184[30] , \ScanLink184[29] , 
        \ScanLink184[28] , \ScanLink184[27] , \ScanLink184[26] , 
        \ScanLink184[25] , \ScanLink184[24] , \ScanLink184[23] , 
        \ScanLink184[22] , \ScanLink184[21] , \ScanLink184[20] , 
        \ScanLink184[19] , \ScanLink184[18] , \ScanLink184[17] , 
        \ScanLink184[16] , \ScanLink184[15] , \ScanLink184[14] , 
        \ScanLink184[13] , \ScanLink184[12] , \ScanLink184[11] , 
        \ScanLink184[10] , \ScanLink184[9] , \ScanLink184[8] , 
        \ScanLink184[7] , \ScanLink184[6] , \ScanLink184[5] , \ScanLink184[4] , 
        \ScanLink184[3] , \ScanLink184[2] , \ScanLink184[1] , \ScanLink184[0] 
        }), .ScanOut({\ScanLink183[31] , \ScanLink183[30] , \ScanLink183[29] , 
        \ScanLink183[28] , \ScanLink183[27] , \ScanLink183[26] , 
        \ScanLink183[25] , \ScanLink183[24] , \ScanLink183[23] , 
        \ScanLink183[22] , \ScanLink183[21] , \ScanLink183[20] , 
        \ScanLink183[19] , \ScanLink183[18] , \ScanLink183[17] , 
        \ScanLink183[16] , \ScanLink183[15] , \ScanLink183[14] , 
        \ScanLink183[13] , \ScanLink183[12] , \ScanLink183[11] , 
        \ScanLink183[10] , \ScanLink183[9] , \ScanLink183[8] , 
        \ScanLink183[7] , \ScanLink183[6] , \ScanLink183[5] , \ScanLink183[4] , 
        \ScanLink183[3] , \ScanLink183[2] , \ScanLink183[1] , \ScanLink183[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_56[31] , 
        \wRegOut_7_56[30] , \wRegOut_7_56[29] , \wRegOut_7_56[28] , 
        \wRegOut_7_56[27] , \wRegOut_7_56[26] , \wRegOut_7_56[25] , 
        \wRegOut_7_56[24] , \wRegOut_7_56[23] , \wRegOut_7_56[22] , 
        \wRegOut_7_56[21] , \wRegOut_7_56[20] , \wRegOut_7_56[19] , 
        \wRegOut_7_56[18] , \wRegOut_7_56[17] , \wRegOut_7_56[16] , 
        \wRegOut_7_56[15] , \wRegOut_7_56[14] , \wRegOut_7_56[13] , 
        \wRegOut_7_56[12] , \wRegOut_7_56[11] , \wRegOut_7_56[10] , 
        \wRegOut_7_56[9] , \wRegOut_7_56[8] , \wRegOut_7_56[7] , 
        \wRegOut_7_56[6] , \wRegOut_7_56[5] , \wRegOut_7_56[4] , 
        \wRegOut_7_56[3] , \wRegOut_7_56[2] , \wRegOut_7_56[1] , 
        \wRegOut_7_56[0] }), .Enable1(\wRegEnTop_7_56[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_56[31] , \wRegInTop_7_56[30] , \wRegInTop_7_56[29] , 
        \wRegInTop_7_56[28] , \wRegInTop_7_56[27] , \wRegInTop_7_56[26] , 
        \wRegInTop_7_56[25] , \wRegInTop_7_56[24] , \wRegInTop_7_56[23] , 
        \wRegInTop_7_56[22] , \wRegInTop_7_56[21] , \wRegInTop_7_56[20] , 
        \wRegInTop_7_56[19] , \wRegInTop_7_56[18] , \wRegInTop_7_56[17] , 
        \wRegInTop_7_56[16] , \wRegInTop_7_56[15] , \wRegInTop_7_56[14] , 
        \wRegInTop_7_56[13] , \wRegInTop_7_56[12] , \wRegInTop_7_56[11] , 
        \wRegInTop_7_56[10] , \wRegInTop_7_56[9] , \wRegInTop_7_56[8] , 
        \wRegInTop_7_56[7] , \wRegInTop_7_56[6] , \wRegInTop_7_56[5] , 
        \wRegInTop_7_56[4] , \wRegInTop_7_56[3] , \wRegInTop_7_56[2] , 
        \wRegInTop_7_56[1] , \wRegInTop_7_56[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_38 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink166[31] , \ScanLink166[30] , \ScanLink166[29] , 
        \ScanLink166[28] , \ScanLink166[27] , \ScanLink166[26] , 
        \ScanLink166[25] , \ScanLink166[24] , \ScanLink166[23] , 
        \ScanLink166[22] , \ScanLink166[21] , \ScanLink166[20] , 
        \ScanLink166[19] , \ScanLink166[18] , \ScanLink166[17] , 
        \ScanLink166[16] , \ScanLink166[15] , \ScanLink166[14] , 
        \ScanLink166[13] , \ScanLink166[12] , \ScanLink166[11] , 
        \ScanLink166[10] , \ScanLink166[9] , \ScanLink166[8] , 
        \ScanLink166[7] , \ScanLink166[6] , \ScanLink166[5] , \ScanLink166[4] , 
        \ScanLink166[3] , \ScanLink166[2] , \ScanLink166[1] , \ScanLink166[0] 
        }), .ScanOut({\ScanLink165[31] , \ScanLink165[30] , \ScanLink165[29] , 
        \ScanLink165[28] , \ScanLink165[27] , \ScanLink165[26] , 
        \ScanLink165[25] , \ScanLink165[24] , \ScanLink165[23] , 
        \ScanLink165[22] , \ScanLink165[21] , \ScanLink165[20] , 
        \ScanLink165[19] , \ScanLink165[18] , \ScanLink165[17] , 
        \ScanLink165[16] , \ScanLink165[15] , \ScanLink165[14] , 
        \ScanLink165[13] , \ScanLink165[12] , \ScanLink165[11] , 
        \ScanLink165[10] , \ScanLink165[9] , \ScanLink165[8] , 
        \ScanLink165[7] , \ScanLink165[6] , \ScanLink165[5] , \ScanLink165[4] , 
        \ScanLink165[3] , \ScanLink165[2] , \ScanLink165[1] , \ScanLink165[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_38[31] , 
        \wRegOut_7_38[30] , \wRegOut_7_38[29] , \wRegOut_7_38[28] , 
        \wRegOut_7_38[27] , \wRegOut_7_38[26] , \wRegOut_7_38[25] , 
        \wRegOut_7_38[24] , \wRegOut_7_38[23] , \wRegOut_7_38[22] , 
        \wRegOut_7_38[21] , \wRegOut_7_38[20] , \wRegOut_7_38[19] , 
        \wRegOut_7_38[18] , \wRegOut_7_38[17] , \wRegOut_7_38[16] , 
        \wRegOut_7_38[15] , \wRegOut_7_38[14] , \wRegOut_7_38[13] , 
        \wRegOut_7_38[12] , \wRegOut_7_38[11] , \wRegOut_7_38[10] , 
        \wRegOut_7_38[9] , \wRegOut_7_38[8] , \wRegOut_7_38[7] , 
        \wRegOut_7_38[6] , \wRegOut_7_38[5] , \wRegOut_7_38[4] , 
        \wRegOut_7_38[3] , \wRegOut_7_38[2] , \wRegOut_7_38[1] , 
        \wRegOut_7_38[0] }), .Enable1(\wRegEnTop_7_38[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_38[31] , \wRegInTop_7_38[30] , \wRegInTop_7_38[29] , 
        \wRegInTop_7_38[28] , \wRegInTop_7_38[27] , \wRegInTop_7_38[26] , 
        \wRegInTop_7_38[25] , \wRegInTop_7_38[24] , \wRegInTop_7_38[23] , 
        \wRegInTop_7_38[22] , \wRegInTop_7_38[21] , \wRegInTop_7_38[20] , 
        \wRegInTop_7_38[19] , \wRegInTop_7_38[18] , \wRegInTop_7_38[17] , 
        \wRegInTop_7_38[16] , \wRegInTop_7_38[15] , \wRegInTop_7_38[14] , 
        \wRegInTop_7_38[13] , \wRegInTop_7_38[12] , \wRegInTop_7_38[11] , 
        \wRegInTop_7_38[10] , \wRegInTop_7_38[9] , \wRegInTop_7_38[8] , 
        \wRegInTop_7_38[7] , \wRegInTop_7_38[6] , \wRegInTop_7_38[5] , 
        \wRegInTop_7_38[4] , \wRegInTop_7_38[3] , \wRegInTop_7_38[2] , 
        \wRegInTop_7_38[1] , \wRegInTop_7_38[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_94 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink222[31] , \ScanLink222[30] , \ScanLink222[29] , 
        \ScanLink222[28] , \ScanLink222[27] , \ScanLink222[26] , 
        \ScanLink222[25] , \ScanLink222[24] , \ScanLink222[23] , 
        \ScanLink222[22] , \ScanLink222[21] , \ScanLink222[20] , 
        \ScanLink222[19] , \ScanLink222[18] , \ScanLink222[17] , 
        \ScanLink222[16] , \ScanLink222[15] , \ScanLink222[14] , 
        \ScanLink222[13] , \ScanLink222[12] , \ScanLink222[11] , 
        \ScanLink222[10] , \ScanLink222[9] , \ScanLink222[8] , 
        \ScanLink222[7] , \ScanLink222[6] , \ScanLink222[5] , \ScanLink222[4] , 
        \ScanLink222[3] , \ScanLink222[2] , \ScanLink222[1] , \ScanLink222[0] 
        }), .ScanOut({\ScanLink221[31] , \ScanLink221[30] , \ScanLink221[29] , 
        \ScanLink221[28] , \ScanLink221[27] , \ScanLink221[26] , 
        \ScanLink221[25] , \ScanLink221[24] , \ScanLink221[23] , 
        \ScanLink221[22] , \ScanLink221[21] , \ScanLink221[20] , 
        \ScanLink221[19] , \ScanLink221[18] , \ScanLink221[17] , 
        \ScanLink221[16] , \ScanLink221[15] , \ScanLink221[14] , 
        \ScanLink221[13] , \ScanLink221[12] , \ScanLink221[11] , 
        \ScanLink221[10] , \ScanLink221[9] , \ScanLink221[8] , 
        \ScanLink221[7] , \ScanLink221[6] , \ScanLink221[5] , \ScanLink221[4] , 
        \ScanLink221[3] , \ScanLink221[2] , \ScanLink221[1] , \ScanLink221[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_94[31] , 
        \wRegOut_7_94[30] , \wRegOut_7_94[29] , \wRegOut_7_94[28] , 
        \wRegOut_7_94[27] , \wRegOut_7_94[26] , \wRegOut_7_94[25] , 
        \wRegOut_7_94[24] , \wRegOut_7_94[23] , \wRegOut_7_94[22] , 
        \wRegOut_7_94[21] , \wRegOut_7_94[20] , \wRegOut_7_94[19] , 
        \wRegOut_7_94[18] , \wRegOut_7_94[17] , \wRegOut_7_94[16] , 
        \wRegOut_7_94[15] , \wRegOut_7_94[14] , \wRegOut_7_94[13] , 
        \wRegOut_7_94[12] , \wRegOut_7_94[11] , \wRegOut_7_94[10] , 
        \wRegOut_7_94[9] , \wRegOut_7_94[8] , \wRegOut_7_94[7] , 
        \wRegOut_7_94[6] , \wRegOut_7_94[5] , \wRegOut_7_94[4] , 
        \wRegOut_7_94[3] , \wRegOut_7_94[2] , \wRegOut_7_94[1] , 
        \wRegOut_7_94[0] }), .Enable1(\wRegEnTop_7_94[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_94[31] , \wRegInTop_7_94[30] , \wRegInTop_7_94[29] , 
        \wRegInTop_7_94[28] , \wRegInTop_7_94[27] , \wRegInTop_7_94[26] , 
        \wRegInTop_7_94[25] , \wRegInTop_7_94[24] , \wRegInTop_7_94[23] , 
        \wRegInTop_7_94[22] , \wRegInTop_7_94[21] , \wRegInTop_7_94[20] , 
        \wRegInTop_7_94[19] , \wRegInTop_7_94[18] , \wRegInTop_7_94[17] , 
        \wRegInTop_7_94[16] , \wRegInTop_7_94[15] , \wRegInTop_7_94[14] , 
        \wRegInTop_7_94[13] , \wRegInTop_7_94[12] , \wRegInTop_7_94[11] , 
        \wRegInTop_7_94[10] , \wRegInTop_7_94[9] , \wRegInTop_7_94[8] , 
        \wRegInTop_7_94[7] , \wRegInTop_7_94[6] , \wRegInTop_7_94[5] , 
        \wRegInTop_7_94[4] , \wRegInTop_7_94[3] , \wRegInTop_7_94[2] , 
        \wRegInTop_7_94[1] , \wRegInTop_7_94[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_43[0] ), .P_In({\wRegOut_6_43[31] , 
        \wRegOut_6_43[30] , \wRegOut_6_43[29] , \wRegOut_6_43[28] , 
        \wRegOut_6_43[27] , \wRegOut_6_43[26] , \wRegOut_6_43[25] , 
        \wRegOut_6_43[24] , \wRegOut_6_43[23] , \wRegOut_6_43[22] , 
        \wRegOut_6_43[21] , \wRegOut_6_43[20] , \wRegOut_6_43[19] , 
        \wRegOut_6_43[18] , \wRegOut_6_43[17] , \wRegOut_6_43[16] , 
        \wRegOut_6_43[15] , \wRegOut_6_43[14] , \wRegOut_6_43[13] , 
        \wRegOut_6_43[12] , \wRegOut_6_43[11] , \wRegOut_6_43[10] , 
        \wRegOut_6_43[9] , \wRegOut_6_43[8] , \wRegOut_6_43[7] , 
        \wRegOut_6_43[6] , \wRegOut_6_43[5] , \wRegOut_6_43[4] , 
        \wRegOut_6_43[3] , \wRegOut_6_43[2] , \wRegOut_6_43[1] , 
        \wRegOut_6_43[0] }), .P_Out({\wRegInBot_6_43[31] , 
        \wRegInBot_6_43[30] , \wRegInBot_6_43[29] , \wRegInBot_6_43[28] , 
        \wRegInBot_6_43[27] , \wRegInBot_6_43[26] , \wRegInBot_6_43[25] , 
        \wRegInBot_6_43[24] , \wRegInBot_6_43[23] , \wRegInBot_6_43[22] , 
        \wRegInBot_6_43[21] , \wRegInBot_6_43[20] , \wRegInBot_6_43[19] , 
        \wRegInBot_6_43[18] , \wRegInBot_6_43[17] , \wRegInBot_6_43[16] , 
        \wRegInBot_6_43[15] , \wRegInBot_6_43[14] , \wRegInBot_6_43[13] , 
        \wRegInBot_6_43[12] , \wRegInBot_6_43[11] , \wRegInBot_6_43[10] , 
        \wRegInBot_6_43[9] , \wRegInBot_6_43[8] , \wRegInBot_6_43[7] , 
        \wRegInBot_6_43[6] , \wRegInBot_6_43[5] , \wRegInBot_6_43[4] , 
        \wRegInBot_6_43[3] , \wRegInBot_6_43[2] , \wRegInBot_6_43[1] , 
        \wRegInBot_6_43[0] }), .L_WR(\wRegEnTop_7_86[0] ), .L_In({
        \wRegOut_7_86[31] , \wRegOut_7_86[30] , \wRegOut_7_86[29] , 
        \wRegOut_7_86[28] , \wRegOut_7_86[27] , \wRegOut_7_86[26] , 
        \wRegOut_7_86[25] , \wRegOut_7_86[24] , \wRegOut_7_86[23] , 
        \wRegOut_7_86[22] , \wRegOut_7_86[21] , \wRegOut_7_86[20] , 
        \wRegOut_7_86[19] , \wRegOut_7_86[18] , \wRegOut_7_86[17] , 
        \wRegOut_7_86[16] , \wRegOut_7_86[15] , \wRegOut_7_86[14] , 
        \wRegOut_7_86[13] , \wRegOut_7_86[12] , \wRegOut_7_86[11] , 
        \wRegOut_7_86[10] , \wRegOut_7_86[9] , \wRegOut_7_86[8] , 
        \wRegOut_7_86[7] , \wRegOut_7_86[6] , \wRegOut_7_86[5] , 
        \wRegOut_7_86[4] , \wRegOut_7_86[3] , \wRegOut_7_86[2] , 
        \wRegOut_7_86[1] , \wRegOut_7_86[0] }), .L_Out({\wRegInTop_7_86[31] , 
        \wRegInTop_7_86[30] , \wRegInTop_7_86[29] , \wRegInTop_7_86[28] , 
        \wRegInTop_7_86[27] , \wRegInTop_7_86[26] , \wRegInTop_7_86[25] , 
        \wRegInTop_7_86[24] , \wRegInTop_7_86[23] , \wRegInTop_7_86[22] , 
        \wRegInTop_7_86[21] , \wRegInTop_7_86[20] , \wRegInTop_7_86[19] , 
        \wRegInTop_7_86[18] , \wRegInTop_7_86[17] , \wRegInTop_7_86[16] , 
        \wRegInTop_7_86[15] , \wRegInTop_7_86[14] , \wRegInTop_7_86[13] , 
        \wRegInTop_7_86[12] , \wRegInTop_7_86[11] , \wRegInTop_7_86[10] , 
        \wRegInTop_7_86[9] , \wRegInTop_7_86[8] , \wRegInTop_7_86[7] , 
        \wRegInTop_7_86[6] , \wRegInTop_7_86[5] , \wRegInTop_7_86[4] , 
        \wRegInTop_7_86[3] , \wRegInTop_7_86[2] , \wRegInTop_7_86[1] , 
        \wRegInTop_7_86[0] }), .R_WR(\wRegEnTop_7_87[0] ), .R_In({
        \wRegOut_7_87[31] , \wRegOut_7_87[30] , \wRegOut_7_87[29] , 
        \wRegOut_7_87[28] , \wRegOut_7_87[27] , \wRegOut_7_87[26] , 
        \wRegOut_7_87[25] , \wRegOut_7_87[24] , \wRegOut_7_87[23] , 
        \wRegOut_7_87[22] , \wRegOut_7_87[21] , \wRegOut_7_87[20] , 
        \wRegOut_7_87[19] , \wRegOut_7_87[18] , \wRegOut_7_87[17] , 
        \wRegOut_7_87[16] , \wRegOut_7_87[15] , \wRegOut_7_87[14] , 
        \wRegOut_7_87[13] , \wRegOut_7_87[12] , \wRegOut_7_87[11] , 
        \wRegOut_7_87[10] , \wRegOut_7_87[9] , \wRegOut_7_87[8] , 
        \wRegOut_7_87[7] , \wRegOut_7_87[6] , \wRegOut_7_87[5] , 
        \wRegOut_7_87[4] , \wRegOut_7_87[3] , \wRegOut_7_87[2] , 
        \wRegOut_7_87[1] , \wRegOut_7_87[0] }), .R_Out({\wRegInTop_7_87[31] , 
        \wRegInTop_7_87[30] , \wRegInTop_7_87[29] , \wRegInTop_7_87[28] , 
        \wRegInTop_7_87[27] , \wRegInTop_7_87[26] , \wRegInTop_7_87[25] , 
        \wRegInTop_7_87[24] , \wRegInTop_7_87[23] , \wRegInTop_7_87[22] , 
        \wRegInTop_7_87[21] , \wRegInTop_7_87[20] , \wRegInTop_7_87[19] , 
        \wRegInTop_7_87[18] , \wRegInTop_7_87[17] , \wRegInTop_7_87[16] , 
        \wRegInTop_7_87[15] , \wRegInTop_7_87[14] , \wRegInTop_7_87[13] , 
        \wRegInTop_7_87[12] , \wRegInTop_7_87[11] , \wRegInTop_7_87[10] , 
        \wRegInTop_7_87[9] , \wRegInTop_7_87[8] , \wRegInTop_7_87[7] , 
        \wRegInTop_7_87[6] , \wRegInTop_7_87[5] , \wRegInTop_7_87[4] , 
        \wRegInTop_7_87[3] , \wRegInTop_7_87[2] , \wRegInTop_7_87[1] , 
        \wRegInTop_7_87[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_110 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink238[31] , \ScanLink238[30] , \ScanLink238[29] , 
        \ScanLink238[28] , \ScanLink238[27] , \ScanLink238[26] , 
        \ScanLink238[25] , \ScanLink238[24] , \ScanLink238[23] , 
        \ScanLink238[22] , \ScanLink238[21] , \ScanLink238[20] , 
        \ScanLink238[19] , \ScanLink238[18] , \ScanLink238[17] , 
        \ScanLink238[16] , \ScanLink238[15] , \ScanLink238[14] , 
        \ScanLink238[13] , \ScanLink238[12] , \ScanLink238[11] , 
        \ScanLink238[10] , \ScanLink238[9] , \ScanLink238[8] , 
        \ScanLink238[7] , \ScanLink238[6] , \ScanLink238[5] , \ScanLink238[4] , 
        \ScanLink238[3] , \ScanLink238[2] , \ScanLink238[1] , \ScanLink238[0] 
        }), .ScanOut({\ScanLink237[31] , \ScanLink237[30] , \ScanLink237[29] , 
        \ScanLink237[28] , \ScanLink237[27] , \ScanLink237[26] , 
        \ScanLink237[25] , \ScanLink237[24] , \ScanLink237[23] , 
        \ScanLink237[22] , \ScanLink237[21] , \ScanLink237[20] , 
        \ScanLink237[19] , \ScanLink237[18] , \ScanLink237[17] , 
        \ScanLink237[16] , \ScanLink237[15] , \ScanLink237[14] , 
        \ScanLink237[13] , \ScanLink237[12] , \ScanLink237[11] , 
        \ScanLink237[10] , \ScanLink237[9] , \ScanLink237[8] , 
        \ScanLink237[7] , \ScanLink237[6] , \ScanLink237[5] , \ScanLink237[4] , 
        \ScanLink237[3] , \ScanLink237[2] , \ScanLink237[1] , \ScanLink237[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_110[31] , 
        \wRegOut_7_110[30] , \wRegOut_7_110[29] , \wRegOut_7_110[28] , 
        \wRegOut_7_110[27] , \wRegOut_7_110[26] , \wRegOut_7_110[25] , 
        \wRegOut_7_110[24] , \wRegOut_7_110[23] , \wRegOut_7_110[22] , 
        \wRegOut_7_110[21] , \wRegOut_7_110[20] , \wRegOut_7_110[19] , 
        \wRegOut_7_110[18] , \wRegOut_7_110[17] , \wRegOut_7_110[16] , 
        \wRegOut_7_110[15] , \wRegOut_7_110[14] , \wRegOut_7_110[13] , 
        \wRegOut_7_110[12] , \wRegOut_7_110[11] , \wRegOut_7_110[10] , 
        \wRegOut_7_110[9] , \wRegOut_7_110[8] , \wRegOut_7_110[7] , 
        \wRegOut_7_110[6] , \wRegOut_7_110[5] , \wRegOut_7_110[4] , 
        \wRegOut_7_110[3] , \wRegOut_7_110[2] , \wRegOut_7_110[1] , 
        \wRegOut_7_110[0] }), .Enable1(\wRegEnTop_7_110[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_110[31] , \wRegInTop_7_110[30] , 
        \wRegInTop_7_110[29] , \wRegInTop_7_110[28] , \wRegInTop_7_110[27] , 
        \wRegInTop_7_110[26] , \wRegInTop_7_110[25] , \wRegInTop_7_110[24] , 
        \wRegInTop_7_110[23] , \wRegInTop_7_110[22] , \wRegInTop_7_110[21] , 
        \wRegInTop_7_110[20] , \wRegInTop_7_110[19] , \wRegInTop_7_110[18] , 
        \wRegInTop_7_110[17] , \wRegInTop_7_110[16] , \wRegInTop_7_110[15] , 
        \wRegInTop_7_110[14] , \wRegInTop_7_110[13] , \wRegInTop_7_110[12] , 
        \wRegInTop_7_110[11] , \wRegInTop_7_110[10] , \wRegInTop_7_110[9] , 
        \wRegInTop_7_110[8] , \wRegInTop_7_110[7] , \wRegInTop_7_110[6] , 
        \wRegInTop_7_110[5] , \wRegInTop_7_110[4] , \wRegInTop_7_110[3] , 
        \wRegInTop_7_110[2] , \wRegInTop_7_110[1] , \wRegInTop_7_110[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_5[0] ), .P_In({\wRegOut_4_5[31] , 
        \wRegOut_4_5[30] , \wRegOut_4_5[29] , \wRegOut_4_5[28] , 
        \wRegOut_4_5[27] , \wRegOut_4_5[26] , \wRegOut_4_5[25] , 
        \wRegOut_4_5[24] , \wRegOut_4_5[23] , \wRegOut_4_5[22] , 
        \wRegOut_4_5[21] , \wRegOut_4_5[20] , \wRegOut_4_5[19] , 
        \wRegOut_4_5[18] , \wRegOut_4_5[17] , \wRegOut_4_5[16] , 
        \wRegOut_4_5[15] , \wRegOut_4_5[14] , \wRegOut_4_5[13] , 
        \wRegOut_4_5[12] , \wRegOut_4_5[11] , \wRegOut_4_5[10] , 
        \wRegOut_4_5[9] , \wRegOut_4_5[8] , \wRegOut_4_5[7] , \wRegOut_4_5[6] , 
        \wRegOut_4_5[5] , \wRegOut_4_5[4] , \wRegOut_4_5[3] , \wRegOut_4_5[2] , 
        \wRegOut_4_5[1] , \wRegOut_4_5[0] }), .P_Out({\wRegInBot_4_5[31] , 
        \wRegInBot_4_5[30] , \wRegInBot_4_5[29] , \wRegInBot_4_5[28] , 
        \wRegInBot_4_5[27] , \wRegInBot_4_5[26] , \wRegInBot_4_5[25] , 
        \wRegInBot_4_5[24] , \wRegInBot_4_5[23] , \wRegInBot_4_5[22] , 
        \wRegInBot_4_5[21] , \wRegInBot_4_5[20] , \wRegInBot_4_5[19] , 
        \wRegInBot_4_5[18] , \wRegInBot_4_5[17] , \wRegInBot_4_5[16] , 
        \wRegInBot_4_5[15] , \wRegInBot_4_5[14] , \wRegInBot_4_5[13] , 
        \wRegInBot_4_5[12] , \wRegInBot_4_5[11] , \wRegInBot_4_5[10] , 
        \wRegInBot_4_5[9] , \wRegInBot_4_5[8] , \wRegInBot_4_5[7] , 
        \wRegInBot_4_5[6] , \wRegInBot_4_5[5] , \wRegInBot_4_5[4] , 
        \wRegInBot_4_5[3] , \wRegInBot_4_5[2] , \wRegInBot_4_5[1] , 
        \wRegInBot_4_5[0] }), .L_WR(\wRegEnTop_5_10[0] ), .L_In({
        \wRegOut_5_10[31] , \wRegOut_5_10[30] , \wRegOut_5_10[29] , 
        \wRegOut_5_10[28] , \wRegOut_5_10[27] , \wRegOut_5_10[26] , 
        \wRegOut_5_10[25] , \wRegOut_5_10[24] , \wRegOut_5_10[23] , 
        \wRegOut_5_10[22] , \wRegOut_5_10[21] , \wRegOut_5_10[20] , 
        \wRegOut_5_10[19] , \wRegOut_5_10[18] , \wRegOut_5_10[17] , 
        \wRegOut_5_10[16] , \wRegOut_5_10[15] , \wRegOut_5_10[14] , 
        \wRegOut_5_10[13] , \wRegOut_5_10[12] , \wRegOut_5_10[11] , 
        \wRegOut_5_10[10] , \wRegOut_5_10[9] , \wRegOut_5_10[8] , 
        \wRegOut_5_10[7] , \wRegOut_5_10[6] , \wRegOut_5_10[5] , 
        \wRegOut_5_10[4] , \wRegOut_5_10[3] , \wRegOut_5_10[2] , 
        \wRegOut_5_10[1] , \wRegOut_5_10[0] }), .L_Out({\wRegInTop_5_10[31] , 
        \wRegInTop_5_10[30] , \wRegInTop_5_10[29] , \wRegInTop_5_10[28] , 
        \wRegInTop_5_10[27] , \wRegInTop_5_10[26] , \wRegInTop_5_10[25] , 
        \wRegInTop_5_10[24] , \wRegInTop_5_10[23] , \wRegInTop_5_10[22] , 
        \wRegInTop_5_10[21] , \wRegInTop_5_10[20] , \wRegInTop_5_10[19] , 
        \wRegInTop_5_10[18] , \wRegInTop_5_10[17] , \wRegInTop_5_10[16] , 
        \wRegInTop_5_10[15] , \wRegInTop_5_10[14] , \wRegInTop_5_10[13] , 
        \wRegInTop_5_10[12] , \wRegInTop_5_10[11] , \wRegInTop_5_10[10] , 
        \wRegInTop_5_10[9] , \wRegInTop_5_10[8] , \wRegInTop_5_10[7] , 
        \wRegInTop_5_10[6] , \wRegInTop_5_10[5] , \wRegInTop_5_10[4] , 
        \wRegInTop_5_10[3] , \wRegInTop_5_10[2] , \wRegInTop_5_10[1] , 
        \wRegInTop_5_10[0] }), .R_WR(\wRegEnTop_5_11[0] ), .R_In({
        \wRegOut_5_11[31] , \wRegOut_5_11[30] , \wRegOut_5_11[29] , 
        \wRegOut_5_11[28] , \wRegOut_5_11[27] , \wRegOut_5_11[26] , 
        \wRegOut_5_11[25] , \wRegOut_5_11[24] , \wRegOut_5_11[23] , 
        \wRegOut_5_11[22] , \wRegOut_5_11[21] , \wRegOut_5_11[20] , 
        \wRegOut_5_11[19] , \wRegOut_5_11[18] , \wRegOut_5_11[17] , 
        \wRegOut_5_11[16] , \wRegOut_5_11[15] , \wRegOut_5_11[14] , 
        \wRegOut_5_11[13] , \wRegOut_5_11[12] , \wRegOut_5_11[11] , 
        \wRegOut_5_11[10] , \wRegOut_5_11[9] , \wRegOut_5_11[8] , 
        \wRegOut_5_11[7] , \wRegOut_5_11[6] , \wRegOut_5_11[5] , 
        \wRegOut_5_11[4] , \wRegOut_5_11[3] , \wRegOut_5_11[2] , 
        \wRegOut_5_11[1] , \wRegOut_5_11[0] }), .R_Out({\wRegInTop_5_11[31] , 
        \wRegInTop_5_11[30] , \wRegInTop_5_11[29] , \wRegInTop_5_11[28] , 
        \wRegInTop_5_11[27] , \wRegInTop_5_11[26] , \wRegInTop_5_11[25] , 
        \wRegInTop_5_11[24] , \wRegInTop_5_11[23] , \wRegInTop_5_11[22] , 
        \wRegInTop_5_11[21] , \wRegInTop_5_11[20] , \wRegInTop_5_11[19] , 
        \wRegInTop_5_11[18] , \wRegInTop_5_11[17] , \wRegInTop_5_11[16] , 
        \wRegInTop_5_11[15] , \wRegInTop_5_11[14] , \wRegInTop_5_11[13] , 
        \wRegInTop_5_11[12] , \wRegInTop_5_11[11] , \wRegInTop_5_11[10] , 
        \wRegInTop_5_11[9] , \wRegInTop_5_11[8] , \wRegInTop_5_11[7] , 
        \wRegInTop_5_11[6] , \wRegInTop_5_11[5] , \wRegInTop_5_11[4] , 
        \wRegInTop_5_11[3] , \wRegInTop_5_11[2] , \wRegInTop_5_11[1] , 
        \wRegInTop_5_11[0] }) );
    BHeap_Node_WIDTH32 BHN_5_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_5[0] ), .P_In({\wRegOut_5_5[31] , 
        \wRegOut_5_5[30] , \wRegOut_5_5[29] , \wRegOut_5_5[28] , 
        \wRegOut_5_5[27] , \wRegOut_5_5[26] , \wRegOut_5_5[25] , 
        \wRegOut_5_5[24] , \wRegOut_5_5[23] , \wRegOut_5_5[22] , 
        \wRegOut_5_5[21] , \wRegOut_5_5[20] , \wRegOut_5_5[19] , 
        \wRegOut_5_5[18] , \wRegOut_5_5[17] , \wRegOut_5_5[16] , 
        \wRegOut_5_5[15] , \wRegOut_5_5[14] , \wRegOut_5_5[13] , 
        \wRegOut_5_5[12] , \wRegOut_5_5[11] , \wRegOut_5_5[10] , 
        \wRegOut_5_5[9] , \wRegOut_5_5[8] , \wRegOut_5_5[7] , \wRegOut_5_5[6] , 
        \wRegOut_5_5[5] , \wRegOut_5_5[4] , \wRegOut_5_5[3] , \wRegOut_5_5[2] , 
        \wRegOut_5_5[1] , \wRegOut_5_5[0] }), .P_Out({\wRegInBot_5_5[31] , 
        \wRegInBot_5_5[30] , \wRegInBot_5_5[29] , \wRegInBot_5_5[28] , 
        \wRegInBot_5_5[27] , \wRegInBot_5_5[26] , \wRegInBot_5_5[25] , 
        \wRegInBot_5_5[24] , \wRegInBot_5_5[23] , \wRegInBot_5_5[22] , 
        \wRegInBot_5_5[21] , \wRegInBot_5_5[20] , \wRegInBot_5_5[19] , 
        \wRegInBot_5_5[18] , \wRegInBot_5_5[17] , \wRegInBot_5_5[16] , 
        \wRegInBot_5_5[15] , \wRegInBot_5_5[14] , \wRegInBot_5_5[13] , 
        \wRegInBot_5_5[12] , \wRegInBot_5_5[11] , \wRegInBot_5_5[10] , 
        \wRegInBot_5_5[9] , \wRegInBot_5_5[8] , \wRegInBot_5_5[7] , 
        \wRegInBot_5_5[6] , \wRegInBot_5_5[5] , \wRegInBot_5_5[4] , 
        \wRegInBot_5_5[3] , \wRegInBot_5_5[2] , \wRegInBot_5_5[1] , 
        \wRegInBot_5_5[0] }), .L_WR(\wRegEnTop_6_10[0] ), .L_In({
        \wRegOut_6_10[31] , \wRegOut_6_10[30] , \wRegOut_6_10[29] , 
        \wRegOut_6_10[28] , \wRegOut_6_10[27] , \wRegOut_6_10[26] , 
        \wRegOut_6_10[25] , \wRegOut_6_10[24] , \wRegOut_6_10[23] , 
        \wRegOut_6_10[22] , \wRegOut_6_10[21] , \wRegOut_6_10[20] , 
        \wRegOut_6_10[19] , \wRegOut_6_10[18] , \wRegOut_6_10[17] , 
        \wRegOut_6_10[16] , \wRegOut_6_10[15] , \wRegOut_6_10[14] , 
        \wRegOut_6_10[13] , \wRegOut_6_10[12] , \wRegOut_6_10[11] , 
        \wRegOut_6_10[10] , \wRegOut_6_10[9] , \wRegOut_6_10[8] , 
        \wRegOut_6_10[7] , \wRegOut_6_10[6] , \wRegOut_6_10[5] , 
        \wRegOut_6_10[4] , \wRegOut_6_10[3] , \wRegOut_6_10[2] , 
        \wRegOut_6_10[1] , \wRegOut_6_10[0] }), .L_Out({\wRegInTop_6_10[31] , 
        \wRegInTop_6_10[30] , \wRegInTop_6_10[29] , \wRegInTop_6_10[28] , 
        \wRegInTop_6_10[27] , \wRegInTop_6_10[26] , \wRegInTop_6_10[25] , 
        \wRegInTop_6_10[24] , \wRegInTop_6_10[23] , \wRegInTop_6_10[22] , 
        \wRegInTop_6_10[21] , \wRegInTop_6_10[20] , \wRegInTop_6_10[19] , 
        \wRegInTop_6_10[18] , \wRegInTop_6_10[17] , \wRegInTop_6_10[16] , 
        \wRegInTop_6_10[15] , \wRegInTop_6_10[14] , \wRegInTop_6_10[13] , 
        \wRegInTop_6_10[12] , \wRegInTop_6_10[11] , \wRegInTop_6_10[10] , 
        \wRegInTop_6_10[9] , \wRegInTop_6_10[8] , \wRegInTop_6_10[7] , 
        \wRegInTop_6_10[6] , \wRegInTop_6_10[5] , \wRegInTop_6_10[4] , 
        \wRegInTop_6_10[3] , \wRegInTop_6_10[2] , \wRegInTop_6_10[1] , 
        \wRegInTop_6_10[0] }), .R_WR(\wRegEnTop_6_11[0] ), .R_In({
        \wRegOut_6_11[31] , \wRegOut_6_11[30] , \wRegOut_6_11[29] , 
        \wRegOut_6_11[28] , \wRegOut_6_11[27] , \wRegOut_6_11[26] , 
        \wRegOut_6_11[25] , \wRegOut_6_11[24] , \wRegOut_6_11[23] , 
        \wRegOut_6_11[22] , \wRegOut_6_11[21] , \wRegOut_6_11[20] , 
        \wRegOut_6_11[19] , \wRegOut_6_11[18] , \wRegOut_6_11[17] , 
        \wRegOut_6_11[16] , \wRegOut_6_11[15] , \wRegOut_6_11[14] , 
        \wRegOut_6_11[13] , \wRegOut_6_11[12] , \wRegOut_6_11[11] , 
        \wRegOut_6_11[10] , \wRegOut_6_11[9] , \wRegOut_6_11[8] , 
        \wRegOut_6_11[7] , \wRegOut_6_11[6] , \wRegOut_6_11[5] , 
        \wRegOut_6_11[4] , \wRegOut_6_11[3] , \wRegOut_6_11[2] , 
        \wRegOut_6_11[1] , \wRegOut_6_11[0] }), .R_Out({\wRegInTop_6_11[31] , 
        \wRegInTop_6_11[30] , \wRegInTop_6_11[29] , \wRegInTop_6_11[28] , 
        \wRegInTop_6_11[27] , \wRegInTop_6_11[26] , \wRegInTop_6_11[25] , 
        \wRegInTop_6_11[24] , \wRegInTop_6_11[23] , \wRegInTop_6_11[22] , 
        \wRegInTop_6_11[21] , \wRegInTop_6_11[20] , \wRegInTop_6_11[19] , 
        \wRegInTop_6_11[18] , \wRegInTop_6_11[17] , \wRegInTop_6_11[16] , 
        \wRegInTop_6_11[15] , \wRegInTop_6_11[14] , \wRegInTop_6_11[13] , 
        \wRegInTop_6_11[12] , \wRegInTop_6_11[11] , \wRegInTop_6_11[10] , 
        \wRegInTop_6_11[9] , \wRegInTop_6_11[8] , \wRegInTop_6_11[7] , 
        \wRegInTop_6_11[6] , \wRegInTop_6_11[5] , \wRegInTop_6_11[4] , 
        \wRegInTop_6_11[3] , \wRegInTop_6_11[2] , \wRegInTop_6_11[1] , 
        \wRegInTop_6_11[0] }) );
    BHeap_Node_WIDTH32 BHN_6_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_9[0] ), .P_In({\wRegOut_6_9[31] , 
        \wRegOut_6_9[30] , \wRegOut_6_9[29] , \wRegOut_6_9[28] , 
        \wRegOut_6_9[27] , \wRegOut_6_9[26] , \wRegOut_6_9[25] , 
        \wRegOut_6_9[24] , \wRegOut_6_9[23] , \wRegOut_6_9[22] , 
        \wRegOut_6_9[21] , \wRegOut_6_9[20] , \wRegOut_6_9[19] , 
        \wRegOut_6_9[18] , \wRegOut_6_9[17] , \wRegOut_6_9[16] , 
        \wRegOut_6_9[15] , \wRegOut_6_9[14] , \wRegOut_6_9[13] , 
        \wRegOut_6_9[12] , \wRegOut_6_9[11] , \wRegOut_6_9[10] , 
        \wRegOut_6_9[9] , \wRegOut_6_9[8] , \wRegOut_6_9[7] , \wRegOut_6_9[6] , 
        \wRegOut_6_9[5] , \wRegOut_6_9[4] , \wRegOut_6_9[3] , \wRegOut_6_9[2] , 
        \wRegOut_6_9[1] , \wRegOut_6_9[0] }), .P_Out({\wRegInBot_6_9[31] , 
        \wRegInBot_6_9[30] , \wRegInBot_6_9[29] , \wRegInBot_6_9[28] , 
        \wRegInBot_6_9[27] , \wRegInBot_6_9[26] , \wRegInBot_6_9[25] , 
        \wRegInBot_6_9[24] , \wRegInBot_6_9[23] , \wRegInBot_6_9[22] , 
        \wRegInBot_6_9[21] , \wRegInBot_6_9[20] , \wRegInBot_6_9[19] , 
        \wRegInBot_6_9[18] , \wRegInBot_6_9[17] , \wRegInBot_6_9[16] , 
        \wRegInBot_6_9[15] , \wRegInBot_6_9[14] , \wRegInBot_6_9[13] , 
        \wRegInBot_6_9[12] , \wRegInBot_6_9[11] , \wRegInBot_6_9[10] , 
        \wRegInBot_6_9[9] , \wRegInBot_6_9[8] , \wRegInBot_6_9[7] , 
        \wRegInBot_6_9[6] , \wRegInBot_6_9[5] , \wRegInBot_6_9[4] , 
        \wRegInBot_6_9[3] , \wRegInBot_6_9[2] , \wRegInBot_6_9[1] , 
        \wRegInBot_6_9[0] }), .L_WR(\wRegEnTop_7_18[0] ), .L_In({
        \wRegOut_7_18[31] , \wRegOut_7_18[30] , \wRegOut_7_18[29] , 
        \wRegOut_7_18[28] , \wRegOut_7_18[27] , \wRegOut_7_18[26] , 
        \wRegOut_7_18[25] , \wRegOut_7_18[24] , \wRegOut_7_18[23] , 
        \wRegOut_7_18[22] , \wRegOut_7_18[21] , \wRegOut_7_18[20] , 
        \wRegOut_7_18[19] , \wRegOut_7_18[18] , \wRegOut_7_18[17] , 
        \wRegOut_7_18[16] , \wRegOut_7_18[15] , \wRegOut_7_18[14] , 
        \wRegOut_7_18[13] , \wRegOut_7_18[12] , \wRegOut_7_18[11] , 
        \wRegOut_7_18[10] , \wRegOut_7_18[9] , \wRegOut_7_18[8] , 
        \wRegOut_7_18[7] , \wRegOut_7_18[6] , \wRegOut_7_18[5] , 
        \wRegOut_7_18[4] , \wRegOut_7_18[3] , \wRegOut_7_18[2] , 
        \wRegOut_7_18[1] , \wRegOut_7_18[0] }), .L_Out({\wRegInTop_7_18[31] , 
        \wRegInTop_7_18[30] , \wRegInTop_7_18[29] , \wRegInTop_7_18[28] , 
        \wRegInTop_7_18[27] , \wRegInTop_7_18[26] , \wRegInTop_7_18[25] , 
        \wRegInTop_7_18[24] , \wRegInTop_7_18[23] , \wRegInTop_7_18[22] , 
        \wRegInTop_7_18[21] , \wRegInTop_7_18[20] , \wRegInTop_7_18[19] , 
        \wRegInTop_7_18[18] , \wRegInTop_7_18[17] , \wRegInTop_7_18[16] , 
        \wRegInTop_7_18[15] , \wRegInTop_7_18[14] , \wRegInTop_7_18[13] , 
        \wRegInTop_7_18[12] , \wRegInTop_7_18[11] , \wRegInTop_7_18[10] , 
        \wRegInTop_7_18[9] , \wRegInTop_7_18[8] , \wRegInTop_7_18[7] , 
        \wRegInTop_7_18[6] , \wRegInTop_7_18[5] , \wRegInTop_7_18[4] , 
        \wRegInTop_7_18[3] , \wRegInTop_7_18[2] , \wRegInTop_7_18[1] , 
        \wRegInTop_7_18[0] }), .R_WR(\wRegEnTop_7_19[0] ), .R_In({
        \wRegOut_7_19[31] , \wRegOut_7_19[30] , \wRegOut_7_19[29] , 
        \wRegOut_7_19[28] , \wRegOut_7_19[27] , \wRegOut_7_19[26] , 
        \wRegOut_7_19[25] , \wRegOut_7_19[24] , \wRegOut_7_19[23] , 
        \wRegOut_7_19[22] , \wRegOut_7_19[21] , \wRegOut_7_19[20] , 
        \wRegOut_7_19[19] , \wRegOut_7_19[18] , \wRegOut_7_19[17] , 
        \wRegOut_7_19[16] , \wRegOut_7_19[15] , \wRegOut_7_19[14] , 
        \wRegOut_7_19[13] , \wRegOut_7_19[12] , \wRegOut_7_19[11] , 
        \wRegOut_7_19[10] , \wRegOut_7_19[9] , \wRegOut_7_19[8] , 
        \wRegOut_7_19[7] , \wRegOut_7_19[6] , \wRegOut_7_19[5] , 
        \wRegOut_7_19[4] , \wRegOut_7_19[3] , \wRegOut_7_19[2] , 
        \wRegOut_7_19[1] , \wRegOut_7_19[0] }), .R_Out({\wRegInTop_7_19[31] , 
        \wRegInTop_7_19[30] , \wRegInTop_7_19[29] , \wRegInTop_7_19[28] , 
        \wRegInTop_7_19[27] , \wRegInTop_7_19[26] , \wRegInTop_7_19[25] , 
        \wRegInTop_7_19[24] , \wRegInTop_7_19[23] , \wRegInTop_7_19[22] , 
        \wRegInTop_7_19[21] , \wRegInTop_7_19[20] , \wRegInTop_7_19[19] , 
        \wRegInTop_7_19[18] , \wRegInTop_7_19[17] , \wRegInTop_7_19[16] , 
        \wRegInTop_7_19[15] , \wRegInTop_7_19[14] , \wRegInTop_7_19[13] , 
        \wRegInTop_7_19[12] , \wRegInTop_7_19[11] , \wRegInTop_7_19[10] , 
        \wRegInTop_7_19[9] , \wRegInTop_7_19[8] , \wRegInTop_7_19[7] , 
        \wRegInTop_7_19[6] , \wRegInTop_7_19[5] , \wRegInTop_7_19[4] , 
        \wRegInTop_7_19[3] , \wRegInTop_7_19[2] , \wRegInTop_7_19[1] , 
        \wRegInTop_7_19[0] }) );
    BHeap_Node_WIDTH32 BHN_6_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_58[0] ), .P_In({\wRegOut_6_58[31] , 
        \wRegOut_6_58[30] , \wRegOut_6_58[29] , \wRegOut_6_58[28] , 
        \wRegOut_6_58[27] , \wRegOut_6_58[26] , \wRegOut_6_58[25] , 
        \wRegOut_6_58[24] , \wRegOut_6_58[23] , \wRegOut_6_58[22] , 
        \wRegOut_6_58[21] , \wRegOut_6_58[20] , \wRegOut_6_58[19] , 
        \wRegOut_6_58[18] , \wRegOut_6_58[17] , \wRegOut_6_58[16] , 
        \wRegOut_6_58[15] , \wRegOut_6_58[14] , \wRegOut_6_58[13] , 
        \wRegOut_6_58[12] , \wRegOut_6_58[11] , \wRegOut_6_58[10] , 
        \wRegOut_6_58[9] , \wRegOut_6_58[8] , \wRegOut_6_58[7] , 
        \wRegOut_6_58[6] , \wRegOut_6_58[5] , \wRegOut_6_58[4] , 
        \wRegOut_6_58[3] , \wRegOut_6_58[2] , \wRegOut_6_58[1] , 
        \wRegOut_6_58[0] }), .P_Out({\wRegInBot_6_58[31] , 
        \wRegInBot_6_58[30] , \wRegInBot_6_58[29] , \wRegInBot_6_58[28] , 
        \wRegInBot_6_58[27] , \wRegInBot_6_58[26] , \wRegInBot_6_58[25] , 
        \wRegInBot_6_58[24] , \wRegInBot_6_58[23] , \wRegInBot_6_58[22] , 
        \wRegInBot_6_58[21] , \wRegInBot_6_58[20] , \wRegInBot_6_58[19] , 
        \wRegInBot_6_58[18] , \wRegInBot_6_58[17] , \wRegInBot_6_58[16] , 
        \wRegInBot_6_58[15] , \wRegInBot_6_58[14] , \wRegInBot_6_58[13] , 
        \wRegInBot_6_58[12] , \wRegInBot_6_58[11] , \wRegInBot_6_58[10] , 
        \wRegInBot_6_58[9] , \wRegInBot_6_58[8] , \wRegInBot_6_58[7] , 
        \wRegInBot_6_58[6] , \wRegInBot_6_58[5] , \wRegInBot_6_58[4] , 
        \wRegInBot_6_58[3] , \wRegInBot_6_58[2] , \wRegInBot_6_58[1] , 
        \wRegInBot_6_58[0] }), .L_WR(\wRegEnTop_7_116[0] ), .L_In({
        \wRegOut_7_116[31] , \wRegOut_7_116[30] , \wRegOut_7_116[29] , 
        \wRegOut_7_116[28] , \wRegOut_7_116[27] , \wRegOut_7_116[26] , 
        \wRegOut_7_116[25] , \wRegOut_7_116[24] , \wRegOut_7_116[23] , 
        \wRegOut_7_116[22] , \wRegOut_7_116[21] , \wRegOut_7_116[20] , 
        \wRegOut_7_116[19] , \wRegOut_7_116[18] , \wRegOut_7_116[17] , 
        \wRegOut_7_116[16] , \wRegOut_7_116[15] , \wRegOut_7_116[14] , 
        \wRegOut_7_116[13] , \wRegOut_7_116[12] , \wRegOut_7_116[11] , 
        \wRegOut_7_116[10] , \wRegOut_7_116[9] , \wRegOut_7_116[8] , 
        \wRegOut_7_116[7] , \wRegOut_7_116[6] , \wRegOut_7_116[5] , 
        \wRegOut_7_116[4] , \wRegOut_7_116[3] , \wRegOut_7_116[2] , 
        \wRegOut_7_116[1] , \wRegOut_7_116[0] }), .L_Out({
        \wRegInTop_7_116[31] , \wRegInTop_7_116[30] , \wRegInTop_7_116[29] , 
        \wRegInTop_7_116[28] , \wRegInTop_7_116[27] , \wRegInTop_7_116[26] , 
        \wRegInTop_7_116[25] , \wRegInTop_7_116[24] , \wRegInTop_7_116[23] , 
        \wRegInTop_7_116[22] , \wRegInTop_7_116[21] , \wRegInTop_7_116[20] , 
        \wRegInTop_7_116[19] , \wRegInTop_7_116[18] , \wRegInTop_7_116[17] , 
        \wRegInTop_7_116[16] , \wRegInTop_7_116[15] , \wRegInTop_7_116[14] , 
        \wRegInTop_7_116[13] , \wRegInTop_7_116[12] , \wRegInTop_7_116[11] , 
        \wRegInTop_7_116[10] , \wRegInTop_7_116[9] , \wRegInTop_7_116[8] , 
        \wRegInTop_7_116[7] , \wRegInTop_7_116[6] , \wRegInTop_7_116[5] , 
        \wRegInTop_7_116[4] , \wRegInTop_7_116[3] , \wRegInTop_7_116[2] , 
        \wRegInTop_7_116[1] , \wRegInTop_7_116[0] }), .R_WR(
        \wRegEnTop_7_117[0] ), .R_In({\wRegOut_7_117[31] , \wRegOut_7_117[30] , 
        \wRegOut_7_117[29] , \wRegOut_7_117[28] , \wRegOut_7_117[27] , 
        \wRegOut_7_117[26] , \wRegOut_7_117[25] , \wRegOut_7_117[24] , 
        \wRegOut_7_117[23] , \wRegOut_7_117[22] , \wRegOut_7_117[21] , 
        \wRegOut_7_117[20] , \wRegOut_7_117[19] , \wRegOut_7_117[18] , 
        \wRegOut_7_117[17] , \wRegOut_7_117[16] , \wRegOut_7_117[15] , 
        \wRegOut_7_117[14] , \wRegOut_7_117[13] , \wRegOut_7_117[12] , 
        \wRegOut_7_117[11] , \wRegOut_7_117[10] , \wRegOut_7_117[9] , 
        \wRegOut_7_117[8] , \wRegOut_7_117[7] , \wRegOut_7_117[6] , 
        \wRegOut_7_117[5] , \wRegOut_7_117[4] , \wRegOut_7_117[3] , 
        \wRegOut_7_117[2] , \wRegOut_7_117[1] , \wRegOut_7_117[0] }), .R_Out({
        \wRegInTop_7_117[31] , \wRegInTop_7_117[30] , \wRegInTop_7_117[29] , 
        \wRegInTop_7_117[28] , \wRegInTop_7_117[27] , \wRegInTop_7_117[26] , 
        \wRegInTop_7_117[25] , \wRegInTop_7_117[24] , \wRegInTop_7_117[23] , 
        \wRegInTop_7_117[22] , \wRegInTop_7_117[21] , \wRegInTop_7_117[20] , 
        \wRegInTop_7_117[19] , \wRegInTop_7_117[18] , \wRegInTop_7_117[17] , 
        \wRegInTop_7_117[16] , \wRegInTop_7_117[15] , \wRegInTop_7_117[14] , 
        \wRegInTop_7_117[13] , \wRegInTop_7_117[12] , \wRegInTop_7_117[11] , 
        \wRegInTop_7_117[10] , \wRegInTop_7_117[9] , \wRegInTop_7_117[8] , 
        \wRegInTop_7_117[7] , \wRegInTop_7_117[6] , \wRegInTop_7_117[5] , 
        \wRegInTop_7_117[4] , \wRegInTop_7_117[3] , \wRegInTop_7_117[2] , 
        \wRegInTop_7_117[1] , \wRegInTop_7_117[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink39[31] , \ScanLink39[30] , \ScanLink39[29] , 
        \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , \ScanLink39[25] , 
        \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , \ScanLink39[21] , 
        \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , \ScanLink39[17] , 
        \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , \ScanLink39[13] , 
        \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , \ScanLink39[9] , 
        \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , \ScanLink39[5] , 
        \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , \ScanLink39[1] , 
        \ScanLink39[0] }), .ScanOut({\ScanLink38[31] , \ScanLink38[30] , 
        \ScanLink38[29] , \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , 
        \ScanLink38[25] , \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , 
        \ScanLink38[21] , \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , 
        \ScanLink38[17] , \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , 
        \ScanLink38[13] , \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , 
        \ScanLink38[9] , \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , 
        \ScanLink38[5] , \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , 
        \ScanLink38[1] , \ScanLink38[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_7[31] , \wRegOut_5_7[30] , \wRegOut_5_7[29] , 
        \wRegOut_5_7[28] , \wRegOut_5_7[27] , \wRegOut_5_7[26] , 
        \wRegOut_5_7[25] , \wRegOut_5_7[24] , \wRegOut_5_7[23] , 
        \wRegOut_5_7[22] , \wRegOut_5_7[21] , \wRegOut_5_7[20] , 
        \wRegOut_5_7[19] , \wRegOut_5_7[18] , \wRegOut_5_7[17] , 
        \wRegOut_5_7[16] , \wRegOut_5_7[15] , \wRegOut_5_7[14] , 
        \wRegOut_5_7[13] , \wRegOut_5_7[12] , \wRegOut_5_7[11] , 
        \wRegOut_5_7[10] , \wRegOut_5_7[9] , \wRegOut_5_7[8] , 
        \wRegOut_5_7[7] , \wRegOut_5_7[6] , \wRegOut_5_7[5] , \wRegOut_5_7[4] , 
        \wRegOut_5_7[3] , \wRegOut_5_7[2] , \wRegOut_5_7[1] , \wRegOut_5_7[0] 
        }), .Enable1(\wRegEnTop_5_7[0] ), .Enable2(\wRegEnBot_5_7[0] ), .In1({
        \wRegInTop_5_7[31] , \wRegInTop_5_7[30] , \wRegInTop_5_7[29] , 
        \wRegInTop_5_7[28] , \wRegInTop_5_7[27] , \wRegInTop_5_7[26] , 
        \wRegInTop_5_7[25] , \wRegInTop_5_7[24] , \wRegInTop_5_7[23] , 
        \wRegInTop_5_7[22] , \wRegInTop_5_7[21] , \wRegInTop_5_7[20] , 
        \wRegInTop_5_7[19] , \wRegInTop_5_7[18] , \wRegInTop_5_7[17] , 
        \wRegInTop_5_7[16] , \wRegInTop_5_7[15] , \wRegInTop_5_7[14] , 
        \wRegInTop_5_7[13] , \wRegInTop_5_7[12] , \wRegInTop_5_7[11] , 
        \wRegInTop_5_7[10] , \wRegInTop_5_7[9] , \wRegInTop_5_7[8] , 
        \wRegInTop_5_7[7] , \wRegInTop_5_7[6] , \wRegInTop_5_7[5] , 
        \wRegInTop_5_7[4] , \wRegInTop_5_7[3] , \wRegInTop_5_7[2] , 
        \wRegInTop_5_7[1] , \wRegInTop_5_7[0] }), .In2({\wRegInBot_5_7[31] , 
        \wRegInBot_5_7[30] , \wRegInBot_5_7[29] , \wRegInBot_5_7[28] , 
        \wRegInBot_5_7[27] , \wRegInBot_5_7[26] , \wRegInBot_5_7[25] , 
        \wRegInBot_5_7[24] , \wRegInBot_5_7[23] , \wRegInBot_5_7[22] , 
        \wRegInBot_5_7[21] , \wRegInBot_5_7[20] , \wRegInBot_5_7[19] , 
        \wRegInBot_5_7[18] , \wRegInBot_5_7[17] , \wRegInBot_5_7[16] , 
        \wRegInBot_5_7[15] , \wRegInBot_5_7[14] , \wRegInBot_5_7[13] , 
        \wRegInBot_5_7[12] , \wRegInBot_5_7[11] , \wRegInBot_5_7[10] , 
        \wRegInBot_5_7[9] , \wRegInBot_5_7[8] , \wRegInBot_5_7[7] , 
        \wRegInBot_5_7[6] , \wRegInBot_5_7[5] , \wRegInBot_5_7[4] , 
        \wRegInBot_5_7[3] , \wRegInBot_5_7[2] , \wRegInBot_5_7[1] , 
        \wRegInBot_5_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_39 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink103[31] , \ScanLink103[30] , \ScanLink103[29] , 
        \ScanLink103[28] , \ScanLink103[27] , \ScanLink103[26] , 
        \ScanLink103[25] , \ScanLink103[24] , \ScanLink103[23] , 
        \ScanLink103[22] , \ScanLink103[21] , \ScanLink103[20] , 
        \ScanLink103[19] , \ScanLink103[18] , \ScanLink103[17] , 
        \ScanLink103[16] , \ScanLink103[15] , \ScanLink103[14] , 
        \ScanLink103[13] , \ScanLink103[12] , \ScanLink103[11] , 
        \ScanLink103[10] , \ScanLink103[9] , \ScanLink103[8] , 
        \ScanLink103[7] , \ScanLink103[6] , \ScanLink103[5] , \ScanLink103[4] , 
        \ScanLink103[3] , \ScanLink103[2] , \ScanLink103[1] , \ScanLink103[0] 
        }), .ScanOut({\ScanLink102[31] , \ScanLink102[30] , \ScanLink102[29] , 
        \ScanLink102[28] , \ScanLink102[27] , \ScanLink102[26] , 
        \ScanLink102[25] , \ScanLink102[24] , \ScanLink102[23] , 
        \ScanLink102[22] , \ScanLink102[21] , \ScanLink102[20] , 
        \ScanLink102[19] , \ScanLink102[18] , \ScanLink102[17] , 
        \ScanLink102[16] , \ScanLink102[15] , \ScanLink102[14] , 
        \ScanLink102[13] , \ScanLink102[12] , \ScanLink102[11] , 
        \ScanLink102[10] , \ScanLink102[9] , \ScanLink102[8] , 
        \ScanLink102[7] , \ScanLink102[6] , \ScanLink102[5] , \ScanLink102[4] , 
        \ScanLink102[3] , \ScanLink102[2] , \ScanLink102[1] , \ScanLink102[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_39[31] , 
        \wRegOut_6_39[30] , \wRegOut_6_39[29] , \wRegOut_6_39[28] , 
        \wRegOut_6_39[27] , \wRegOut_6_39[26] , \wRegOut_6_39[25] , 
        \wRegOut_6_39[24] , \wRegOut_6_39[23] , \wRegOut_6_39[22] , 
        \wRegOut_6_39[21] , \wRegOut_6_39[20] , \wRegOut_6_39[19] , 
        \wRegOut_6_39[18] , \wRegOut_6_39[17] , \wRegOut_6_39[16] , 
        \wRegOut_6_39[15] , \wRegOut_6_39[14] , \wRegOut_6_39[13] , 
        \wRegOut_6_39[12] , \wRegOut_6_39[11] , \wRegOut_6_39[10] , 
        \wRegOut_6_39[9] , \wRegOut_6_39[8] , \wRegOut_6_39[7] , 
        \wRegOut_6_39[6] , \wRegOut_6_39[5] , \wRegOut_6_39[4] , 
        \wRegOut_6_39[3] , \wRegOut_6_39[2] , \wRegOut_6_39[1] , 
        \wRegOut_6_39[0] }), .Enable1(\wRegEnTop_6_39[0] ), .Enable2(
        \wRegEnBot_6_39[0] ), .In1({\wRegInTop_6_39[31] , \wRegInTop_6_39[30] , 
        \wRegInTop_6_39[29] , \wRegInTop_6_39[28] , \wRegInTop_6_39[27] , 
        \wRegInTop_6_39[26] , \wRegInTop_6_39[25] , \wRegInTop_6_39[24] , 
        \wRegInTop_6_39[23] , \wRegInTop_6_39[22] , \wRegInTop_6_39[21] , 
        \wRegInTop_6_39[20] , \wRegInTop_6_39[19] , \wRegInTop_6_39[18] , 
        \wRegInTop_6_39[17] , \wRegInTop_6_39[16] , \wRegInTop_6_39[15] , 
        \wRegInTop_6_39[14] , \wRegInTop_6_39[13] , \wRegInTop_6_39[12] , 
        \wRegInTop_6_39[11] , \wRegInTop_6_39[10] , \wRegInTop_6_39[9] , 
        \wRegInTop_6_39[8] , \wRegInTop_6_39[7] , \wRegInTop_6_39[6] , 
        \wRegInTop_6_39[5] , \wRegInTop_6_39[4] , \wRegInTop_6_39[3] , 
        \wRegInTop_6_39[2] , \wRegInTop_6_39[1] , \wRegInTop_6_39[0] }), .In2(
        {\wRegInBot_6_39[31] , \wRegInBot_6_39[30] , \wRegInBot_6_39[29] , 
        \wRegInBot_6_39[28] , \wRegInBot_6_39[27] , \wRegInBot_6_39[26] , 
        \wRegInBot_6_39[25] , \wRegInBot_6_39[24] , \wRegInBot_6_39[23] , 
        \wRegInBot_6_39[22] , \wRegInBot_6_39[21] , \wRegInBot_6_39[20] , 
        \wRegInBot_6_39[19] , \wRegInBot_6_39[18] , \wRegInBot_6_39[17] , 
        \wRegInBot_6_39[16] , \wRegInBot_6_39[15] , \wRegInBot_6_39[14] , 
        \wRegInBot_6_39[13] , \wRegInBot_6_39[12] , \wRegInBot_6_39[11] , 
        \wRegInBot_6_39[10] , \wRegInBot_6_39[9] , \wRegInBot_6_39[8] , 
        \wRegInBot_6_39[7] , \wRegInBot_6_39[6] , \wRegInBot_6_39[5] , 
        \wRegInBot_6_39[4] , \wRegInBot_6_39[3] , \wRegInBot_6_39[2] , 
        \wRegInBot_6_39[1] , \wRegInBot_6_39[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_57 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink121[31] , \ScanLink121[30] , \ScanLink121[29] , 
        \ScanLink121[28] , \ScanLink121[27] , \ScanLink121[26] , 
        \ScanLink121[25] , \ScanLink121[24] , \ScanLink121[23] , 
        \ScanLink121[22] , \ScanLink121[21] , \ScanLink121[20] , 
        \ScanLink121[19] , \ScanLink121[18] , \ScanLink121[17] , 
        \ScanLink121[16] , \ScanLink121[15] , \ScanLink121[14] , 
        \ScanLink121[13] , \ScanLink121[12] , \ScanLink121[11] , 
        \ScanLink121[10] , \ScanLink121[9] , \ScanLink121[8] , 
        \ScanLink121[7] , \ScanLink121[6] , \ScanLink121[5] , \ScanLink121[4] , 
        \ScanLink121[3] , \ScanLink121[2] , \ScanLink121[1] , \ScanLink121[0] 
        }), .ScanOut({\ScanLink120[31] , \ScanLink120[30] , \ScanLink120[29] , 
        \ScanLink120[28] , \ScanLink120[27] , \ScanLink120[26] , 
        \ScanLink120[25] , \ScanLink120[24] , \ScanLink120[23] , 
        \ScanLink120[22] , \ScanLink120[21] , \ScanLink120[20] , 
        \ScanLink120[19] , \ScanLink120[18] , \ScanLink120[17] , 
        \ScanLink120[16] , \ScanLink120[15] , \ScanLink120[14] , 
        \ScanLink120[13] , \ScanLink120[12] , \ScanLink120[11] , 
        \ScanLink120[10] , \ScanLink120[9] , \ScanLink120[8] , 
        \ScanLink120[7] , \ScanLink120[6] , \ScanLink120[5] , \ScanLink120[4] , 
        \ScanLink120[3] , \ScanLink120[2] , \ScanLink120[1] , \ScanLink120[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_57[31] , 
        \wRegOut_6_57[30] , \wRegOut_6_57[29] , \wRegOut_6_57[28] , 
        \wRegOut_6_57[27] , \wRegOut_6_57[26] , \wRegOut_6_57[25] , 
        \wRegOut_6_57[24] , \wRegOut_6_57[23] , \wRegOut_6_57[22] , 
        \wRegOut_6_57[21] , \wRegOut_6_57[20] , \wRegOut_6_57[19] , 
        \wRegOut_6_57[18] , \wRegOut_6_57[17] , \wRegOut_6_57[16] , 
        \wRegOut_6_57[15] , \wRegOut_6_57[14] , \wRegOut_6_57[13] , 
        \wRegOut_6_57[12] , \wRegOut_6_57[11] , \wRegOut_6_57[10] , 
        \wRegOut_6_57[9] , \wRegOut_6_57[8] , \wRegOut_6_57[7] , 
        \wRegOut_6_57[6] , \wRegOut_6_57[5] , \wRegOut_6_57[4] , 
        \wRegOut_6_57[3] , \wRegOut_6_57[2] , \wRegOut_6_57[1] , 
        \wRegOut_6_57[0] }), .Enable1(\wRegEnTop_6_57[0] ), .Enable2(
        \wRegEnBot_6_57[0] ), .In1({\wRegInTop_6_57[31] , \wRegInTop_6_57[30] , 
        \wRegInTop_6_57[29] , \wRegInTop_6_57[28] , \wRegInTop_6_57[27] , 
        \wRegInTop_6_57[26] , \wRegInTop_6_57[25] , \wRegInTop_6_57[24] , 
        \wRegInTop_6_57[23] , \wRegInTop_6_57[22] , \wRegInTop_6_57[21] , 
        \wRegInTop_6_57[20] , \wRegInTop_6_57[19] , \wRegInTop_6_57[18] , 
        \wRegInTop_6_57[17] , \wRegInTop_6_57[16] , \wRegInTop_6_57[15] , 
        \wRegInTop_6_57[14] , \wRegInTop_6_57[13] , \wRegInTop_6_57[12] , 
        \wRegInTop_6_57[11] , \wRegInTop_6_57[10] , \wRegInTop_6_57[9] , 
        \wRegInTop_6_57[8] , \wRegInTop_6_57[7] , \wRegInTop_6_57[6] , 
        \wRegInTop_6_57[5] , \wRegInTop_6_57[4] , \wRegInTop_6_57[3] , 
        \wRegInTop_6_57[2] , \wRegInTop_6_57[1] , \wRegInTop_6_57[0] }), .In2(
        {\wRegInBot_6_57[31] , \wRegInBot_6_57[30] , \wRegInBot_6_57[29] , 
        \wRegInBot_6_57[28] , \wRegInBot_6_57[27] , \wRegInBot_6_57[26] , 
        \wRegInBot_6_57[25] , \wRegInBot_6_57[24] , \wRegInBot_6_57[23] , 
        \wRegInBot_6_57[22] , \wRegInBot_6_57[21] , \wRegInBot_6_57[20] , 
        \wRegInBot_6_57[19] , \wRegInBot_6_57[18] , \wRegInBot_6_57[17] , 
        \wRegInBot_6_57[16] , \wRegInBot_6_57[15] , \wRegInBot_6_57[14] , 
        \wRegInBot_6_57[13] , \wRegInBot_6_57[12] , \wRegInBot_6_57[11] , 
        \wRegInBot_6_57[10] , \wRegInBot_6_57[9] , \wRegInBot_6_57[8] , 
        \wRegInBot_6_57[7] , \wRegInBot_6_57[6] , \wRegInBot_6_57[5] , 
        \wRegInBot_6_57[4] , \wRegInBot_6_57[3] , \wRegInBot_6_57[2] , 
        \wRegInBot_6_57[1] , \wRegInBot_6_57[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_23 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink151[31] , \ScanLink151[30] , \ScanLink151[29] , 
        \ScanLink151[28] , \ScanLink151[27] , \ScanLink151[26] , 
        \ScanLink151[25] , \ScanLink151[24] , \ScanLink151[23] , 
        \ScanLink151[22] , \ScanLink151[21] , \ScanLink151[20] , 
        \ScanLink151[19] , \ScanLink151[18] , \ScanLink151[17] , 
        \ScanLink151[16] , \ScanLink151[15] , \ScanLink151[14] , 
        \ScanLink151[13] , \ScanLink151[12] , \ScanLink151[11] , 
        \ScanLink151[10] , \ScanLink151[9] , \ScanLink151[8] , 
        \ScanLink151[7] , \ScanLink151[6] , \ScanLink151[5] , \ScanLink151[4] , 
        \ScanLink151[3] , \ScanLink151[2] , \ScanLink151[1] , \ScanLink151[0] 
        }), .ScanOut({\ScanLink150[31] , \ScanLink150[30] , \ScanLink150[29] , 
        \ScanLink150[28] , \ScanLink150[27] , \ScanLink150[26] , 
        \ScanLink150[25] , \ScanLink150[24] , \ScanLink150[23] , 
        \ScanLink150[22] , \ScanLink150[21] , \ScanLink150[20] , 
        \ScanLink150[19] , \ScanLink150[18] , \ScanLink150[17] , 
        \ScanLink150[16] , \ScanLink150[15] , \ScanLink150[14] , 
        \ScanLink150[13] , \ScanLink150[12] , \ScanLink150[11] , 
        \ScanLink150[10] , \ScanLink150[9] , \ScanLink150[8] , 
        \ScanLink150[7] , \ScanLink150[6] , \ScanLink150[5] , \ScanLink150[4] , 
        \ScanLink150[3] , \ScanLink150[2] , \ScanLink150[1] , \ScanLink150[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_23[31] , 
        \wRegOut_7_23[30] , \wRegOut_7_23[29] , \wRegOut_7_23[28] , 
        \wRegOut_7_23[27] , \wRegOut_7_23[26] , \wRegOut_7_23[25] , 
        \wRegOut_7_23[24] , \wRegOut_7_23[23] , \wRegOut_7_23[22] , 
        \wRegOut_7_23[21] , \wRegOut_7_23[20] , \wRegOut_7_23[19] , 
        \wRegOut_7_23[18] , \wRegOut_7_23[17] , \wRegOut_7_23[16] , 
        \wRegOut_7_23[15] , \wRegOut_7_23[14] , \wRegOut_7_23[13] , 
        \wRegOut_7_23[12] , \wRegOut_7_23[11] , \wRegOut_7_23[10] , 
        \wRegOut_7_23[9] , \wRegOut_7_23[8] , \wRegOut_7_23[7] , 
        \wRegOut_7_23[6] , \wRegOut_7_23[5] , \wRegOut_7_23[4] , 
        \wRegOut_7_23[3] , \wRegOut_7_23[2] , \wRegOut_7_23[1] , 
        \wRegOut_7_23[0] }), .Enable1(\wRegEnTop_7_23[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_23[31] , \wRegInTop_7_23[30] , \wRegInTop_7_23[29] , 
        \wRegInTop_7_23[28] , \wRegInTop_7_23[27] , \wRegInTop_7_23[26] , 
        \wRegInTop_7_23[25] , \wRegInTop_7_23[24] , \wRegInTop_7_23[23] , 
        \wRegInTop_7_23[22] , \wRegInTop_7_23[21] , \wRegInTop_7_23[20] , 
        \wRegInTop_7_23[19] , \wRegInTop_7_23[18] , \wRegInTop_7_23[17] , 
        \wRegInTop_7_23[16] , \wRegInTop_7_23[15] , \wRegInTop_7_23[14] , 
        \wRegInTop_7_23[13] , \wRegInTop_7_23[12] , \wRegInTop_7_23[11] , 
        \wRegInTop_7_23[10] , \wRegInTop_7_23[9] , \wRegInTop_7_23[8] , 
        \wRegInTop_7_23[7] , \wRegInTop_7_23[6] , \wRegInTop_7_23[5] , 
        \wRegInTop_7_23[4] , \wRegInTop_7_23[3] , \wRegInTop_7_23[2] , 
        \wRegInTop_7_23[1] , \wRegInTop_7_23[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_21[0] ), .P_In({\wRegOut_5_21[31] , 
        \wRegOut_5_21[30] , \wRegOut_5_21[29] , \wRegOut_5_21[28] , 
        \wRegOut_5_21[27] , \wRegOut_5_21[26] , \wRegOut_5_21[25] , 
        \wRegOut_5_21[24] , \wRegOut_5_21[23] , \wRegOut_5_21[22] , 
        \wRegOut_5_21[21] , \wRegOut_5_21[20] , \wRegOut_5_21[19] , 
        \wRegOut_5_21[18] , \wRegOut_5_21[17] , \wRegOut_5_21[16] , 
        \wRegOut_5_21[15] , \wRegOut_5_21[14] , \wRegOut_5_21[13] , 
        \wRegOut_5_21[12] , \wRegOut_5_21[11] , \wRegOut_5_21[10] , 
        \wRegOut_5_21[9] , \wRegOut_5_21[8] , \wRegOut_5_21[7] , 
        \wRegOut_5_21[6] , \wRegOut_5_21[5] , \wRegOut_5_21[4] , 
        \wRegOut_5_21[3] , \wRegOut_5_21[2] , \wRegOut_5_21[1] , 
        \wRegOut_5_21[0] }), .P_Out({\wRegInBot_5_21[31] , 
        \wRegInBot_5_21[30] , \wRegInBot_5_21[29] , \wRegInBot_5_21[28] , 
        \wRegInBot_5_21[27] , \wRegInBot_5_21[26] , \wRegInBot_5_21[25] , 
        \wRegInBot_5_21[24] , \wRegInBot_5_21[23] , \wRegInBot_5_21[22] , 
        \wRegInBot_5_21[21] , \wRegInBot_5_21[20] , \wRegInBot_5_21[19] , 
        \wRegInBot_5_21[18] , \wRegInBot_5_21[17] , \wRegInBot_5_21[16] , 
        \wRegInBot_5_21[15] , \wRegInBot_5_21[14] , \wRegInBot_5_21[13] , 
        \wRegInBot_5_21[12] , \wRegInBot_5_21[11] , \wRegInBot_5_21[10] , 
        \wRegInBot_5_21[9] , \wRegInBot_5_21[8] , \wRegInBot_5_21[7] , 
        \wRegInBot_5_21[6] , \wRegInBot_5_21[5] , \wRegInBot_5_21[4] , 
        \wRegInBot_5_21[3] , \wRegInBot_5_21[2] , \wRegInBot_5_21[1] , 
        \wRegInBot_5_21[0] }), .L_WR(\wRegEnTop_6_42[0] ), .L_In({
        \wRegOut_6_42[31] , \wRegOut_6_42[30] , \wRegOut_6_42[29] , 
        \wRegOut_6_42[28] , \wRegOut_6_42[27] , \wRegOut_6_42[26] , 
        \wRegOut_6_42[25] , \wRegOut_6_42[24] , \wRegOut_6_42[23] , 
        \wRegOut_6_42[22] , \wRegOut_6_42[21] , \wRegOut_6_42[20] , 
        \wRegOut_6_42[19] , \wRegOut_6_42[18] , \wRegOut_6_42[17] , 
        \wRegOut_6_42[16] , \wRegOut_6_42[15] , \wRegOut_6_42[14] , 
        \wRegOut_6_42[13] , \wRegOut_6_42[12] , \wRegOut_6_42[11] , 
        \wRegOut_6_42[10] , \wRegOut_6_42[9] , \wRegOut_6_42[8] , 
        \wRegOut_6_42[7] , \wRegOut_6_42[6] , \wRegOut_6_42[5] , 
        \wRegOut_6_42[4] , \wRegOut_6_42[3] , \wRegOut_6_42[2] , 
        \wRegOut_6_42[1] , \wRegOut_6_42[0] }), .L_Out({\wRegInTop_6_42[31] , 
        \wRegInTop_6_42[30] , \wRegInTop_6_42[29] , \wRegInTop_6_42[28] , 
        \wRegInTop_6_42[27] , \wRegInTop_6_42[26] , \wRegInTop_6_42[25] , 
        \wRegInTop_6_42[24] , \wRegInTop_6_42[23] , \wRegInTop_6_42[22] , 
        \wRegInTop_6_42[21] , \wRegInTop_6_42[20] , \wRegInTop_6_42[19] , 
        \wRegInTop_6_42[18] , \wRegInTop_6_42[17] , \wRegInTop_6_42[16] , 
        \wRegInTop_6_42[15] , \wRegInTop_6_42[14] , \wRegInTop_6_42[13] , 
        \wRegInTop_6_42[12] , \wRegInTop_6_42[11] , \wRegInTop_6_42[10] , 
        \wRegInTop_6_42[9] , \wRegInTop_6_42[8] , \wRegInTop_6_42[7] , 
        \wRegInTop_6_42[6] , \wRegInTop_6_42[5] , \wRegInTop_6_42[4] , 
        \wRegInTop_6_42[3] , \wRegInTop_6_42[2] , \wRegInTop_6_42[1] , 
        \wRegInTop_6_42[0] }), .R_WR(\wRegEnTop_6_43[0] ), .R_In({
        \wRegOut_6_43[31] , \wRegOut_6_43[30] , \wRegOut_6_43[29] , 
        \wRegOut_6_43[28] , \wRegOut_6_43[27] , \wRegOut_6_43[26] , 
        \wRegOut_6_43[25] , \wRegOut_6_43[24] , \wRegOut_6_43[23] , 
        \wRegOut_6_43[22] , \wRegOut_6_43[21] , \wRegOut_6_43[20] , 
        \wRegOut_6_43[19] , \wRegOut_6_43[18] , \wRegOut_6_43[17] , 
        \wRegOut_6_43[16] , \wRegOut_6_43[15] , \wRegOut_6_43[14] , 
        \wRegOut_6_43[13] , \wRegOut_6_43[12] , \wRegOut_6_43[11] , 
        \wRegOut_6_43[10] , \wRegOut_6_43[9] , \wRegOut_6_43[8] , 
        \wRegOut_6_43[7] , \wRegOut_6_43[6] , \wRegOut_6_43[5] , 
        \wRegOut_6_43[4] , \wRegOut_6_43[3] , \wRegOut_6_43[2] , 
        \wRegOut_6_43[1] , \wRegOut_6_43[0] }), .R_Out({\wRegInTop_6_43[31] , 
        \wRegInTop_6_43[30] , \wRegInTop_6_43[29] , \wRegInTop_6_43[28] , 
        \wRegInTop_6_43[27] , \wRegInTop_6_43[26] , \wRegInTop_6_43[25] , 
        \wRegInTop_6_43[24] , \wRegInTop_6_43[23] , \wRegInTop_6_43[22] , 
        \wRegInTop_6_43[21] , \wRegInTop_6_43[20] , \wRegInTop_6_43[19] , 
        \wRegInTop_6_43[18] , \wRegInTop_6_43[17] , \wRegInTop_6_43[16] , 
        \wRegInTop_6_43[15] , \wRegInTop_6_43[14] , \wRegInTop_6_43[13] , 
        \wRegInTop_6_43[12] , \wRegInTop_6_43[11] , \wRegInTop_6_43[10] , 
        \wRegInTop_6_43[9] , \wRegInTop_6_43[8] , \wRegInTop_6_43[7] , 
        \wRegInTop_6_43[6] , \wRegInTop_6_43[5] , \wRegInTop_6_43[4] , 
        \wRegInTop_6_43[3] , \wRegInTop_6_43[2] , \wRegInTop_6_43[1] , 
        \wRegInTop_6_43[0] }) );
    BHeap_Node_WIDTH32 BHN_6_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_11[0] ), .P_In({\wRegOut_6_11[31] , 
        \wRegOut_6_11[30] , \wRegOut_6_11[29] , \wRegOut_6_11[28] , 
        \wRegOut_6_11[27] , \wRegOut_6_11[26] , \wRegOut_6_11[25] , 
        \wRegOut_6_11[24] , \wRegOut_6_11[23] , \wRegOut_6_11[22] , 
        \wRegOut_6_11[21] , \wRegOut_6_11[20] , \wRegOut_6_11[19] , 
        \wRegOut_6_11[18] , \wRegOut_6_11[17] , \wRegOut_6_11[16] , 
        \wRegOut_6_11[15] , \wRegOut_6_11[14] , \wRegOut_6_11[13] , 
        \wRegOut_6_11[12] , \wRegOut_6_11[11] , \wRegOut_6_11[10] , 
        \wRegOut_6_11[9] , \wRegOut_6_11[8] , \wRegOut_6_11[7] , 
        \wRegOut_6_11[6] , \wRegOut_6_11[5] , \wRegOut_6_11[4] , 
        \wRegOut_6_11[3] , \wRegOut_6_11[2] , \wRegOut_6_11[1] , 
        \wRegOut_6_11[0] }), .P_Out({\wRegInBot_6_11[31] , 
        \wRegInBot_6_11[30] , \wRegInBot_6_11[29] , \wRegInBot_6_11[28] , 
        \wRegInBot_6_11[27] , \wRegInBot_6_11[26] , \wRegInBot_6_11[25] , 
        \wRegInBot_6_11[24] , \wRegInBot_6_11[23] , \wRegInBot_6_11[22] , 
        \wRegInBot_6_11[21] , \wRegInBot_6_11[20] , \wRegInBot_6_11[19] , 
        \wRegInBot_6_11[18] , \wRegInBot_6_11[17] , \wRegInBot_6_11[16] , 
        \wRegInBot_6_11[15] , \wRegInBot_6_11[14] , \wRegInBot_6_11[13] , 
        \wRegInBot_6_11[12] , \wRegInBot_6_11[11] , \wRegInBot_6_11[10] , 
        \wRegInBot_6_11[9] , \wRegInBot_6_11[8] , \wRegInBot_6_11[7] , 
        \wRegInBot_6_11[6] , \wRegInBot_6_11[5] , \wRegInBot_6_11[4] , 
        \wRegInBot_6_11[3] , \wRegInBot_6_11[2] , \wRegInBot_6_11[1] , 
        \wRegInBot_6_11[0] }), .L_WR(\wRegEnTop_7_22[0] ), .L_In({
        \wRegOut_7_22[31] , \wRegOut_7_22[30] , \wRegOut_7_22[29] , 
        \wRegOut_7_22[28] , \wRegOut_7_22[27] , \wRegOut_7_22[26] , 
        \wRegOut_7_22[25] , \wRegOut_7_22[24] , \wRegOut_7_22[23] , 
        \wRegOut_7_22[22] , \wRegOut_7_22[21] , \wRegOut_7_22[20] , 
        \wRegOut_7_22[19] , \wRegOut_7_22[18] , \wRegOut_7_22[17] , 
        \wRegOut_7_22[16] , \wRegOut_7_22[15] , \wRegOut_7_22[14] , 
        \wRegOut_7_22[13] , \wRegOut_7_22[12] , \wRegOut_7_22[11] , 
        \wRegOut_7_22[10] , \wRegOut_7_22[9] , \wRegOut_7_22[8] , 
        \wRegOut_7_22[7] , \wRegOut_7_22[6] , \wRegOut_7_22[5] , 
        \wRegOut_7_22[4] , \wRegOut_7_22[3] , \wRegOut_7_22[2] , 
        \wRegOut_7_22[1] , \wRegOut_7_22[0] }), .L_Out({\wRegInTop_7_22[31] , 
        \wRegInTop_7_22[30] , \wRegInTop_7_22[29] , \wRegInTop_7_22[28] , 
        \wRegInTop_7_22[27] , \wRegInTop_7_22[26] , \wRegInTop_7_22[25] , 
        \wRegInTop_7_22[24] , \wRegInTop_7_22[23] , \wRegInTop_7_22[22] , 
        \wRegInTop_7_22[21] , \wRegInTop_7_22[20] , \wRegInTop_7_22[19] , 
        \wRegInTop_7_22[18] , \wRegInTop_7_22[17] , \wRegInTop_7_22[16] , 
        \wRegInTop_7_22[15] , \wRegInTop_7_22[14] , \wRegInTop_7_22[13] , 
        \wRegInTop_7_22[12] , \wRegInTop_7_22[11] , \wRegInTop_7_22[10] , 
        \wRegInTop_7_22[9] , \wRegInTop_7_22[8] , \wRegInTop_7_22[7] , 
        \wRegInTop_7_22[6] , \wRegInTop_7_22[5] , \wRegInTop_7_22[4] , 
        \wRegInTop_7_22[3] , \wRegInTop_7_22[2] , \wRegInTop_7_22[1] , 
        \wRegInTop_7_22[0] }), .R_WR(\wRegEnTop_7_23[0] ), .R_In({
        \wRegOut_7_23[31] , \wRegOut_7_23[30] , \wRegOut_7_23[29] , 
        \wRegOut_7_23[28] , \wRegOut_7_23[27] , \wRegOut_7_23[26] , 
        \wRegOut_7_23[25] , \wRegOut_7_23[24] , \wRegOut_7_23[23] , 
        \wRegOut_7_23[22] , \wRegOut_7_23[21] , \wRegOut_7_23[20] , 
        \wRegOut_7_23[19] , \wRegOut_7_23[18] , \wRegOut_7_23[17] , 
        \wRegOut_7_23[16] , \wRegOut_7_23[15] , \wRegOut_7_23[14] , 
        \wRegOut_7_23[13] , \wRegOut_7_23[12] , \wRegOut_7_23[11] , 
        \wRegOut_7_23[10] , \wRegOut_7_23[9] , \wRegOut_7_23[8] , 
        \wRegOut_7_23[7] , \wRegOut_7_23[6] , \wRegOut_7_23[5] , 
        \wRegOut_7_23[4] , \wRegOut_7_23[3] , \wRegOut_7_23[2] , 
        \wRegOut_7_23[1] , \wRegOut_7_23[0] }), .R_Out({\wRegInTop_7_23[31] , 
        \wRegInTop_7_23[30] , \wRegInTop_7_23[29] , \wRegInTop_7_23[28] , 
        \wRegInTop_7_23[27] , \wRegInTop_7_23[26] , \wRegInTop_7_23[25] , 
        \wRegInTop_7_23[24] , \wRegInTop_7_23[23] , \wRegInTop_7_23[22] , 
        \wRegInTop_7_23[21] , \wRegInTop_7_23[20] , \wRegInTop_7_23[19] , 
        \wRegInTop_7_23[18] , \wRegInTop_7_23[17] , \wRegInTop_7_23[16] , 
        \wRegInTop_7_23[15] , \wRegInTop_7_23[14] , \wRegInTop_7_23[13] , 
        \wRegInTop_7_23[12] , \wRegInTop_7_23[11] , \wRegInTop_7_23[10] , 
        \wRegInTop_7_23[9] , \wRegInTop_7_23[8] , \wRegInTop_7_23[7] , 
        \wRegInTop_7_23[6] , \wRegInTop_7_23[5] , \wRegInTop_7_23[4] , 
        \wRegInTop_7_23[3] , \wRegInTop_7_23[2] , \wRegInTop_7_23[1] , 
        \wRegInTop_7_23[0] }) );
    BHeap_Node_WIDTH32 BHN_6_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_36[0] ), .P_In({\wRegOut_6_36[31] , 
        \wRegOut_6_36[30] , \wRegOut_6_36[29] , \wRegOut_6_36[28] , 
        \wRegOut_6_36[27] , \wRegOut_6_36[26] , \wRegOut_6_36[25] , 
        \wRegOut_6_36[24] , \wRegOut_6_36[23] , \wRegOut_6_36[22] , 
        \wRegOut_6_36[21] , \wRegOut_6_36[20] , \wRegOut_6_36[19] , 
        \wRegOut_6_36[18] , \wRegOut_6_36[17] , \wRegOut_6_36[16] , 
        \wRegOut_6_36[15] , \wRegOut_6_36[14] , \wRegOut_6_36[13] , 
        \wRegOut_6_36[12] , \wRegOut_6_36[11] , \wRegOut_6_36[10] , 
        \wRegOut_6_36[9] , \wRegOut_6_36[8] , \wRegOut_6_36[7] , 
        \wRegOut_6_36[6] , \wRegOut_6_36[5] , \wRegOut_6_36[4] , 
        \wRegOut_6_36[3] , \wRegOut_6_36[2] , \wRegOut_6_36[1] , 
        \wRegOut_6_36[0] }), .P_Out({\wRegInBot_6_36[31] , 
        \wRegInBot_6_36[30] , \wRegInBot_6_36[29] , \wRegInBot_6_36[28] , 
        \wRegInBot_6_36[27] , \wRegInBot_6_36[26] , \wRegInBot_6_36[25] , 
        \wRegInBot_6_36[24] , \wRegInBot_6_36[23] , \wRegInBot_6_36[22] , 
        \wRegInBot_6_36[21] , \wRegInBot_6_36[20] , \wRegInBot_6_36[19] , 
        \wRegInBot_6_36[18] , \wRegInBot_6_36[17] , \wRegInBot_6_36[16] , 
        \wRegInBot_6_36[15] , \wRegInBot_6_36[14] , \wRegInBot_6_36[13] , 
        \wRegInBot_6_36[12] , \wRegInBot_6_36[11] , \wRegInBot_6_36[10] , 
        \wRegInBot_6_36[9] , \wRegInBot_6_36[8] , \wRegInBot_6_36[7] , 
        \wRegInBot_6_36[6] , \wRegInBot_6_36[5] , \wRegInBot_6_36[4] , 
        \wRegInBot_6_36[3] , \wRegInBot_6_36[2] , \wRegInBot_6_36[1] , 
        \wRegInBot_6_36[0] }), .L_WR(\wRegEnTop_7_72[0] ), .L_In({
        \wRegOut_7_72[31] , \wRegOut_7_72[30] , \wRegOut_7_72[29] , 
        \wRegOut_7_72[28] , \wRegOut_7_72[27] , \wRegOut_7_72[26] , 
        \wRegOut_7_72[25] , \wRegOut_7_72[24] , \wRegOut_7_72[23] , 
        \wRegOut_7_72[22] , \wRegOut_7_72[21] , \wRegOut_7_72[20] , 
        \wRegOut_7_72[19] , \wRegOut_7_72[18] , \wRegOut_7_72[17] , 
        \wRegOut_7_72[16] , \wRegOut_7_72[15] , \wRegOut_7_72[14] , 
        \wRegOut_7_72[13] , \wRegOut_7_72[12] , \wRegOut_7_72[11] , 
        \wRegOut_7_72[10] , \wRegOut_7_72[9] , \wRegOut_7_72[8] , 
        \wRegOut_7_72[7] , \wRegOut_7_72[6] , \wRegOut_7_72[5] , 
        \wRegOut_7_72[4] , \wRegOut_7_72[3] , \wRegOut_7_72[2] , 
        \wRegOut_7_72[1] , \wRegOut_7_72[0] }), .L_Out({\wRegInTop_7_72[31] , 
        \wRegInTop_7_72[30] , \wRegInTop_7_72[29] , \wRegInTop_7_72[28] , 
        \wRegInTop_7_72[27] , \wRegInTop_7_72[26] , \wRegInTop_7_72[25] , 
        \wRegInTop_7_72[24] , \wRegInTop_7_72[23] , \wRegInTop_7_72[22] , 
        \wRegInTop_7_72[21] , \wRegInTop_7_72[20] , \wRegInTop_7_72[19] , 
        \wRegInTop_7_72[18] , \wRegInTop_7_72[17] , \wRegInTop_7_72[16] , 
        \wRegInTop_7_72[15] , \wRegInTop_7_72[14] , \wRegInTop_7_72[13] , 
        \wRegInTop_7_72[12] , \wRegInTop_7_72[11] , \wRegInTop_7_72[10] , 
        \wRegInTop_7_72[9] , \wRegInTop_7_72[8] , \wRegInTop_7_72[7] , 
        \wRegInTop_7_72[6] , \wRegInTop_7_72[5] , \wRegInTop_7_72[4] , 
        \wRegInTop_7_72[3] , \wRegInTop_7_72[2] , \wRegInTop_7_72[1] , 
        \wRegInTop_7_72[0] }), .R_WR(\wRegEnTop_7_73[0] ), .R_In({
        \wRegOut_7_73[31] , \wRegOut_7_73[30] , \wRegOut_7_73[29] , 
        \wRegOut_7_73[28] , \wRegOut_7_73[27] , \wRegOut_7_73[26] , 
        \wRegOut_7_73[25] , \wRegOut_7_73[24] , \wRegOut_7_73[23] , 
        \wRegOut_7_73[22] , \wRegOut_7_73[21] , \wRegOut_7_73[20] , 
        \wRegOut_7_73[19] , \wRegOut_7_73[18] , \wRegOut_7_73[17] , 
        \wRegOut_7_73[16] , \wRegOut_7_73[15] , \wRegOut_7_73[14] , 
        \wRegOut_7_73[13] , \wRegOut_7_73[12] , \wRegOut_7_73[11] , 
        \wRegOut_7_73[10] , \wRegOut_7_73[9] , \wRegOut_7_73[8] , 
        \wRegOut_7_73[7] , \wRegOut_7_73[6] , \wRegOut_7_73[5] , 
        \wRegOut_7_73[4] , \wRegOut_7_73[3] , \wRegOut_7_73[2] , 
        \wRegOut_7_73[1] , \wRegOut_7_73[0] }), .R_Out({\wRegInTop_7_73[31] , 
        \wRegInTop_7_73[30] , \wRegInTop_7_73[29] , \wRegInTop_7_73[28] , 
        \wRegInTop_7_73[27] , \wRegInTop_7_73[26] , \wRegInTop_7_73[25] , 
        \wRegInTop_7_73[24] , \wRegInTop_7_73[23] , \wRegInTop_7_73[22] , 
        \wRegInTop_7_73[21] , \wRegInTop_7_73[20] , \wRegInTop_7_73[19] , 
        \wRegInTop_7_73[18] , \wRegInTop_7_73[17] , \wRegInTop_7_73[16] , 
        \wRegInTop_7_73[15] , \wRegInTop_7_73[14] , \wRegInTop_7_73[13] , 
        \wRegInTop_7_73[12] , \wRegInTop_7_73[11] , \wRegInTop_7_73[10] , 
        \wRegInTop_7_73[9] , \wRegInTop_7_73[8] , \wRegInTop_7_73[7] , 
        \wRegInTop_7_73[6] , \wRegInTop_7_73[5] , \wRegInTop_7_73[4] , 
        \wRegInTop_7_73[3] , \wRegInTop_7_73[2] , \wRegInTop_7_73[1] , 
        \wRegInTop_7_73[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_19 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink51[31] , \ScanLink51[30] , \ScanLink51[29] , 
        \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , \ScanLink51[25] , 
        \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , \ScanLink51[21] , 
        \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , \ScanLink51[17] , 
        \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , \ScanLink51[13] , 
        \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , \ScanLink51[9] , 
        \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , \ScanLink51[5] , 
        \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , \ScanLink51[1] , 
        \ScanLink51[0] }), .ScanOut({\ScanLink50[31] , \ScanLink50[30] , 
        \ScanLink50[29] , \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , 
        \ScanLink50[25] , \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , 
        \ScanLink50[21] , \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , 
        \ScanLink50[17] , \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , 
        \ScanLink50[13] , \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , 
        \ScanLink50[9] , \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , 
        \ScanLink50[5] , \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , 
        \ScanLink50[1] , \ScanLink50[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_19[31] , \wRegOut_5_19[30] , 
        \wRegOut_5_19[29] , \wRegOut_5_19[28] , \wRegOut_5_19[27] , 
        \wRegOut_5_19[26] , \wRegOut_5_19[25] , \wRegOut_5_19[24] , 
        \wRegOut_5_19[23] , \wRegOut_5_19[22] , \wRegOut_5_19[21] , 
        \wRegOut_5_19[20] , \wRegOut_5_19[19] , \wRegOut_5_19[18] , 
        \wRegOut_5_19[17] , \wRegOut_5_19[16] , \wRegOut_5_19[15] , 
        \wRegOut_5_19[14] , \wRegOut_5_19[13] , \wRegOut_5_19[12] , 
        \wRegOut_5_19[11] , \wRegOut_5_19[10] , \wRegOut_5_19[9] , 
        \wRegOut_5_19[8] , \wRegOut_5_19[7] , \wRegOut_5_19[6] , 
        \wRegOut_5_19[5] , \wRegOut_5_19[4] , \wRegOut_5_19[3] , 
        \wRegOut_5_19[2] , \wRegOut_5_19[1] , \wRegOut_5_19[0] }), .Enable1(
        \wRegEnTop_5_19[0] ), .Enable2(\wRegEnBot_5_19[0] ), .In1({
        \wRegInTop_5_19[31] , \wRegInTop_5_19[30] , \wRegInTop_5_19[29] , 
        \wRegInTop_5_19[28] , \wRegInTop_5_19[27] , \wRegInTop_5_19[26] , 
        \wRegInTop_5_19[25] , \wRegInTop_5_19[24] , \wRegInTop_5_19[23] , 
        \wRegInTop_5_19[22] , \wRegInTop_5_19[21] , \wRegInTop_5_19[20] , 
        \wRegInTop_5_19[19] , \wRegInTop_5_19[18] , \wRegInTop_5_19[17] , 
        \wRegInTop_5_19[16] , \wRegInTop_5_19[15] , \wRegInTop_5_19[14] , 
        \wRegInTop_5_19[13] , \wRegInTop_5_19[12] , \wRegInTop_5_19[11] , 
        \wRegInTop_5_19[10] , \wRegInTop_5_19[9] , \wRegInTop_5_19[8] , 
        \wRegInTop_5_19[7] , \wRegInTop_5_19[6] , \wRegInTop_5_19[5] , 
        \wRegInTop_5_19[4] , \wRegInTop_5_19[3] , \wRegInTop_5_19[2] , 
        \wRegInTop_5_19[1] , \wRegInTop_5_19[0] }), .In2({\wRegInBot_5_19[31] , 
        \wRegInBot_5_19[30] , \wRegInBot_5_19[29] , \wRegInBot_5_19[28] , 
        \wRegInBot_5_19[27] , \wRegInBot_5_19[26] , \wRegInBot_5_19[25] , 
        \wRegInBot_5_19[24] , \wRegInBot_5_19[23] , \wRegInBot_5_19[22] , 
        \wRegInBot_5_19[21] , \wRegInBot_5_19[20] , \wRegInBot_5_19[19] , 
        \wRegInBot_5_19[18] , \wRegInBot_5_19[17] , \wRegInBot_5_19[16] , 
        \wRegInBot_5_19[15] , \wRegInBot_5_19[14] , \wRegInBot_5_19[13] , 
        \wRegInBot_5_19[12] , \wRegInBot_5_19[11] , \wRegInBot_5_19[10] , 
        \wRegInBot_5_19[9] , \wRegInBot_5_19[8] , \wRegInBot_5_19[7] , 
        \wRegInBot_5_19[6] , \wRegInBot_5_19[5] , \wRegInBot_5_19[4] , 
        \wRegInBot_5_19[3] , \wRegInBot_5_19[2] , \wRegInBot_5_19[1] , 
        \wRegInBot_5_19[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_25 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink57[31] , \ScanLink57[30] , \ScanLink57[29] , 
        \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , \ScanLink57[25] , 
        \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , \ScanLink57[21] , 
        \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , \ScanLink57[17] , 
        \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , \ScanLink57[13] , 
        \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , \ScanLink57[9] , 
        \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , \ScanLink57[5] , 
        \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , \ScanLink57[1] , 
        \ScanLink57[0] }), .ScanOut({\ScanLink56[31] , \ScanLink56[30] , 
        \ScanLink56[29] , \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , 
        \ScanLink56[25] , \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , 
        \ScanLink56[21] , \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , 
        \ScanLink56[17] , \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , 
        \ScanLink56[13] , \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , 
        \ScanLink56[9] , \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , 
        \ScanLink56[5] , \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , 
        \ScanLink56[1] , \ScanLink56[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_25[31] , \wRegOut_5_25[30] , 
        \wRegOut_5_25[29] , \wRegOut_5_25[28] , \wRegOut_5_25[27] , 
        \wRegOut_5_25[26] , \wRegOut_5_25[25] , \wRegOut_5_25[24] , 
        \wRegOut_5_25[23] , \wRegOut_5_25[22] , \wRegOut_5_25[21] , 
        \wRegOut_5_25[20] , \wRegOut_5_25[19] , \wRegOut_5_25[18] , 
        \wRegOut_5_25[17] , \wRegOut_5_25[16] , \wRegOut_5_25[15] , 
        \wRegOut_5_25[14] , \wRegOut_5_25[13] , \wRegOut_5_25[12] , 
        \wRegOut_5_25[11] , \wRegOut_5_25[10] , \wRegOut_5_25[9] , 
        \wRegOut_5_25[8] , \wRegOut_5_25[7] , \wRegOut_5_25[6] , 
        \wRegOut_5_25[5] , \wRegOut_5_25[4] , \wRegOut_5_25[3] , 
        \wRegOut_5_25[2] , \wRegOut_5_25[1] , \wRegOut_5_25[0] }), .Enable1(
        \wRegEnTop_5_25[0] ), .Enable2(\wRegEnBot_5_25[0] ), .In1({
        \wRegInTop_5_25[31] , \wRegInTop_5_25[30] , \wRegInTop_5_25[29] , 
        \wRegInTop_5_25[28] , \wRegInTop_5_25[27] , \wRegInTop_5_25[26] , 
        \wRegInTop_5_25[25] , \wRegInTop_5_25[24] , \wRegInTop_5_25[23] , 
        \wRegInTop_5_25[22] , \wRegInTop_5_25[21] , \wRegInTop_5_25[20] , 
        \wRegInTop_5_25[19] , \wRegInTop_5_25[18] , \wRegInTop_5_25[17] , 
        \wRegInTop_5_25[16] , \wRegInTop_5_25[15] , \wRegInTop_5_25[14] , 
        \wRegInTop_5_25[13] , \wRegInTop_5_25[12] , \wRegInTop_5_25[11] , 
        \wRegInTop_5_25[10] , \wRegInTop_5_25[9] , \wRegInTop_5_25[8] , 
        \wRegInTop_5_25[7] , \wRegInTop_5_25[6] , \wRegInTop_5_25[5] , 
        \wRegInTop_5_25[4] , \wRegInTop_5_25[3] , \wRegInTop_5_25[2] , 
        \wRegInTop_5_25[1] , \wRegInTop_5_25[0] }), .In2({\wRegInBot_5_25[31] , 
        \wRegInBot_5_25[30] , \wRegInBot_5_25[29] , \wRegInBot_5_25[28] , 
        \wRegInBot_5_25[27] , \wRegInBot_5_25[26] , \wRegInBot_5_25[25] , 
        \wRegInBot_5_25[24] , \wRegInBot_5_25[23] , \wRegInBot_5_25[22] , 
        \wRegInBot_5_25[21] , \wRegInBot_5_25[20] , \wRegInBot_5_25[19] , 
        \wRegInBot_5_25[18] , \wRegInBot_5_25[17] , \wRegInBot_5_25[16] , 
        \wRegInBot_5_25[15] , \wRegInBot_5_25[14] , \wRegInBot_5_25[13] , 
        \wRegInBot_5_25[12] , \wRegInBot_5_25[11] , \wRegInBot_5_25[10] , 
        \wRegInBot_5_25[9] , \wRegInBot_5_25[8] , \wRegInBot_5_25[7] , 
        \wRegInBot_5_25[6] , \wRegInBot_5_25[5] , \wRegInBot_5_25[4] , 
        \wRegInBot_5_25[3] , \wRegInBot_5_25[2] , \wRegInBot_5_25[1] , 
        \wRegInBot_5_25[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink79[31] , \ScanLink79[30] , \ScanLink79[29] , 
        \ScanLink79[28] , \ScanLink79[27] , \ScanLink79[26] , \ScanLink79[25] , 
        \ScanLink79[24] , \ScanLink79[23] , \ScanLink79[22] , \ScanLink79[21] , 
        \ScanLink79[20] , \ScanLink79[19] , \ScanLink79[18] , \ScanLink79[17] , 
        \ScanLink79[16] , \ScanLink79[15] , \ScanLink79[14] , \ScanLink79[13] , 
        \ScanLink79[12] , \ScanLink79[11] , \ScanLink79[10] , \ScanLink79[9] , 
        \ScanLink79[8] , \ScanLink79[7] , \ScanLink79[6] , \ScanLink79[5] , 
        \ScanLink79[4] , \ScanLink79[3] , \ScanLink79[2] , \ScanLink79[1] , 
        \ScanLink79[0] }), .ScanOut({\ScanLink78[31] , \ScanLink78[30] , 
        \ScanLink78[29] , \ScanLink78[28] , \ScanLink78[27] , \ScanLink78[26] , 
        \ScanLink78[25] , \ScanLink78[24] , \ScanLink78[23] , \ScanLink78[22] , 
        \ScanLink78[21] , \ScanLink78[20] , \ScanLink78[19] , \ScanLink78[18] , 
        \ScanLink78[17] , \ScanLink78[16] , \ScanLink78[15] , \ScanLink78[14] , 
        \ScanLink78[13] , \ScanLink78[12] , \ScanLink78[11] , \ScanLink78[10] , 
        \ScanLink78[9] , \ScanLink78[8] , \ScanLink78[7] , \ScanLink78[6] , 
        \ScanLink78[5] , \ScanLink78[4] , \ScanLink78[3] , \ScanLink78[2] , 
        \ScanLink78[1] , \ScanLink78[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_15[31] , \wRegOut_6_15[30] , 
        \wRegOut_6_15[29] , \wRegOut_6_15[28] , \wRegOut_6_15[27] , 
        \wRegOut_6_15[26] , \wRegOut_6_15[25] , \wRegOut_6_15[24] , 
        \wRegOut_6_15[23] , \wRegOut_6_15[22] , \wRegOut_6_15[21] , 
        \wRegOut_6_15[20] , \wRegOut_6_15[19] , \wRegOut_6_15[18] , 
        \wRegOut_6_15[17] , \wRegOut_6_15[16] , \wRegOut_6_15[15] , 
        \wRegOut_6_15[14] , \wRegOut_6_15[13] , \wRegOut_6_15[12] , 
        \wRegOut_6_15[11] , \wRegOut_6_15[10] , \wRegOut_6_15[9] , 
        \wRegOut_6_15[8] , \wRegOut_6_15[7] , \wRegOut_6_15[6] , 
        \wRegOut_6_15[5] , \wRegOut_6_15[4] , \wRegOut_6_15[3] , 
        \wRegOut_6_15[2] , \wRegOut_6_15[1] , \wRegOut_6_15[0] }), .Enable1(
        \wRegEnTop_6_15[0] ), .Enable2(\wRegEnBot_6_15[0] ), .In1({
        \wRegInTop_6_15[31] , \wRegInTop_6_15[30] , \wRegInTop_6_15[29] , 
        \wRegInTop_6_15[28] , \wRegInTop_6_15[27] , \wRegInTop_6_15[26] , 
        \wRegInTop_6_15[25] , \wRegInTop_6_15[24] , \wRegInTop_6_15[23] , 
        \wRegInTop_6_15[22] , \wRegInTop_6_15[21] , \wRegInTop_6_15[20] , 
        \wRegInTop_6_15[19] , \wRegInTop_6_15[18] , \wRegInTop_6_15[17] , 
        \wRegInTop_6_15[16] , \wRegInTop_6_15[15] , \wRegInTop_6_15[14] , 
        \wRegInTop_6_15[13] , \wRegInTop_6_15[12] , \wRegInTop_6_15[11] , 
        \wRegInTop_6_15[10] , \wRegInTop_6_15[9] , \wRegInTop_6_15[8] , 
        \wRegInTop_6_15[7] , \wRegInTop_6_15[6] , \wRegInTop_6_15[5] , 
        \wRegInTop_6_15[4] , \wRegInTop_6_15[3] , \wRegInTop_6_15[2] , 
        \wRegInTop_6_15[1] , \wRegInTop_6_15[0] }), .In2({\wRegInBot_6_15[31] , 
        \wRegInBot_6_15[30] , \wRegInBot_6_15[29] , \wRegInBot_6_15[28] , 
        \wRegInBot_6_15[27] , \wRegInBot_6_15[26] , \wRegInBot_6_15[25] , 
        \wRegInBot_6_15[24] , \wRegInBot_6_15[23] , \wRegInBot_6_15[22] , 
        \wRegInBot_6_15[21] , \wRegInBot_6_15[20] , \wRegInBot_6_15[19] , 
        \wRegInBot_6_15[18] , \wRegInBot_6_15[17] , \wRegInBot_6_15[16] , 
        \wRegInBot_6_15[15] , \wRegInBot_6_15[14] , \wRegInBot_6_15[13] , 
        \wRegInBot_6_15[12] , \wRegInBot_6_15[11] , \wRegInBot_6_15[10] , 
        \wRegInBot_6_15[9] , \wRegInBot_6_15[8] , \wRegInBot_6_15[7] , 
        \wRegInBot_6_15[6] , \wRegInBot_6_15[5] , \wRegInBot_6_15[4] , 
        \wRegInBot_6_15[3] , \wRegInBot_6_15[2] , \wRegInBot_6_15[1] , 
        \wRegInBot_6_15[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_32 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink96[31] , \ScanLink96[30] , \ScanLink96[29] , 
        \ScanLink96[28] , \ScanLink96[27] , \ScanLink96[26] , \ScanLink96[25] , 
        \ScanLink96[24] , \ScanLink96[23] , \ScanLink96[22] , \ScanLink96[21] , 
        \ScanLink96[20] , \ScanLink96[19] , \ScanLink96[18] , \ScanLink96[17] , 
        \ScanLink96[16] , \ScanLink96[15] , \ScanLink96[14] , \ScanLink96[13] , 
        \ScanLink96[12] , \ScanLink96[11] , \ScanLink96[10] , \ScanLink96[9] , 
        \ScanLink96[8] , \ScanLink96[7] , \ScanLink96[6] , \ScanLink96[5] , 
        \ScanLink96[4] , \ScanLink96[3] , \ScanLink96[2] , \ScanLink96[1] , 
        \ScanLink96[0] }), .ScanOut({\ScanLink95[31] , \ScanLink95[30] , 
        \ScanLink95[29] , \ScanLink95[28] , \ScanLink95[27] , \ScanLink95[26] , 
        \ScanLink95[25] , \ScanLink95[24] , \ScanLink95[23] , \ScanLink95[22] , 
        \ScanLink95[21] , \ScanLink95[20] , \ScanLink95[19] , \ScanLink95[18] , 
        \ScanLink95[17] , \ScanLink95[16] , \ScanLink95[15] , \ScanLink95[14] , 
        \ScanLink95[13] , \ScanLink95[12] , \ScanLink95[11] , \ScanLink95[10] , 
        \ScanLink95[9] , \ScanLink95[8] , \ScanLink95[7] , \ScanLink95[6] , 
        \ScanLink95[5] , \ScanLink95[4] , \ScanLink95[3] , \ScanLink95[2] , 
        \ScanLink95[1] , \ScanLink95[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_32[31] , \wRegOut_6_32[30] , 
        \wRegOut_6_32[29] , \wRegOut_6_32[28] , \wRegOut_6_32[27] , 
        \wRegOut_6_32[26] , \wRegOut_6_32[25] , \wRegOut_6_32[24] , 
        \wRegOut_6_32[23] , \wRegOut_6_32[22] , \wRegOut_6_32[21] , 
        \wRegOut_6_32[20] , \wRegOut_6_32[19] , \wRegOut_6_32[18] , 
        \wRegOut_6_32[17] , \wRegOut_6_32[16] , \wRegOut_6_32[15] , 
        \wRegOut_6_32[14] , \wRegOut_6_32[13] , \wRegOut_6_32[12] , 
        \wRegOut_6_32[11] , \wRegOut_6_32[10] , \wRegOut_6_32[9] , 
        \wRegOut_6_32[8] , \wRegOut_6_32[7] , \wRegOut_6_32[6] , 
        \wRegOut_6_32[5] , \wRegOut_6_32[4] , \wRegOut_6_32[3] , 
        \wRegOut_6_32[2] , \wRegOut_6_32[1] , \wRegOut_6_32[0] }), .Enable1(
        \wRegEnTop_6_32[0] ), .Enable2(\wRegEnBot_6_32[0] ), .In1({
        \wRegInTop_6_32[31] , \wRegInTop_6_32[30] , \wRegInTop_6_32[29] , 
        \wRegInTop_6_32[28] , \wRegInTop_6_32[27] , \wRegInTop_6_32[26] , 
        \wRegInTop_6_32[25] , \wRegInTop_6_32[24] , \wRegInTop_6_32[23] , 
        \wRegInTop_6_32[22] , \wRegInTop_6_32[21] , \wRegInTop_6_32[20] , 
        \wRegInTop_6_32[19] , \wRegInTop_6_32[18] , \wRegInTop_6_32[17] , 
        \wRegInTop_6_32[16] , \wRegInTop_6_32[15] , \wRegInTop_6_32[14] , 
        \wRegInTop_6_32[13] , \wRegInTop_6_32[12] , \wRegInTop_6_32[11] , 
        \wRegInTop_6_32[10] , \wRegInTop_6_32[9] , \wRegInTop_6_32[8] , 
        \wRegInTop_6_32[7] , \wRegInTop_6_32[6] , \wRegInTop_6_32[5] , 
        \wRegInTop_6_32[4] , \wRegInTop_6_32[3] , \wRegInTop_6_32[2] , 
        \wRegInTop_6_32[1] , \wRegInTop_6_32[0] }), .In2({\wRegInBot_6_32[31] , 
        \wRegInBot_6_32[30] , \wRegInBot_6_32[29] , \wRegInBot_6_32[28] , 
        \wRegInBot_6_32[27] , \wRegInBot_6_32[26] , \wRegInBot_6_32[25] , 
        \wRegInBot_6_32[24] , \wRegInBot_6_32[23] , \wRegInBot_6_32[22] , 
        \wRegInBot_6_32[21] , \wRegInBot_6_32[20] , \wRegInBot_6_32[19] , 
        \wRegInBot_6_32[18] , \wRegInBot_6_32[17] , \wRegInBot_6_32[16] , 
        \wRegInBot_6_32[15] , \wRegInBot_6_32[14] , \wRegInBot_6_32[13] , 
        \wRegInBot_6_32[12] , \wRegInBot_6_32[11] , \wRegInBot_6_32[10] , 
        \wRegInBot_6_32[9] , \wRegInBot_6_32[8] , \wRegInBot_6_32[7] , 
        \wRegInBot_6_32[6] , \wRegInBot_6_32[5] , \wRegInBot_6_32[4] , 
        \wRegInBot_6_32[3] , \wRegInBot_6_32[2] , \wRegInBot_6_32[1] , 
        \wRegInBot_6_32[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink128[31] , \ScanLink128[30] , \ScanLink128[29] , 
        \ScanLink128[28] , \ScanLink128[27] , \ScanLink128[26] , 
        \ScanLink128[25] , \ScanLink128[24] , \ScanLink128[23] , 
        \ScanLink128[22] , \ScanLink128[21] , \ScanLink128[20] , 
        \ScanLink128[19] , \ScanLink128[18] , \ScanLink128[17] , 
        \ScanLink128[16] , \ScanLink128[15] , \ScanLink128[14] , 
        \ScanLink128[13] , \ScanLink128[12] , \ScanLink128[11] , 
        \ScanLink128[10] , \ScanLink128[9] , \ScanLink128[8] , 
        \ScanLink128[7] , \ScanLink128[6] , \ScanLink128[5] , \ScanLink128[4] , 
        \ScanLink128[3] , \ScanLink128[2] , \ScanLink128[1] , \ScanLink128[0] 
        }), .ScanOut({\ScanLink127[31] , \ScanLink127[30] , \ScanLink127[29] , 
        \ScanLink127[28] , \ScanLink127[27] , \ScanLink127[26] , 
        \ScanLink127[25] , \ScanLink127[24] , \ScanLink127[23] , 
        \ScanLink127[22] , \ScanLink127[21] , \ScanLink127[20] , 
        \ScanLink127[19] , \ScanLink127[18] , \ScanLink127[17] , 
        \ScanLink127[16] , \ScanLink127[15] , \ScanLink127[14] , 
        \ScanLink127[13] , \ScanLink127[12] , \ScanLink127[11] , 
        \ScanLink127[10] , \ScanLink127[9] , \ScanLink127[8] , 
        \ScanLink127[7] , \ScanLink127[6] , \ScanLink127[5] , \ScanLink127[4] , 
        \ScanLink127[3] , \ScanLink127[2] , \ScanLink127[1] , \ScanLink127[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_0[31] , 
        \wRegOut_7_0[30] , \wRegOut_7_0[29] , \wRegOut_7_0[28] , 
        \wRegOut_7_0[27] , \wRegOut_7_0[26] , \wRegOut_7_0[25] , 
        \wRegOut_7_0[24] , \wRegOut_7_0[23] , \wRegOut_7_0[22] , 
        \wRegOut_7_0[21] , \wRegOut_7_0[20] , \wRegOut_7_0[19] , 
        \wRegOut_7_0[18] , \wRegOut_7_0[17] , \wRegOut_7_0[16] , 
        \wRegOut_7_0[15] , \wRegOut_7_0[14] , \wRegOut_7_0[13] , 
        \wRegOut_7_0[12] , \wRegOut_7_0[11] , \wRegOut_7_0[10] , 
        \wRegOut_7_0[9] , \wRegOut_7_0[8] , \wRegOut_7_0[7] , \wRegOut_7_0[6] , 
        \wRegOut_7_0[5] , \wRegOut_7_0[4] , \wRegOut_7_0[3] , \wRegOut_7_0[2] , 
        \wRegOut_7_0[1] , \wRegOut_7_0[0] }), .Enable1(\wRegEnTop_7_0[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_0[31] , \wRegInTop_7_0[30] , 
        \wRegInTop_7_0[29] , \wRegInTop_7_0[28] , \wRegInTop_7_0[27] , 
        \wRegInTop_7_0[26] , \wRegInTop_7_0[25] , \wRegInTop_7_0[24] , 
        \wRegInTop_7_0[23] , \wRegInTop_7_0[22] , \wRegInTop_7_0[21] , 
        \wRegInTop_7_0[20] , \wRegInTop_7_0[19] , \wRegInTop_7_0[18] , 
        \wRegInTop_7_0[17] , \wRegInTop_7_0[16] , \wRegInTop_7_0[15] , 
        \wRegInTop_7_0[14] , \wRegInTop_7_0[13] , \wRegInTop_7_0[12] , 
        \wRegInTop_7_0[11] , \wRegInTop_7_0[10] , \wRegInTop_7_0[9] , 
        \wRegInTop_7_0[8] , \wRegInTop_7_0[7] , \wRegInTop_7_0[6] , 
        \wRegInTop_7_0[5] , \wRegInTop_7_0[4] , \wRegInTop_7_0[3] , 
        \wRegInTop_7_0[2] , \wRegInTop_7_0[1] , \wRegInTop_7_0[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_46 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink174[31] , \ScanLink174[30] , \ScanLink174[29] , 
        \ScanLink174[28] , \ScanLink174[27] , \ScanLink174[26] , 
        \ScanLink174[25] , \ScanLink174[24] , \ScanLink174[23] , 
        \ScanLink174[22] , \ScanLink174[21] , \ScanLink174[20] , 
        \ScanLink174[19] , \ScanLink174[18] , \ScanLink174[17] , 
        \ScanLink174[16] , \ScanLink174[15] , \ScanLink174[14] , 
        \ScanLink174[13] , \ScanLink174[12] , \ScanLink174[11] , 
        \ScanLink174[10] , \ScanLink174[9] , \ScanLink174[8] , 
        \ScanLink174[7] , \ScanLink174[6] , \ScanLink174[5] , \ScanLink174[4] , 
        \ScanLink174[3] , \ScanLink174[2] , \ScanLink174[1] , \ScanLink174[0] 
        }), .ScanOut({\ScanLink173[31] , \ScanLink173[30] , \ScanLink173[29] , 
        \ScanLink173[28] , \ScanLink173[27] , \ScanLink173[26] , 
        \ScanLink173[25] , \ScanLink173[24] , \ScanLink173[23] , 
        \ScanLink173[22] , \ScanLink173[21] , \ScanLink173[20] , 
        \ScanLink173[19] , \ScanLink173[18] , \ScanLink173[17] , 
        \ScanLink173[16] , \ScanLink173[15] , \ScanLink173[14] , 
        \ScanLink173[13] , \ScanLink173[12] , \ScanLink173[11] , 
        \ScanLink173[10] , \ScanLink173[9] , \ScanLink173[8] , 
        \ScanLink173[7] , \ScanLink173[6] , \ScanLink173[5] , \ScanLink173[4] , 
        \ScanLink173[3] , \ScanLink173[2] , \ScanLink173[1] , \ScanLink173[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_46[31] , 
        \wRegOut_7_46[30] , \wRegOut_7_46[29] , \wRegOut_7_46[28] , 
        \wRegOut_7_46[27] , \wRegOut_7_46[26] , \wRegOut_7_46[25] , 
        \wRegOut_7_46[24] , \wRegOut_7_46[23] , \wRegOut_7_46[22] , 
        \wRegOut_7_46[21] , \wRegOut_7_46[20] , \wRegOut_7_46[19] , 
        \wRegOut_7_46[18] , \wRegOut_7_46[17] , \wRegOut_7_46[16] , 
        \wRegOut_7_46[15] , \wRegOut_7_46[14] , \wRegOut_7_46[13] , 
        \wRegOut_7_46[12] , \wRegOut_7_46[11] , \wRegOut_7_46[10] , 
        \wRegOut_7_46[9] , \wRegOut_7_46[8] , \wRegOut_7_46[7] , 
        \wRegOut_7_46[6] , \wRegOut_7_46[5] , \wRegOut_7_46[4] , 
        \wRegOut_7_46[3] , \wRegOut_7_46[2] , \wRegOut_7_46[1] , 
        \wRegOut_7_46[0] }), .Enable1(\wRegEnTop_7_46[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_46[31] , \wRegInTop_7_46[30] , \wRegInTop_7_46[29] , 
        \wRegInTop_7_46[28] , \wRegInTop_7_46[27] , \wRegInTop_7_46[26] , 
        \wRegInTop_7_46[25] , \wRegInTop_7_46[24] , \wRegInTop_7_46[23] , 
        \wRegInTop_7_46[22] , \wRegInTop_7_46[21] , \wRegInTop_7_46[20] , 
        \wRegInTop_7_46[19] , \wRegInTop_7_46[18] , \wRegInTop_7_46[17] , 
        \wRegInTop_7_46[16] , \wRegInTop_7_46[15] , \wRegInTop_7_46[14] , 
        \wRegInTop_7_46[13] , \wRegInTop_7_46[12] , \wRegInTop_7_46[11] , 
        \wRegInTop_7_46[10] , \wRegInTop_7_46[9] , \wRegInTop_7_46[8] , 
        \wRegInTop_7_46[7] , \wRegInTop_7_46[6] , \wRegInTop_7_46[5] , 
        \wRegInTop_7_46[4] , \wRegInTop_7_46[3] , \wRegInTop_7_46[2] , 
        \wRegInTop_7_46[1] , \wRegInTop_7_46[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_47 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink111[31] , \ScanLink111[30] , \ScanLink111[29] , 
        \ScanLink111[28] , \ScanLink111[27] , \ScanLink111[26] , 
        \ScanLink111[25] , \ScanLink111[24] , \ScanLink111[23] , 
        \ScanLink111[22] , \ScanLink111[21] , \ScanLink111[20] , 
        \ScanLink111[19] , \ScanLink111[18] , \ScanLink111[17] , 
        \ScanLink111[16] , \ScanLink111[15] , \ScanLink111[14] , 
        \ScanLink111[13] , \ScanLink111[12] , \ScanLink111[11] , 
        \ScanLink111[10] , \ScanLink111[9] , \ScanLink111[8] , 
        \ScanLink111[7] , \ScanLink111[6] , \ScanLink111[5] , \ScanLink111[4] , 
        \ScanLink111[3] , \ScanLink111[2] , \ScanLink111[1] , \ScanLink111[0] 
        }), .ScanOut({\ScanLink110[31] , \ScanLink110[30] , \ScanLink110[29] , 
        \ScanLink110[28] , \ScanLink110[27] , \ScanLink110[26] , 
        \ScanLink110[25] , \ScanLink110[24] , \ScanLink110[23] , 
        \ScanLink110[22] , \ScanLink110[21] , \ScanLink110[20] , 
        \ScanLink110[19] , \ScanLink110[18] , \ScanLink110[17] , 
        \ScanLink110[16] , \ScanLink110[15] , \ScanLink110[14] , 
        \ScanLink110[13] , \ScanLink110[12] , \ScanLink110[11] , 
        \ScanLink110[10] , \ScanLink110[9] , \ScanLink110[8] , 
        \ScanLink110[7] , \ScanLink110[6] , \ScanLink110[5] , \ScanLink110[4] , 
        \ScanLink110[3] , \ScanLink110[2] , \ScanLink110[1] , \ScanLink110[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_47[31] , 
        \wRegOut_6_47[30] , \wRegOut_6_47[29] , \wRegOut_6_47[28] , 
        \wRegOut_6_47[27] , \wRegOut_6_47[26] , \wRegOut_6_47[25] , 
        \wRegOut_6_47[24] , \wRegOut_6_47[23] , \wRegOut_6_47[22] , 
        \wRegOut_6_47[21] , \wRegOut_6_47[20] , \wRegOut_6_47[19] , 
        \wRegOut_6_47[18] , \wRegOut_6_47[17] , \wRegOut_6_47[16] , 
        \wRegOut_6_47[15] , \wRegOut_6_47[14] , \wRegOut_6_47[13] , 
        \wRegOut_6_47[12] , \wRegOut_6_47[11] , \wRegOut_6_47[10] , 
        \wRegOut_6_47[9] , \wRegOut_6_47[8] , \wRegOut_6_47[7] , 
        \wRegOut_6_47[6] , \wRegOut_6_47[5] , \wRegOut_6_47[4] , 
        \wRegOut_6_47[3] , \wRegOut_6_47[2] , \wRegOut_6_47[1] , 
        \wRegOut_6_47[0] }), .Enable1(\wRegEnTop_6_47[0] ), .Enable2(
        \wRegEnBot_6_47[0] ), .In1({\wRegInTop_6_47[31] , \wRegInTop_6_47[30] , 
        \wRegInTop_6_47[29] , \wRegInTop_6_47[28] , \wRegInTop_6_47[27] , 
        \wRegInTop_6_47[26] , \wRegInTop_6_47[25] , \wRegInTop_6_47[24] , 
        \wRegInTop_6_47[23] , \wRegInTop_6_47[22] , \wRegInTop_6_47[21] , 
        \wRegInTop_6_47[20] , \wRegInTop_6_47[19] , \wRegInTop_6_47[18] , 
        \wRegInTop_6_47[17] , \wRegInTop_6_47[16] , \wRegInTop_6_47[15] , 
        \wRegInTop_6_47[14] , \wRegInTop_6_47[13] , \wRegInTop_6_47[12] , 
        \wRegInTop_6_47[11] , \wRegInTop_6_47[10] , \wRegInTop_6_47[9] , 
        \wRegInTop_6_47[8] , \wRegInTop_6_47[7] , \wRegInTop_6_47[6] , 
        \wRegInTop_6_47[5] , \wRegInTop_6_47[4] , \wRegInTop_6_47[3] , 
        \wRegInTop_6_47[2] , \wRegInTop_6_47[1] , \wRegInTop_6_47[0] }), .In2(
        {\wRegInBot_6_47[31] , \wRegInBot_6_47[30] , \wRegInBot_6_47[29] , 
        \wRegInBot_6_47[28] , \wRegInBot_6_47[27] , \wRegInBot_6_47[26] , 
        \wRegInBot_6_47[25] , \wRegInBot_6_47[24] , \wRegInBot_6_47[23] , 
        \wRegInBot_6_47[22] , \wRegInBot_6_47[21] , \wRegInBot_6_47[20] , 
        \wRegInBot_6_47[19] , \wRegInBot_6_47[18] , \wRegInBot_6_47[17] , 
        \wRegInBot_6_47[16] , \wRegInBot_6_47[15] , \wRegInBot_6_47[14] , 
        \wRegInBot_6_47[13] , \wRegInBot_6_47[12] , \wRegInBot_6_47[11] , 
        \wRegInBot_6_47[10] , \wRegInBot_6_47[9] , \wRegInBot_6_47[8] , 
        \wRegInBot_6_47[7] , \wRegInBot_6_47[6] , \wRegInBot_6_47[5] , 
        \wRegInBot_6_47[4] , \wRegInBot_6_47[3] , \wRegInBot_6_47[2] , 
        \wRegInBot_6_47[1] , \wRegInBot_6_47[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_28 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink156[31] , \ScanLink156[30] , \ScanLink156[29] , 
        \ScanLink156[28] , \ScanLink156[27] , \ScanLink156[26] , 
        \ScanLink156[25] , \ScanLink156[24] , \ScanLink156[23] , 
        \ScanLink156[22] , \ScanLink156[21] , \ScanLink156[20] , 
        \ScanLink156[19] , \ScanLink156[18] , \ScanLink156[17] , 
        \ScanLink156[16] , \ScanLink156[15] , \ScanLink156[14] , 
        \ScanLink156[13] , \ScanLink156[12] , \ScanLink156[11] , 
        \ScanLink156[10] , \ScanLink156[9] , \ScanLink156[8] , 
        \ScanLink156[7] , \ScanLink156[6] , \ScanLink156[5] , \ScanLink156[4] , 
        \ScanLink156[3] , \ScanLink156[2] , \ScanLink156[1] , \ScanLink156[0] 
        }), .ScanOut({\ScanLink155[31] , \ScanLink155[30] , \ScanLink155[29] , 
        \ScanLink155[28] , \ScanLink155[27] , \ScanLink155[26] , 
        \ScanLink155[25] , \ScanLink155[24] , \ScanLink155[23] , 
        \ScanLink155[22] , \ScanLink155[21] , \ScanLink155[20] , 
        \ScanLink155[19] , \ScanLink155[18] , \ScanLink155[17] , 
        \ScanLink155[16] , \ScanLink155[15] , \ScanLink155[14] , 
        \ScanLink155[13] , \ScanLink155[12] , \ScanLink155[11] , 
        \ScanLink155[10] , \ScanLink155[9] , \ScanLink155[8] , 
        \ScanLink155[7] , \ScanLink155[6] , \ScanLink155[5] , \ScanLink155[4] , 
        \ScanLink155[3] , \ScanLink155[2] , \ScanLink155[1] , \ScanLink155[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_28[31] , 
        \wRegOut_7_28[30] , \wRegOut_7_28[29] , \wRegOut_7_28[28] , 
        \wRegOut_7_28[27] , \wRegOut_7_28[26] , \wRegOut_7_28[25] , 
        \wRegOut_7_28[24] , \wRegOut_7_28[23] , \wRegOut_7_28[22] , 
        \wRegOut_7_28[21] , \wRegOut_7_28[20] , \wRegOut_7_28[19] , 
        \wRegOut_7_28[18] , \wRegOut_7_28[17] , \wRegOut_7_28[16] , 
        \wRegOut_7_28[15] , \wRegOut_7_28[14] , \wRegOut_7_28[13] , 
        \wRegOut_7_28[12] , \wRegOut_7_28[11] , \wRegOut_7_28[10] , 
        \wRegOut_7_28[9] , \wRegOut_7_28[8] , \wRegOut_7_28[7] , 
        \wRegOut_7_28[6] , \wRegOut_7_28[5] , \wRegOut_7_28[4] , 
        \wRegOut_7_28[3] , \wRegOut_7_28[2] , \wRegOut_7_28[1] , 
        \wRegOut_7_28[0] }), .Enable1(\wRegEnTop_7_28[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_28[31] , \wRegInTop_7_28[30] , \wRegInTop_7_28[29] , 
        \wRegInTop_7_28[28] , \wRegInTop_7_28[27] , \wRegInTop_7_28[26] , 
        \wRegInTop_7_28[25] , \wRegInTop_7_28[24] , \wRegInTop_7_28[23] , 
        \wRegInTop_7_28[22] , \wRegInTop_7_28[21] , \wRegInTop_7_28[20] , 
        \wRegInTop_7_28[19] , \wRegInTop_7_28[18] , \wRegInTop_7_28[17] , 
        \wRegInTop_7_28[16] , \wRegInTop_7_28[15] , \wRegInTop_7_28[14] , 
        \wRegInTop_7_28[13] , \wRegInTop_7_28[12] , \wRegInTop_7_28[11] , 
        \wRegInTop_7_28[10] , \wRegInTop_7_28[9] , \wRegInTop_7_28[8] , 
        \wRegInTop_7_28[7] , \wRegInTop_7_28[6] , \wRegInTop_7_28[5] , 
        \wRegInTop_7_28[4] , \wRegInTop_7_28[3] , \wRegInTop_7_28[2] , 
        \wRegInTop_7_28[1] , \wRegInTop_7_28[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_61 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink189[31] , \ScanLink189[30] , \ScanLink189[29] , 
        \ScanLink189[28] , \ScanLink189[27] , \ScanLink189[26] , 
        \ScanLink189[25] , \ScanLink189[24] , \ScanLink189[23] , 
        \ScanLink189[22] , \ScanLink189[21] , \ScanLink189[20] , 
        \ScanLink189[19] , \ScanLink189[18] , \ScanLink189[17] , 
        \ScanLink189[16] , \ScanLink189[15] , \ScanLink189[14] , 
        \ScanLink189[13] , \ScanLink189[12] , \ScanLink189[11] , 
        \ScanLink189[10] , \ScanLink189[9] , \ScanLink189[8] , 
        \ScanLink189[7] , \ScanLink189[6] , \ScanLink189[5] , \ScanLink189[4] , 
        \ScanLink189[3] , \ScanLink189[2] , \ScanLink189[1] , \ScanLink189[0] 
        }), .ScanOut({\ScanLink188[31] , \ScanLink188[30] , \ScanLink188[29] , 
        \ScanLink188[28] , \ScanLink188[27] , \ScanLink188[26] , 
        \ScanLink188[25] , \ScanLink188[24] , \ScanLink188[23] , 
        \ScanLink188[22] , \ScanLink188[21] , \ScanLink188[20] , 
        \ScanLink188[19] , \ScanLink188[18] , \ScanLink188[17] , 
        \ScanLink188[16] , \ScanLink188[15] , \ScanLink188[14] , 
        \ScanLink188[13] , \ScanLink188[12] , \ScanLink188[11] , 
        \ScanLink188[10] , \ScanLink188[9] , \ScanLink188[8] , 
        \ScanLink188[7] , \ScanLink188[6] , \ScanLink188[5] , \ScanLink188[4] , 
        \ScanLink188[3] , \ScanLink188[2] , \ScanLink188[1] , \ScanLink188[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_61[31] , 
        \wRegOut_7_61[30] , \wRegOut_7_61[29] , \wRegOut_7_61[28] , 
        \wRegOut_7_61[27] , \wRegOut_7_61[26] , \wRegOut_7_61[25] , 
        \wRegOut_7_61[24] , \wRegOut_7_61[23] , \wRegOut_7_61[22] , 
        \wRegOut_7_61[21] , \wRegOut_7_61[20] , \wRegOut_7_61[19] , 
        \wRegOut_7_61[18] , \wRegOut_7_61[17] , \wRegOut_7_61[16] , 
        \wRegOut_7_61[15] , \wRegOut_7_61[14] , \wRegOut_7_61[13] , 
        \wRegOut_7_61[12] , \wRegOut_7_61[11] , \wRegOut_7_61[10] , 
        \wRegOut_7_61[9] , \wRegOut_7_61[8] , \wRegOut_7_61[7] , 
        \wRegOut_7_61[6] , \wRegOut_7_61[5] , \wRegOut_7_61[4] , 
        \wRegOut_7_61[3] , \wRegOut_7_61[2] , \wRegOut_7_61[1] , 
        \wRegOut_7_61[0] }), .Enable1(\wRegEnTop_7_61[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_61[31] , \wRegInTop_7_61[30] , \wRegInTop_7_61[29] , 
        \wRegInTop_7_61[28] , \wRegInTop_7_61[27] , \wRegInTop_7_61[26] , 
        \wRegInTop_7_61[25] , \wRegInTop_7_61[24] , \wRegInTop_7_61[23] , 
        \wRegInTop_7_61[22] , \wRegInTop_7_61[21] , \wRegInTop_7_61[20] , 
        \wRegInTop_7_61[19] , \wRegInTop_7_61[18] , \wRegInTop_7_61[17] , 
        \wRegInTop_7_61[16] , \wRegInTop_7_61[15] , \wRegInTop_7_61[14] , 
        \wRegInTop_7_61[13] , \wRegInTop_7_61[12] , \wRegInTop_7_61[11] , 
        \wRegInTop_7_61[10] , \wRegInTop_7_61[9] , \wRegInTop_7_61[8] , 
        \wRegInTop_7_61[7] , \wRegInTop_7_61[6] , \wRegInTop_7_61[5] , 
        \wRegInTop_7_61[4] , \wRegInTop_7_61[3] , \wRegInTop_7_61[2] , 
        \wRegInTop_7_61[1] , \wRegInTop_7_61[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_53[0] ), .P_In({\wRegOut_6_53[31] , 
        \wRegOut_6_53[30] , \wRegOut_6_53[29] , \wRegOut_6_53[28] , 
        \wRegOut_6_53[27] , \wRegOut_6_53[26] , \wRegOut_6_53[25] , 
        \wRegOut_6_53[24] , \wRegOut_6_53[23] , \wRegOut_6_53[22] , 
        \wRegOut_6_53[21] , \wRegOut_6_53[20] , \wRegOut_6_53[19] , 
        \wRegOut_6_53[18] , \wRegOut_6_53[17] , \wRegOut_6_53[16] , 
        \wRegOut_6_53[15] , \wRegOut_6_53[14] , \wRegOut_6_53[13] , 
        \wRegOut_6_53[12] , \wRegOut_6_53[11] , \wRegOut_6_53[10] , 
        \wRegOut_6_53[9] , \wRegOut_6_53[8] , \wRegOut_6_53[7] , 
        \wRegOut_6_53[6] , \wRegOut_6_53[5] , \wRegOut_6_53[4] , 
        \wRegOut_6_53[3] , \wRegOut_6_53[2] , \wRegOut_6_53[1] , 
        \wRegOut_6_53[0] }), .P_Out({\wRegInBot_6_53[31] , 
        \wRegInBot_6_53[30] , \wRegInBot_6_53[29] , \wRegInBot_6_53[28] , 
        \wRegInBot_6_53[27] , \wRegInBot_6_53[26] , \wRegInBot_6_53[25] , 
        \wRegInBot_6_53[24] , \wRegInBot_6_53[23] , \wRegInBot_6_53[22] , 
        \wRegInBot_6_53[21] , \wRegInBot_6_53[20] , \wRegInBot_6_53[19] , 
        \wRegInBot_6_53[18] , \wRegInBot_6_53[17] , \wRegInBot_6_53[16] , 
        \wRegInBot_6_53[15] , \wRegInBot_6_53[14] , \wRegInBot_6_53[13] , 
        \wRegInBot_6_53[12] , \wRegInBot_6_53[11] , \wRegInBot_6_53[10] , 
        \wRegInBot_6_53[9] , \wRegInBot_6_53[8] , \wRegInBot_6_53[7] , 
        \wRegInBot_6_53[6] , \wRegInBot_6_53[5] , \wRegInBot_6_53[4] , 
        \wRegInBot_6_53[3] , \wRegInBot_6_53[2] , \wRegInBot_6_53[1] , 
        \wRegInBot_6_53[0] }), .L_WR(\wRegEnTop_7_106[0] ), .L_In({
        \wRegOut_7_106[31] , \wRegOut_7_106[30] , \wRegOut_7_106[29] , 
        \wRegOut_7_106[28] , \wRegOut_7_106[27] , \wRegOut_7_106[26] , 
        \wRegOut_7_106[25] , \wRegOut_7_106[24] , \wRegOut_7_106[23] , 
        \wRegOut_7_106[22] , \wRegOut_7_106[21] , \wRegOut_7_106[20] , 
        \wRegOut_7_106[19] , \wRegOut_7_106[18] , \wRegOut_7_106[17] , 
        \wRegOut_7_106[16] , \wRegOut_7_106[15] , \wRegOut_7_106[14] , 
        \wRegOut_7_106[13] , \wRegOut_7_106[12] , \wRegOut_7_106[11] , 
        \wRegOut_7_106[10] , \wRegOut_7_106[9] , \wRegOut_7_106[8] , 
        \wRegOut_7_106[7] , \wRegOut_7_106[6] , \wRegOut_7_106[5] , 
        \wRegOut_7_106[4] , \wRegOut_7_106[3] , \wRegOut_7_106[2] , 
        \wRegOut_7_106[1] , \wRegOut_7_106[0] }), .L_Out({
        \wRegInTop_7_106[31] , \wRegInTop_7_106[30] , \wRegInTop_7_106[29] , 
        \wRegInTop_7_106[28] , \wRegInTop_7_106[27] , \wRegInTop_7_106[26] , 
        \wRegInTop_7_106[25] , \wRegInTop_7_106[24] , \wRegInTop_7_106[23] , 
        \wRegInTop_7_106[22] , \wRegInTop_7_106[21] , \wRegInTop_7_106[20] , 
        \wRegInTop_7_106[19] , \wRegInTop_7_106[18] , \wRegInTop_7_106[17] , 
        \wRegInTop_7_106[16] , \wRegInTop_7_106[15] , \wRegInTop_7_106[14] , 
        \wRegInTop_7_106[13] , \wRegInTop_7_106[12] , \wRegInTop_7_106[11] , 
        \wRegInTop_7_106[10] , \wRegInTop_7_106[9] , \wRegInTop_7_106[8] , 
        \wRegInTop_7_106[7] , \wRegInTop_7_106[6] , \wRegInTop_7_106[5] , 
        \wRegInTop_7_106[4] , \wRegInTop_7_106[3] , \wRegInTop_7_106[2] , 
        \wRegInTop_7_106[1] , \wRegInTop_7_106[0] }), .R_WR(
        \wRegEnTop_7_107[0] ), .R_In({\wRegOut_7_107[31] , \wRegOut_7_107[30] , 
        \wRegOut_7_107[29] , \wRegOut_7_107[28] , \wRegOut_7_107[27] , 
        \wRegOut_7_107[26] , \wRegOut_7_107[25] , \wRegOut_7_107[24] , 
        \wRegOut_7_107[23] , \wRegOut_7_107[22] , \wRegOut_7_107[21] , 
        \wRegOut_7_107[20] , \wRegOut_7_107[19] , \wRegOut_7_107[18] , 
        \wRegOut_7_107[17] , \wRegOut_7_107[16] , \wRegOut_7_107[15] , 
        \wRegOut_7_107[14] , \wRegOut_7_107[13] , \wRegOut_7_107[12] , 
        \wRegOut_7_107[11] , \wRegOut_7_107[10] , \wRegOut_7_107[9] , 
        \wRegOut_7_107[8] , \wRegOut_7_107[7] , \wRegOut_7_107[6] , 
        \wRegOut_7_107[5] , \wRegOut_7_107[4] , \wRegOut_7_107[3] , 
        \wRegOut_7_107[2] , \wRegOut_7_107[1] , \wRegOut_7_107[0] }), .R_Out({
        \wRegInTop_7_107[31] , \wRegInTop_7_107[30] , \wRegInTop_7_107[29] , 
        \wRegInTop_7_107[28] , \wRegInTop_7_107[27] , \wRegInTop_7_107[26] , 
        \wRegInTop_7_107[25] , \wRegInTop_7_107[24] , \wRegInTop_7_107[23] , 
        \wRegInTop_7_107[22] , \wRegInTop_7_107[21] , \wRegInTop_7_107[20] , 
        \wRegInTop_7_107[19] , \wRegInTop_7_107[18] , \wRegInTop_7_107[17] , 
        \wRegInTop_7_107[16] , \wRegInTop_7_107[15] , \wRegInTop_7_107[14] , 
        \wRegInTop_7_107[13] , \wRegInTop_7_107[12] , \wRegInTop_7_107[11] , 
        \wRegInTop_7_107[10] , \wRegInTop_7_107[9] , \wRegInTop_7_107[8] , 
        \wRegInTop_7_107[7] , \wRegInTop_7_107[6] , \wRegInTop_7_107[5] , 
        \wRegInTop_7_107[4] , \wRegInTop_7_107[3] , \wRegInTop_7_107[2] , 
        \wRegInTop_7_107[1] , \wRegInTop_7_107[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_33 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink161[31] , \ScanLink161[30] , \ScanLink161[29] , 
        \ScanLink161[28] , \ScanLink161[27] , \ScanLink161[26] , 
        \ScanLink161[25] , \ScanLink161[24] , \ScanLink161[23] , 
        \ScanLink161[22] , \ScanLink161[21] , \ScanLink161[20] , 
        \ScanLink161[19] , \ScanLink161[18] , \ScanLink161[17] , 
        \ScanLink161[16] , \ScanLink161[15] , \ScanLink161[14] , 
        \ScanLink161[13] , \ScanLink161[12] , \ScanLink161[11] , 
        \ScanLink161[10] , \ScanLink161[9] , \ScanLink161[8] , 
        \ScanLink161[7] , \ScanLink161[6] , \ScanLink161[5] , \ScanLink161[4] , 
        \ScanLink161[3] , \ScanLink161[2] , \ScanLink161[1] , \ScanLink161[0] 
        }), .ScanOut({\ScanLink160[31] , \ScanLink160[30] , \ScanLink160[29] , 
        \ScanLink160[28] , \ScanLink160[27] , \ScanLink160[26] , 
        \ScanLink160[25] , \ScanLink160[24] , \ScanLink160[23] , 
        \ScanLink160[22] , \ScanLink160[21] , \ScanLink160[20] , 
        \ScanLink160[19] , \ScanLink160[18] , \ScanLink160[17] , 
        \ScanLink160[16] , \ScanLink160[15] , \ScanLink160[14] , 
        \ScanLink160[13] , \ScanLink160[12] , \ScanLink160[11] , 
        \ScanLink160[10] , \ScanLink160[9] , \ScanLink160[8] , 
        \ScanLink160[7] , \ScanLink160[6] , \ScanLink160[5] , \ScanLink160[4] , 
        \ScanLink160[3] , \ScanLink160[2] , \ScanLink160[1] , \ScanLink160[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_33[31] , 
        \wRegOut_7_33[30] , \wRegOut_7_33[29] , \wRegOut_7_33[28] , 
        \wRegOut_7_33[27] , \wRegOut_7_33[26] , \wRegOut_7_33[25] , 
        \wRegOut_7_33[24] , \wRegOut_7_33[23] , \wRegOut_7_33[22] , 
        \wRegOut_7_33[21] , \wRegOut_7_33[20] , \wRegOut_7_33[19] , 
        \wRegOut_7_33[18] , \wRegOut_7_33[17] , \wRegOut_7_33[16] , 
        \wRegOut_7_33[15] , \wRegOut_7_33[14] , \wRegOut_7_33[13] , 
        \wRegOut_7_33[12] , \wRegOut_7_33[11] , \wRegOut_7_33[10] , 
        \wRegOut_7_33[9] , \wRegOut_7_33[8] , \wRegOut_7_33[7] , 
        \wRegOut_7_33[6] , \wRegOut_7_33[5] , \wRegOut_7_33[4] , 
        \wRegOut_7_33[3] , \wRegOut_7_33[2] , \wRegOut_7_33[1] , 
        \wRegOut_7_33[0] }), .Enable1(\wRegEnTop_7_33[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_33[31] , \wRegInTop_7_33[30] , \wRegInTop_7_33[29] , 
        \wRegInTop_7_33[28] , \wRegInTop_7_33[27] , \wRegInTop_7_33[26] , 
        \wRegInTop_7_33[25] , \wRegInTop_7_33[24] , \wRegInTop_7_33[23] , 
        \wRegInTop_7_33[22] , \wRegInTop_7_33[21] , \wRegInTop_7_33[20] , 
        \wRegInTop_7_33[19] , \wRegInTop_7_33[18] , \wRegInTop_7_33[17] , 
        \wRegInTop_7_33[16] , \wRegInTop_7_33[15] , \wRegInTop_7_33[14] , 
        \wRegInTop_7_33[13] , \wRegInTop_7_33[12] , \wRegInTop_7_33[11] , 
        \wRegInTop_7_33[10] , \wRegInTop_7_33[9] , \wRegInTop_7_33[8] , 
        \wRegInTop_7_33[7] , \wRegInTop_7_33[6] , \wRegInTop_7_33[5] , 
        \wRegInTop_7_33[4] , \wRegInTop_7_33[3] , \wRegInTop_7_33[2] , 
        \wRegInTop_7_33[1] , \wRegInTop_7_33[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_84 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink212[31] , \ScanLink212[30] , \ScanLink212[29] , 
        \ScanLink212[28] , \ScanLink212[27] , \ScanLink212[26] , 
        \ScanLink212[25] , \ScanLink212[24] , \ScanLink212[23] , 
        \ScanLink212[22] , \ScanLink212[21] , \ScanLink212[20] , 
        \ScanLink212[19] , \ScanLink212[18] , \ScanLink212[17] , 
        \ScanLink212[16] , \ScanLink212[15] , \ScanLink212[14] , 
        \ScanLink212[13] , \ScanLink212[12] , \ScanLink212[11] , 
        \ScanLink212[10] , \ScanLink212[9] , \ScanLink212[8] , 
        \ScanLink212[7] , \ScanLink212[6] , \ScanLink212[5] , \ScanLink212[4] , 
        \ScanLink212[3] , \ScanLink212[2] , \ScanLink212[1] , \ScanLink212[0] 
        }), .ScanOut({\ScanLink211[31] , \ScanLink211[30] , \ScanLink211[29] , 
        \ScanLink211[28] , \ScanLink211[27] , \ScanLink211[26] , 
        \ScanLink211[25] , \ScanLink211[24] , \ScanLink211[23] , 
        \ScanLink211[22] , \ScanLink211[21] , \ScanLink211[20] , 
        \ScanLink211[19] , \ScanLink211[18] , \ScanLink211[17] , 
        \ScanLink211[16] , \ScanLink211[15] , \ScanLink211[14] , 
        \ScanLink211[13] , \ScanLink211[12] , \ScanLink211[11] , 
        \ScanLink211[10] , \ScanLink211[9] , \ScanLink211[8] , 
        \ScanLink211[7] , \ScanLink211[6] , \ScanLink211[5] , \ScanLink211[4] , 
        \ScanLink211[3] , \ScanLink211[2] , \ScanLink211[1] , \ScanLink211[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_84[31] , 
        \wRegOut_7_84[30] , \wRegOut_7_84[29] , \wRegOut_7_84[28] , 
        \wRegOut_7_84[27] , \wRegOut_7_84[26] , \wRegOut_7_84[25] , 
        \wRegOut_7_84[24] , \wRegOut_7_84[23] , \wRegOut_7_84[22] , 
        \wRegOut_7_84[21] , \wRegOut_7_84[20] , \wRegOut_7_84[19] , 
        \wRegOut_7_84[18] , \wRegOut_7_84[17] , \wRegOut_7_84[16] , 
        \wRegOut_7_84[15] , \wRegOut_7_84[14] , \wRegOut_7_84[13] , 
        \wRegOut_7_84[12] , \wRegOut_7_84[11] , \wRegOut_7_84[10] , 
        \wRegOut_7_84[9] , \wRegOut_7_84[8] , \wRegOut_7_84[7] , 
        \wRegOut_7_84[6] , \wRegOut_7_84[5] , \wRegOut_7_84[4] , 
        \wRegOut_7_84[3] , \wRegOut_7_84[2] , \wRegOut_7_84[1] , 
        \wRegOut_7_84[0] }), .Enable1(\wRegEnTop_7_84[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_84[31] , \wRegInTop_7_84[30] , \wRegInTop_7_84[29] , 
        \wRegInTop_7_84[28] , \wRegInTop_7_84[27] , \wRegInTop_7_84[26] , 
        \wRegInTop_7_84[25] , \wRegInTop_7_84[24] , \wRegInTop_7_84[23] , 
        \wRegInTop_7_84[22] , \wRegInTop_7_84[21] , \wRegInTop_7_84[20] , 
        \wRegInTop_7_84[19] , \wRegInTop_7_84[18] , \wRegInTop_7_84[17] , 
        \wRegInTop_7_84[16] , \wRegInTop_7_84[15] , \wRegInTop_7_84[14] , 
        \wRegInTop_7_84[13] , \wRegInTop_7_84[12] , \wRegInTop_7_84[11] , 
        \wRegInTop_7_84[10] , \wRegInTop_7_84[9] , \wRegInTop_7_84[8] , 
        \wRegInTop_7_84[7] , \wRegInTop_7_84[6] , \wRegInTop_7_84[5] , 
        \wRegInTop_7_84[4] , \wRegInTop_7_84[3] , \wRegInTop_7_84[2] , 
        \wRegInTop_7_84[1] , \wRegInTop_7_84[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_4[0] ), .P_In({\wRegOut_3_4[31] , 
        \wRegOut_3_4[30] , \wRegOut_3_4[29] , \wRegOut_3_4[28] , 
        \wRegOut_3_4[27] , \wRegOut_3_4[26] , \wRegOut_3_4[25] , 
        \wRegOut_3_4[24] , \wRegOut_3_4[23] , \wRegOut_3_4[22] , 
        \wRegOut_3_4[21] , \wRegOut_3_4[20] , \wRegOut_3_4[19] , 
        \wRegOut_3_4[18] , \wRegOut_3_4[17] , \wRegOut_3_4[16] , 
        \wRegOut_3_4[15] , \wRegOut_3_4[14] , \wRegOut_3_4[13] , 
        \wRegOut_3_4[12] , \wRegOut_3_4[11] , \wRegOut_3_4[10] , 
        \wRegOut_3_4[9] , \wRegOut_3_4[8] , \wRegOut_3_4[7] , \wRegOut_3_4[6] , 
        \wRegOut_3_4[5] , \wRegOut_3_4[4] , \wRegOut_3_4[3] , \wRegOut_3_4[2] , 
        \wRegOut_3_4[1] , \wRegOut_3_4[0] }), .P_Out({\wRegInBot_3_4[31] , 
        \wRegInBot_3_4[30] , \wRegInBot_3_4[29] , \wRegInBot_3_4[28] , 
        \wRegInBot_3_4[27] , \wRegInBot_3_4[26] , \wRegInBot_3_4[25] , 
        \wRegInBot_3_4[24] , \wRegInBot_3_4[23] , \wRegInBot_3_4[22] , 
        \wRegInBot_3_4[21] , \wRegInBot_3_4[20] , \wRegInBot_3_4[19] , 
        \wRegInBot_3_4[18] , \wRegInBot_3_4[17] , \wRegInBot_3_4[16] , 
        \wRegInBot_3_4[15] , \wRegInBot_3_4[14] , \wRegInBot_3_4[13] , 
        \wRegInBot_3_4[12] , \wRegInBot_3_4[11] , \wRegInBot_3_4[10] , 
        \wRegInBot_3_4[9] , \wRegInBot_3_4[8] , \wRegInBot_3_4[7] , 
        \wRegInBot_3_4[6] , \wRegInBot_3_4[5] , \wRegInBot_3_4[4] , 
        \wRegInBot_3_4[3] , \wRegInBot_3_4[2] , \wRegInBot_3_4[1] , 
        \wRegInBot_3_4[0] }), .L_WR(\wRegEnTop_4_8[0] ), .L_In({
        \wRegOut_4_8[31] , \wRegOut_4_8[30] , \wRegOut_4_8[29] , 
        \wRegOut_4_8[28] , \wRegOut_4_8[27] , \wRegOut_4_8[26] , 
        \wRegOut_4_8[25] , \wRegOut_4_8[24] , \wRegOut_4_8[23] , 
        \wRegOut_4_8[22] , \wRegOut_4_8[21] , \wRegOut_4_8[20] , 
        \wRegOut_4_8[19] , \wRegOut_4_8[18] , \wRegOut_4_8[17] , 
        \wRegOut_4_8[16] , \wRegOut_4_8[15] , \wRegOut_4_8[14] , 
        \wRegOut_4_8[13] , \wRegOut_4_8[12] , \wRegOut_4_8[11] , 
        \wRegOut_4_8[10] , \wRegOut_4_8[9] , \wRegOut_4_8[8] , 
        \wRegOut_4_8[7] , \wRegOut_4_8[6] , \wRegOut_4_8[5] , \wRegOut_4_8[4] , 
        \wRegOut_4_8[3] , \wRegOut_4_8[2] , \wRegOut_4_8[1] , \wRegOut_4_8[0] 
        }), .L_Out({\wRegInTop_4_8[31] , \wRegInTop_4_8[30] , 
        \wRegInTop_4_8[29] , \wRegInTop_4_8[28] , \wRegInTop_4_8[27] , 
        \wRegInTop_4_8[26] , \wRegInTop_4_8[25] , \wRegInTop_4_8[24] , 
        \wRegInTop_4_8[23] , \wRegInTop_4_8[22] , \wRegInTop_4_8[21] , 
        \wRegInTop_4_8[20] , \wRegInTop_4_8[19] , \wRegInTop_4_8[18] , 
        \wRegInTop_4_8[17] , \wRegInTop_4_8[16] , \wRegInTop_4_8[15] , 
        \wRegInTop_4_8[14] , \wRegInTop_4_8[13] , \wRegInTop_4_8[12] , 
        \wRegInTop_4_8[11] , \wRegInTop_4_8[10] , \wRegInTop_4_8[9] , 
        \wRegInTop_4_8[8] , \wRegInTop_4_8[7] , \wRegInTop_4_8[6] , 
        \wRegInTop_4_8[5] , \wRegInTop_4_8[4] , \wRegInTop_4_8[3] , 
        \wRegInTop_4_8[2] , \wRegInTop_4_8[1] , \wRegInTop_4_8[0] }), .R_WR(
        \wRegEnTop_4_9[0] ), .R_In({\wRegOut_4_9[31] , \wRegOut_4_9[30] , 
        \wRegOut_4_9[29] , \wRegOut_4_9[28] , \wRegOut_4_9[27] , 
        \wRegOut_4_9[26] , \wRegOut_4_9[25] , \wRegOut_4_9[24] , 
        \wRegOut_4_9[23] , \wRegOut_4_9[22] , \wRegOut_4_9[21] , 
        \wRegOut_4_9[20] , \wRegOut_4_9[19] , \wRegOut_4_9[18] , 
        \wRegOut_4_9[17] , \wRegOut_4_9[16] , \wRegOut_4_9[15] , 
        \wRegOut_4_9[14] , \wRegOut_4_9[13] , \wRegOut_4_9[12] , 
        \wRegOut_4_9[11] , \wRegOut_4_9[10] , \wRegOut_4_9[9] , 
        \wRegOut_4_9[8] , \wRegOut_4_9[7] , \wRegOut_4_9[6] , \wRegOut_4_9[5] , 
        \wRegOut_4_9[4] , \wRegOut_4_9[3] , \wRegOut_4_9[2] , \wRegOut_4_9[1] , 
        \wRegOut_4_9[0] }), .R_Out({\wRegInTop_4_9[31] , \wRegInTop_4_9[30] , 
        \wRegInTop_4_9[29] , \wRegInTop_4_9[28] , \wRegInTop_4_9[27] , 
        \wRegInTop_4_9[26] , \wRegInTop_4_9[25] , \wRegInTop_4_9[24] , 
        \wRegInTop_4_9[23] , \wRegInTop_4_9[22] , \wRegInTop_4_9[21] , 
        \wRegInTop_4_9[20] , \wRegInTop_4_9[19] , \wRegInTop_4_9[18] , 
        \wRegInTop_4_9[17] , \wRegInTop_4_9[16] , \wRegInTop_4_9[15] , 
        \wRegInTop_4_9[14] , \wRegInTop_4_9[13] , \wRegInTop_4_9[12] , 
        \wRegInTop_4_9[11] , \wRegInTop_4_9[10] , \wRegInTop_4_9[9] , 
        \wRegInTop_4_9[8] , \wRegInTop_4_9[7] , \wRegInTop_4_9[6] , 
        \wRegInTop_4_9[5] , \wRegInTop_4_9[4] , \wRegInTop_4_9[3] , 
        \wRegInTop_4_9[2] , \wRegInTop_4_9[1] , \wRegInTop_4_9[0] }) );
    BHeap_Node_WIDTH32 BHN_6_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_2[0] ), .P_In({\wRegOut_6_2[31] , 
        \wRegOut_6_2[30] , \wRegOut_6_2[29] , \wRegOut_6_2[28] , 
        \wRegOut_6_2[27] , \wRegOut_6_2[26] , \wRegOut_6_2[25] , 
        \wRegOut_6_2[24] , \wRegOut_6_2[23] , \wRegOut_6_2[22] , 
        \wRegOut_6_2[21] , \wRegOut_6_2[20] , \wRegOut_6_2[19] , 
        \wRegOut_6_2[18] , \wRegOut_6_2[17] , \wRegOut_6_2[16] , 
        \wRegOut_6_2[15] , \wRegOut_6_2[14] , \wRegOut_6_2[13] , 
        \wRegOut_6_2[12] , \wRegOut_6_2[11] , \wRegOut_6_2[10] , 
        \wRegOut_6_2[9] , \wRegOut_6_2[8] , \wRegOut_6_2[7] , \wRegOut_6_2[6] , 
        \wRegOut_6_2[5] , \wRegOut_6_2[4] , \wRegOut_6_2[3] , \wRegOut_6_2[2] , 
        \wRegOut_6_2[1] , \wRegOut_6_2[0] }), .P_Out({\wRegInBot_6_2[31] , 
        \wRegInBot_6_2[30] , \wRegInBot_6_2[29] , \wRegInBot_6_2[28] , 
        \wRegInBot_6_2[27] , \wRegInBot_6_2[26] , \wRegInBot_6_2[25] , 
        \wRegInBot_6_2[24] , \wRegInBot_6_2[23] , \wRegInBot_6_2[22] , 
        \wRegInBot_6_2[21] , \wRegInBot_6_2[20] , \wRegInBot_6_2[19] , 
        \wRegInBot_6_2[18] , \wRegInBot_6_2[17] , \wRegInBot_6_2[16] , 
        \wRegInBot_6_2[15] , \wRegInBot_6_2[14] , \wRegInBot_6_2[13] , 
        \wRegInBot_6_2[12] , \wRegInBot_6_2[11] , \wRegInBot_6_2[10] , 
        \wRegInBot_6_2[9] , \wRegInBot_6_2[8] , \wRegInBot_6_2[7] , 
        \wRegInBot_6_2[6] , \wRegInBot_6_2[5] , \wRegInBot_6_2[4] , 
        \wRegInBot_6_2[3] , \wRegInBot_6_2[2] , \wRegInBot_6_2[1] , 
        \wRegInBot_6_2[0] }), .L_WR(\wRegEnTop_7_4[0] ), .L_In({
        \wRegOut_7_4[31] , \wRegOut_7_4[30] , \wRegOut_7_4[29] , 
        \wRegOut_7_4[28] , \wRegOut_7_4[27] , \wRegOut_7_4[26] , 
        \wRegOut_7_4[25] , \wRegOut_7_4[24] , \wRegOut_7_4[23] , 
        \wRegOut_7_4[22] , \wRegOut_7_4[21] , \wRegOut_7_4[20] , 
        \wRegOut_7_4[19] , \wRegOut_7_4[18] , \wRegOut_7_4[17] , 
        \wRegOut_7_4[16] , \wRegOut_7_4[15] , \wRegOut_7_4[14] , 
        \wRegOut_7_4[13] , \wRegOut_7_4[12] , \wRegOut_7_4[11] , 
        \wRegOut_7_4[10] , \wRegOut_7_4[9] , \wRegOut_7_4[8] , 
        \wRegOut_7_4[7] , \wRegOut_7_4[6] , \wRegOut_7_4[5] , \wRegOut_7_4[4] , 
        \wRegOut_7_4[3] , \wRegOut_7_4[2] , \wRegOut_7_4[1] , \wRegOut_7_4[0] 
        }), .L_Out({\wRegInTop_7_4[31] , \wRegInTop_7_4[30] , 
        \wRegInTop_7_4[29] , \wRegInTop_7_4[28] , \wRegInTop_7_4[27] , 
        \wRegInTop_7_4[26] , \wRegInTop_7_4[25] , \wRegInTop_7_4[24] , 
        \wRegInTop_7_4[23] , \wRegInTop_7_4[22] , \wRegInTop_7_4[21] , 
        \wRegInTop_7_4[20] , \wRegInTop_7_4[19] , \wRegInTop_7_4[18] , 
        \wRegInTop_7_4[17] , \wRegInTop_7_4[16] , \wRegInTop_7_4[15] , 
        \wRegInTop_7_4[14] , \wRegInTop_7_4[13] , \wRegInTop_7_4[12] , 
        \wRegInTop_7_4[11] , \wRegInTop_7_4[10] , \wRegInTop_7_4[9] , 
        \wRegInTop_7_4[8] , \wRegInTop_7_4[7] , \wRegInTop_7_4[6] , 
        \wRegInTop_7_4[5] , \wRegInTop_7_4[4] , \wRegInTop_7_4[3] , 
        \wRegInTop_7_4[2] , \wRegInTop_7_4[1] , \wRegInTop_7_4[0] }), .R_WR(
        \wRegEnTop_7_5[0] ), .R_In({\wRegOut_7_5[31] , \wRegOut_7_5[30] , 
        \wRegOut_7_5[29] , \wRegOut_7_5[28] , \wRegOut_7_5[27] , 
        \wRegOut_7_5[26] , \wRegOut_7_5[25] , \wRegOut_7_5[24] , 
        \wRegOut_7_5[23] , \wRegOut_7_5[22] , \wRegOut_7_5[21] , 
        \wRegOut_7_5[20] , \wRegOut_7_5[19] , \wRegOut_7_5[18] , 
        \wRegOut_7_5[17] , \wRegOut_7_5[16] , \wRegOut_7_5[15] , 
        \wRegOut_7_5[14] , \wRegOut_7_5[13] , \wRegOut_7_5[12] , 
        \wRegOut_7_5[11] , \wRegOut_7_5[10] , \wRegOut_7_5[9] , 
        \wRegOut_7_5[8] , \wRegOut_7_5[7] , \wRegOut_7_5[6] , \wRegOut_7_5[5] , 
        \wRegOut_7_5[4] , \wRegOut_7_5[3] , \wRegOut_7_5[2] , \wRegOut_7_5[1] , 
        \wRegOut_7_5[0] }), .R_Out({\wRegInTop_7_5[31] , \wRegInTop_7_5[30] , 
        \wRegInTop_7_5[29] , \wRegInTop_7_5[28] , \wRegInTop_7_5[27] , 
        \wRegInTop_7_5[26] , \wRegInTop_7_5[25] , \wRegInTop_7_5[24] , 
        \wRegInTop_7_5[23] , \wRegInTop_7_5[22] , \wRegInTop_7_5[21] , 
        \wRegInTop_7_5[20] , \wRegInTop_7_5[19] , \wRegInTop_7_5[18] , 
        \wRegInTop_7_5[17] , \wRegInTop_7_5[16] , \wRegInTop_7_5[15] , 
        \wRegInTop_7_5[14] , \wRegInTop_7_5[13] , \wRegInTop_7_5[12] , 
        \wRegInTop_7_5[11] , \wRegInTop_7_5[10] , \wRegInTop_7_5[9] , 
        \wRegInTop_7_5[8] , \wRegInTop_7_5[7] , \wRegInTop_7_5[6] , 
        \wRegInTop_7_5[5] , \wRegInTop_7_5[4] , \wRegInTop_7_5[3] , 
        \wRegInTop_7_5[2] , \wRegInTop_7_5[1] , \wRegInTop_7_5[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_60 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink124[31] , \ScanLink124[30] , \ScanLink124[29] , 
        \ScanLink124[28] , \ScanLink124[27] , \ScanLink124[26] , 
        \ScanLink124[25] , \ScanLink124[24] , \ScanLink124[23] , 
        \ScanLink124[22] , \ScanLink124[21] , \ScanLink124[20] , 
        \ScanLink124[19] , \ScanLink124[18] , \ScanLink124[17] , 
        \ScanLink124[16] , \ScanLink124[15] , \ScanLink124[14] , 
        \ScanLink124[13] , \ScanLink124[12] , \ScanLink124[11] , 
        \ScanLink124[10] , \ScanLink124[9] , \ScanLink124[8] , 
        \ScanLink124[7] , \ScanLink124[6] , \ScanLink124[5] , \ScanLink124[4] , 
        \ScanLink124[3] , \ScanLink124[2] , \ScanLink124[1] , \ScanLink124[0] 
        }), .ScanOut({\ScanLink123[31] , \ScanLink123[30] , \ScanLink123[29] , 
        \ScanLink123[28] , \ScanLink123[27] , \ScanLink123[26] , 
        \ScanLink123[25] , \ScanLink123[24] , \ScanLink123[23] , 
        \ScanLink123[22] , \ScanLink123[21] , \ScanLink123[20] , 
        \ScanLink123[19] , \ScanLink123[18] , \ScanLink123[17] , 
        \ScanLink123[16] , \ScanLink123[15] , \ScanLink123[14] , 
        \ScanLink123[13] , \ScanLink123[12] , \ScanLink123[11] , 
        \ScanLink123[10] , \ScanLink123[9] , \ScanLink123[8] , 
        \ScanLink123[7] , \ScanLink123[6] , \ScanLink123[5] , \ScanLink123[4] , 
        \ScanLink123[3] , \ScanLink123[2] , \ScanLink123[1] , \ScanLink123[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_60[31] , 
        \wRegOut_6_60[30] , \wRegOut_6_60[29] , \wRegOut_6_60[28] , 
        \wRegOut_6_60[27] , \wRegOut_6_60[26] , \wRegOut_6_60[25] , 
        \wRegOut_6_60[24] , \wRegOut_6_60[23] , \wRegOut_6_60[22] , 
        \wRegOut_6_60[21] , \wRegOut_6_60[20] , \wRegOut_6_60[19] , 
        \wRegOut_6_60[18] , \wRegOut_6_60[17] , \wRegOut_6_60[16] , 
        \wRegOut_6_60[15] , \wRegOut_6_60[14] , \wRegOut_6_60[13] , 
        \wRegOut_6_60[12] , \wRegOut_6_60[11] , \wRegOut_6_60[10] , 
        \wRegOut_6_60[9] , \wRegOut_6_60[8] , \wRegOut_6_60[7] , 
        \wRegOut_6_60[6] , \wRegOut_6_60[5] , \wRegOut_6_60[4] , 
        \wRegOut_6_60[3] , \wRegOut_6_60[2] , \wRegOut_6_60[1] , 
        \wRegOut_6_60[0] }), .Enable1(\wRegEnTop_6_60[0] ), .Enable2(
        \wRegEnBot_6_60[0] ), .In1({\wRegInTop_6_60[31] , \wRegInTop_6_60[30] , 
        \wRegInTop_6_60[29] , \wRegInTop_6_60[28] , \wRegInTop_6_60[27] , 
        \wRegInTop_6_60[26] , \wRegInTop_6_60[25] , \wRegInTop_6_60[24] , 
        \wRegInTop_6_60[23] , \wRegInTop_6_60[22] , \wRegInTop_6_60[21] , 
        \wRegInTop_6_60[20] , \wRegInTop_6_60[19] , \wRegInTop_6_60[18] , 
        \wRegInTop_6_60[17] , \wRegInTop_6_60[16] , \wRegInTop_6_60[15] , 
        \wRegInTop_6_60[14] , \wRegInTop_6_60[13] , \wRegInTop_6_60[12] , 
        \wRegInTop_6_60[11] , \wRegInTop_6_60[10] , \wRegInTop_6_60[9] , 
        \wRegInTop_6_60[8] , \wRegInTop_6_60[7] , \wRegInTop_6_60[6] , 
        \wRegInTop_6_60[5] , \wRegInTop_6_60[4] , \wRegInTop_6_60[3] , 
        \wRegInTop_6_60[2] , \wRegInTop_6_60[1] , \wRegInTop_6_60[0] }), .In2(
        {\wRegInBot_6_60[31] , \wRegInBot_6_60[30] , \wRegInBot_6_60[29] , 
        \wRegInBot_6_60[28] , \wRegInBot_6_60[27] , \wRegInBot_6_60[26] , 
        \wRegInBot_6_60[25] , \wRegInBot_6_60[24] , \wRegInBot_6_60[23] , 
        \wRegInBot_6_60[22] , \wRegInBot_6_60[21] , \wRegInBot_6_60[20] , 
        \wRegInBot_6_60[19] , \wRegInBot_6_60[18] , \wRegInBot_6_60[17] , 
        \wRegInBot_6_60[16] , \wRegInBot_6_60[15] , \wRegInBot_6_60[14] , 
        \wRegInBot_6_60[13] , \wRegInBot_6_60[12] , \wRegInBot_6_60[11] , 
        \wRegInBot_6_60[10] , \wRegInBot_6_60[9] , \wRegInBot_6_60[8] , 
        \wRegInBot_6_60[7] , \wRegInBot_6_60[6] , \wRegInBot_6_60[5] , 
        \wRegInBot_6_60[4] , \wRegInBot_6_60[3] , \wRegInBot_6_60[2] , 
        \wRegInBot_6_60[1] , \wRegInBot_6_60[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink142[31] , \ScanLink142[30] , \ScanLink142[29] , 
        \ScanLink142[28] , \ScanLink142[27] , \ScanLink142[26] , 
        \ScanLink142[25] , \ScanLink142[24] , \ScanLink142[23] , 
        \ScanLink142[22] , \ScanLink142[21] , \ScanLink142[20] , 
        \ScanLink142[19] , \ScanLink142[18] , \ScanLink142[17] , 
        \ScanLink142[16] , \ScanLink142[15] , \ScanLink142[14] , 
        \ScanLink142[13] , \ScanLink142[12] , \ScanLink142[11] , 
        \ScanLink142[10] , \ScanLink142[9] , \ScanLink142[8] , 
        \ScanLink142[7] , \ScanLink142[6] , \ScanLink142[5] , \ScanLink142[4] , 
        \ScanLink142[3] , \ScanLink142[2] , \ScanLink142[1] , \ScanLink142[0] 
        }), .ScanOut({\ScanLink141[31] , \ScanLink141[30] , \ScanLink141[29] , 
        \ScanLink141[28] , \ScanLink141[27] , \ScanLink141[26] , 
        \ScanLink141[25] , \ScanLink141[24] , \ScanLink141[23] , 
        \ScanLink141[22] , \ScanLink141[21] , \ScanLink141[20] , 
        \ScanLink141[19] , \ScanLink141[18] , \ScanLink141[17] , 
        \ScanLink141[16] , \ScanLink141[15] , \ScanLink141[14] , 
        \ScanLink141[13] , \ScanLink141[12] , \ScanLink141[11] , 
        \ScanLink141[10] , \ScanLink141[9] , \ScanLink141[8] , 
        \ScanLink141[7] , \ScanLink141[6] , \ScanLink141[5] , \ScanLink141[4] , 
        \ScanLink141[3] , \ScanLink141[2] , \ScanLink141[1] , \ScanLink141[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_14[31] , 
        \wRegOut_7_14[30] , \wRegOut_7_14[29] , \wRegOut_7_14[28] , 
        \wRegOut_7_14[27] , \wRegOut_7_14[26] , \wRegOut_7_14[25] , 
        \wRegOut_7_14[24] , \wRegOut_7_14[23] , \wRegOut_7_14[22] , 
        \wRegOut_7_14[21] , \wRegOut_7_14[20] , \wRegOut_7_14[19] , 
        \wRegOut_7_14[18] , \wRegOut_7_14[17] , \wRegOut_7_14[16] , 
        \wRegOut_7_14[15] , \wRegOut_7_14[14] , \wRegOut_7_14[13] , 
        \wRegOut_7_14[12] , \wRegOut_7_14[11] , \wRegOut_7_14[10] , 
        \wRegOut_7_14[9] , \wRegOut_7_14[8] , \wRegOut_7_14[7] , 
        \wRegOut_7_14[6] , \wRegOut_7_14[5] , \wRegOut_7_14[4] , 
        \wRegOut_7_14[3] , \wRegOut_7_14[2] , \wRegOut_7_14[1] , 
        \wRegOut_7_14[0] }), .Enable1(\wRegEnTop_7_14[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_14[31] , \wRegInTop_7_14[30] , \wRegInTop_7_14[29] , 
        \wRegInTop_7_14[28] , \wRegInTop_7_14[27] , \wRegInTop_7_14[26] , 
        \wRegInTop_7_14[25] , \wRegInTop_7_14[24] , \wRegInTop_7_14[23] , 
        \wRegInTop_7_14[22] , \wRegInTop_7_14[21] , \wRegInTop_7_14[20] , 
        \wRegInTop_7_14[19] , \wRegInTop_7_14[18] , \wRegInTop_7_14[17] , 
        \wRegInTop_7_14[16] , \wRegInTop_7_14[15] , \wRegInTop_7_14[14] , 
        \wRegInTop_7_14[13] , \wRegInTop_7_14[12] , \wRegInTop_7_14[11] , 
        \wRegInTop_7_14[10] , \wRegInTop_7_14[9] , \wRegInTop_7_14[8] , 
        \wRegInTop_7_14[7] , \wRegInTop_7_14[6] , \wRegInTop_7_14[5] , 
        \wRegInTop_7_14[4] , \wRegInTop_7_14[3] , \wRegInTop_7_14[2] , 
        \wRegInTop_7_14[1] , \wRegInTop_7_14[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_127 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink255[31] , \ScanLink255[30] , \ScanLink255[29] , 
        \ScanLink255[28] , \ScanLink255[27] , \ScanLink255[26] , 
        \ScanLink255[25] , \ScanLink255[24] , \ScanLink255[23] , 
        \ScanLink255[22] , \ScanLink255[21] , \ScanLink255[20] , 
        \ScanLink255[19] , \ScanLink255[18] , \ScanLink255[17] , 
        \ScanLink255[16] , \ScanLink255[15] , \ScanLink255[14] , 
        \ScanLink255[13] , \ScanLink255[12] , \ScanLink255[11] , 
        \ScanLink255[10] , \ScanLink255[9] , \ScanLink255[8] , 
        \ScanLink255[7] , \ScanLink255[6] , \ScanLink255[5] , \ScanLink255[4] , 
        \ScanLink255[3] , \ScanLink255[2] , \ScanLink255[1] , \ScanLink255[0] 
        }), .ScanOut({\ScanLink254[31] , \ScanLink254[30] , \ScanLink254[29] , 
        \ScanLink254[28] , \ScanLink254[27] , \ScanLink254[26] , 
        \ScanLink254[25] , \ScanLink254[24] , \ScanLink254[23] , 
        \ScanLink254[22] , \ScanLink254[21] , \ScanLink254[20] , 
        \ScanLink254[19] , \ScanLink254[18] , \ScanLink254[17] , 
        \ScanLink254[16] , \ScanLink254[15] , \ScanLink254[14] , 
        \ScanLink254[13] , \ScanLink254[12] , \ScanLink254[11] , 
        \ScanLink254[10] , \ScanLink254[9] , \ScanLink254[8] , 
        \ScanLink254[7] , \ScanLink254[6] , \ScanLink254[5] , \ScanLink254[4] , 
        \ScanLink254[3] , \ScanLink254[2] , \ScanLink254[1] , \ScanLink254[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_127[31] , 
        \wRegOut_7_127[30] , \wRegOut_7_127[29] , \wRegOut_7_127[28] , 
        \wRegOut_7_127[27] , \wRegOut_7_127[26] , \wRegOut_7_127[25] , 
        \wRegOut_7_127[24] , \wRegOut_7_127[23] , \wRegOut_7_127[22] , 
        \wRegOut_7_127[21] , \wRegOut_7_127[20] , \wRegOut_7_127[19] , 
        \wRegOut_7_127[18] , \wRegOut_7_127[17] , \wRegOut_7_127[16] , 
        \wRegOut_7_127[15] , \wRegOut_7_127[14] , \wRegOut_7_127[13] , 
        \wRegOut_7_127[12] , \wRegOut_7_127[11] , \wRegOut_7_127[10] , 
        \wRegOut_7_127[9] , \wRegOut_7_127[8] , \wRegOut_7_127[7] , 
        \wRegOut_7_127[6] , \wRegOut_7_127[5] , \wRegOut_7_127[4] , 
        \wRegOut_7_127[3] , \wRegOut_7_127[2] , \wRegOut_7_127[1] , 
        \wRegOut_7_127[0] }), .Enable1(\wRegEnTop_7_127[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_127[31] , \wRegInTop_7_127[30] , 
        \wRegInTop_7_127[29] , \wRegInTop_7_127[28] , \wRegInTop_7_127[27] , 
        \wRegInTop_7_127[26] , \wRegInTop_7_127[25] , \wRegInTop_7_127[24] , 
        \wRegInTop_7_127[23] , \wRegInTop_7_127[22] , \wRegInTop_7_127[21] , 
        \wRegInTop_7_127[20] , \wRegInTop_7_127[19] , \wRegInTop_7_127[18] , 
        \wRegInTop_7_127[17] , \wRegInTop_7_127[16] , \wRegInTop_7_127[15] , 
        \wRegInTop_7_127[14] , \wRegInTop_7_127[13] , \wRegInTop_7_127[12] , 
        \wRegInTop_7_127[11] , \wRegInTop_7_127[10] , \wRegInTop_7_127[9] , 
        \wRegInTop_7_127[8] , \wRegInTop_7_127[7] , \wRegInTop_7_127[6] , 
        \wRegInTop_7_127[5] , \wRegInTop_7_127[4] , \wRegInTop_7_127[3] , 
        \wRegInTop_7_127[2] , \wRegInTop_7_127[1] , \wRegInTop_7_127[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_48[0] ), .P_In({\wRegOut_6_48[31] , 
        \wRegOut_6_48[30] , \wRegOut_6_48[29] , \wRegOut_6_48[28] , 
        \wRegOut_6_48[27] , \wRegOut_6_48[26] , \wRegOut_6_48[25] , 
        \wRegOut_6_48[24] , \wRegOut_6_48[23] , \wRegOut_6_48[22] , 
        \wRegOut_6_48[21] , \wRegOut_6_48[20] , \wRegOut_6_48[19] , 
        \wRegOut_6_48[18] , \wRegOut_6_48[17] , \wRegOut_6_48[16] , 
        \wRegOut_6_48[15] , \wRegOut_6_48[14] , \wRegOut_6_48[13] , 
        \wRegOut_6_48[12] , \wRegOut_6_48[11] , \wRegOut_6_48[10] , 
        \wRegOut_6_48[9] , \wRegOut_6_48[8] , \wRegOut_6_48[7] , 
        \wRegOut_6_48[6] , \wRegOut_6_48[5] , \wRegOut_6_48[4] , 
        \wRegOut_6_48[3] , \wRegOut_6_48[2] , \wRegOut_6_48[1] , 
        \wRegOut_6_48[0] }), .P_Out({\wRegInBot_6_48[31] , 
        \wRegInBot_6_48[30] , \wRegInBot_6_48[29] , \wRegInBot_6_48[28] , 
        \wRegInBot_6_48[27] , \wRegInBot_6_48[26] , \wRegInBot_6_48[25] , 
        \wRegInBot_6_48[24] , \wRegInBot_6_48[23] , \wRegInBot_6_48[22] , 
        \wRegInBot_6_48[21] , \wRegInBot_6_48[20] , \wRegInBot_6_48[19] , 
        \wRegInBot_6_48[18] , \wRegInBot_6_48[17] , \wRegInBot_6_48[16] , 
        \wRegInBot_6_48[15] , \wRegInBot_6_48[14] , \wRegInBot_6_48[13] , 
        \wRegInBot_6_48[12] , \wRegInBot_6_48[11] , \wRegInBot_6_48[10] , 
        \wRegInBot_6_48[9] , \wRegInBot_6_48[8] , \wRegInBot_6_48[7] , 
        \wRegInBot_6_48[6] , \wRegInBot_6_48[5] , \wRegInBot_6_48[4] , 
        \wRegInBot_6_48[3] , \wRegInBot_6_48[2] , \wRegInBot_6_48[1] , 
        \wRegInBot_6_48[0] }), .L_WR(\wRegEnTop_7_96[0] ), .L_In({
        \wRegOut_7_96[31] , \wRegOut_7_96[30] , \wRegOut_7_96[29] , 
        \wRegOut_7_96[28] , \wRegOut_7_96[27] , \wRegOut_7_96[26] , 
        \wRegOut_7_96[25] , \wRegOut_7_96[24] , \wRegOut_7_96[23] , 
        \wRegOut_7_96[22] , \wRegOut_7_96[21] , \wRegOut_7_96[20] , 
        \wRegOut_7_96[19] , \wRegOut_7_96[18] , \wRegOut_7_96[17] , 
        \wRegOut_7_96[16] , \wRegOut_7_96[15] , \wRegOut_7_96[14] , 
        \wRegOut_7_96[13] , \wRegOut_7_96[12] , \wRegOut_7_96[11] , 
        \wRegOut_7_96[10] , \wRegOut_7_96[9] , \wRegOut_7_96[8] , 
        \wRegOut_7_96[7] , \wRegOut_7_96[6] , \wRegOut_7_96[5] , 
        \wRegOut_7_96[4] , \wRegOut_7_96[3] , \wRegOut_7_96[2] , 
        \wRegOut_7_96[1] , \wRegOut_7_96[0] }), .L_Out({\wRegInTop_7_96[31] , 
        \wRegInTop_7_96[30] , \wRegInTop_7_96[29] , \wRegInTop_7_96[28] , 
        \wRegInTop_7_96[27] , \wRegInTop_7_96[26] , \wRegInTop_7_96[25] , 
        \wRegInTop_7_96[24] , \wRegInTop_7_96[23] , \wRegInTop_7_96[22] , 
        \wRegInTop_7_96[21] , \wRegInTop_7_96[20] , \wRegInTop_7_96[19] , 
        \wRegInTop_7_96[18] , \wRegInTop_7_96[17] , \wRegInTop_7_96[16] , 
        \wRegInTop_7_96[15] , \wRegInTop_7_96[14] , \wRegInTop_7_96[13] , 
        \wRegInTop_7_96[12] , \wRegInTop_7_96[11] , \wRegInTop_7_96[10] , 
        \wRegInTop_7_96[9] , \wRegInTop_7_96[8] , \wRegInTop_7_96[7] , 
        \wRegInTop_7_96[6] , \wRegInTop_7_96[5] , \wRegInTop_7_96[4] , 
        \wRegInTop_7_96[3] , \wRegInTop_7_96[2] , \wRegInTop_7_96[1] , 
        \wRegInTop_7_96[0] }), .R_WR(\wRegEnTop_7_97[0] ), .R_In({
        \wRegOut_7_97[31] , \wRegOut_7_97[30] , \wRegOut_7_97[29] , 
        \wRegOut_7_97[28] , \wRegOut_7_97[27] , \wRegOut_7_97[26] , 
        \wRegOut_7_97[25] , \wRegOut_7_97[24] , \wRegOut_7_97[23] , 
        \wRegOut_7_97[22] , \wRegOut_7_97[21] , \wRegOut_7_97[20] , 
        \wRegOut_7_97[19] , \wRegOut_7_97[18] , \wRegOut_7_97[17] , 
        \wRegOut_7_97[16] , \wRegOut_7_97[15] , \wRegOut_7_97[14] , 
        \wRegOut_7_97[13] , \wRegOut_7_97[12] , \wRegOut_7_97[11] , 
        \wRegOut_7_97[10] , \wRegOut_7_97[9] , \wRegOut_7_97[8] , 
        \wRegOut_7_97[7] , \wRegOut_7_97[6] , \wRegOut_7_97[5] , 
        \wRegOut_7_97[4] , \wRegOut_7_97[3] , \wRegOut_7_97[2] , 
        \wRegOut_7_97[1] , \wRegOut_7_97[0] }), .R_Out({\wRegInTop_7_97[31] , 
        \wRegInTop_7_97[30] , \wRegInTop_7_97[29] , \wRegInTop_7_97[28] , 
        \wRegInTop_7_97[27] , \wRegInTop_7_97[26] , \wRegInTop_7_97[25] , 
        \wRegInTop_7_97[24] , \wRegInTop_7_97[23] , \wRegInTop_7_97[22] , 
        \wRegInTop_7_97[21] , \wRegInTop_7_97[20] , \wRegInTop_7_97[19] , 
        \wRegInTop_7_97[18] , \wRegInTop_7_97[17] , \wRegInTop_7_97[16] , 
        \wRegInTop_7_97[15] , \wRegInTop_7_97[14] , \wRegInTop_7_97[13] , 
        \wRegInTop_7_97[12] , \wRegInTop_7_97[11] , \wRegInTop_7_97[10] , 
        \wRegInTop_7_97[9] , \wRegInTop_7_97[8] , \wRegInTop_7_97[7] , 
        \wRegInTop_7_97[6] , \wRegInTop_7_97[5] , \wRegInTop_7_97[4] , 
        \wRegInTop_7_97[3] , \wRegInTop_7_97[2] , \wRegInTop_7_97[1] , 
        \wRegInTop_7_97[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_100 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink228[31] , \ScanLink228[30] , \ScanLink228[29] , 
        \ScanLink228[28] , \ScanLink228[27] , \ScanLink228[26] , 
        \ScanLink228[25] , \ScanLink228[24] , \ScanLink228[23] , 
        \ScanLink228[22] , \ScanLink228[21] , \ScanLink228[20] , 
        \ScanLink228[19] , \ScanLink228[18] , \ScanLink228[17] , 
        \ScanLink228[16] , \ScanLink228[15] , \ScanLink228[14] , 
        \ScanLink228[13] , \ScanLink228[12] , \ScanLink228[11] , 
        \ScanLink228[10] , \ScanLink228[9] , \ScanLink228[8] , 
        \ScanLink228[7] , \ScanLink228[6] , \ScanLink228[5] , \ScanLink228[4] , 
        \ScanLink228[3] , \ScanLink228[2] , \ScanLink228[1] , \ScanLink228[0] 
        }), .ScanOut({\ScanLink227[31] , \ScanLink227[30] , \ScanLink227[29] , 
        \ScanLink227[28] , \ScanLink227[27] , \ScanLink227[26] , 
        \ScanLink227[25] , \ScanLink227[24] , \ScanLink227[23] , 
        \ScanLink227[22] , \ScanLink227[21] , \ScanLink227[20] , 
        \ScanLink227[19] , \ScanLink227[18] , \ScanLink227[17] , 
        \ScanLink227[16] , \ScanLink227[15] , \ScanLink227[14] , 
        \ScanLink227[13] , \ScanLink227[12] , \ScanLink227[11] , 
        \ScanLink227[10] , \ScanLink227[9] , \ScanLink227[8] , 
        \ScanLink227[7] , \ScanLink227[6] , \ScanLink227[5] , \ScanLink227[4] , 
        \ScanLink227[3] , \ScanLink227[2] , \ScanLink227[1] , \ScanLink227[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_100[31] , 
        \wRegOut_7_100[30] , \wRegOut_7_100[29] , \wRegOut_7_100[28] , 
        \wRegOut_7_100[27] , \wRegOut_7_100[26] , \wRegOut_7_100[25] , 
        \wRegOut_7_100[24] , \wRegOut_7_100[23] , \wRegOut_7_100[22] , 
        \wRegOut_7_100[21] , \wRegOut_7_100[20] , \wRegOut_7_100[19] , 
        \wRegOut_7_100[18] , \wRegOut_7_100[17] , \wRegOut_7_100[16] , 
        \wRegOut_7_100[15] , \wRegOut_7_100[14] , \wRegOut_7_100[13] , 
        \wRegOut_7_100[12] , \wRegOut_7_100[11] , \wRegOut_7_100[10] , 
        \wRegOut_7_100[9] , \wRegOut_7_100[8] , \wRegOut_7_100[7] , 
        \wRegOut_7_100[6] , \wRegOut_7_100[5] , \wRegOut_7_100[4] , 
        \wRegOut_7_100[3] , \wRegOut_7_100[2] , \wRegOut_7_100[1] , 
        \wRegOut_7_100[0] }), .Enable1(\wRegEnTop_7_100[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_100[31] , \wRegInTop_7_100[30] , 
        \wRegInTop_7_100[29] , \wRegInTop_7_100[28] , \wRegInTop_7_100[27] , 
        \wRegInTop_7_100[26] , \wRegInTop_7_100[25] , \wRegInTop_7_100[24] , 
        \wRegInTop_7_100[23] , \wRegInTop_7_100[22] , \wRegInTop_7_100[21] , 
        \wRegInTop_7_100[20] , \wRegInTop_7_100[19] , \wRegInTop_7_100[18] , 
        \wRegInTop_7_100[17] , \wRegInTop_7_100[16] , \wRegInTop_7_100[15] , 
        \wRegInTop_7_100[14] , \wRegInTop_7_100[13] , \wRegInTop_7_100[12] , 
        \wRegInTop_7_100[11] , \wRegInTop_7_100[10] , \wRegInTop_7_100[9] , 
        \wRegInTop_7_100[8] , \wRegInTop_7_100[7] , \wRegInTop_7_100[6] , 
        \wRegInTop_7_100[5] , \wRegInTop_7_100[4] , \wRegInTop_7_100[3] , 
        \wRegInTop_7_100[2] , \wRegInTop_7_100[1] , \wRegInTop_7_100[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_CtrlReg_WIDTH32 BHCR_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_1[0] ), 
        .Out(\wCtrlOut_0[0] ), .Enable(\wEnable_0[0] ) );
    BHeap_Node_WIDTH32 BHN_5_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_16[0] ), .P_In({\wRegOut_5_16[31] , 
        \wRegOut_5_16[30] , \wRegOut_5_16[29] , \wRegOut_5_16[28] , 
        \wRegOut_5_16[27] , \wRegOut_5_16[26] , \wRegOut_5_16[25] , 
        \wRegOut_5_16[24] , \wRegOut_5_16[23] , \wRegOut_5_16[22] , 
        \wRegOut_5_16[21] , \wRegOut_5_16[20] , \wRegOut_5_16[19] , 
        \wRegOut_5_16[18] , \wRegOut_5_16[17] , \wRegOut_5_16[16] , 
        \wRegOut_5_16[15] , \wRegOut_5_16[14] , \wRegOut_5_16[13] , 
        \wRegOut_5_16[12] , \wRegOut_5_16[11] , \wRegOut_5_16[10] , 
        \wRegOut_5_16[9] , \wRegOut_5_16[8] , \wRegOut_5_16[7] , 
        \wRegOut_5_16[6] , \wRegOut_5_16[5] , \wRegOut_5_16[4] , 
        \wRegOut_5_16[3] , \wRegOut_5_16[2] , \wRegOut_5_16[1] , 
        \wRegOut_5_16[0] }), .P_Out({\wRegInBot_5_16[31] , 
        \wRegInBot_5_16[30] , \wRegInBot_5_16[29] , \wRegInBot_5_16[28] , 
        \wRegInBot_5_16[27] , \wRegInBot_5_16[26] , \wRegInBot_5_16[25] , 
        \wRegInBot_5_16[24] , \wRegInBot_5_16[23] , \wRegInBot_5_16[22] , 
        \wRegInBot_5_16[21] , \wRegInBot_5_16[20] , \wRegInBot_5_16[19] , 
        \wRegInBot_5_16[18] , \wRegInBot_5_16[17] , \wRegInBot_5_16[16] , 
        \wRegInBot_5_16[15] , \wRegInBot_5_16[14] , \wRegInBot_5_16[13] , 
        \wRegInBot_5_16[12] , \wRegInBot_5_16[11] , \wRegInBot_5_16[10] , 
        \wRegInBot_5_16[9] , \wRegInBot_5_16[8] , \wRegInBot_5_16[7] , 
        \wRegInBot_5_16[6] , \wRegInBot_5_16[5] , \wRegInBot_5_16[4] , 
        \wRegInBot_5_16[3] , \wRegInBot_5_16[2] , \wRegInBot_5_16[1] , 
        \wRegInBot_5_16[0] }), .L_WR(\wRegEnTop_6_32[0] ), .L_In({
        \wRegOut_6_32[31] , \wRegOut_6_32[30] , \wRegOut_6_32[29] , 
        \wRegOut_6_32[28] , \wRegOut_6_32[27] , \wRegOut_6_32[26] , 
        \wRegOut_6_32[25] , \wRegOut_6_32[24] , \wRegOut_6_32[23] , 
        \wRegOut_6_32[22] , \wRegOut_6_32[21] , \wRegOut_6_32[20] , 
        \wRegOut_6_32[19] , \wRegOut_6_32[18] , \wRegOut_6_32[17] , 
        \wRegOut_6_32[16] , \wRegOut_6_32[15] , \wRegOut_6_32[14] , 
        \wRegOut_6_32[13] , \wRegOut_6_32[12] , \wRegOut_6_32[11] , 
        \wRegOut_6_32[10] , \wRegOut_6_32[9] , \wRegOut_6_32[8] , 
        \wRegOut_6_32[7] , \wRegOut_6_32[6] , \wRegOut_6_32[5] , 
        \wRegOut_6_32[4] , \wRegOut_6_32[3] , \wRegOut_6_32[2] , 
        \wRegOut_6_32[1] , \wRegOut_6_32[0] }), .L_Out({\wRegInTop_6_32[31] , 
        \wRegInTop_6_32[30] , \wRegInTop_6_32[29] , \wRegInTop_6_32[28] , 
        \wRegInTop_6_32[27] , \wRegInTop_6_32[26] , \wRegInTop_6_32[25] , 
        \wRegInTop_6_32[24] , \wRegInTop_6_32[23] , \wRegInTop_6_32[22] , 
        \wRegInTop_6_32[21] , \wRegInTop_6_32[20] , \wRegInTop_6_32[19] , 
        \wRegInTop_6_32[18] , \wRegInTop_6_32[17] , \wRegInTop_6_32[16] , 
        \wRegInTop_6_32[15] , \wRegInTop_6_32[14] , \wRegInTop_6_32[13] , 
        \wRegInTop_6_32[12] , \wRegInTop_6_32[11] , \wRegInTop_6_32[10] , 
        \wRegInTop_6_32[9] , \wRegInTop_6_32[8] , \wRegInTop_6_32[7] , 
        \wRegInTop_6_32[6] , \wRegInTop_6_32[5] , \wRegInTop_6_32[4] , 
        \wRegInTop_6_32[3] , \wRegInTop_6_32[2] , \wRegInTop_6_32[1] , 
        \wRegInTop_6_32[0] }), .R_WR(\wRegEnTop_6_33[0] ), .R_In({
        \wRegOut_6_33[31] , \wRegOut_6_33[30] , \wRegOut_6_33[29] , 
        \wRegOut_6_33[28] , \wRegOut_6_33[27] , \wRegOut_6_33[26] , 
        \wRegOut_6_33[25] , \wRegOut_6_33[24] , \wRegOut_6_33[23] , 
        \wRegOut_6_33[22] , \wRegOut_6_33[21] , \wRegOut_6_33[20] , 
        \wRegOut_6_33[19] , \wRegOut_6_33[18] , \wRegOut_6_33[17] , 
        \wRegOut_6_33[16] , \wRegOut_6_33[15] , \wRegOut_6_33[14] , 
        \wRegOut_6_33[13] , \wRegOut_6_33[12] , \wRegOut_6_33[11] , 
        \wRegOut_6_33[10] , \wRegOut_6_33[9] , \wRegOut_6_33[8] , 
        \wRegOut_6_33[7] , \wRegOut_6_33[6] , \wRegOut_6_33[5] , 
        \wRegOut_6_33[4] , \wRegOut_6_33[3] , \wRegOut_6_33[2] , 
        \wRegOut_6_33[1] , \wRegOut_6_33[0] }), .R_Out({\wRegInTop_6_33[31] , 
        \wRegInTop_6_33[30] , \wRegInTop_6_33[29] , \wRegInTop_6_33[28] , 
        \wRegInTop_6_33[27] , \wRegInTop_6_33[26] , \wRegInTop_6_33[25] , 
        \wRegInTop_6_33[24] , \wRegInTop_6_33[23] , \wRegInTop_6_33[22] , 
        \wRegInTop_6_33[21] , \wRegInTop_6_33[20] , \wRegInTop_6_33[19] , 
        \wRegInTop_6_33[18] , \wRegInTop_6_33[17] , \wRegInTop_6_33[16] , 
        \wRegInTop_6_33[15] , \wRegInTop_6_33[14] , \wRegInTop_6_33[13] , 
        \wRegInTop_6_33[12] , \wRegInTop_6_33[11] , \wRegInTop_6_33[10] , 
        \wRegInTop_6_33[9] , \wRegInTop_6_33[8] , \wRegInTop_6_33[7] , 
        \wRegInTop_6_33[6] , \wRegInTop_6_33[5] , \wRegInTop_6_33[4] , 
        \wRegInTop_6_33[3] , \wRegInTop_6_33[2] , \wRegInTop_6_33[1] , 
        \wRegInTop_6_33[0] }) );
    BHeap_Node_WIDTH32 BHN_6_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_26[0] ), .P_In({\wRegOut_6_26[31] , 
        \wRegOut_6_26[30] , \wRegOut_6_26[29] , \wRegOut_6_26[28] , 
        \wRegOut_6_26[27] , \wRegOut_6_26[26] , \wRegOut_6_26[25] , 
        \wRegOut_6_26[24] , \wRegOut_6_26[23] , \wRegOut_6_26[22] , 
        \wRegOut_6_26[21] , \wRegOut_6_26[20] , \wRegOut_6_26[19] , 
        \wRegOut_6_26[18] , \wRegOut_6_26[17] , \wRegOut_6_26[16] , 
        \wRegOut_6_26[15] , \wRegOut_6_26[14] , \wRegOut_6_26[13] , 
        \wRegOut_6_26[12] , \wRegOut_6_26[11] , \wRegOut_6_26[10] , 
        \wRegOut_6_26[9] , \wRegOut_6_26[8] , \wRegOut_6_26[7] , 
        \wRegOut_6_26[6] , \wRegOut_6_26[5] , \wRegOut_6_26[4] , 
        \wRegOut_6_26[3] , \wRegOut_6_26[2] , \wRegOut_6_26[1] , 
        \wRegOut_6_26[0] }), .P_Out({\wRegInBot_6_26[31] , 
        \wRegInBot_6_26[30] , \wRegInBot_6_26[29] , \wRegInBot_6_26[28] , 
        \wRegInBot_6_26[27] , \wRegInBot_6_26[26] , \wRegInBot_6_26[25] , 
        \wRegInBot_6_26[24] , \wRegInBot_6_26[23] , \wRegInBot_6_26[22] , 
        \wRegInBot_6_26[21] , \wRegInBot_6_26[20] , \wRegInBot_6_26[19] , 
        \wRegInBot_6_26[18] , \wRegInBot_6_26[17] , \wRegInBot_6_26[16] , 
        \wRegInBot_6_26[15] , \wRegInBot_6_26[14] , \wRegInBot_6_26[13] , 
        \wRegInBot_6_26[12] , \wRegInBot_6_26[11] , \wRegInBot_6_26[10] , 
        \wRegInBot_6_26[9] , \wRegInBot_6_26[8] , \wRegInBot_6_26[7] , 
        \wRegInBot_6_26[6] , \wRegInBot_6_26[5] , \wRegInBot_6_26[4] , 
        \wRegInBot_6_26[3] , \wRegInBot_6_26[2] , \wRegInBot_6_26[1] , 
        \wRegInBot_6_26[0] }), .L_WR(\wRegEnTop_7_52[0] ), .L_In({
        \wRegOut_7_52[31] , \wRegOut_7_52[30] , \wRegOut_7_52[29] , 
        \wRegOut_7_52[28] , \wRegOut_7_52[27] , \wRegOut_7_52[26] , 
        \wRegOut_7_52[25] , \wRegOut_7_52[24] , \wRegOut_7_52[23] , 
        \wRegOut_7_52[22] , \wRegOut_7_52[21] , \wRegOut_7_52[20] , 
        \wRegOut_7_52[19] , \wRegOut_7_52[18] , \wRegOut_7_52[17] , 
        \wRegOut_7_52[16] , \wRegOut_7_52[15] , \wRegOut_7_52[14] , 
        \wRegOut_7_52[13] , \wRegOut_7_52[12] , \wRegOut_7_52[11] , 
        \wRegOut_7_52[10] , \wRegOut_7_52[9] , \wRegOut_7_52[8] , 
        \wRegOut_7_52[7] , \wRegOut_7_52[6] , \wRegOut_7_52[5] , 
        \wRegOut_7_52[4] , \wRegOut_7_52[3] , \wRegOut_7_52[2] , 
        \wRegOut_7_52[1] , \wRegOut_7_52[0] }), .L_Out({\wRegInTop_7_52[31] , 
        \wRegInTop_7_52[30] , \wRegInTop_7_52[29] , \wRegInTop_7_52[28] , 
        \wRegInTop_7_52[27] , \wRegInTop_7_52[26] , \wRegInTop_7_52[25] , 
        \wRegInTop_7_52[24] , \wRegInTop_7_52[23] , \wRegInTop_7_52[22] , 
        \wRegInTop_7_52[21] , \wRegInTop_7_52[20] , \wRegInTop_7_52[19] , 
        \wRegInTop_7_52[18] , \wRegInTop_7_52[17] , \wRegInTop_7_52[16] , 
        \wRegInTop_7_52[15] , \wRegInTop_7_52[14] , \wRegInTop_7_52[13] , 
        \wRegInTop_7_52[12] , \wRegInTop_7_52[11] , \wRegInTop_7_52[10] , 
        \wRegInTop_7_52[9] , \wRegInTop_7_52[8] , \wRegInTop_7_52[7] , 
        \wRegInTop_7_52[6] , \wRegInTop_7_52[5] , \wRegInTop_7_52[4] , 
        \wRegInTop_7_52[3] , \wRegInTop_7_52[2] , \wRegInTop_7_52[1] , 
        \wRegInTop_7_52[0] }), .R_WR(\wRegEnTop_7_53[0] ), .R_In({
        \wRegOut_7_53[31] , \wRegOut_7_53[30] , \wRegOut_7_53[29] , 
        \wRegOut_7_53[28] , \wRegOut_7_53[27] , \wRegOut_7_53[26] , 
        \wRegOut_7_53[25] , \wRegOut_7_53[24] , \wRegOut_7_53[23] , 
        \wRegOut_7_53[22] , \wRegOut_7_53[21] , \wRegOut_7_53[20] , 
        \wRegOut_7_53[19] , \wRegOut_7_53[18] , \wRegOut_7_53[17] , 
        \wRegOut_7_53[16] , \wRegOut_7_53[15] , \wRegOut_7_53[14] , 
        \wRegOut_7_53[13] , \wRegOut_7_53[12] , \wRegOut_7_53[11] , 
        \wRegOut_7_53[10] , \wRegOut_7_53[9] , \wRegOut_7_53[8] , 
        \wRegOut_7_53[7] , \wRegOut_7_53[6] , \wRegOut_7_53[5] , 
        \wRegOut_7_53[4] , \wRegOut_7_53[3] , \wRegOut_7_53[2] , 
        \wRegOut_7_53[1] , \wRegOut_7_53[0] }), .R_Out({\wRegInTop_7_53[31] , 
        \wRegInTop_7_53[30] , \wRegInTop_7_53[29] , \wRegInTop_7_53[28] , 
        \wRegInTop_7_53[27] , \wRegInTop_7_53[26] , \wRegInTop_7_53[25] , 
        \wRegInTop_7_53[24] , \wRegInTop_7_53[23] , \wRegInTop_7_53[22] , 
        \wRegInTop_7_53[21] , \wRegInTop_7_53[20] , \wRegInTop_7_53[19] , 
        \wRegInTop_7_53[18] , \wRegInTop_7_53[17] , \wRegInTop_7_53[16] , 
        \wRegInTop_7_53[15] , \wRegInTop_7_53[14] , \wRegInTop_7_53[13] , 
        \wRegInTop_7_53[12] , \wRegInTop_7_53[11] , \wRegInTop_7_53[10] , 
        \wRegInTop_7_53[9] , \wRegInTop_7_53[8] , \wRegInTop_7_53[7] , 
        \wRegInTop_7_53[6] , \wRegInTop_7_53[5] , \wRegInTop_7_53[4] , 
        \wRegInTop_7_53[3] , \wRegInTop_7_53[2] , \wRegInTop_7_53[1] , 
        \wRegInTop_7_53[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_29 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink93[31] , \ScanLink93[30] , \ScanLink93[29] , 
        \ScanLink93[28] , \ScanLink93[27] , \ScanLink93[26] , \ScanLink93[25] , 
        \ScanLink93[24] , \ScanLink93[23] , \ScanLink93[22] , \ScanLink93[21] , 
        \ScanLink93[20] , \ScanLink93[19] , \ScanLink93[18] , \ScanLink93[17] , 
        \ScanLink93[16] , \ScanLink93[15] , \ScanLink93[14] , \ScanLink93[13] , 
        \ScanLink93[12] , \ScanLink93[11] , \ScanLink93[10] , \ScanLink93[9] , 
        \ScanLink93[8] , \ScanLink93[7] , \ScanLink93[6] , \ScanLink93[5] , 
        \ScanLink93[4] , \ScanLink93[3] , \ScanLink93[2] , \ScanLink93[1] , 
        \ScanLink93[0] }), .ScanOut({\ScanLink92[31] , \ScanLink92[30] , 
        \ScanLink92[29] , \ScanLink92[28] , \ScanLink92[27] , \ScanLink92[26] , 
        \ScanLink92[25] , \ScanLink92[24] , \ScanLink92[23] , \ScanLink92[22] , 
        \ScanLink92[21] , \ScanLink92[20] , \ScanLink92[19] , \ScanLink92[18] , 
        \ScanLink92[17] , \ScanLink92[16] , \ScanLink92[15] , \ScanLink92[14] , 
        \ScanLink92[13] , \ScanLink92[12] , \ScanLink92[11] , \ScanLink92[10] , 
        \ScanLink92[9] , \ScanLink92[8] , \ScanLink92[7] , \ScanLink92[6] , 
        \ScanLink92[5] , \ScanLink92[4] , \ScanLink92[3] , \ScanLink92[2] , 
        \ScanLink92[1] , \ScanLink92[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_29[31] , \wRegOut_6_29[30] , 
        \wRegOut_6_29[29] , \wRegOut_6_29[28] , \wRegOut_6_29[27] , 
        \wRegOut_6_29[26] , \wRegOut_6_29[25] , \wRegOut_6_29[24] , 
        \wRegOut_6_29[23] , \wRegOut_6_29[22] , \wRegOut_6_29[21] , 
        \wRegOut_6_29[20] , \wRegOut_6_29[19] , \wRegOut_6_29[18] , 
        \wRegOut_6_29[17] , \wRegOut_6_29[16] , \wRegOut_6_29[15] , 
        \wRegOut_6_29[14] , \wRegOut_6_29[13] , \wRegOut_6_29[12] , 
        \wRegOut_6_29[11] , \wRegOut_6_29[10] , \wRegOut_6_29[9] , 
        \wRegOut_6_29[8] , \wRegOut_6_29[7] , \wRegOut_6_29[6] , 
        \wRegOut_6_29[5] , \wRegOut_6_29[4] , \wRegOut_6_29[3] , 
        \wRegOut_6_29[2] , \wRegOut_6_29[1] , \wRegOut_6_29[0] }), .Enable1(
        \wRegEnTop_6_29[0] ), .Enable2(\wRegEnBot_6_29[0] ), .In1({
        \wRegInTop_6_29[31] , \wRegInTop_6_29[30] , \wRegInTop_6_29[29] , 
        \wRegInTop_6_29[28] , \wRegInTop_6_29[27] , \wRegInTop_6_29[26] , 
        \wRegInTop_6_29[25] , \wRegInTop_6_29[24] , \wRegInTop_6_29[23] , 
        \wRegInTop_6_29[22] , \wRegInTop_6_29[21] , \wRegInTop_6_29[20] , 
        \wRegInTop_6_29[19] , \wRegInTop_6_29[18] , \wRegInTop_6_29[17] , 
        \wRegInTop_6_29[16] , \wRegInTop_6_29[15] , \wRegInTop_6_29[14] , 
        \wRegInTop_6_29[13] , \wRegInTop_6_29[12] , \wRegInTop_6_29[11] , 
        \wRegInTop_6_29[10] , \wRegInTop_6_29[9] , \wRegInTop_6_29[8] , 
        \wRegInTop_6_29[7] , \wRegInTop_6_29[6] , \wRegInTop_6_29[5] , 
        \wRegInTop_6_29[4] , \wRegInTop_6_29[3] , \wRegInTop_6_29[2] , 
        \wRegInTop_6_29[1] , \wRegInTop_6_29[0] }), .In2({\wRegInBot_6_29[31] , 
        \wRegInBot_6_29[30] , \wRegInBot_6_29[29] , \wRegInBot_6_29[28] , 
        \wRegInBot_6_29[27] , \wRegInBot_6_29[26] , \wRegInBot_6_29[25] , 
        \wRegInBot_6_29[24] , \wRegInBot_6_29[23] , \wRegInBot_6_29[22] , 
        \wRegInBot_6_29[21] , \wRegInBot_6_29[20] , \wRegInBot_6_29[19] , 
        \wRegInBot_6_29[18] , \wRegInBot_6_29[17] , \wRegInBot_6_29[16] , 
        \wRegInBot_6_29[15] , \wRegInBot_6_29[14] , \wRegInBot_6_29[13] , 
        \wRegInBot_6_29[12] , \wRegInBot_6_29[11] , \wRegInBot_6_29[10] , 
        \wRegInBot_6_29[9] , \wRegInBot_6_29[8] , \wRegInBot_6_29[7] , 
        \wRegInBot_6_29[6] , \wRegInBot_6_29[5] , \wRegInBot_6_29[4] , 
        \wRegInBot_6_29[3] , \wRegInBot_6_29[2] , \wRegInBot_6_29[1] , 
        \wRegInBot_6_29[0] }) );
    BHeap_Node_WIDTH32 BHN_5_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_31[0] ), .P_In({\wRegOut_5_31[31] , 
        \wRegOut_5_31[30] , \wRegOut_5_31[29] , \wRegOut_5_31[28] , 
        \wRegOut_5_31[27] , \wRegOut_5_31[26] , \wRegOut_5_31[25] , 
        \wRegOut_5_31[24] , \wRegOut_5_31[23] , \wRegOut_5_31[22] , 
        \wRegOut_5_31[21] , \wRegOut_5_31[20] , \wRegOut_5_31[19] , 
        \wRegOut_5_31[18] , \wRegOut_5_31[17] , \wRegOut_5_31[16] , 
        \wRegOut_5_31[15] , \wRegOut_5_31[14] , \wRegOut_5_31[13] , 
        \wRegOut_5_31[12] , \wRegOut_5_31[11] , \wRegOut_5_31[10] , 
        \wRegOut_5_31[9] , \wRegOut_5_31[8] , \wRegOut_5_31[7] , 
        \wRegOut_5_31[6] , \wRegOut_5_31[5] , \wRegOut_5_31[4] , 
        \wRegOut_5_31[3] , \wRegOut_5_31[2] , \wRegOut_5_31[1] , 
        \wRegOut_5_31[0] }), .P_Out({\wRegInBot_5_31[31] , 
        \wRegInBot_5_31[30] , \wRegInBot_5_31[29] , \wRegInBot_5_31[28] , 
        \wRegInBot_5_31[27] , \wRegInBot_5_31[26] , \wRegInBot_5_31[25] , 
        \wRegInBot_5_31[24] , \wRegInBot_5_31[23] , \wRegInBot_5_31[22] , 
        \wRegInBot_5_31[21] , \wRegInBot_5_31[20] , \wRegInBot_5_31[19] , 
        \wRegInBot_5_31[18] , \wRegInBot_5_31[17] , \wRegInBot_5_31[16] , 
        \wRegInBot_5_31[15] , \wRegInBot_5_31[14] , \wRegInBot_5_31[13] , 
        \wRegInBot_5_31[12] , \wRegInBot_5_31[11] , \wRegInBot_5_31[10] , 
        \wRegInBot_5_31[9] , \wRegInBot_5_31[8] , \wRegInBot_5_31[7] , 
        \wRegInBot_5_31[6] , \wRegInBot_5_31[5] , \wRegInBot_5_31[4] , 
        \wRegInBot_5_31[3] , \wRegInBot_5_31[2] , \wRegInBot_5_31[1] , 
        \wRegInBot_5_31[0] }), .L_WR(\wRegEnTop_6_62[0] ), .L_In({
        \wRegOut_6_62[31] , \wRegOut_6_62[30] , \wRegOut_6_62[29] , 
        \wRegOut_6_62[28] , \wRegOut_6_62[27] , \wRegOut_6_62[26] , 
        \wRegOut_6_62[25] , \wRegOut_6_62[24] , \wRegOut_6_62[23] , 
        \wRegOut_6_62[22] , \wRegOut_6_62[21] , \wRegOut_6_62[20] , 
        \wRegOut_6_62[19] , \wRegOut_6_62[18] , \wRegOut_6_62[17] , 
        \wRegOut_6_62[16] , \wRegOut_6_62[15] , \wRegOut_6_62[14] , 
        \wRegOut_6_62[13] , \wRegOut_6_62[12] , \wRegOut_6_62[11] , 
        \wRegOut_6_62[10] , \wRegOut_6_62[9] , \wRegOut_6_62[8] , 
        \wRegOut_6_62[7] , \wRegOut_6_62[6] , \wRegOut_6_62[5] , 
        \wRegOut_6_62[4] , \wRegOut_6_62[3] , \wRegOut_6_62[2] , 
        \wRegOut_6_62[1] , \wRegOut_6_62[0] }), .L_Out({\wRegInTop_6_62[31] , 
        \wRegInTop_6_62[30] , \wRegInTop_6_62[29] , \wRegInTop_6_62[28] , 
        \wRegInTop_6_62[27] , \wRegInTop_6_62[26] , \wRegInTop_6_62[25] , 
        \wRegInTop_6_62[24] , \wRegInTop_6_62[23] , \wRegInTop_6_62[22] , 
        \wRegInTop_6_62[21] , \wRegInTop_6_62[20] , \wRegInTop_6_62[19] , 
        \wRegInTop_6_62[18] , \wRegInTop_6_62[17] , \wRegInTop_6_62[16] , 
        \wRegInTop_6_62[15] , \wRegInTop_6_62[14] , \wRegInTop_6_62[13] , 
        \wRegInTop_6_62[12] , \wRegInTop_6_62[11] , \wRegInTop_6_62[10] , 
        \wRegInTop_6_62[9] , \wRegInTop_6_62[8] , \wRegInTop_6_62[7] , 
        \wRegInTop_6_62[6] , \wRegInTop_6_62[5] , \wRegInTop_6_62[4] , 
        \wRegInTop_6_62[3] , \wRegInTop_6_62[2] , \wRegInTop_6_62[1] , 
        \wRegInTop_6_62[0] }), .R_WR(\wRegEnTop_6_63[0] ), .R_In({
        \wRegOut_6_63[31] , \wRegOut_6_63[30] , \wRegOut_6_63[29] , 
        \wRegOut_6_63[28] , \wRegOut_6_63[27] , \wRegOut_6_63[26] , 
        \wRegOut_6_63[25] , \wRegOut_6_63[24] , \wRegOut_6_63[23] , 
        \wRegOut_6_63[22] , \wRegOut_6_63[21] , \wRegOut_6_63[20] , 
        \wRegOut_6_63[19] , \wRegOut_6_63[18] , \wRegOut_6_63[17] , 
        \wRegOut_6_63[16] , \wRegOut_6_63[15] , \wRegOut_6_63[14] , 
        \wRegOut_6_63[13] , \wRegOut_6_63[12] , \wRegOut_6_63[11] , 
        \wRegOut_6_63[10] , \wRegOut_6_63[9] , \wRegOut_6_63[8] , 
        \wRegOut_6_63[7] , \wRegOut_6_63[6] , \wRegOut_6_63[5] , 
        \wRegOut_6_63[4] , \wRegOut_6_63[3] , \wRegOut_6_63[2] , 
        \wRegOut_6_63[1] , \wRegOut_6_63[0] }), .R_Out({\wRegInTop_6_63[31] , 
        \wRegInTop_6_63[30] , \wRegInTop_6_63[29] , \wRegInTop_6_63[28] , 
        \wRegInTop_6_63[27] , \wRegInTop_6_63[26] , \wRegInTop_6_63[25] , 
        \wRegInTop_6_63[24] , \wRegInTop_6_63[23] , \wRegInTop_6_63[22] , 
        \wRegInTop_6_63[21] , \wRegInTop_6_63[20] , \wRegInTop_6_63[19] , 
        \wRegInTop_6_63[18] , \wRegInTop_6_63[17] , \wRegInTop_6_63[16] , 
        \wRegInTop_6_63[15] , \wRegInTop_6_63[14] , \wRegInTop_6_63[13] , 
        \wRegInTop_6_63[12] , \wRegInTop_6_63[11] , \wRegInTop_6_63[10] , 
        \wRegInTop_6_63[9] , \wRegInTop_6_63[8] , \wRegInTop_6_63[7] , 
        \wRegInTop_6_63[6] , \wRegInTop_6_63[5] , \wRegInTop_6_63[4] , 
        \wRegInTop_6_63[3] , \wRegInTop_6_63[2] , \wRegInTop_6_63[1] , 
        \wRegInTop_6_63[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink18[31] , \ScanLink18[30] , \ScanLink18[29] , 
        \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , \ScanLink18[25] , 
        \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , \ScanLink18[21] , 
        \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , \ScanLink18[17] , 
        \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , \ScanLink18[13] , 
        \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , \ScanLink18[9] , 
        \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , \ScanLink18[5] , 
        \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , \ScanLink18[1] , 
        \ScanLink18[0] }), .ScanOut({\ScanLink17[31] , \ScanLink17[30] , 
        \ScanLink17[29] , \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , 
        \ScanLink17[25] , \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , 
        \ScanLink17[21] , \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , 
        \ScanLink17[17] , \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , 
        \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , 
        \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , 
        \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , 
        \ScanLink17[1] , \ScanLink17[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_2[31] , \wRegOut_4_2[30] , \wRegOut_4_2[29] , 
        \wRegOut_4_2[28] , \wRegOut_4_2[27] , \wRegOut_4_2[26] , 
        \wRegOut_4_2[25] , \wRegOut_4_2[24] , \wRegOut_4_2[23] , 
        \wRegOut_4_2[22] , \wRegOut_4_2[21] , \wRegOut_4_2[20] , 
        \wRegOut_4_2[19] , \wRegOut_4_2[18] , \wRegOut_4_2[17] , 
        \wRegOut_4_2[16] , \wRegOut_4_2[15] , \wRegOut_4_2[14] , 
        \wRegOut_4_2[13] , \wRegOut_4_2[12] , \wRegOut_4_2[11] , 
        \wRegOut_4_2[10] , \wRegOut_4_2[9] , \wRegOut_4_2[8] , 
        \wRegOut_4_2[7] , \wRegOut_4_2[6] , \wRegOut_4_2[5] , \wRegOut_4_2[4] , 
        \wRegOut_4_2[3] , \wRegOut_4_2[2] , \wRegOut_4_2[1] , \wRegOut_4_2[0] 
        }), .Enable1(\wRegEnTop_4_2[0] ), .Enable2(\wRegEnBot_4_2[0] ), .In1({
        \wRegInTop_4_2[31] , \wRegInTop_4_2[30] , \wRegInTop_4_2[29] , 
        \wRegInTop_4_2[28] , \wRegInTop_4_2[27] , \wRegInTop_4_2[26] , 
        \wRegInTop_4_2[25] , \wRegInTop_4_2[24] , \wRegInTop_4_2[23] , 
        \wRegInTop_4_2[22] , \wRegInTop_4_2[21] , \wRegInTop_4_2[20] , 
        \wRegInTop_4_2[19] , \wRegInTop_4_2[18] , \wRegInTop_4_2[17] , 
        \wRegInTop_4_2[16] , \wRegInTop_4_2[15] , \wRegInTop_4_2[14] , 
        \wRegInTop_4_2[13] , \wRegInTop_4_2[12] , \wRegInTop_4_2[11] , 
        \wRegInTop_4_2[10] , \wRegInTop_4_2[9] , \wRegInTop_4_2[8] , 
        \wRegInTop_4_2[7] , \wRegInTop_4_2[6] , \wRegInTop_4_2[5] , 
        \wRegInTop_4_2[4] , \wRegInTop_4_2[3] , \wRegInTop_4_2[2] , 
        \wRegInTop_4_2[1] , \wRegInTop_4_2[0] }), .In2({\wRegInBot_4_2[31] , 
        \wRegInBot_4_2[30] , \wRegInBot_4_2[29] , \wRegInBot_4_2[28] , 
        \wRegInBot_4_2[27] , \wRegInBot_4_2[26] , \wRegInBot_4_2[25] , 
        \wRegInBot_4_2[24] , \wRegInBot_4_2[23] , \wRegInBot_4_2[22] , 
        \wRegInBot_4_2[21] , \wRegInBot_4_2[20] , \wRegInBot_4_2[19] , 
        \wRegInBot_4_2[18] , \wRegInBot_4_2[17] , \wRegInBot_4_2[16] , 
        \wRegInBot_4_2[15] , \wRegInBot_4_2[14] , \wRegInBot_4_2[13] , 
        \wRegInBot_4_2[12] , \wRegInBot_4_2[11] , \wRegInBot_4_2[10] , 
        \wRegInBot_4_2[9] , \wRegInBot_4_2[8] , \wRegInBot_4_2[7] , 
        \wRegInBot_4_2[6] , \wRegInBot_4_2[5] , \wRegInBot_4_2[4] , 
        \wRegInBot_4_2[3] , \wRegInBot_4_2[2] , \wRegInBot_4_2[1] , 
        \wRegInBot_4_2[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink21[31] , \ScanLink21[30] , \ScanLink21[29] , 
        \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , \ScanLink21[25] , 
        \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , \ScanLink21[21] , 
        \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , \ScanLink21[17] , 
        \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , \ScanLink21[13] , 
        \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , \ScanLink21[9] , 
        \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , \ScanLink21[5] , 
        \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , \ScanLink21[1] , 
        \ScanLink21[0] }), .ScanOut({\ScanLink20[31] , \ScanLink20[30] , 
        \ScanLink20[29] , \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , 
        \ScanLink20[25] , \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , 
        \ScanLink20[21] , \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , 
        \ScanLink20[17] , \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , 
        \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , 
        \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , 
        \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , 
        \ScanLink20[1] , \ScanLink20[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_5[31] , \wRegOut_4_5[30] , \wRegOut_4_5[29] , 
        \wRegOut_4_5[28] , \wRegOut_4_5[27] , \wRegOut_4_5[26] , 
        \wRegOut_4_5[25] , \wRegOut_4_5[24] , \wRegOut_4_5[23] , 
        \wRegOut_4_5[22] , \wRegOut_4_5[21] , \wRegOut_4_5[20] , 
        \wRegOut_4_5[19] , \wRegOut_4_5[18] , \wRegOut_4_5[17] , 
        \wRegOut_4_5[16] , \wRegOut_4_5[15] , \wRegOut_4_5[14] , 
        \wRegOut_4_5[13] , \wRegOut_4_5[12] , \wRegOut_4_5[11] , 
        \wRegOut_4_5[10] , \wRegOut_4_5[9] , \wRegOut_4_5[8] , 
        \wRegOut_4_5[7] , \wRegOut_4_5[6] , \wRegOut_4_5[5] , \wRegOut_4_5[4] , 
        \wRegOut_4_5[3] , \wRegOut_4_5[2] , \wRegOut_4_5[1] , \wRegOut_4_5[0] 
        }), .Enable1(\wRegEnTop_4_5[0] ), .Enable2(\wRegEnBot_4_5[0] ), .In1({
        \wRegInTop_4_5[31] , \wRegInTop_4_5[30] , \wRegInTop_4_5[29] , 
        \wRegInTop_4_5[28] , \wRegInTop_4_5[27] , \wRegInTop_4_5[26] , 
        \wRegInTop_4_5[25] , \wRegInTop_4_5[24] , \wRegInTop_4_5[23] , 
        \wRegInTop_4_5[22] , \wRegInTop_4_5[21] , \wRegInTop_4_5[20] , 
        \wRegInTop_4_5[19] , \wRegInTop_4_5[18] , \wRegInTop_4_5[17] , 
        \wRegInTop_4_5[16] , \wRegInTop_4_5[15] , \wRegInTop_4_5[14] , 
        \wRegInTop_4_5[13] , \wRegInTop_4_5[12] , \wRegInTop_4_5[11] , 
        \wRegInTop_4_5[10] , \wRegInTop_4_5[9] , \wRegInTop_4_5[8] , 
        \wRegInTop_4_5[7] , \wRegInTop_4_5[6] , \wRegInTop_4_5[5] , 
        \wRegInTop_4_5[4] , \wRegInTop_4_5[3] , \wRegInTop_4_5[2] , 
        \wRegInTop_4_5[1] , \wRegInTop_4_5[0] }), .In2({\wRegInBot_4_5[31] , 
        \wRegInBot_4_5[30] , \wRegInBot_4_5[29] , \wRegInBot_4_5[28] , 
        \wRegInBot_4_5[27] , \wRegInBot_4_5[26] , \wRegInBot_4_5[25] , 
        \wRegInBot_4_5[24] , \wRegInBot_4_5[23] , \wRegInBot_4_5[22] , 
        \wRegInBot_4_5[21] , \wRegInBot_4_5[20] , \wRegInBot_4_5[19] , 
        \wRegInBot_4_5[18] , \wRegInBot_4_5[17] , \wRegInBot_4_5[16] , 
        \wRegInBot_4_5[15] , \wRegInBot_4_5[14] , \wRegInBot_4_5[13] , 
        \wRegInBot_4_5[12] , \wRegInBot_4_5[11] , \wRegInBot_4_5[10] , 
        \wRegInBot_4_5[9] , \wRegInBot_4_5[8] , \wRegInBot_4_5[7] , 
        \wRegInBot_4_5[6] , \wRegInBot_4_5[5] , \wRegInBot_4_5[4] , 
        \wRegInBot_4_5[3] , \wRegInBot_4_5[2] , \wRegInBot_4_5[1] , 
        \wRegInBot_4_5[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink27[31] , \ScanLink27[30] , \ScanLink27[29] , 
        \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , \ScanLink27[25] , 
        \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , \ScanLink27[21] , 
        \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , \ScanLink27[17] , 
        \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , \ScanLink27[13] , 
        \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , \ScanLink27[9] , 
        \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , \ScanLink27[5] , 
        \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , \ScanLink27[1] , 
        \ScanLink27[0] }), .ScanOut({\ScanLink26[31] , \ScanLink26[30] , 
        \ScanLink26[29] , \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , 
        \ScanLink26[25] , \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , 
        \ScanLink26[21] , \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , 
        \ScanLink26[17] , \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , 
        \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , 
        \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , 
        \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , 
        \ScanLink26[1] , \ScanLink26[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_11[31] , \wRegOut_4_11[30] , 
        \wRegOut_4_11[29] , \wRegOut_4_11[28] , \wRegOut_4_11[27] , 
        \wRegOut_4_11[26] , \wRegOut_4_11[25] , \wRegOut_4_11[24] , 
        \wRegOut_4_11[23] , \wRegOut_4_11[22] , \wRegOut_4_11[21] , 
        \wRegOut_4_11[20] , \wRegOut_4_11[19] , \wRegOut_4_11[18] , 
        \wRegOut_4_11[17] , \wRegOut_4_11[16] , \wRegOut_4_11[15] , 
        \wRegOut_4_11[14] , \wRegOut_4_11[13] , \wRegOut_4_11[12] , 
        \wRegOut_4_11[11] , \wRegOut_4_11[10] , \wRegOut_4_11[9] , 
        \wRegOut_4_11[8] , \wRegOut_4_11[7] , \wRegOut_4_11[6] , 
        \wRegOut_4_11[5] , \wRegOut_4_11[4] , \wRegOut_4_11[3] , 
        \wRegOut_4_11[2] , \wRegOut_4_11[1] , \wRegOut_4_11[0] }), .Enable1(
        \wRegEnTop_4_11[0] ), .Enable2(\wRegEnBot_4_11[0] ), .In1({
        \wRegInTop_4_11[31] , \wRegInTop_4_11[30] , \wRegInTop_4_11[29] , 
        \wRegInTop_4_11[28] , \wRegInTop_4_11[27] , \wRegInTop_4_11[26] , 
        \wRegInTop_4_11[25] , \wRegInTop_4_11[24] , \wRegInTop_4_11[23] , 
        \wRegInTop_4_11[22] , \wRegInTop_4_11[21] , \wRegInTop_4_11[20] , 
        \wRegInTop_4_11[19] , \wRegInTop_4_11[18] , \wRegInTop_4_11[17] , 
        \wRegInTop_4_11[16] , \wRegInTop_4_11[15] , \wRegInTop_4_11[14] , 
        \wRegInTop_4_11[13] , \wRegInTop_4_11[12] , \wRegInTop_4_11[11] , 
        \wRegInTop_4_11[10] , \wRegInTop_4_11[9] , \wRegInTop_4_11[8] , 
        \wRegInTop_4_11[7] , \wRegInTop_4_11[6] , \wRegInTop_4_11[5] , 
        \wRegInTop_4_11[4] , \wRegInTop_4_11[3] , \wRegInTop_4_11[2] , 
        \wRegInTop_4_11[1] , \wRegInTop_4_11[0] }), .In2({\wRegInBot_4_11[31] , 
        \wRegInBot_4_11[30] , \wRegInBot_4_11[29] , \wRegInBot_4_11[28] , 
        \wRegInBot_4_11[27] , \wRegInBot_4_11[26] , \wRegInBot_4_11[25] , 
        \wRegInBot_4_11[24] , \wRegInBot_4_11[23] , \wRegInBot_4_11[22] , 
        \wRegInBot_4_11[21] , \wRegInBot_4_11[20] , \wRegInBot_4_11[19] , 
        \wRegInBot_4_11[18] , \wRegInBot_4_11[17] , \wRegInBot_4_11[16] , 
        \wRegInBot_4_11[15] , \wRegInBot_4_11[14] , \wRegInBot_4_11[13] , 
        \wRegInBot_4_11[12] , \wRegInBot_4_11[11] , \wRegInBot_4_11[10] , 
        \wRegInBot_4_11[9] , \wRegInBot_4_11[8] , \wRegInBot_4_11[7] , 
        \wRegInBot_4_11[6] , \wRegInBot_4_11[5] , \wRegInBot_4_11[4] , 
        \wRegInBot_4_11[3] , \wRegInBot_4_11[2] , \wRegInBot_4_11[1] , 
        \wRegInBot_4_11[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink37[31] , \ScanLink37[30] , \ScanLink37[29] , 
        \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , \ScanLink37[25] , 
        \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , \ScanLink37[21] , 
        \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , \ScanLink37[17] , 
        \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , \ScanLink37[13] , 
        \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , \ScanLink37[9] , 
        \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , \ScanLink37[5] , 
        \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , \ScanLink37[1] , 
        \ScanLink37[0] }), .ScanOut({\ScanLink36[31] , \ScanLink36[30] , 
        \ScanLink36[29] , \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , 
        \ScanLink36[25] , \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , 
        \ScanLink36[21] , \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , 
        \ScanLink36[17] , \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , 
        \ScanLink36[13] , \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , 
        \ScanLink36[9] , \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , 
        \ScanLink36[5] , \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , 
        \ScanLink36[1] , \ScanLink36[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_5[31] , \wRegOut_5_5[30] , \wRegOut_5_5[29] , 
        \wRegOut_5_5[28] , \wRegOut_5_5[27] , \wRegOut_5_5[26] , 
        \wRegOut_5_5[25] , \wRegOut_5_5[24] , \wRegOut_5_5[23] , 
        \wRegOut_5_5[22] , \wRegOut_5_5[21] , \wRegOut_5_5[20] , 
        \wRegOut_5_5[19] , \wRegOut_5_5[18] , \wRegOut_5_5[17] , 
        \wRegOut_5_5[16] , \wRegOut_5_5[15] , \wRegOut_5_5[14] , 
        \wRegOut_5_5[13] , \wRegOut_5_5[12] , \wRegOut_5_5[11] , 
        \wRegOut_5_5[10] , \wRegOut_5_5[9] , \wRegOut_5_5[8] , 
        \wRegOut_5_5[7] , \wRegOut_5_5[6] , \wRegOut_5_5[5] , \wRegOut_5_5[4] , 
        \wRegOut_5_5[3] , \wRegOut_5_5[2] , \wRegOut_5_5[1] , \wRegOut_5_5[0] 
        }), .Enable1(\wRegEnTop_5_5[0] ), .Enable2(\wRegEnBot_5_5[0] ), .In1({
        \wRegInTop_5_5[31] , \wRegInTop_5_5[30] , \wRegInTop_5_5[29] , 
        \wRegInTop_5_5[28] , \wRegInTop_5_5[27] , \wRegInTop_5_5[26] , 
        \wRegInTop_5_5[25] , \wRegInTop_5_5[24] , \wRegInTop_5_5[23] , 
        \wRegInTop_5_5[22] , \wRegInTop_5_5[21] , \wRegInTop_5_5[20] , 
        \wRegInTop_5_5[19] , \wRegInTop_5_5[18] , \wRegInTop_5_5[17] , 
        \wRegInTop_5_5[16] , \wRegInTop_5_5[15] , \wRegInTop_5_5[14] , 
        \wRegInTop_5_5[13] , \wRegInTop_5_5[12] , \wRegInTop_5_5[11] , 
        \wRegInTop_5_5[10] , \wRegInTop_5_5[9] , \wRegInTop_5_5[8] , 
        \wRegInTop_5_5[7] , \wRegInTop_5_5[6] , \wRegInTop_5_5[5] , 
        \wRegInTop_5_5[4] , \wRegInTop_5_5[3] , \wRegInTop_5_5[2] , 
        \wRegInTop_5_5[1] , \wRegInTop_5_5[0] }), .In2({\wRegInBot_5_5[31] , 
        \wRegInBot_5_5[30] , \wRegInBot_5_5[29] , \wRegInBot_5_5[28] , 
        \wRegInBot_5_5[27] , \wRegInBot_5_5[26] , \wRegInBot_5_5[25] , 
        \wRegInBot_5_5[24] , \wRegInBot_5_5[23] , \wRegInBot_5_5[22] , 
        \wRegInBot_5_5[21] , \wRegInBot_5_5[20] , \wRegInBot_5_5[19] , 
        \wRegInBot_5_5[18] , \wRegInBot_5_5[17] , \wRegInBot_5_5[16] , 
        \wRegInBot_5_5[15] , \wRegInBot_5_5[14] , \wRegInBot_5_5[13] , 
        \wRegInBot_5_5[12] , \wRegInBot_5_5[11] , \wRegInBot_5_5[10] , 
        \wRegInBot_5_5[9] , \wRegInBot_5_5[8] , \wRegInBot_5_5[7] , 
        \wRegInBot_5_5[6] , \wRegInBot_5_5[5] , \wRegInBot_5_5[4] , 
        \wRegInBot_5_5[3] , \wRegInBot_5_5[2] , \wRegInBot_5_5[1] , 
        \wRegInBot_5_5[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink64[31] , \ScanLink64[30] , \ScanLink64[29] , 
        \ScanLink64[28] , \ScanLink64[27] , \ScanLink64[26] , \ScanLink64[25] , 
        \ScanLink64[24] , \ScanLink64[23] , \ScanLink64[22] , \ScanLink64[21] , 
        \ScanLink64[20] , \ScanLink64[19] , \ScanLink64[18] , \ScanLink64[17] , 
        \ScanLink64[16] , \ScanLink64[15] , \ScanLink64[14] , \ScanLink64[13] , 
        \ScanLink64[12] , \ScanLink64[11] , \ScanLink64[10] , \ScanLink64[9] , 
        \ScanLink64[8] , \ScanLink64[7] , \ScanLink64[6] , \ScanLink64[5] , 
        \ScanLink64[4] , \ScanLink64[3] , \ScanLink64[2] , \ScanLink64[1] , 
        \ScanLink64[0] }), .ScanOut({\ScanLink63[31] , \ScanLink63[30] , 
        \ScanLink63[29] , \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , 
        \ScanLink63[25] , \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , 
        \ScanLink63[21] , \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , 
        \ScanLink63[17] , \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , 
        \ScanLink63[13] , \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , 
        \ScanLink63[9] , \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , 
        \ScanLink63[5] , \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , 
        \ScanLink63[1] , \ScanLink63[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_0[31] , \wRegOut_6_0[30] , \wRegOut_6_0[29] , 
        \wRegOut_6_0[28] , \wRegOut_6_0[27] , \wRegOut_6_0[26] , 
        \wRegOut_6_0[25] , \wRegOut_6_0[24] , \wRegOut_6_0[23] , 
        \wRegOut_6_0[22] , \wRegOut_6_0[21] , \wRegOut_6_0[20] , 
        \wRegOut_6_0[19] , \wRegOut_6_0[18] , \wRegOut_6_0[17] , 
        \wRegOut_6_0[16] , \wRegOut_6_0[15] , \wRegOut_6_0[14] , 
        \wRegOut_6_0[13] , \wRegOut_6_0[12] , \wRegOut_6_0[11] , 
        \wRegOut_6_0[10] , \wRegOut_6_0[9] , \wRegOut_6_0[8] , 
        \wRegOut_6_0[7] , \wRegOut_6_0[6] , \wRegOut_6_0[5] , \wRegOut_6_0[4] , 
        \wRegOut_6_0[3] , \wRegOut_6_0[2] , \wRegOut_6_0[1] , \wRegOut_6_0[0] 
        }), .Enable1(\wRegEnTop_6_0[0] ), .Enable2(\wRegEnBot_6_0[0] ), .In1({
        \wRegInTop_6_0[31] , \wRegInTop_6_0[30] , \wRegInTop_6_0[29] , 
        \wRegInTop_6_0[28] , \wRegInTop_6_0[27] , \wRegInTop_6_0[26] , 
        \wRegInTop_6_0[25] , \wRegInTop_6_0[24] , \wRegInTop_6_0[23] , 
        \wRegInTop_6_0[22] , \wRegInTop_6_0[21] , \wRegInTop_6_0[20] , 
        \wRegInTop_6_0[19] , \wRegInTop_6_0[18] , \wRegInTop_6_0[17] , 
        \wRegInTop_6_0[16] , \wRegInTop_6_0[15] , \wRegInTop_6_0[14] , 
        \wRegInTop_6_0[13] , \wRegInTop_6_0[12] , \wRegInTop_6_0[11] , 
        \wRegInTop_6_0[10] , \wRegInTop_6_0[9] , \wRegInTop_6_0[8] , 
        \wRegInTop_6_0[7] , \wRegInTop_6_0[6] , \wRegInTop_6_0[5] , 
        \wRegInTop_6_0[4] , \wRegInTop_6_0[3] , \wRegInTop_6_0[2] , 
        \wRegInTop_6_0[1] , \wRegInTop_6_0[0] }), .In2({\wRegInBot_6_0[31] , 
        \wRegInBot_6_0[30] , \wRegInBot_6_0[29] , \wRegInBot_6_0[28] , 
        \wRegInBot_6_0[27] , \wRegInBot_6_0[26] , \wRegInBot_6_0[25] , 
        \wRegInBot_6_0[24] , \wRegInBot_6_0[23] , \wRegInBot_6_0[22] , 
        \wRegInBot_6_0[21] , \wRegInBot_6_0[20] , \wRegInBot_6_0[19] , 
        \wRegInBot_6_0[18] , \wRegInBot_6_0[17] , \wRegInBot_6_0[16] , 
        \wRegInBot_6_0[15] , \wRegInBot_6_0[14] , \wRegInBot_6_0[13] , 
        \wRegInBot_6_0[12] , \wRegInBot_6_0[11] , \wRegInBot_6_0[10] , 
        \wRegInBot_6_0[9] , \wRegInBot_6_0[8] , \wRegInBot_6_0[7] , 
        \wRegInBot_6_0[6] , \wRegInBot_6_0[5] , \wRegInBot_6_0[4] , 
        \wRegInBot_6_0[3] , \wRegInBot_6_0[2] , \wRegInBot_6_0[1] , 
        \wRegInBot_6_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_55 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink119[31] , \ScanLink119[30] , \ScanLink119[29] , 
        \ScanLink119[28] , \ScanLink119[27] , \ScanLink119[26] , 
        \ScanLink119[25] , \ScanLink119[24] , \ScanLink119[23] , 
        \ScanLink119[22] , \ScanLink119[21] , \ScanLink119[20] , 
        \ScanLink119[19] , \ScanLink119[18] , \ScanLink119[17] , 
        \ScanLink119[16] , \ScanLink119[15] , \ScanLink119[14] , 
        \ScanLink119[13] , \ScanLink119[12] , \ScanLink119[11] , 
        \ScanLink119[10] , \ScanLink119[9] , \ScanLink119[8] , 
        \ScanLink119[7] , \ScanLink119[6] , \ScanLink119[5] , \ScanLink119[4] , 
        \ScanLink119[3] , \ScanLink119[2] , \ScanLink119[1] , \ScanLink119[0] 
        }), .ScanOut({\ScanLink118[31] , \ScanLink118[30] , \ScanLink118[29] , 
        \ScanLink118[28] , \ScanLink118[27] , \ScanLink118[26] , 
        \ScanLink118[25] , \ScanLink118[24] , \ScanLink118[23] , 
        \ScanLink118[22] , \ScanLink118[21] , \ScanLink118[20] , 
        \ScanLink118[19] , \ScanLink118[18] , \ScanLink118[17] , 
        \ScanLink118[16] , \ScanLink118[15] , \ScanLink118[14] , 
        \ScanLink118[13] , \ScanLink118[12] , \ScanLink118[11] , 
        \ScanLink118[10] , \ScanLink118[9] , \ScanLink118[8] , 
        \ScanLink118[7] , \ScanLink118[6] , \ScanLink118[5] , \ScanLink118[4] , 
        \ScanLink118[3] , \ScanLink118[2] , \ScanLink118[1] , \ScanLink118[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_55[31] , 
        \wRegOut_6_55[30] , \wRegOut_6_55[29] , \wRegOut_6_55[28] , 
        \wRegOut_6_55[27] , \wRegOut_6_55[26] , \wRegOut_6_55[25] , 
        \wRegOut_6_55[24] , \wRegOut_6_55[23] , \wRegOut_6_55[22] , 
        \wRegOut_6_55[21] , \wRegOut_6_55[20] , \wRegOut_6_55[19] , 
        \wRegOut_6_55[18] , \wRegOut_6_55[17] , \wRegOut_6_55[16] , 
        \wRegOut_6_55[15] , \wRegOut_6_55[14] , \wRegOut_6_55[13] , 
        \wRegOut_6_55[12] , \wRegOut_6_55[11] , \wRegOut_6_55[10] , 
        \wRegOut_6_55[9] , \wRegOut_6_55[8] , \wRegOut_6_55[7] , 
        \wRegOut_6_55[6] , \wRegOut_6_55[5] , \wRegOut_6_55[4] , 
        \wRegOut_6_55[3] , \wRegOut_6_55[2] , \wRegOut_6_55[1] , 
        \wRegOut_6_55[0] }), .Enable1(\wRegEnTop_6_55[0] ), .Enable2(
        \wRegEnBot_6_55[0] ), .In1({\wRegInTop_6_55[31] , \wRegInTop_6_55[30] , 
        \wRegInTop_6_55[29] , \wRegInTop_6_55[28] , \wRegInTop_6_55[27] , 
        \wRegInTop_6_55[26] , \wRegInTop_6_55[25] , \wRegInTop_6_55[24] , 
        \wRegInTop_6_55[23] , \wRegInTop_6_55[22] , \wRegInTop_6_55[21] , 
        \wRegInTop_6_55[20] , \wRegInTop_6_55[19] , \wRegInTop_6_55[18] , 
        \wRegInTop_6_55[17] , \wRegInTop_6_55[16] , \wRegInTop_6_55[15] , 
        \wRegInTop_6_55[14] , \wRegInTop_6_55[13] , \wRegInTop_6_55[12] , 
        \wRegInTop_6_55[11] , \wRegInTop_6_55[10] , \wRegInTop_6_55[9] , 
        \wRegInTop_6_55[8] , \wRegInTop_6_55[7] , \wRegInTop_6_55[6] , 
        \wRegInTop_6_55[5] , \wRegInTop_6_55[4] , \wRegInTop_6_55[3] , 
        \wRegInTop_6_55[2] , \wRegInTop_6_55[1] , \wRegInTop_6_55[0] }), .In2(
        {\wRegInBot_6_55[31] , \wRegInBot_6_55[30] , \wRegInBot_6_55[29] , 
        \wRegInBot_6_55[28] , \wRegInBot_6_55[27] , \wRegInBot_6_55[26] , 
        \wRegInBot_6_55[25] , \wRegInBot_6_55[24] , \wRegInBot_6_55[23] , 
        \wRegInBot_6_55[22] , \wRegInBot_6_55[21] , \wRegInBot_6_55[20] , 
        \wRegInBot_6_55[19] , \wRegInBot_6_55[18] , \wRegInBot_6_55[17] , 
        \wRegInBot_6_55[16] , \wRegInBot_6_55[15] , \wRegInBot_6_55[14] , 
        \wRegInBot_6_55[13] , \wRegInBot_6_55[12] , \wRegInBot_6_55[11] , 
        \wRegInBot_6_55[10] , \wRegInBot_6_55[9] , \wRegInBot_6_55[8] , 
        \wRegInBot_6_55[7] , \wRegInBot_6_55[6] , \wRegInBot_6_55[5] , 
        \wRegInBot_6_55[4] , \wRegInBot_6_55[3] , \wRegInBot_6_55[2] , 
        \wRegInBot_6_55[1] , \wRegInBot_6_55[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink137[31] , \ScanLink137[30] , \ScanLink137[29] , 
        \ScanLink137[28] , \ScanLink137[27] , \ScanLink137[26] , 
        \ScanLink137[25] , \ScanLink137[24] , \ScanLink137[23] , 
        \ScanLink137[22] , \ScanLink137[21] , \ScanLink137[20] , 
        \ScanLink137[19] , \ScanLink137[18] , \ScanLink137[17] , 
        \ScanLink137[16] , \ScanLink137[15] , \ScanLink137[14] , 
        \ScanLink137[13] , \ScanLink137[12] , \ScanLink137[11] , 
        \ScanLink137[10] , \ScanLink137[9] , \ScanLink137[8] , 
        \ScanLink137[7] , \ScanLink137[6] , \ScanLink137[5] , \ScanLink137[4] , 
        \ScanLink137[3] , \ScanLink137[2] , \ScanLink137[1] , \ScanLink137[0] 
        }), .ScanOut({\ScanLink136[31] , \ScanLink136[30] , \ScanLink136[29] , 
        \ScanLink136[28] , \ScanLink136[27] , \ScanLink136[26] , 
        \ScanLink136[25] , \ScanLink136[24] , \ScanLink136[23] , 
        \ScanLink136[22] , \ScanLink136[21] , \ScanLink136[20] , 
        \ScanLink136[19] , \ScanLink136[18] , \ScanLink136[17] , 
        \ScanLink136[16] , \ScanLink136[15] , \ScanLink136[14] , 
        \ScanLink136[13] , \ScanLink136[12] , \ScanLink136[11] , 
        \ScanLink136[10] , \ScanLink136[9] , \ScanLink136[8] , 
        \ScanLink136[7] , \ScanLink136[6] , \ScanLink136[5] , \ScanLink136[4] , 
        \ScanLink136[3] , \ScanLink136[2] , \ScanLink136[1] , \ScanLink136[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_9[31] , 
        \wRegOut_7_9[30] , \wRegOut_7_9[29] , \wRegOut_7_9[28] , 
        \wRegOut_7_9[27] , \wRegOut_7_9[26] , \wRegOut_7_9[25] , 
        \wRegOut_7_9[24] , \wRegOut_7_9[23] , \wRegOut_7_9[22] , 
        \wRegOut_7_9[21] , \wRegOut_7_9[20] , \wRegOut_7_9[19] , 
        \wRegOut_7_9[18] , \wRegOut_7_9[17] , \wRegOut_7_9[16] , 
        \wRegOut_7_9[15] , \wRegOut_7_9[14] , \wRegOut_7_9[13] , 
        \wRegOut_7_9[12] , \wRegOut_7_9[11] , \wRegOut_7_9[10] , 
        \wRegOut_7_9[9] , \wRegOut_7_9[8] , \wRegOut_7_9[7] , \wRegOut_7_9[6] , 
        \wRegOut_7_9[5] , \wRegOut_7_9[4] , \wRegOut_7_9[3] , \wRegOut_7_9[2] , 
        \wRegOut_7_9[1] , \wRegOut_7_9[0] }), .Enable1(\wRegEnTop_7_9[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_9[31] , \wRegInTop_7_9[30] , 
        \wRegInTop_7_9[29] , \wRegInTop_7_9[28] , \wRegInTop_7_9[27] , 
        \wRegInTop_7_9[26] , \wRegInTop_7_9[25] , \wRegInTop_7_9[24] , 
        \wRegInTop_7_9[23] , \wRegInTop_7_9[22] , \wRegInTop_7_9[21] , 
        \wRegInTop_7_9[20] , \wRegInTop_7_9[19] , \wRegInTop_7_9[18] , 
        \wRegInTop_7_9[17] , \wRegInTop_7_9[16] , \wRegInTop_7_9[15] , 
        \wRegInTop_7_9[14] , \wRegInTop_7_9[13] , \wRegInTop_7_9[12] , 
        \wRegInTop_7_9[11] , \wRegInTop_7_9[10] , \wRegInTop_7_9[9] , 
        \wRegInTop_7_9[8] , \wRegInTop_7_9[7] , \wRegInTop_7_9[6] , 
        \wRegInTop_7_9[5] , \wRegInTop_7_9[4] , \wRegInTop_7_9[3] , 
        \wRegInTop_7_9[2] , \wRegInTop_7_9[1] , \wRegInTop_7_9[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_68 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink196[31] , \ScanLink196[30] , \ScanLink196[29] , 
        \ScanLink196[28] , \ScanLink196[27] , \ScanLink196[26] , 
        \ScanLink196[25] , \ScanLink196[24] , \ScanLink196[23] , 
        \ScanLink196[22] , \ScanLink196[21] , \ScanLink196[20] , 
        \ScanLink196[19] , \ScanLink196[18] , \ScanLink196[17] , 
        \ScanLink196[16] , \ScanLink196[15] , \ScanLink196[14] , 
        \ScanLink196[13] , \ScanLink196[12] , \ScanLink196[11] , 
        \ScanLink196[10] , \ScanLink196[9] , \ScanLink196[8] , 
        \ScanLink196[7] , \ScanLink196[6] , \ScanLink196[5] , \ScanLink196[4] , 
        \ScanLink196[3] , \ScanLink196[2] , \ScanLink196[1] , \ScanLink196[0] 
        }), .ScanOut({\ScanLink195[31] , \ScanLink195[30] , \ScanLink195[29] , 
        \ScanLink195[28] , \ScanLink195[27] , \ScanLink195[26] , 
        \ScanLink195[25] , \ScanLink195[24] , \ScanLink195[23] , 
        \ScanLink195[22] , \ScanLink195[21] , \ScanLink195[20] , 
        \ScanLink195[19] , \ScanLink195[18] , \ScanLink195[17] , 
        \ScanLink195[16] , \ScanLink195[15] , \ScanLink195[14] , 
        \ScanLink195[13] , \ScanLink195[12] , \ScanLink195[11] , 
        \ScanLink195[10] , \ScanLink195[9] , \ScanLink195[8] , 
        \ScanLink195[7] , \ScanLink195[6] , \ScanLink195[5] , \ScanLink195[4] , 
        \ScanLink195[3] , \ScanLink195[2] , \ScanLink195[1] , \ScanLink195[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_68[31] , 
        \wRegOut_7_68[30] , \wRegOut_7_68[29] , \wRegOut_7_68[28] , 
        \wRegOut_7_68[27] , \wRegOut_7_68[26] , \wRegOut_7_68[25] , 
        \wRegOut_7_68[24] , \wRegOut_7_68[23] , \wRegOut_7_68[22] , 
        \wRegOut_7_68[21] , \wRegOut_7_68[20] , \wRegOut_7_68[19] , 
        \wRegOut_7_68[18] , \wRegOut_7_68[17] , \wRegOut_7_68[16] , 
        \wRegOut_7_68[15] , \wRegOut_7_68[14] , \wRegOut_7_68[13] , 
        \wRegOut_7_68[12] , \wRegOut_7_68[11] , \wRegOut_7_68[10] , 
        \wRegOut_7_68[9] , \wRegOut_7_68[8] , \wRegOut_7_68[7] , 
        \wRegOut_7_68[6] , \wRegOut_7_68[5] , \wRegOut_7_68[4] , 
        \wRegOut_7_68[3] , \wRegOut_7_68[2] , \wRegOut_7_68[1] , 
        \wRegOut_7_68[0] }), .Enable1(\wRegEnTop_7_68[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_68[31] , \wRegInTop_7_68[30] , \wRegInTop_7_68[29] , 
        \wRegInTop_7_68[28] , \wRegInTop_7_68[27] , \wRegInTop_7_68[26] , 
        \wRegInTop_7_68[25] , \wRegInTop_7_68[24] , \wRegInTop_7_68[23] , 
        \wRegInTop_7_68[22] , \wRegInTop_7_68[21] , \wRegInTop_7_68[20] , 
        \wRegInTop_7_68[19] , \wRegInTop_7_68[18] , \wRegInTop_7_68[17] , 
        \wRegInTop_7_68[16] , \wRegInTop_7_68[15] , \wRegInTop_7_68[14] , 
        \wRegInTop_7_68[13] , \wRegInTop_7_68[12] , \wRegInTop_7_68[11] , 
        \wRegInTop_7_68[10] , \wRegInTop_7_68[9] , \wRegInTop_7_68[8] , 
        \wRegInTop_7_68[7] , \wRegInTop_7_68[6] , \wRegInTop_7_68[5] , 
        \wRegInTop_7_68[4] , \wRegInTop_7_68[3] , \wRegInTop_7_68[2] , 
        \wRegInTop_7_68[1] , \wRegInTop_7_68[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_34[0] ), .P_In({\wRegOut_6_34[31] , 
        \wRegOut_6_34[30] , \wRegOut_6_34[29] , \wRegOut_6_34[28] , 
        \wRegOut_6_34[27] , \wRegOut_6_34[26] , \wRegOut_6_34[25] , 
        \wRegOut_6_34[24] , \wRegOut_6_34[23] , \wRegOut_6_34[22] , 
        \wRegOut_6_34[21] , \wRegOut_6_34[20] , \wRegOut_6_34[19] , 
        \wRegOut_6_34[18] , \wRegOut_6_34[17] , \wRegOut_6_34[16] , 
        \wRegOut_6_34[15] , \wRegOut_6_34[14] , \wRegOut_6_34[13] , 
        \wRegOut_6_34[12] , \wRegOut_6_34[11] , \wRegOut_6_34[10] , 
        \wRegOut_6_34[9] , \wRegOut_6_34[8] , \wRegOut_6_34[7] , 
        \wRegOut_6_34[6] , \wRegOut_6_34[5] , \wRegOut_6_34[4] , 
        \wRegOut_6_34[3] , \wRegOut_6_34[2] , \wRegOut_6_34[1] , 
        \wRegOut_6_34[0] }), .P_Out({\wRegInBot_6_34[31] , 
        \wRegInBot_6_34[30] , \wRegInBot_6_34[29] , \wRegInBot_6_34[28] , 
        \wRegInBot_6_34[27] , \wRegInBot_6_34[26] , \wRegInBot_6_34[25] , 
        \wRegInBot_6_34[24] , \wRegInBot_6_34[23] , \wRegInBot_6_34[22] , 
        \wRegInBot_6_34[21] , \wRegInBot_6_34[20] , \wRegInBot_6_34[19] , 
        \wRegInBot_6_34[18] , \wRegInBot_6_34[17] , \wRegInBot_6_34[16] , 
        \wRegInBot_6_34[15] , \wRegInBot_6_34[14] , \wRegInBot_6_34[13] , 
        \wRegInBot_6_34[12] , \wRegInBot_6_34[11] , \wRegInBot_6_34[10] , 
        \wRegInBot_6_34[9] , \wRegInBot_6_34[8] , \wRegInBot_6_34[7] , 
        \wRegInBot_6_34[6] , \wRegInBot_6_34[5] , \wRegInBot_6_34[4] , 
        \wRegInBot_6_34[3] , \wRegInBot_6_34[2] , \wRegInBot_6_34[1] , 
        \wRegInBot_6_34[0] }), .L_WR(\wRegEnTop_7_68[0] ), .L_In({
        \wRegOut_7_68[31] , \wRegOut_7_68[30] , \wRegOut_7_68[29] , 
        \wRegOut_7_68[28] , \wRegOut_7_68[27] , \wRegOut_7_68[26] , 
        \wRegOut_7_68[25] , \wRegOut_7_68[24] , \wRegOut_7_68[23] , 
        \wRegOut_7_68[22] , \wRegOut_7_68[21] , \wRegOut_7_68[20] , 
        \wRegOut_7_68[19] , \wRegOut_7_68[18] , \wRegOut_7_68[17] , 
        \wRegOut_7_68[16] , \wRegOut_7_68[15] , \wRegOut_7_68[14] , 
        \wRegOut_7_68[13] , \wRegOut_7_68[12] , \wRegOut_7_68[11] , 
        \wRegOut_7_68[10] , \wRegOut_7_68[9] , \wRegOut_7_68[8] , 
        \wRegOut_7_68[7] , \wRegOut_7_68[6] , \wRegOut_7_68[5] , 
        \wRegOut_7_68[4] , \wRegOut_7_68[3] , \wRegOut_7_68[2] , 
        \wRegOut_7_68[1] , \wRegOut_7_68[0] }), .L_Out({\wRegInTop_7_68[31] , 
        \wRegInTop_7_68[30] , \wRegInTop_7_68[29] , \wRegInTop_7_68[28] , 
        \wRegInTop_7_68[27] , \wRegInTop_7_68[26] , \wRegInTop_7_68[25] , 
        \wRegInTop_7_68[24] , \wRegInTop_7_68[23] , \wRegInTop_7_68[22] , 
        \wRegInTop_7_68[21] , \wRegInTop_7_68[20] , \wRegInTop_7_68[19] , 
        \wRegInTop_7_68[18] , \wRegInTop_7_68[17] , \wRegInTop_7_68[16] , 
        \wRegInTop_7_68[15] , \wRegInTop_7_68[14] , \wRegInTop_7_68[13] , 
        \wRegInTop_7_68[12] , \wRegInTop_7_68[11] , \wRegInTop_7_68[10] , 
        \wRegInTop_7_68[9] , \wRegInTop_7_68[8] , \wRegInTop_7_68[7] , 
        \wRegInTop_7_68[6] , \wRegInTop_7_68[5] , \wRegInTop_7_68[4] , 
        \wRegInTop_7_68[3] , \wRegInTop_7_68[2] , \wRegInTop_7_68[1] , 
        \wRegInTop_7_68[0] }), .R_WR(\wRegEnTop_7_69[0] ), .R_In({
        \wRegOut_7_69[31] , \wRegOut_7_69[30] , \wRegOut_7_69[29] , 
        \wRegOut_7_69[28] , \wRegOut_7_69[27] , \wRegOut_7_69[26] , 
        \wRegOut_7_69[25] , \wRegOut_7_69[24] , \wRegOut_7_69[23] , 
        \wRegOut_7_69[22] , \wRegOut_7_69[21] , \wRegOut_7_69[20] , 
        \wRegOut_7_69[19] , \wRegOut_7_69[18] , \wRegOut_7_69[17] , 
        \wRegOut_7_69[16] , \wRegOut_7_69[15] , \wRegOut_7_69[14] , 
        \wRegOut_7_69[13] , \wRegOut_7_69[12] , \wRegOut_7_69[11] , 
        \wRegOut_7_69[10] , \wRegOut_7_69[9] , \wRegOut_7_69[8] , 
        \wRegOut_7_69[7] , \wRegOut_7_69[6] , \wRegOut_7_69[5] , 
        \wRegOut_7_69[4] , \wRegOut_7_69[3] , \wRegOut_7_69[2] , 
        \wRegOut_7_69[1] , \wRegOut_7_69[0] }), .R_Out({\wRegInTop_7_69[31] , 
        \wRegInTop_7_69[30] , \wRegInTop_7_69[29] , \wRegInTop_7_69[28] , 
        \wRegInTop_7_69[27] , \wRegInTop_7_69[26] , \wRegInTop_7_69[25] , 
        \wRegInTop_7_69[24] , \wRegInTop_7_69[23] , \wRegInTop_7_69[22] , 
        \wRegInTop_7_69[21] , \wRegInTop_7_69[20] , \wRegInTop_7_69[19] , 
        \wRegInTop_7_69[18] , \wRegInTop_7_69[17] , \wRegInTop_7_69[16] , 
        \wRegInTop_7_69[15] , \wRegInTop_7_69[14] , \wRegInTop_7_69[13] , 
        \wRegInTop_7_69[12] , \wRegInTop_7_69[11] , \wRegInTop_7_69[10] , 
        \wRegInTop_7_69[9] , \wRegInTop_7_69[8] , \wRegInTop_7_69[7] , 
        \wRegInTop_7_69[6] , \wRegInTop_7_69[5] , \wRegInTop_7_69[4] , 
        \wRegInTop_7_69[3] , \wRegInTop_7_69[2] , \wRegInTop_7_69[1] , 
        \wRegInTop_7_69[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_21 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink149[31] , \ScanLink149[30] , \ScanLink149[29] , 
        \ScanLink149[28] , \ScanLink149[27] , \ScanLink149[26] , 
        \ScanLink149[25] , \ScanLink149[24] , \ScanLink149[23] , 
        \ScanLink149[22] , \ScanLink149[21] , \ScanLink149[20] , 
        \ScanLink149[19] , \ScanLink149[18] , \ScanLink149[17] , 
        \ScanLink149[16] , \ScanLink149[15] , \ScanLink149[14] , 
        \ScanLink149[13] , \ScanLink149[12] , \ScanLink149[11] , 
        \ScanLink149[10] , \ScanLink149[9] , \ScanLink149[8] , 
        \ScanLink149[7] , \ScanLink149[6] , \ScanLink149[5] , \ScanLink149[4] , 
        \ScanLink149[3] , \ScanLink149[2] , \ScanLink149[1] , \ScanLink149[0] 
        }), .ScanOut({\ScanLink148[31] , \ScanLink148[30] , \ScanLink148[29] , 
        \ScanLink148[28] , \ScanLink148[27] , \ScanLink148[26] , 
        \ScanLink148[25] , \ScanLink148[24] , \ScanLink148[23] , 
        \ScanLink148[22] , \ScanLink148[21] , \ScanLink148[20] , 
        \ScanLink148[19] , \ScanLink148[18] , \ScanLink148[17] , 
        \ScanLink148[16] , \ScanLink148[15] , \ScanLink148[14] , 
        \ScanLink148[13] , \ScanLink148[12] , \ScanLink148[11] , 
        \ScanLink148[10] , \ScanLink148[9] , \ScanLink148[8] , 
        \ScanLink148[7] , \ScanLink148[6] , \ScanLink148[5] , \ScanLink148[4] , 
        \ScanLink148[3] , \ScanLink148[2] , \ScanLink148[1] , \ScanLink148[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_21[31] , 
        \wRegOut_7_21[30] , \wRegOut_7_21[29] , \wRegOut_7_21[28] , 
        \wRegOut_7_21[27] , \wRegOut_7_21[26] , \wRegOut_7_21[25] , 
        \wRegOut_7_21[24] , \wRegOut_7_21[23] , \wRegOut_7_21[22] , 
        \wRegOut_7_21[21] , \wRegOut_7_21[20] , \wRegOut_7_21[19] , 
        \wRegOut_7_21[18] , \wRegOut_7_21[17] , \wRegOut_7_21[16] , 
        \wRegOut_7_21[15] , \wRegOut_7_21[14] , \wRegOut_7_21[13] , 
        \wRegOut_7_21[12] , \wRegOut_7_21[11] , \wRegOut_7_21[10] , 
        \wRegOut_7_21[9] , \wRegOut_7_21[8] , \wRegOut_7_21[7] , 
        \wRegOut_7_21[6] , \wRegOut_7_21[5] , \wRegOut_7_21[4] , 
        \wRegOut_7_21[3] , \wRegOut_7_21[2] , \wRegOut_7_21[1] , 
        \wRegOut_7_21[0] }), .Enable1(\wRegEnTop_7_21[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_21[31] , \wRegInTop_7_21[30] , \wRegInTop_7_21[29] , 
        \wRegInTop_7_21[28] , \wRegInTop_7_21[27] , \wRegInTop_7_21[26] , 
        \wRegInTop_7_21[25] , \wRegInTop_7_21[24] , \wRegInTop_7_21[23] , 
        \wRegInTop_7_21[22] , \wRegInTop_7_21[21] , \wRegInTop_7_21[20] , 
        \wRegInTop_7_21[19] , \wRegInTop_7_21[18] , \wRegInTop_7_21[17] , 
        \wRegInTop_7_21[16] , \wRegInTop_7_21[15] , \wRegInTop_7_21[14] , 
        \wRegInTop_7_21[13] , \wRegInTop_7_21[12] , \wRegInTop_7_21[11] , 
        \wRegInTop_7_21[10] , \wRegInTop_7_21[9] , \wRegInTop_7_21[8] , 
        \wRegInTop_7_21[7] , \wRegInTop_7_21[6] , \wRegInTop_7_21[5] , 
        \wRegInTop_7_21[4] , \wRegInTop_7_21[3] , \wRegInTop_7_21[2] , 
        \wRegInTop_7_21[1] , \wRegInTop_7_21[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_1[0] ), .P_WR(\wRegEnBot_1_1[0] ), .P_In({\wRegOut_1_1[31] , 
        \wRegOut_1_1[30] , \wRegOut_1_1[29] , \wRegOut_1_1[28] , 
        \wRegOut_1_1[27] , \wRegOut_1_1[26] , \wRegOut_1_1[25] , 
        \wRegOut_1_1[24] , \wRegOut_1_1[23] , \wRegOut_1_1[22] , 
        \wRegOut_1_1[21] , \wRegOut_1_1[20] , \wRegOut_1_1[19] , 
        \wRegOut_1_1[18] , \wRegOut_1_1[17] , \wRegOut_1_1[16] , 
        \wRegOut_1_1[15] , \wRegOut_1_1[14] , \wRegOut_1_1[13] , 
        \wRegOut_1_1[12] , \wRegOut_1_1[11] , \wRegOut_1_1[10] , 
        \wRegOut_1_1[9] , \wRegOut_1_1[8] , \wRegOut_1_1[7] , \wRegOut_1_1[6] , 
        \wRegOut_1_1[5] , \wRegOut_1_1[4] , \wRegOut_1_1[3] , \wRegOut_1_1[2] , 
        \wRegOut_1_1[1] , \wRegOut_1_1[0] }), .P_Out({\wRegInBot_1_1[31] , 
        \wRegInBot_1_1[30] , \wRegInBot_1_1[29] , \wRegInBot_1_1[28] , 
        \wRegInBot_1_1[27] , \wRegInBot_1_1[26] , \wRegInBot_1_1[25] , 
        \wRegInBot_1_1[24] , \wRegInBot_1_1[23] , \wRegInBot_1_1[22] , 
        \wRegInBot_1_1[21] , \wRegInBot_1_1[20] , \wRegInBot_1_1[19] , 
        \wRegInBot_1_1[18] , \wRegInBot_1_1[17] , \wRegInBot_1_1[16] , 
        \wRegInBot_1_1[15] , \wRegInBot_1_1[14] , \wRegInBot_1_1[13] , 
        \wRegInBot_1_1[12] , \wRegInBot_1_1[11] , \wRegInBot_1_1[10] , 
        \wRegInBot_1_1[9] , \wRegInBot_1_1[8] , \wRegInBot_1_1[7] , 
        \wRegInBot_1_1[6] , \wRegInBot_1_1[5] , \wRegInBot_1_1[4] , 
        \wRegInBot_1_1[3] , \wRegInBot_1_1[2] , \wRegInBot_1_1[1] , 
        \wRegInBot_1_1[0] }), .L_WR(\wRegEnTop_2_2[0] ), .L_In({
        \wRegOut_2_2[31] , \wRegOut_2_2[30] , \wRegOut_2_2[29] , 
        \wRegOut_2_2[28] , \wRegOut_2_2[27] , \wRegOut_2_2[26] , 
        \wRegOut_2_2[25] , \wRegOut_2_2[24] , \wRegOut_2_2[23] , 
        \wRegOut_2_2[22] , \wRegOut_2_2[21] , \wRegOut_2_2[20] , 
        \wRegOut_2_2[19] , \wRegOut_2_2[18] , \wRegOut_2_2[17] , 
        \wRegOut_2_2[16] , \wRegOut_2_2[15] , \wRegOut_2_2[14] , 
        \wRegOut_2_2[13] , \wRegOut_2_2[12] , \wRegOut_2_2[11] , 
        \wRegOut_2_2[10] , \wRegOut_2_2[9] , \wRegOut_2_2[8] , 
        \wRegOut_2_2[7] , \wRegOut_2_2[6] , \wRegOut_2_2[5] , \wRegOut_2_2[4] , 
        \wRegOut_2_2[3] , \wRegOut_2_2[2] , \wRegOut_2_2[1] , \wRegOut_2_2[0] 
        }), .L_Out({\wRegInTop_2_2[31] , \wRegInTop_2_2[30] , 
        \wRegInTop_2_2[29] , \wRegInTop_2_2[28] , \wRegInTop_2_2[27] , 
        \wRegInTop_2_2[26] , \wRegInTop_2_2[25] , \wRegInTop_2_2[24] , 
        \wRegInTop_2_2[23] , \wRegInTop_2_2[22] , \wRegInTop_2_2[21] , 
        \wRegInTop_2_2[20] , \wRegInTop_2_2[19] , \wRegInTop_2_2[18] , 
        \wRegInTop_2_2[17] , \wRegInTop_2_2[16] , \wRegInTop_2_2[15] , 
        \wRegInTop_2_2[14] , \wRegInTop_2_2[13] , \wRegInTop_2_2[12] , 
        \wRegInTop_2_2[11] , \wRegInTop_2_2[10] , \wRegInTop_2_2[9] , 
        \wRegInTop_2_2[8] , \wRegInTop_2_2[7] , \wRegInTop_2_2[6] , 
        \wRegInTop_2_2[5] , \wRegInTop_2_2[4] , \wRegInTop_2_2[3] , 
        \wRegInTop_2_2[2] , \wRegInTop_2_2[1] , \wRegInTop_2_2[0] }), .R_WR(
        \wRegEnTop_2_3[0] ), .R_In({\wRegOut_2_3[31] , \wRegOut_2_3[30] , 
        \wRegOut_2_3[29] , \wRegOut_2_3[28] , \wRegOut_2_3[27] , 
        \wRegOut_2_3[26] , \wRegOut_2_3[25] , \wRegOut_2_3[24] , 
        \wRegOut_2_3[23] , \wRegOut_2_3[22] , \wRegOut_2_3[21] , 
        \wRegOut_2_3[20] , \wRegOut_2_3[19] , \wRegOut_2_3[18] , 
        \wRegOut_2_3[17] , \wRegOut_2_3[16] , \wRegOut_2_3[15] , 
        \wRegOut_2_3[14] , \wRegOut_2_3[13] , \wRegOut_2_3[12] , 
        \wRegOut_2_3[11] , \wRegOut_2_3[10] , \wRegOut_2_3[9] , 
        \wRegOut_2_3[8] , \wRegOut_2_3[7] , \wRegOut_2_3[6] , \wRegOut_2_3[5] , 
        \wRegOut_2_3[4] , \wRegOut_2_3[3] , \wRegOut_2_3[2] , \wRegOut_2_3[1] , 
        \wRegOut_2_3[0] }), .R_Out({\wRegInTop_2_3[31] , \wRegInTop_2_3[30] , 
        \wRegInTop_2_3[29] , \wRegInTop_2_3[28] , \wRegInTop_2_3[27] , 
        \wRegInTop_2_3[26] , \wRegInTop_2_3[25] , \wRegInTop_2_3[24] , 
        \wRegInTop_2_3[23] , \wRegInTop_2_3[22] , \wRegInTop_2_3[21] , 
        \wRegInTop_2_3[20] , \wRegInTop_2_3[19] , \wRegInTop_2_3[18] , 
        \wRegInTop_2_3[17] , \wRegInTop_2_3[16] , \wRegInTop_2_3[15] , 
        \wRegInTop_2_3[14] , \wRegInTop_2_3[13] , \wRegInTop_2_3[12] , 
        \wRegInTop_2_3[11] , \wRegInTop_2_3[10] , \wRegInTop_2_3[9] , 
        \wRegInTop_2_3[8] , \wRegInTop_2_3[7] , \wRegInTop_2_3[6] , 
        \wRegInTop_2_3[5] , \wRegInTop_2_3[4] , \wRegInTop_2_3[3] , 
        \wRegInTop_2_3[2] , \wRegInTop_2_3[1] , \wRegInTop_2_3[0] }) );
    BHeap_Node_WIDTH32 BHN_5_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_23[0] ), .P_In({\wRegOut_5_23[31] , 
        \wRegOut_5_23[30] , \wRegOut_5_23[29] , \wRegOut_5_23[28] , 
        \wRegOut_5_23[27] , \wRegOut_5_23[26] , \wRegOut_5_23[25] , 
        \wRegOut_5_23[24] , \wRegOut_5_23[23] , \wRegOut_5_23[22] , 
        \wRegOut_5_23[21] , \wRegOut_5_23[20] , \wRegOut_5_23[19] , 
        \wRegOut_5_23[18] , \wRegOut_5_23[17] , \wRegOut_5_23[16] , 
        \wRegOut_5_23[15] , \wRegOut_5_23[14] , \wRegOut_5_23[13] , 
        \wRegOut_5_23[12] , \wRegOut_5_23[11] , \wRegOut_5_23[10] , 
        \wRegOut_5_23[9] , \wRegOut_5_23[8] , \wRegOut_5_23[7] , 
        \wRegOut_5_23[6] , \wRegOut_5_23[5] , \wRegOut_5_23[4] , 
        \wRegOut_5_23[3] , \wRegOut_5_23[2] , \wRegOut_5_23[1] , 
        \wRegOut_5_23[0] }), .P_Out({\wRegInBot_5_23[31] , 
        \wRegInBot_5_23[30] , \wRegInBot_5_23[29] , \wRegInBot_5_23[28] , 
        \wRegInBot_5_23[27] , \wRegInBot_5_23[26] , \wRegInBot_5_23[25] , 
        \wRegInBot_5_23[24] , \wRegInBot_5_23[23] , \wRegInBot_5_23[22] , 
        \wRegInBot_5_23[21] , \wRegInBot_5_23[20] , \wRegInBot_5_23[19] , 
        \wRegInBot_5_23[18] , \wRegInBot_5_23[17] , \wRegInBot_5_23[16] , 
        \wRegInBot_5_23[15] , \wRegInBot_5_23[14] , \wRegInBot_5_23[13] , 
        \wRegInBot_5_23[12] , \wRegInBot_5_23[11] , \wRegInBot_5_23[10] , 
        \wRegInBot_5_23[9] , \wRegInBot_5_23[8] , \wRegInBot_5_23[7] , 
        \wRegInBot_5_23[6] , \wRegInBot_5_23[5] , \wRegInBot_5_23[4] , 
        \wRegInBot_5_23[3] , \wRegInBot_5_23[2] , \wRegInBot_5_23[1] , 
        \wRegInBot_5_23[0] }), .L_WR(\wRegEnTop_6_46[0] ), .L_In({
        \wRegOut_6_46[31] , \wRegOut_6_46[30] , \wRegOut_6_46[29] , 
        \wRegOut_6_46[28] , \wRegOut_6_46[27] , \wRegOut_6_46[26] , 
        \wRegOut_6_46[25] , \wRegOut_6_46[24] , \wRegOut_6_46[23] , 
        \wRegOut_6_46[22] , \wRegOut_6_46[21] , \wRegOut_6_46[20] , 
        \wRegOut_6_46[19] , \wRegOut_6_46[18] , \wRegOut_6_46[17] , 
        \wRegOut_6_46[16] , \wRegOut_6_46[15] , \wRegOut_6_46[14] , 
        \wRegOut_6_46[13] , \wRegOut_6_46[12] , \wRegOut_6_46[11] , 
        \wRegOut_6_46[10] , \wRegOut_6_46[9] , \wRegOut_6_46[8] , 
        \wRegOut_6_46[7] , \wRegOut_6_46[6] , \wRegOut_6_46[5] , 
        \wRegOut_6_46[4] , \wRegOut_6_46[3] , \wRegOut_6_46[2] , 
        \wRegOut_6_46[1] , \wRegOut_6_46[0] }), .L_Out({\wRegInTop_6_46[31] , 
        \wRegInTop_6_46[30] , \wRegInTop_6_46[29] , \wRegInTop_6_46[28] , 
        \wRegInTop_6_46[27] , \wRegInTop_6_46[26] , \wRegInTop_6_46[25] , 
        \wRegInTop_6_46[24] , \wRegInTop_6_46[23] , \wRegInTop_6_46[22] , 
        \wRegInTop_6_46[21] , \wRegInTop_6_46[20] , \wRegInTop_6_46[19] , 
        \wRegInTop_6_46[18] , \wRegInTop_6_46[17] , \wRegInTop_6_46[16] , 
        \wRegInTop_6_46[15] , \wRegInTop_6_46[14] , \wRegInTop_6_46[13] , 
        \wRegInTop_6_46[12] , \wRegInTop_6_46[11] , \wRegInTop_6_46[10] , 
        \wRegInTop_6_46[9] , \wRegInTop_6_46[8] , \wRegInTop_6_46[7] , 
        \wRegInTop_6_46[6] , \wRegInTop_6_46[5] , \wRegInTop_6_46[4] , 
        \wRegInTop_6_46[3] , \wRegInTop_6_46[2] , \wRegInTop_6_46[1] , 
        \wRegInTop_6_46[0] }), .R_WR(\wRegEnTop_6_47[0] ), .R_In({
        \wRegOut_6_47[31] , \wRegOut_6_47[30] , \wRegOut_6_47[29] , 
        \wRegOut_6_47[28] , \wRegOut_6_47[27] , \wRegOut_6_47[26] , 
        \wRegOut_6_47[25] , \wRegOut_6_47[24] , \wRegOut_6_47[23] , 
        \wRegOut_6_47[22] , \wRegOut_6_47[21] , \wRegOut_6_47[20] , 
        \wRegOut_6_47[19] , \wRegOut_6_47[18] , \wRegOut_6_47[17] , 
        \wRegOut_6_47[16] , \wRegOut_6_47[15] , \wRegOut_6_47[14] , 
        \wRegOut_6_47[13] , \wRegOut_6_47[12] , \wRegOut_6_47[11] , 
        \wRegOut_6_47[10] , \wRegOut_6_47[9] , \wRegOut_6_47[8] , 
        \wRegOut_6_47[7] , \wRegOut_6_47[6] , \wRegOut_6_47[5] , 
        \wRegOut_6_47[4] , \wRegOut_6_47[3] , \wRegOut_6_47[2] , 
        \wRegOut_6_47[1] , \wRegOut_6_47[0] }), .R_Out({\wRegInTop_6_47[31] , 
        \wRegInTop_6_47[30] , \wRegInTop_6_47[29] , \wRegInTop_6_47[28] , 
        \wRegInTop_6_47[27] , \wRegInTop_6_47[26] , \wRegInTop_6_47[25] , 
        \wRegInTop_6_47[24] , \wRegInTop_6_47[23] , \wRegInTop_6_47[22] , 
        \wRegInTop_6_47[21] , \wRegInTop_6_47[20] , \wRegInTop_6_47[19] , 
        \wRegInTop_6_47[18] , \wRegInTop_6_47[17] , \wRegInTop_6_47[16] , 
        \wRegInTop_6_47[15] , \wRegInTop_6_47[14] , \wRegInTop_6_47[13] , 
        \wRegInTop_6_47[12] , \wRegInTop_6_47[11] , \wRegInTop_6_47[10] , 
        \wRegInTop_6_47[9] , \wRegInTop_6_47[8] , \wRegInTop_6_47[7] , 
        \wRegInTop_6_47[6] , \wRegInTop_6_47[5] , \wRegInTop_6_47[4] , 
        \wRegInTop_6_47[3] , \wRegInTop_6_47[2] , \wRegInTop_6_47[1] , 
        \wRegInTop_6_47[0] }) );
    BHeap_Node_WIDTH32 BHN_6_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_13[0] ), .P_In({\wRegOut_6_13[31] , 
        \wRegOut_6_13[30] , \wRegOut_6_13[29] , \wRegOut_6_13[28] , 
        \wRegOut_6_13[27] , \wRegOut_6_13[26] , \wRegOut_6_13[25] , 
        \wRegOut_6_13[24] , \wRegOut_6_13[23] , \wRegOut_6_13[22] , 
        \wRegOut_6_13[21] , \wRegOut_6_13[20] , \wRegOut_6_13[19] , 
        \wRegOut_6_13[18] , \wRegOut_6_13[17] , \wRegOut_6_13[16] , 
        \wRegOut_6_13[15] , \wRegOut_6_13[14] , \wRegOut_6_13[13] , 
        \wRegOut_6_13[12] , \wRegOut_6_13[11] , \wRegOut_6_13[10] , 
        \wRegOut_6_13[9] , \wRegOut_6_13[8] , \wRegOut_6_13[7] , 
        \wRegOut_6_13[6] , \wRegOut_6_13[5] , \wRegOut_6_13[4] , 
        \wRegOut_6_13[3] , \wRegOut_6_13[2] , \wRegOut_6_13[1] , 
        \wRegOut_6_13[0] }), .P_Out({\wRegInBot_6_13[31] , 
        \wRegInBot_6_13[30] , \wRegInBot_6_13[29] , \wRegInBot_6_13[28] , 
        \wRegInBot_6_13[27] , \wRegInBot_6_13[26] , \wRegInBot_6_13[25] , 
        \wRegInBot_6_13[24] , \wRegInBot_6_13[23] , \wRegInBot_6_13[22] , 
        \wRegInBot_6_13[21] , \wRegInBot_6_13[20] , \wRegInBot_6_13[19] , 
        \wRegInBot_6_13[18] , \wRegInBot_6_13[17] , \wRegInBot_6_13[16] , 
        \wRegInBot_6_13[15] , \wRegInBot_6_13[14] , \wRegInBot_6_13[13] , 
        \wRegInBot_6_13[12] , \wRegInBot_6_13[11] , \wRegInBot_6_13[10] , 
        \wRegInBot_6_13[9] , \wRegInBot_6_13[8] , \wRegInBot_6_13[7] , 
        \wRegInBot_6_13[6] , \wRegInBot_6_13[5] , \wRegInBot_6_13[4] , 
        \wRegInBot_6_13[3] , \wRegInBot_6_13[2] , \wRegInBot_6_13[1] , 
        \wRegInBot_6_13[0] }), .L_WR(\wRegEnTop_7_26[0] ), .L_In({
        \wRegOut_7_26[31] , \wRegOut_7_26[30] , \wRegOut_7_26[29] , 
        \wRegOut_7_26[28] , \wRegOut_7_26[27] , \wRegOut_7_26[26] , 
        \wRegOut_7_26[25] , \wRegOut_7_26[24] , \wRegOut_7_26[23] , 
        \wRegOut_7_26[22] , \wRegOut_7_26[21] , \wRegOut_7_26[20] , 
        \wRegOut_7_26[19] , \wRegOut_7_26[18] , \wRegOut_7_26[17] , 
        \wRegOut_7_26[16] , \wRegOut_7_26[15] , \wRegOut_7_26[14] , 
        \wRegOut_7_26[13] , \wRegOut_7_26[12] , \wRegOut_7_26[11] , 
        \wRegOut_7_26[10] , \wRegOut_7_26[9] , \wRegOut_7_26[8] , 
        \wRegOut_7_26[7] , \wRegOut_7_26[6] , \wRegOut_7_26[5] , 
        \wRegOut_7_26[4] , \wRegOut_7_26[3] , \wRegOut_7_26[2] , 
        \wRegOut_7_26[1] , \wRegOut_7_26[0] }), .L_Out({\wRegInTop_7_26[31] , 
        \wRegInTop_7_26[30] , \wRegInTop_7_26[29] , \wRegInTop_7_26[28] , 
        \wRegInTop_7_26[27] , \wRegInTop_7_26[26] , \wRegInTop_7_26[25] , 
        \wRegInTop_7_26[24] , \wRegInTop_7_26[23] , \wRegInTop_7_26[22] , 
        \wRegInTop_7_26[21] , \wRegInTop_7_26[20] , \wRegInTop_7_26[19] , 
        \wRegInTop_7_26[18] , \wRegInTop_7_26[17] , \wRegInTop_7_26[16] , 
        \wRegInTop_7_26[15] , \wRegInTop_7_26[14] , \wRegInTop_7_26[13] , 
        \wRegInTop_7_26[12] , \wRegInTop_7_26[11] , \wRegInTop_7_26[10] , 
        \wRegInTop_7_26[9] , \wRegInTop_7_26[8] , \wRegInTop_7_26[7] , 
        \wRegInTop_7_26[6] , \wRegInTop_7_26[5] , \wRegInTop_7_26[4] , 
        \wRegInTop_7_26[3] , \wRegInTop_7_26[2] , \wRegInTop_7_26[1] , 
        \wRegInTop_7_26[0] }), .R_WR(\wRegEnTop_7_27[0] ), .R_In({
        \wRegOut_7_27[31] , \wRegOut_7_27[30] , \wRegOut_7_27[29] , 
        \wRegOut_7_27[28] , \wRegOut_7_27[27] , \wRegOut_7_27[26] , 
        \wRegOut_7_27[25] , \wRegOut_7_27[24] , \wRegOut_7_27[23] , 
        \wRegOut_7_27[22] , \wRegOut_7_27[21] , \wRegOut_7_27[20] , 
        \wRegOut_7_27[19] , \wRegOut_7_27[18] , \wRegOut_7_27[17] , 
        \wRegOut_7_27[16] , \wRegOut_7_27[15] , \wRegOut_7_27[14] , 
        \wRegOut_7_27[13] , \wRegOut_7_27[12] , \wRegOut_7_27[11] , 
        \wRegOut_7_27[10] , \wRegOut_7_27[9] , \wRegOut_7_27[8] , 
        \wRegOut_7_27[7] , \wRegOut_7_27[6] , \wRegOut_7_27[5] , 
        \wRegOut_7_27[4] , \wRegOut_7_27[3] , \wRegOut_7_27[2] , 
        \wRegOut_7_27[1] , \wRegOut_7_27[0] }), .R_Out({\wRegInTop_7_27[31] , 
        \wRegInTop_7_27[30] , \wRegInTop_7_27[29] , \wRegInTop_7_27[28] , 
        \wRegInTop_7_27[27] , \wRegInTop_7_27[26] , \wRegInTop_7_27[25] , 
        \wRegInTop_7_27[24] , \wRegInTop_7_27[23] , \wRegInTop_7_27[22] , 
        \wRegInTop_7_27[21] , \wRegInTop_7_27[20] , \wRegInTop_7_27[19] , 
        \wRegInTop_7_27[18] , \wRegInTop_7_27[17] , \wRegInTop_7_27[16] , 
        \wRegInTop_7_27[15] , \wRegInTop_7_27[14] , \wRegInTop_7_27[13] , 
        \wRegInTop_7_27[12] , \wRegInTop_7_27[11] , \wRegInTop_7_27[10] , 
        \wRegInTop_7_27[9] , \wRegInTop_7_27[8] , \wRegInTop_7_27[7] , 
        \wRegInTop_7_27[6] , \wRegInTop_7_27[5] , \wRegInTop_7_27[4] , 
        \wRegInTop_7_27[3] , \wRegInTop_7_27[2] , \wRegInTop_7_27[1] , 
        \wRegInTop_7_27[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink42[31] , \ScanLink42[30] , \ScanLink42[29] , 
        \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , \ScanLink42[25] , 
        \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , \ScanLink42[21] , 
        \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , \ScanLink42[17] , 
        \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , \ScanLink42[13] , 
        \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , \ScanLink42[9] , 
        \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , \ScanLink42[5] , 
        \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , \ScanLink42[1] , 
        \ScanLink42[0] }), .ScanOut({\ScanLink41[31] , \ScanLink41[30] , 
        \ScanLink41[29] , \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , 
        \ScanLink41[25] , \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , 
        \ScanLink41[21] , \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , 
        \ScanLink41[17] , \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , 
        \ScanLink41[13] , \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , 
        \ScanLink41[9] , \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , 
        \ScanLink41[5] , \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , 
        \ScanLink41[1] , \ScanLink41[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_10[31] , \wRegOut_5_10[30] , 
        \wRegOut_5_10[29] , \wRegOut_5_10[28] , \wRegOut_5_10[27] , 
        \wRegOut_5_10[26] , \wRegOut_5_10[25] , \wRegOut_5_10[24] , 
        \wRegOut_5_10[23] , \wRegOut_5_10[22] , \wRegOut_5_10[21] , 
        \wRegOut_5_10[20] , \wRegOut_5_10[19] , \wRegOut_5_10[18] , 
        \wRegOut_5_10[17] , \wRegOut_5_10[16] , \wRegOut_5_10[15] , 
        \wRegOut_5_10[14] , \wRegOut_5_10[13] , \wRegOut_5_10[12] , 
        \wRegOut_5_10[11] , \wRegOut_5_10[10] , \wRegOut_5_10[9] , 
        \wRegOut_5_10[8] , \wRegOut_5_10[7] , \wRegOut_5_10[6] , 
        \wRegOut_5_10[5] , \wRegOut_5_10[4] , \wRegOut_5_10[3] , 
        \wRegOut_5_10[2] , \wRegOut_5_10[1] , \wRegOut_5_10[0] }), .Enable1(
        \wRegEnTop_5_10[0] ), .Enable2(\wRegEnBot_5_10[0] ), .In1({
        \wRegInTop_5_10[31] , \wRegInTop_5_10[30] , \wRegInTop_5_10[29] , 
        \wRegInTop_5_10[28] , \wRegInTop_5_10[27] , \wRegInTop_5_10[26] , 
        \wRegInTop_5_10[25] , \wRegInTop_5_10[24] , \wRegInTop_5_10[23] , 
        \wRegInTop_5_10[22] , \wRegInTop_5_10[21] , \wRegInTop_5_10[20] , 
        \wRegInTop_5_10[19] , \wRegInTop_5_10[18] , \wRegInTop_5_10[17] , 
        \wRegInTop_5_10[16] , \wRegInTop_5_10[15] , \wRegInTop_5_10[14] , 
        \wRegInTop_5_10[13] , \wRegInTop_5_10[12] , \wRegInTop_5_10[11] , 
        \wRegInTop_5_10[10] , \wRegInTop_5_10[9] , \wRegInTop_5_10[8] , 
        \wRegInTop_5_10[7] , \wRegInTop_5_10[6] , \wRegInTop_5_10[5] , 
        \wRegInTop_5_10[4] , \wRegInTop_5_10[3] , \wRegInTop_5_10[2] , 
        \wRegInTop_5_10[1] , \wRegInTop_5_10[0] }), .In2({\wRegInBot_5_10[31] , 
        \wRegInBot_5_10[30] , \wRegInBot_5_10[29] , \wRegInBot_5_10[28] , 
        \wRegInBot_5_10[27] , \wRegInBot_5_10[26] , \wRegInBot_5_10[25] , 
        \wRegInBot_5_10[24] , \wRegInBot_5_10[23] , \wRegInBot_5_10[22] , 
        \wRegInBot_5_10[21] , \wRegInBot_5_10[20] , \wRegInBot_5_10[19] , 
        \wRegInBot_5_10[18] , \wRegInBot_5_10[17] , \wRegInBot_5_10[16] , 
        \wRegInBot_5_10[15] , \wRegInBot_5_10[14] , \wRegInBot_5_10[13] , 
        \wRegInBot_5_10[12] , \wRegInBot_5_10[11] , \wRegInBot_5_10[10] , 
        \wRegInBot_5_10[9] , \wRegInBot_5_10[8] , \wRegInBot_5_10[7] , 
        \wRegInBot_5_10[6] , \wRegInBot_5_10[5] , \wRegInBot_5_10[4] , 
        \wRegInBot_5_10[3] , \wRegInBot_5_10[2] , \wRegInBot_5_10[1] , 
        \wRegInBot_5_10[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_20 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink84[31] , \ScanLink84[30] , \ScanLink84[29] , 
        \ScanLink84[28] , \ScanLink84[27] , \ScanLink84[26] , \ScanLink84[25] , 
        \ScanLink84[24] , \ScanLink84[23] , \ScanLink84[22] , \ScanLink84[21] , 
        \ScanLink84[20] , \ScanLink84[19] , \ScanLink84[18] , \ScanLink84[17] , 
        \ScanLink84[16] , \ScanLink84[15] , \ScanLink84[14] , \ScanLink84[13] , 
        \ScanLink84[12] , \ScanLink84[11] , \ScanLink84[10] , \ScanLink84[9] , 
        \ScanLink84[8] , \ScanLink84[7] , \ScanLink84[6] , \ScanLink84[5] , 
        \ScanLink84[4] , \ScanLink84[3] , \ScanLink84[2] , \ScanLink84[1] , 
        \ScanLink84[0] }), .ScanOut({\ScanLink83[31] , \ScanLink83[30] , 
        \ScanLink83[29] , \ScanLink83[28] , \ScanLink83[27] , \ScanLink83[26] , 
        \ScanLink83[25] , \ScanLink83[24] , \ScanLink83[23] , \ScanLink83[22] , 
        \ScanLink83[21] , \ScanLink83[20] , \ScanLink83[19] , \ScanLink83[18] , 
        \ScanLink83[17] , \ScanLink83[16] , \ScanLink83[15] , \ScanLink83[14] , 
        \ScanLink83[13] , \ScanLink83[12] , \ScanLink83[11] , \ScanLink83[10] , 
        \ScanLink83[9] , \ScanLink83[8] , \ScanLink83[7] , \ScanLink83[6] , 
        \ScanLink83[5] , \ScanLink83[4] , \ScanLink83[3] , \ScanLink83[2] , 
        \ScanLink83[1] , \ScanLink83[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_20[31] , \wRegOut_6_20[30] , 
        \wRegOut_6_20[29] , \wRegOut_6_20[28] , \wRegOut_6_20[27] , 
        \wRegOut_6_20[26] , \wRegOut_6_20[25] , \wRegOut_6_20[24] , 
        \wRegOut_6_20[23] , \wRegOut_6_20[22] , \wRegOut_6_20[21] , 
        \wRegOut_6_20[20] , \wRegOut_6_20[19] , \wRegOut_6_20[18] , 
        \wRegOut_6_20[17] , \wRegOut_6_20[16] , \wRegOut_6_20[15] , 
        \wRegOut_6_20[14] , \wRegOut_6_20[13] , \wRegOut_6_20[12] , 
        \wRegOut_6_20[11] , \wRegOut_6_20[10] , \wRegOut_6_20[9] , 
        \wRegOut_6_20[8] , \wRegOut_6_20[7] , \wRegOut_6_20[6] , 
        \wRegOut_6_20[5] , \wRegOut_6_20[4] , \wRegOut_6_20[3] , 
        \wRegOut_6_20[2] , \wRegOut_6_20[1] , \wRegOut_6_20[0] }), .Enable1(
        \wRegEnTop_6_20[0] ), .Enable2(\wRegEnBot_6_20[0] ), .In1({
        \wRegInTop_6_20[31] , \wRegInTop_6_20[30] , \wRegInTop_6_20[29] , 
        \wRegInTop_6_20[28] , \wRegInTop_6_20[27] , \wRegInTop_6_20[26] , 
        \wRegInTop_6_20[25] , \wRegInTop_6_20[24] , \wRegInTop_6_20[23] , 
        \wRegInTop_6_20[22] , \wRegInTop_6_20[21] , \wRegInTop_6_20[20] , 
        \wRegInTop_6_20[19] , \wRegInTop_6_20[18] , \wRegInTop_6_20[17] , 
        \wRegInTop_6_20[16] , \wRegInTop_6_20[15] , \wRegInTop_6_20[14] , 
        \wRegInTop_6_20[13] , \wRegInTop_6_20[12] , \wRegInTop_6_20[11] , 
        \wRegInTop_6_20[10] , \wRegInTop_6_20[9] , \wRegInTop_6_20[8] , 
        \wRegInTop_6_20[7] , \wRegInTop_6_20[6] , \wRegInTop_6_20[5] , 
        \wRegInTop_6_20[4] , \wRegInTop_6_20[3] , \wRegInTop_6_20[2] , 
        \wRegInTop_6_20[1] , \wRegInTop_6_20[0] }), .In2({\wRegInBot_6_20[31] , 
        \wRegInBot_6_20[30] , \wRegInBot_6_20[29] , \wRegInBot_6_20[28] , 
        \wRegInBot_6_20[27] , \wRegInBot_6_20[26] , \wRegInBot_6_20[25] , 
        \wRegInBot_6_20[24] , \wRegInBot_6_20[23] , \wRegInBot_6_20[22] , 
        \wRegInBot_6_20[21] , \wRegInBot_6_20[20] , \wRegInBot_6_20[19] , 
        \wRegInBot_6_20[18] , \wRegInBot_6_20[17] , \wRegInBot_6_20[16] , 
        \wRegInBot_6_20[15] , \wRegInBot_6_20[14] , \wRegInBot_6_20[13] , 
        \wRegInBot_6_20[12] , \wRegInBot_6_20[11] , \wRegInBot_6_20[10] , 
        \wRegInBot_6_20[9] , \wRegInBot_6_20[8] , \wRegInBot_6_20[7] , 
        \wRegInBot_6_20[6] , \wRegInBot_6_20[5] , \wRegInBot_6_20[4] , 
        \wRegInBot_6_20[3] , \wRegInBot_6_20[2] , \wRegInBot_6_20[1] , 
        \wRegInBot_6_20[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_96 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink224[31] , \ScanLink224[30] , \ScanLink224[29] , 
        \ScanLink224[28] , \ScanLink224[27] , \ScanLink224[26] , 
        \ScanLink224[25] , \ScanLink224[24] , \ScanLink224[23] , 
        \ScanLink224[22] , \ScanLink224[21] , \ScanLink224[20] , 
        \ScanLink224[19] , \ScanLink224[18] , \ScanLink224[17] , 
        \ScanLink224[16] , \ScanLink224[15] , \ScanLink224[14] , 
        \ScanLink224[13] , \ScanLink224[12] , \ScanLink224[11] , 
        \ScanLink224[10] , \ScanLink224[9] , \ScanLink224[8] , 
        \ScanLink224[7] , \ScanLink224[6] , \ScanLink224[5] , \ScanLink224[4] , 
        \ScanLink224[3] , \ScanLink224[2] , \ScanLink224[1] , \ScanLink224[0] 
        }), .ScanOut({\ScanLink223[31] , \ScanLink223[30] , \ScanLink223[29] , 
        \ScanLink223[28] , \ScanLink223[27] , \ScanLink223[26] , 
        \ScanLink223[25] , \ScanLink223[24] , \ScanLink223[23] , 
        \ScanLink223[22] , \ScanLink223[21] , \ScanLink223[20] , 
        \ScanLink223[19] , \ScanLink223[18] , \ScanLink223[17] , 
        \ScanLink223[16] , \ScanLink223[15] , \ScanLink223[14] , 
        \ScanLink223[13] , \ScanLink223[12] , \ScanLink223[11] , 
        \ScanLink223[10] , \ScanLink223[9] , \ScanLink223[8] , 
        \ScanLink223[7] , \ScanLink223[6] , \ScanLink223[5] , \ScanLink223[4] , 
        \ScanLink223[3] , \ScanLink223[2] , \ScanLink223[1] , \ScanLink223[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_96[31] , 
        \wRegOut_7_96[30] , \wRegOut_7_96[29] , \wRegOut_7_96[28] , 
        \wRegOut_7_96[27] , \wRegOut_7_96[26] , \wRegOut_7_96[25] , 
        \wRegOut_7_96[24] , \wRegOut_7_96[23] , \wRegOut_7_96[22] , 
        \wRegOut_7_96[21] , \wRegOut_7_96[20] , \wRegOut_7_96[19] , 
        \wRegOut_7_96[18] , \wRegOut_7_96[17] , \wRegOut_7_96[16] , 
        \wRegOut_7_96[15] , \wRegOut_7_96[14] , \wRegOut_7_96[13] , 
        \wRegOut_7_96[12] , \wRegOut_7_96[11] , \wRegOut_7_96[10] , 
        \wRegOut_7_96[9] , \wRegOut_7_96[8] , \wRegOut_7_96[7] , 
        \wRegOut_7_96[6] , \wRegOut_7_96[5] , \wRegOut_7_96[4] , 
        \wRegOut_7_96[3] , \wRegOut_7_96[2] , \wRegOut_7_96[1] , 
        \wRegOut_7_96[0] }), .Enable1(\wRegEnTop_7_96[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_96[31] , \wRegInTop_7_96[30] , \wRegInTop_7_96[29] , 
        \wRegInTop_7_96[28] , \wRegInTop_7_96[27] , \wRegInTop_7_96[26] , 
        \wRegInTop_7_96[25] , \wRegInTop_7_96[24] , \wRegInTop_7_96[23] , 
        \wRegInTop_7_96[22] , \wRegInTop_7_96[21] , \wRegInTop_7_96[20] , 
        \wRegInTop_7_96[19] , \wRegInTop_7_96[18] , \wRegInTop_7_96[17] , 
        \wRegInTop_7_96[16] , \wRegInTop_7_96[15] , \wRegInTop_7_96[14] , 
        \wRegInTop_7_96[13] , \wRegInTop_7_96[12] , \wRegInTop_7_96[11] , 
        \wRegInTop_7_96[10] , \wRegInTop_7_96[9] , \wRegInTop_7_96[8] , 
        \wRegInTop_7_96[7] , \wRegInTop_7_96[6] , \wRegInTop_7_96[5] , 
        \wRegInTop_7_96[4] , \wRegInTop_7_96[3] , \wRegInTop_7_96[2] , 
        \wRegInTop_7_96[1] , \wRegInTop_7_96[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_112 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink240[31] , \ScanLink240[30] , \ScanLink240[29] , 
        \ScanLink240[28] , \ScanLink240[27] , \ScanLink240[26] , 
        \ScanLink240[25] , \ScanLink240[24] , \ScanLink240[23] , 
        \ScanLink240[22] , \ScanLink240[21] , \ScanLink240[20] , 
        \ScanLink240[19] , \ScanLink240[18] , \ScanLink240[17] , 
        \ScanLink240[16] , \ScanLink240[15] , \ScanLink240[14] , 
        \ScanLink240[13] , \ScanLink240[12] , \ScanLink240[11] , 
        \ScanLink240[10] , \ScanLink240[9] , \ScanLink240[8] , 
        \ScanLink240[7] , \ScanLink240[6] , \ScanLink240[5] , \ScanLink240[4] , 
        \ScanLink240[3] , \ScanLink240[2] , \ScanLink240[1] , \ScanLink240[0] 
        }), .ScanOut({\ScanLink239[31] , \ScanLink239[30] , \ScanLink239[29] , 
        \ScanLink239[28] , \ScanLink239[27] , \ScanLink239[26] , 
        \ScanLink239[25] , \ScanLink239[24] , \ScanLink239[23] , 
        \ScanLink239[22] , \ScanLink239[21] , \ScanLink239[20] , 
        \ScanLink239[19] , \ScanLink239[18] , \ScanLink239[17] , 
        \ScanLink239[16] , \ScanLink239[15] , \ScanLink239[14] , 
        \ScanLink239[13] , \ScanLink239[12] , \ScanLink239[11] , 
        \ScanLink239[10] , \ScanLink239[9] , \ScanLink239[8] , 
        \ScanLink239[7] , \ScanLink239[6] , \ScanLink239[5] , \ScanLink239[4] , 
        \ScanLink239[3] , \ScanLink239[2] , \ScanLink239[1] , \ScanLink239[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_112[31] , 
        \wRegOut_7_112[30] , \wRegOut_7_112[29] , \wRegOut_7_112[28] , 
        \wRegOut_7_112[27] , \wRegOut_7_112[26] , \wRegOut_7_112[25] , 
        \wRegOut_7_112[24] , \wRegOut_7_112[23] , \wRegOut_7_112[22] , 
        \wRegOut_7_112[21] , \wRegOut_7_112[20] , \wRegOut_7_112[19] , 
        \wRegOut_7_112[18] , \wRegOut_7_112[17] , \wRegOut_7_112[16] , 
        \wRegOut_7_112[15] , \wRegOut_7_112[14] , \wRegOut_7_112[13] , 
        \wRegOut_7_112[12] , \wRegOut_7_112[11] , \wRegOut_7_112[10] , 
        \wRegOut_7_112[9] , \wRegOut_7_112[8] , \wRegOut_7_112[7] , 
        \wRegOut_7_112[6] , \wRegOut_7_112[5] , \wRegOut_7_112[4] , 
        \wRegOut_7_112[3] , \wRegOut_7_112[2] , \wRegOut_7_112[1] , 
        \wRegOut_7_112[0] }), .Enable1(\wRegEnTop_7_112[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_112[31] , \wRegInTop_7_112[30] , 
        \wRegInTop_7_112[29] , \wRegInTop_7_112[28] , \wRegInTop_7_112[27] , 
        \wRegInTop_7_112[26] , \wRegInTop_7_112[25] , \wRegInTop_7_112[24] , 
        \wRegInTop_7_112[23] , \wRegInTop_7_112[22] , \wRegInTop_7_112[21] , 
        \wRegInTop_7_112[20] , \wRegInTop_7_112[19] , \wRegInTop_7_112[18] , 
        \wRegInTop_7_112[17] , \wRegInTop_7_112[16] , \wRegInTop_7_112[15] , 
        \wRegInTop_7_112[14] , \wRegInTop_7_112[13] , \wRegInTop_7_112[12] , 
        \wRegInTop_7_112[11] , \wRegInTop_7_112[10] , \wRegInTop_7_112[9] , 
        \wRegInTop_7_112[8] , \wRegInTop_7_112[7] , \wRegInTop_7_112[6] , 
        \wRegInTop_7_112[5] , \wRegInTop_7_112[4] , \wRegInTop_7_112[3] , 
        \wRegInTop_7_112[2] , \wRegInTop_7_112[1] , \wRegInTop_7_112[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_7[0] ), .P_In({\wRegOut_4_7[31] , 
        \wRegOut_4_7[30] , \wRegOut_4_7[29] , \wRegOut_4_7[28] , 
        \wRegOut_4_7[27] , \wRegOut_4_7[26] , \wRegOut_4_7[25] , 
        \wRegOut_4_7[24] , \wRegOut_4_7[23] , \wRegOut_4_7[22] , 
        \wRegOut_4_7[21] , \wRegOut_4_7[20] , \wRegOut_4_7[19] , 
        \wRegOut_4_7[18] , \wRegOut_4_7[17] , \wRegOut_4_7[16] , 
        \wRegOut_4_7[15] , \wRegOut_4_7[14] , \wRegOut_4_7[13] , 
        \wRegOut_4_7[12] , \wRegOut_4_7[11] , \wRegOut_4_7[10] , 
        \wRegOut_4_7[9] , \wRegOut_4_7[8] , \wRegOut_4_7[7] , \wRegOut_4_7[6] , 
        \wRegOut_4_7[5] , \wRegOut_4_7[4] , \wRegOut_4_7[3] , \wRegOut_4_7[2] , 
        \wRegOut_4_7[1] , \wRegOut_4_7[0] }), .P_Out({\wRegInBot_4_7[31] , 
        \wRegInBot_4_7[30] , \wRegInBot_4_7[29] , \wRegInBot_4_7[28] , 
        \wRegInBot_4_7[27] , \wRegInBot_4_7[26] , \wRegInBot_4_7[25] , 
        \wRegInBot_4_7[24] , \wRegInBot_4_7[23] , \wRegInBot_4_7[22] , 
        \wRegInBot_4_7[21] , \wRegInBot_4_7[20] , \wRegInBot_4_7[19] , 
        \wRegInBot_4_7[18] , \wRegInBot_4_7[17] , \wRegInBot_4_7[16] , 
        \wRegInBot_4_7[15] , \wRegInBot_4_7[14] , \wRegInBot_4_7[13] , 
        \wRegInBot_4_7[12] , \wRegInBot_4_7[11] , \wRegInBot_4_7[10] , 
        \wRegInBot_4_7[9] , \wRegInBot_4_7[8] , \wRegInBot_4_7[7] , 
        \wRegInBot_4_7[6] , \wRegInBot_4_7[5] , \wRegInBot_4_7[4] , 
        \wRegInBot_4_7[3] , \wRegInBot_4_7[2] , \wRegInBot_4_7[1] , 
        \wRegInBot_4_7[0] }), .L_WR(\wRegEnTop_5_14[0] ), .L_In({
        \wRegOut_5_14[31] , \wRegOut_5_14[30] , \wRegOut_5_14[29] , 
        \wRegOut_5_14[28] , \wRegOut_5_14[27] , \wRegOut_5_14[26] , 
        \wRegOut_5_14[25] , \wRegOut_5_14[24] , \wRegOut_5_14[23] , 
        \wRegOut_5_14[22] , \wRegOut_5_14[21] , \wRegOut_5_14[20] , 
        \wRegOut_5_14[19] , \wRegOut_5_14[18] , \wRegOut_5_14[17] , 
        \wRegOut_5_14[16] , \wRegOut_5_14[15] , \wRegOut_5_14[14] , 
        \wRegOut_5_14[13] , \wRegOut_5_14[12] , \wRegOut_5_14[11] , 
        \wRegOut_5_14[10] , \wRegOut_5_14[9] , \wRegOut_5_14[8] , 
        \wRegOut_5_14[7] , \wRegOut_5_14[6] , \wRegOut_5_14[5] , 
        \wRegOut_5_14[4] , \wRegOut_5_14[3] , \wRegOut_5_14[2] , 
        \wRegOut_5_14[1] , \wRegOut_5_14[0] }), .L_Out({\wRegInTop_5_14[31] , 
        \wRegInTop_5_14[30] , \wRegInTop_5_14[29] , \wRegInTop_5_14[28] , 
        \wRegInTop_5_14[27] , \wRegInTop_5_14[26] , \wRegInTop_5_14[25] , 
        \wRegInTop_5_14[24] , \wRegInTop_5_14[23] , \wRegInTop_5_14[22] , 
        \wRegInTop_5_14[21] , \wRegInTop_5_14[20] , \wRegInTop_5_14[19] , 
        \wRegInTop_5_14[18] , \wRegInTop_5_14[17] , \wRegInTop_5_14[16] , 
        \wRegInTop_5_14[15] , \wRegInTop_5_14[14] , \wRegInTop_5_14[13] , 
        \wRegInTop_5_14[12] , \wRegInTop_5_14[11] , \wRegInTop_5_14[10] , 
        \wRegInTop_5_14[9] , \wRegInTop_5_14[8] , \wRegInTop_5_14[7] , 
        \wRegInTop_5_14[6] , \wRegInTop_5_14[5] , \wRegInTop_5_14[4] , 
        \wRegInTop_5_14[3] , \wRegInTop_5_14[2] , \wRegInTop_5_14[1] , 
        \wRegInTop_5_14[0] }), .R_WR(\wRegEnTop_5_15[0] ), .R_In({
        \wRegOut_5_15[31] , \wRegOut_5_15[30] , \wRegOut_5_15[29] , 
        \wRegOut_5_15[28] , \wRegOut_5_15[27] , \wRegOut_5_15[26] , 
        \wRegOut_5_15[25] , \wRegOut_5_15[24] , \wRegOut_5_15[23] , 
        \wRegOut_5_15[22] , \wRegOut_5_15[21] , \wRegOut_5_15[20] , 
        \wRegOut_5_15[19] , \wRegOut_5_15[18] , \wRegOut_5_15[17] , 
        \wRegOut_5_15[16] , \wRegOut_5_15[15] , \wRegOut_5_15[14] , 
        \wRegOut_5_15[13] , \wRegOut_5_15[12] , \wRegOut_5_15[11] , 
        \wRegOut_5_15[10] , \wRegOut_5_15[9] , \wRegOut_5_15[8] , 
        \wRegOut_5_15[7] , \wRegOut_5_15[6] , \wRegOut_5_15[5] , 
        \wRegOut_5_15[4] , \wRegOut_5_15[3] , \wRegOut_5_15[2] , 
        \wRegOut_5_15[1] , \wRegOut_5_15[0] }), .R_Out({\wRegInTop_5_15[31] , 
        \wRegInTop_5_15[30] , \wRegInTop_5_15[29] , \wRegInTop_5_15[28] , 
        \wRegInTop_5_15[27] , \wRegInTop_5_15[26] , \wRegInTop_5_15[25] , 
        \wRegInTop_5_15[24] , \wRegInTop_5_15[23] , \wRegInTop_5_15[22] , 
        \wRegInTop_5_15[21] , \wRegInTop_5_15[20] , \wRegInTop_5_15[19] , 
        \wRegInTop_5_15[18] , \wRegInTop_5_15[17] , \wRegInTop_5_15[16] , 
        \wRegInTop_5_15[15] , \wRegInTop_5_15[14] , \wRegInTop_5_15[13] , 
        \wRegInTop_5_15[12] , \wRegInTop_5_15[11] , \wRegInTop_5_15[10] , 
        \wRegInTop_5_15[9] , \wRegInTop_5_15[8] , \wRegInTop_5_15[7] , 
        \wRegInTop_5_15[6] , \wRegInTop_5_15[5] , \wRegInTop_5_15[4] , 
        \wRegInTop_5_15[3] , \wRegInTop_5_15[2] , \wRegInTop_5_15[1] , 
        \wRegInTop_5_15[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_109 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink237[31] , \ScanLink237[30] , \ScanLink237[29] , 
        \ScanLink237[28] , \ScanLink237[27] , \ScanLink237[26] , 
        \ScanLink237[25] , \ScanLink237[24] , \ScanLink237[23] , 
        \ScanLink237[22] , \ScanLink237[21] , \ScanLink237[20] , 
        \ScanLink237[19] , \ScanLink237[18] , \ScanLink237[17] , 
        \ScanLink237[16] , \ScanLink237[15] , \ScanLink237[14] , 
        \ScanLink237[13] , \ScanLink237[12] , \ScanLink237[11] , 
        \ScanLink237[10] , \ScanLink237[9] , \ScanLink237[8] , 
        \ScanLink237[7] , \ScanLink237[6] , \ScanLink237[5] , \ScanLink237[4] , 
        \ScanLink237[3] , \ScanLink237[2] , \ScanLink237[1] , \ScanLink237[0] 
        }), .ScanOut({\ScanLink236[31] , \ScanLink236[30] , \ScanLink236[29] , 
        \ScanLink236[28] , \ScanLink236[27] , \ScanLink236[26] , 
        \ScanLink236[25] , \ScanLink236[24] , \ScanLink236[23] , 
        \ScanLink236[22] , \ScanLink236[21] , \ScanLink236[20] , 
        \ScanLink236[19] , \ScanLink236[18] , \ScanLink236[17] , 
        \ScanLink236[16] , \ScanLink236[15] , \ScanLink236[14] , 
        \ScanLink236[13] , \ScanLink236[12] , \ScanLink236[11] , 
        \ScanLink236[10] , \ScanLink236[9] , \ScanLink236[8] , 
        \ScanLink236[7] , \ScanLink236[6] , \ScanLink236[5] , \ScanLink236[4] , 
        \ScanLink236[3] , \ScanLink236[2] , \ScanLink236[1] , \ScanLink236[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_109[31] , 
        \wRegOut_7_109[30] , \wRegOut_7_109[29] , \wRegOut_7_109[28] , 
        \wRegOut_7_109[27] , \wRegOut_7_109[26] , \wRegOut_7_109[25] , 
        \wRegOut_7_109[24] , \wRegOut_7_109[23] , \wRegOut_7_109[22] , 
        \wRegOut_7_109[21] , \wRegOut_7_109[20] , \wRegOut_7_109[19] , 
        \wRegOut_7_109[18] , \wRegOut_7_109[17] , \wRegOut_7_109[16] , 
        \wRegOut_7_109[15] , \wRegOut_7_109[14] , \wRegOut_7_109[13] , 
        \wRegOut_7_109[12] , \wRegOut_7_109[11] , \wRegOut_7_109[10] , 
        \wRegOut_7_109[9] , \wRegOut_7_109[8] , \wRegOut_7_109[7] , 
        \wRegOut_7_109[6] , \wRegOut_7_109[5] , \wRegOut_7_109[4] , 
        \wRegOut_7_109[3] , \wRegOut_7_109[2] , \wRegOut_7_109[1] , 
        \wRegOut_7_109[0] }), .Enable1(\wRegEnTop_7_109[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_109[31] , \wRegInTop_7_109[30] , 
        \wRegInTop_7_109[29] , \wRegInTop_7_109[28] , \wRegInTop_7_109[27] , 
        \wRegInTop_7_109[26] , \wRegInTop_7_109[25] , \wRegInTop_7_109[24] , 
        \wRegInTop_7_109[23] , \wRegInTop_7_109[22] , \wRegInTop_7_109[21] , 
        \wRegInTop_7_109[20] , \wRegInTop_7_109[19] , \wRegInTop_7_109[18] , 
        \wRegInTop_7_109[17] , \wRegInTop_7_109[16] , \wRegInTop_7_109[15] , 
        \wRegInTop_7_109[14] , \wRegInTop_7_109[13] , \wRegInTop_7_109[12] , 
        \wRegInTop_7_109[11] , \wRegInTop_7_109[10] , \wRegInTop_7_109[9] , 
        \wRegInTop_7_109[8] , \wRegInTop_7_109[7] , \wRegInTop_7_109[6] , 
        \wRegInTop_7_109[5] , \wRegInTop_7_109[4] , \wRegInTop_7_109[3] , 
        \wRegInTop_7_109[2] , \wRegInTop_7_109[1] , \wRegInTop_7_109[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_7[0] ), .P_In({\wRegOut_5_7[31] , 
        \wRegOut_5_7[30] , \wRegOut_5_7[29] , \wRegOut_5_7[28] , 
        \wRegOut_5_7[27] , \wRegOut_5_7[26] , \wRegOut_5_7[25] , 
        \wRegOut_5_7[24] , \wRegOut_5_7[23] , \wRegOut_5_7[22] , 
        \wRegOut_5_7[21] , \wRegOut_5_7[20] , \wRegOut_5_7[19] , 
        \wRegOut_5_7[18] , \wRegOut_5_7[17] , \wRegOut_5_7[16] , 
        \wRegOut_5_7[15] , \wRegOut_5_7[14] , \wRegOut_5_7[13] , 
        \wRegOut_5_7[12] , \wRegOut_5_7[11] , \wRegOut_5_7[10] , 
        \wRegOut_5_7[9] , \wRegOut_5_7[8] , \wRegOut_5_7[7] , \wRegOut_5_7[6] , 
        \wRegOut_5_7[5] , \wRegOut_5_7[4] , \wRegOut_5_7[3] , \wRegOut_5_7[2] , 
        \wRegOut_5_7[1] , \wRegOut_5_7[0] }), .P_Out({\wRegInBot_5_7[31] , 
        \wRegInBot_5_7[30] , \wRegInBot_5_7[29] , \wRegInBot_5_7[28] , 
        \wRegInBot_5_7[27] , \wRegInBot_5_7[26] , \wRegInBot_5_7[25] , 
        \wRegInBot_5_7[24] , \wRegInBot_5_7[23] , \wRegInBot_5_7[22] , 
        \wRegInBot_5_7[21] , \wRegInBot_5_7[20] , \wRegInBot_5_7[19] , 
        \wRegInBot_5_7[18] , \wRegInBot_5_7[17] , \wRegInBot_5_7[16] , 
        \wRegInBot_5_7[15] , \wRegInBot_5_7[14] , \wRegInBot_5_7[13] , 
        \wRegInBot_5_7[12] , \wRegInBot_5_7[11] , \wRegInBot_5_7[10] , 
        \wRegInBot_5_7[9] , \wRegInBot_5_7[8] , \wRegInBot_5_7[7] , 
        \wRegInBot_5_7[6] , \wRegInBot_5_7[5] , \wRegInBot_5_7[4] , 
        \wRegInBot_5_7[3] , \wRegInBot_5_7[2] , \wRegInBot_5_7[1] , 
        \wRegInBot_5_7[0] }), .L_WR(\wRegEnTop_6_14[0] ), .L_In({
        \wRegOut_6_14[31] , \wRegOut_6_14[30] , \wRegOut_6_14[29] , 
        \wRegOut_6_14[28] , \wRegOut_6_14[27] , \wRegOut_6_14[26] , 
        \wRegOut_6_14[25] , \wRegOut_6_14[24] , \wRegOut_6_14[23] , 
        \wRegOut_6_14[22] , \wRegOut_6_14[21] , \wRegOut_6_14[20] , 
        \wRegOut_6_14[19] , \wRegOut_6_14[18] , \wRegOut_6_14[17] , 
        \wRegOut_6_14[16] , \wRegOut_6_14[15] , \wRegOut_6_14[14] , 
        \wRegOut_6_14[13] , \wRegOut_6_14[12] , \wRegOut_6_14[11] , 
        \wRegOut_6_14[10] , \wRegOut_6_14[9] , \wRegOut_6_14[8] , 
        \wRegOut_6_14[7] , \wRegOut_6_14[6] , \wRegOut_6_14[5] , 
        \wRegOut_6_14[4] , \wRegOut_6_14[3] , \wRegOut_6_14[2] , 
        \wRegOut_6_14[1] , \wRegOut_6_14[0] }), .L_Out({\wRegInTop_6_14[31] , 
        \wRegInTop_6_14[30] , \wRegInTop_6_14[29] , \wRegInTop_6_14[28] , 
        \wRegInTop_6_14[27] , \wRegInTop_6_14[26] , \wRegInTop_6_14[25] , 
        \wRegInTop_6_14[24] , \wRegInTop_6_14[23] , \wRegInTop_6_14[22] , 
        \wRegInTop_6_14[21] , \wRegInTop_6_14[20] , \wRegInTop_6_14[19] , 
        \wRegInTop_6_14[18] , \wRegInTop_6_14[17] , \wRegInTop_6_14[16] , 
        \wRegInTop_6_14[15] , \wRegInTop_6_14[14] , \wRegInTop_6_14[13] , 
        \wRegInTop_6_14[12] , \wRegInTop_6_14[11] , \wRegInTop_6_14[10] , 
        \wRegInTop_6_14[9] , \wRegInTop_6_14[8] , \wRegInTop_6_14[7] , 
        \wRegInTop_6_14[6] , \wRegInTop_6_14[5] , \wRegInTop_6_14[4] , 
        \wRegInTop_6_14[3] , \wRegInTop_6_14[2] , \wRegInTop_6_14[1] , 
        \wRegInTop_6_14[0] }), .R_WR(\wRegEnTop_6_15[0] ), .R_In({
        \wRegOut_6_15[31] , \wRegOut_6_15[30] , \wRegOut_6_15[29] , 
        \wRegOut_6_15[28] , \wRegOut_6_15[27] , \wRegOut_6_15[26] , 
        \wRegOut_6_15[25] , \wRegOut_6_15[24] , \wRegOut_6_15[23] , 
        \wRegOut_6_15[22] , \wRegOut_6_15[21] , \wRegOut_6_15[20] , 
        \wRegOut_6_15[19] , \wRegOut_6_15[18] , \wRegOut_6_15[17] , 
        \wRegOut_6_15[16] , \wRegOut_6_15[15] , \wRegOut_6_15[14] , 
        \wRegOut_6_15[13] , \wRegOut_6_15[12] , \wRegOut_6_15[11] , 
        \wRegOut_6_15[10] , \wRegOut_6_15[9] , \wRegOut_6_15[8] , 
        \wRegOut_6_15[7] , \wRegOut_6_15[6] , \wRegOut_6_15[5] , 
        \wRegOut_6_15[4] , \wRegOut_6_15[3] , \wRegOut_6_15[2] , 
        \wRegOut_6_15[1] , \wRegOut_6_15[0] }), .R_Out({\wRegInTop_6_15[31] , 
        \wRegInTop_6_15[30] , \wRegInTop_6_15[29] , \wRegInTop_6_15[28] , 
        \wRegInTop_6_15[27] , \wRegInTop_6_15[26] , \wRegInTop_6_15[25] , 
        \wRegInTop_6_15[24] , \wRegInTop_6_15[23] , \wRegInTop_6_15[22] , 
        \wRegInTop_6_15[21] , \wRegInTop_6_15[20] , \wRegInTop_6_15[19] , 
        \wRegInTop_6_15[18] , \wRegInTop_6_15[17] , \wRegInTop_6_15[16] , 
        \wRegInTop_6_15[15] , \wRegInTop_6_15[14] , \wRegInTop_6_15[13] , 
        \wRegInTop_6_15[12] , \wRegInTop_6_15[11] , \wRegInTop_6_15[10] , 
        \wRegInTop_6_15[9] , \wRegInTop_6_15[8] , \wRegInTop_6_15[7] , 
        \wRegInTop_6_15[6] , \wRegInTop_6_15[5] , \wRegInTop_6_15[4] , 
        \wRegInTop_6_15[3] , \wRegInTop_6_15[2] , \wRegInTop_6_15[1] , 
        \wRegInTop_6_15[0] }) );
    BHeap_Node_WIDTH32 BHN_6_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_41[0] ), .P_In({\wRegOut_6_41[31] , 
        \wRegOut_6_41[30] , \wRegOut_6_41[29] , \wRegOut_6_41[28] , 
        \wRegOut_6_41[27] , \wRegOut_6_41[26] , \wRegOut_6_41[25] , 
        \wRegOut_6_41[24] , \wRegOut_6_41[23] , \wRegOut_6_41[22] , 
        \wRegOut_6_41[21] , \wRegOut_6_41[20] , \wRegOut_6_41[19] , 
        \wRegOut_6_41[18] , \wRegOut_6_41[17] , \wRegOut_6_41[16] , 
        \wRegOut_6_41[15] , \wRegOut_6_41[14] , \wRegOut_6_41[13] , 
        \wRegOut_6_41[12] , \wRegOut_6_41[11] , \wRegOut_6_41[10] , 
        \wRegOut_6_41[9] , \wRegOut_6_41[8] , \wRegOut_6_41[7] , 
        \wRegOut_6_41[6] , \wRegOut_6_41[5] , \wRegOut_6_41[4] , 
        \wRegOut_6_41[3] , \wRegOut_6_41[2] , \wRegOut_6_41[1] , 
        \wRegOut_6_41[0] }), .P_Out({\wRegInBot_6_41[31] , 
        \wRegInBot_6_41[30] , \wRegInBot_6_41[29] , \wRegInBot_6_41[28] , 
        \wRegInBot_6_41[27] , \wRegInBot_6_41[26] , \wRegInBot_6_41[25] , 
        \wRegInBot_6_41[24] , \wRegInBot_6_41[23] , \wRegInBot_6_41[22] , 
        \wRegInBot_6_41[21] , \wRegInBot_6_41[20] , \wRegInBot_6_41[19] , 
        \wRegInBot_6_41[18] , \wRegInBot_6_41[17] , \wRegInBot_6_41[16] , 
        \wRegInBot_6_41[15] , \wRegInBot_6_41[14] , \wRegInBot_6_41[13] , 
        \wRegInBot_6_41[12] , \wRegInBot_6_41[11] , \wRegInBot_6_41[10] , 
        \wRegInBot_6_41[9] , \wRegInBot_6_41[8] , \wRegInBot_6_41[7] , 
        \wRegInBot_6_41[6] , \wRegInBot_6_41[5] , \wRegInBot_6_41[4] , 
        \wRegInBot_6_41[3] , \wRegInBot_6_41[2] , \wRegInBot_6_41[1] , 
        \wRegInBot_6_41[0] }), .L_WR(\wRegEnTop_7_82[0] ), .L_In({
        \wRegOut_7_82[31] , \wRegOut_7_82[30] , \wRegOut_7_82[29] , 
        \wRegOut_7_82[28] , \wRegOut_7_82[27] , \wRegOut_7_82[26] , 
        \wRegOut_7_82[25] , \wRegOut_7_82[24] , \wRegOut_7_82[23] , 
        \wRegOut_7_82[22] , \wRegOut_7_82[21] , \wRegOut_7_82[20] , 
        \wRegOut_7_82[19] , \wRegOut_7_82[18] , \wRegOut_7_82[17] , 
        \wRegOut_7_82[16] , \wRegOut_7_82[15] , \wRegOut_7_82[14] , 
        \wRegOut_7_82[13] , \wRegOut_7_82[12] , \wRegOut_7_82[11] , 
        \wRegOut_7_82[10] , \wRegOut_7_82[9] , \wRegOut_7_82[8] , 
        \wRegOut_7_82[7] , \wRegOut_7_82[6] , \wRegOut_7_82[5] , 
        \wRegOut_7_82[4] , \wRegOut_7_82[3] , \wRegOut_7_82[2] , 
        \wRegOut_7_82[1] , \wRegOut_7_82[0] }), .L_Out({\wRegInTop_7_82[31] , 
        \wRegInTop_7_82[30] , \wRegInTop_7_82[29] , \wRegInTop_7_82[28] , 
        \wRegInTop_7_82[27] , \wRegInTop_7_82[26] , \wRegInTop_7_82[25] , 
        \wRegInTop_7_82[24] , \wRegInTop_7_82[23] , \wRegInTop_7_82[22] , 
        \wRegInTop_7_82[21] , \wRegInTop_7_82[20] , \wRegInTop_7_82[19] , 
        \wRegInTop_7_82[18] , \wRegInTop_7_82[17] , \wRegInTop_7_82[16] , 
        \wRegInTop_7_82[15] , \wRegInTop_7_82[14] , \wRegInTop_7_82[13] , 
        \wRegInTop_7_82[12] , \wRegInTop_7_82[11] , \wRegInTop_7_82[10] , 
        \wRegInTop_7_82[9] , \wRegInTop_7_82[8] , \wRegInTop_7_82[7] , 
        \wRegInTop_7_82[6] , \wRegInTop_7_82[5] , \wRegInTop_7_82[4] , 
        \wRegInTop_7_82[3] , \wRegInTop_7_82[2] , \wRegInTop_7_82[1] , 
        \wRegInTop_7_82[0] }), .R_WR(\wRegEnTop_7_83[0] ), .R_In({
        \wRegOut_7_83[31] , \wRegOut_7_83[30] , \wRegOut_7_83[29] , 
        \wRegOut_7_83[28] , \wRegOut_7_83[27] , \wRegOut_7_83[26] , 
        \wRegOut_7_83[25] , \wRegOut_7_83[24] , \wRegOut_7_83[23] , 
        \wRegOut_7_83[22] , \wRegOut_7_83[21] , \wRegOut_7_83[20] , 
        \wRegOut_7_83[19] , \wRegOut_7_83[18] , \wRegOut_7_83[17] , 
        \wRegOut_7_83[16] , \wRegOut_7_83[15] , \wRegOut_7_83[14] , 
        \wRegOut_7_83[13] , \wRegOut_7_83[12] , \wRegOut_7_83[11] , 
        \wRegOut_7_83[10] , \wRegOut_7_83[9] , \wRegOut_7_83[8] , 
        \wRegOut_7_83[7] , \wRegOut_7_83[6] , \wRegOut_7_83[5] , 
        \wRegOut_7_83[4] , \wRegOut_7_83[3] , \wRegOut_7_83[2] , 
        \wRegOut_7_83[1] , \wRegOut_7_83[0] }), .R_Out({\wRegInTop_7_83[31] , 
        \wRegInTop_7_83[30] , \wRegInTop_7_83[29] , \wRegInTop_7_83[28] , 
        \wRegInTop_7_83[27] , \wRegInTop_7_83[26] , \wRegInTop_7_83[25] , 
        \wRegInTop_7_83[24] , \wRegInTop_7_83[23] , \wRegInTop_7_83[22] , 
        \wRegInTop_7_83[21] , \wRegInTop_7_83[20] , \wRegInTop_7_83[19] , 
        \wRegInTop_7_83[18] , \wRegInTop_7_83[17] , \wRegInTop_7_83[16] , 
        \wRegInTop_7_83[15] , \wRegInTop_7_83[14] , \wRegInTop_7_83[13] , 
        \wRegInTop_7_83[12] , \wRegInTop_7_83[11] , \wRegInTop_7_83[10] , 
        \wRegInTop_7_83[9] , \wRegInTop_7_83[8] , \wRegInTop_7_83[7] , 
        \wRegInTop_7_83[6] , \wRegInTop_7_83[5] , \wRegInTop_7_83[4] , 
        \wRegInTop_7_83[3] , \wRegInTop_7_83[2] , \wRegInTop_7_83[1] , 
        \wRegInTop_7_83[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_54 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink182[31] , \ScanLink182[30] , \ScanLink182[29] , 
        \ScanLink182[28] , \ScanLink182[27] , \ScanLink182[26] , 
        \ScanLink182[25] , \ScanLink182[24] , \ScanLink182[23] , 
        \ScanLink182[22] , \ScanLink182[21] , \ScanLink182[20] , 
        \ScanLink182[19] , \ScanLink182[18] , \ScanLink182[17] , 
        \ScanLink182[16] , \ScanLink182[15] , \ScanLink182[14] , 
        \ScanLink182[13] , \ScanLink182[12] , \ScanLink182[11] , 
        \ScanLink182[10] , \ScanLink182[9] , \ScanLink182[8] , 
        \ScanLink182[7] , \ScanLink182[6] , \ScanLink182[5] , \ScanLink182[4] , 
        \ScanLink182[3] , \ScanLink182[2] , \ScanLink182[1] , \ScanLink182[0] 
        }), .ScanOut({\ScanLink181[31] , \ScanLink181[30] , \ScanLink181[29] , 
        \ScanLink181[28] , \ScanLink181[27] , \ScanLink181[26] , 
        \ScanLink181[25] , \ScanLink181[24] , \ScanLink181[23] , 
        \ScanLink181[22] , \ScanLink181[21] , \ScanLink181[20] , 
        \ScanLink181[19] , \ScanLink181[18] , \ScanLink181[17] , 
        \ScanLink181[16] , \ScanLink181[15] , \ScanLink181[14] , 
        \ScanLink181[13] , \ScanLink181[12] , \ScanLink181[11] , 
        \ScanLink181[10] , \ScanLink181[9] , \ScanLink181[8] , 
        \ScanLink181[7] , \ScanLink181[6] , \ScanLink181[5] , \ScanLink181[4] , 
        \ScanLink181[3] , \ScanLink181[2] , \ScanLink181[1] , \ScanLink181[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_54[31] , 
        \wRegOut_7_54[30] , \wRegOut_7_54[29] , \wRegOut_7_54[28] , 
        \wRegOut_7_54[27] , \wRegOut_7_54[26] , \wRegOut_7_54[25] , 
        \wRegOut_7_54[24] , \wRegOut_7_54[23] , \wRegOut_7_54[22] , 
        \wRegOut_7_54[21] , \wRegOut_7_54[20] , \wRegOut_7_54[19] , 
        \wRegOut_7_54[18] , \wRegOut_7_54[17] , \wRegOut_7_54[16] , 
        \wRegOut_7_54[15] , \wRegOut_7_54[14] , \wRegOut_7_54[13] , 
        \wRegOut_7_54[12] , \wRegOut_7_54[11] , \wRegOut_7_54[10] , 
        \wRegOut_7_54[9] , \wRegOut_7_54[8] , \wRegOut_7_54[7] , 
        \wRegOut_7_54[6] , \wRegOut_7_54[5] , \wRegOut_7_54[4] , 
        \wRegOut_7_54[3] , \wRegOut_7_54[2] , \wRegOut_7_54[1] , 
        \wRegOut_7_54[0] }), .Enable1(\wRegEnTop_7_54[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_54[31] , \wRegInTop_7_54[30] , \wRegInTop_7_54[29] , 
        \wRegInTop_7_54[28] , \wRegInTop_7_54[27] , \wRegInTop_7_54[26] , 
        \wRegInTop_7_54[25] , \wRegInTop_7_54[24] , \wRegInTop_7_54[23] , 
        \wRegInTop_7_54[22] , \wRegInTop_7_54[21] , \wRegInTop_7_54[20] , 
        \wRegInTop_7_54[19] , \wRegInTop_7_54[18] , \wRegInTop_7_54[17] , 
        \wRegInTop_7_54[16] , \wRegInTop_7_54[15] , \wRegInTop_7_54[14] , 
        \wRegInTop_7_54[13] , \wRegInTop_7_54[12] , \wRegInTop_7_54[11] , 
        \wRegInTop_7_54[10] , \wRegInTop_7_54[9] , \wRegInTop_7_54[8] , 
        \wRegInTop_7_54[7] , \wRegInTop_7_54[6] , \wRegInTop_7_54[5] , 
        \wRegInTop_7_54[4] , \wRegInTop_7_54[3] , \wRegInTop_7_54[2] , 
        \wRegInTop_7_54[1] , \wRegInTop_7_54[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_73 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink201[31] , \ScanLink201[30] , \ScanLink201[29] , 
        \ScanLink201[28] , \ScanLink201[27] , \ScanLink201[26] , 
        \ScanLink201[25] , \ScanLink201[24] , \ScanLink201[23] , 
        \ScanLink201[22] , \ScanLink201[21] , \ScanLink201[20] , 
        \ScanLink201[19] , \ScanLink201[18] , \ScanLink201[17] , 
        \ScanLink201[16] , \ScanLink201[15] , \ScanLink201[14] , 
        \ScanLink201[13] , \ScanLink201[12] , \ScanLink201[11] , 
        \ScanLink201[10] , \ScanLink201[9] , \ScanLink201[8] , 
        \ScanLink201[7] , \ScanLink201[6] , \ScanLink201[5] , \ScanLink201[4] , 
        \ScanLink201[3] , \ScanLink201[2] , \ScanLink201[1] , \ScanLink201[0] 
        }), .ScanOut({\ScanLink200[31] , \ScanLink200[30] , \ScanLink200[29] , 
        \ScanLink200[28] , \ScanLink200[27] , \ScanLink200[26] , 
        \ScanLink200[25] , \ScanLink200[24] , \ScanLink200[23] , 
        \ScanLink200[22] , \ScanLink200[21] , \ScanLink200[20] , 
        \ScanLink200[19] , \ScanLink200[18] , \ScanLink200[17] , 
        \ScanLink200[16] , \ScanLink200[15] , \ScanLink200[14] , 
        \ScanLink200[13] , \ScanLink200[12] , \ScanLink200[11] , 
        \ScanLink200[10] , \ScanLink200[9] , \ScanLink200[8] , 
        \ScanLink200[7] , \ScanLink200[6] , \ScanLink200[5] , \ScanLink200[4] , 
        \ScanLink200[3] , \ScanLink200[2] , \ScanLink200[1] , \ScanLink200[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_73[31] , 
        \wRegOut_7_73[30] , \wRegOut_7_73[29] , \wRegOut_7_73[28] , 
        \wRegOut_7_73[27] , \wRegOut_7_73[26] , \wRegOut_7_73[25] , 
        \wRegOut_7_73[24] , \wRegOut_7_73[23] , \wRegOut_7_73[22] , 
        \wRegOut_7_73[21] , \wRegOut_7_73[20] , \wRegOut_7_73[19] , 
        \wRegOut_7_73[18] , \wRegOut_7_73[17] , \wRegOut_7_73[16] , 
        \wRegOut_7_73[15] , \wRegOut_7_73[14] , \wRegOut_7_73[13] , 
        \wRegOut_7_73[12] , \wRegOut_7_73[11] , \wRegOut_7_73[10] , 
        \wRegOut_7_73[9] , \wRegOut_7_73[8] , \wRegOut_7_73[7] , 
        \wRegOut_7_73[6] , \wRegOut_7_73[5] , \wRegOut_7_73[4] , 
        \wRegOut_7_73[3] , \wRegOut_7_73[2] , \wRegOut_7_73[1] , 
        \wRegOut_7_73[0] }), .Enable1(\wRegEnTop_7_73[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_73[31] , \wRegInTop_7_73[30] , \wRegInTop_7_73[29] , 
        \wRegInTop_7_73[28] , \wRegInTop_7_73[27] , \wRegInTop_7_73[26] , 
        \wRegInTop_7_73[25] , \wRegInTop_7_73[24] , \wRegInTop_7_73[23] , 
        \wRegInTop_7_73[22] , \wRegInTop_7_73[21] , \wRegInTop_7_73[20] , 
        \wRegInTop_7_73[19] , \wRegInTop_7_73[18] , \wRegInTop_7_73[17] , 
        \wRegInTop_7_73[16] , \wRegInTop_7_73[15] , \wRegInTop_7_73[14] , 
        \wRegInTop_7_73[13] , \wRegInTop_7_73[12] , \wRegInTop_7_73[11] , 
        \wRegInTop_7_73[10] , \wRegInTop_7_73[9] , \wRegInTop_7_73[8] , 
        \wRegInTop_7_73[7] , \wRegInTop_7_73[6] , \wRegInTop_7_73[5] , 
        \wRegInTop_7_73[4] , \wRegInTop_7_73[3] , \wRegInTop_7_73[2] , 
        \wRegInTop_7_73[1] , \wRegInTop_7_73[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink73[31] , \ScanLink73[30] , \ScanLink73[29] , 
        \ScanLink73[28] , \ScanLink73[27] , \ScanLink73[26] , \ScanLink73[25] , 
        \ScanLink73[24] , \ScanLink73[23] , \ScanLink73[22] , \ScanLink73[21] , 
        \ScanLink73[20] , \ScanLink73[19] , \ScanLink73[18] , \ScanLink73[17] , 
        \ScanLink73[16] , \ScanLink73[15] , \ScanLink73[14] , \ScanLink73[13] , 
        \ScanLink73[12] , \ScanLink73[11] , \ScanLink73[10] , \ScanLink73[9] , 
        \ScanLink73[8] , \ScanLink73[7] , \ScanLink73[6] , \ScanLink73[5] , 
        \ScanLink73[4] , \ScanLink73[3] , \ScanLink73[2] , \ScanLink73[1] , 
        \ScanLink73[0] }), .ScanOut({\ScanLink72[31] , \ScanLink72[30] , 
        \ScanLink72[29] , \ScanLink72[28] , \ScanLink72[27] , \ScanLink72[26] , 
        \ScanLink72[25] , \ScanLink72[24] , \ScanLink72[23] , \ScanLink72[22] , 
        \ScanLink72[21] , \ScanLink72[20] , \ScanLink72[19] , \ScanLink72[18] , 
        \ScanLink72[17] , \ScanLink72[16] , \ScanLink72[15] , \ScanLink72[14] , 
        \ScanLink72[13] , \ScanLink72[12] , \ScanLink72[11] , \ScanLink72[10] , 
        \ScanLink72[9] , \ScanLink72[8] , \ScanLink72[7] , \ScanLink72[6] , 
        \ScanLink72[5] , \ScanLink72[4] , \ScanLink72[3] , \ScanLink72[2] , 
        \ScanLink72[1] , \ScanLink72[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_9[31] , \wRegOut_6_9[30] , \wRegOut_6_9[29] , 
        \wRegOut_6_9[28] , \wRegOut_6_9[27] , \wRegOut_6_9[26] , 
        \wRegOut_6_9[25] , \wRegOut_6_9[24] , \wRegOut_6_9[23] , 
        \wRegOut_6_9[22] , \wRegOut_6_9[21] , \wRegOut_6_9[20] , 
        \wRegOut_6_9[19] , \wRegOut_6_9[18] , \wRegOut_6_9[17] , 
        \wRegOut_6_9[16] , \wRegOut_6_9[15] , \wRegOut_6_9[14] , 
        \wRegOut_6_9[13] , \wRegOut_6_9[12] , \wRegOut_6_9[11] , 
        \wRegOut_6_9[10] , \wRegOut_6_9[9] , \wRegOut_6_9[8] , 
        \wRegOut_6_9[7] , \wRegOut_6_9[6] , \wRegOut_6_9[5] , \wRegOut_6_9[4] , 
        \wRegOut_6_9[3] , \wRegOut_6_9[2] , \wRegOut_6_9[1] , \wRegOut_6_9[0] 
        }), .Enable1(\wRegEnTop_6_9[0] ), .Enable2(\wRegEnBot_6_9[0] ), .In1({
        \wRegInTop_6_9[31] , \wRegInTop_6_9[30] , \wRegInTop_6_9[29] , 
        \wRegInTop_6_9[28] , \wRegInTop_6_9[27] , \wRegInTop_6_9[26] , 
        \wRegInTop_6_9[25] , \wRegInTop_6_9[24] , \wRegInTop_6_9[23] , 
        \wRegInTop_6_9[22] , \wRegInTop_6_9[21] , \wRegInTop_6_9[20] , 
        \wRegInTop_6_9[19] , \wRegInTop_6_9[18] , \wRegInTop_6_9[17] , 
        \wRegInTop_6_9[16] , \wRegInTop_6_9[15] , \wRegInTop_6_9[14] , 
        \wRegInTop_6_9[13] , \wRegInTop_6_9[12] , \wRegInTop_6_9[11] , 
        \wRegInTop_6_9[10] , \wRegInTop_6_9[9] , \wRegInTop_6_9[8] , 
        \wRegInTop_6_9[7] , \wRegInTop_6_9[6] , \wRegInTop_6_9[5] , 
        \wRegInTop_6_9[4] , \wRegInTop_6_9[3] , \wRegInTop_6_9[2] , 
        \wRegInTop_6_9[1] , \wRegInTop_6_9[0] }), .In2({\wRegInBot_6_9[31] , 
        \wRegInBot_6_9[30] , \wRegInBot_6_9[29] , \wRegInBot_6_9[28] , 
        \wRegInBot_6_9[27] , \wRegInBot_6_9[26] , \wRegInBot_6_9[25] , 
        \wRegInBot_6_9[24] , \wRegInBot_6_9[23] , \wRegInBot_6_9[22] , 
        \wRegInBot_6_9[21] , \wRegInBot_6_9[20] , \wRegInBot_6_9[19] , 
        \wRegInBot_6_9[18] , \wRegInBot_6_9[17] , \wRegInBot_6_9[16] , 
        \wRegInBot_6_9[15] , \wRegInBot_6_9[14] , \wRegInBot_6_9[13] , 
        \wRegInBot_6_9[12] , \wRegInBot_6_9[11] , \wRegInBot_6_9[10] , 
        \wRegInBot_6_9[9] , \wRegInBot_6_9[8] , \wRegInBot_6_9[7] , 
        \wRegInBot_6_9[6] , \wRegInBot_6_9[5] , \wRegInBot_6_9[4] , 
        \wRegInBot_6_9[3] , \wRegInBot_6_9[2] , \wRegInBot_6_9[1] , 
        \wRegInBot_6_9[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink34[31] , \ScanLink34[30] , \ScanLink34[29] , 
        \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , \ScanLink34[25] , 
        \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , \ScanLink34[21] , 
        \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , \ScanLink34[17] , 
        \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , \ScanLink34[13] , 
        \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , \ScanLink34[9] , 
        \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , \ScanLink34[5] , 
        \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , \ScanLink34[1] , 
        \ScanLink34[0] }), .ScanOut({\ScanLink33[31] , \ScanLink33[30] , 
        \ScanLink33[29] , \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , 
        \ScanLink33[25] , \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , 
        \ScanLink33[21] , \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , 
        \ScanLink33[17] , \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , 
        \ScanLink33[13] , \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , 
        \ScanLink33[9] , \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , 
        \ScanLink33[5] , \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , 
        \ScanLink33[1] , \ScanLink33[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_2[31] , \wRegOut_5_2[30] , \wRegOut_5_2[29] , 
        \wRegOut_5_2[28] , \wRegOut_5_2[27] , \wRegOut_5_2[26] , 
        \wRegOut_5_2[25] , \wRegOut_5_2[24] , \wRegOut_5_2[23] , 
        \wRegOut_5_2[22] , \wRegOut_5_2[21] , \wRegOut_5_2[20] , 
        \wRegOut_5_2[19] , \wRegOut_5_2[18] , \wRegOut_5_2[17] , 
        \wRegOut_5_2[16] , \wRegOut_5_2[15] , \wRegOut_5_2[14] , 
        \wRegOut_5_2[13] , \wRegOut_5_2[12] , \wRegOut_5_2[11] , 
        \wRegOut_5_2[10] , \wRegOut_5_2[9] , \wRegOut_5_2[8] , 
        \wRegOut_5_2[7] , \wRegOut_5_2[6] , \wRegOut_5_2[5] , \wRegOut_5_2[4] , 
        \wRegOut_5_2[3] , \wRegOut_5_2[2] , \wRegOut_5_2[1] , \wRegOut_5_2[0] 
        }), .Enable1(\wRegEnTop_5_2[0] ), .Enable2(\wRegEnBot_5_2[0] ), .In1({
        \wRegInTop_5_2[31] , \wRegInTop_5_2[30] , \wRegInTop_5_2[29] , 
        \wRegInTop_5_2[28] , \wRegInTop_5_2[27] , \wRegInTop_5_2[26] , 
        \wRegInTop_5_2[25] , \wRegInTop_5_2[24] , \wRegInTop_5_2[23] , 
        \wRegInTop_5_2[22] , \wRegInTop_5_2[21] , \wRegInTop_5_2[20] , 
        \wRegInTop_5_2[19] , \wRegInTop_5_2[18] , \wRegInTop_5_2[17] , 
        \wRegInTop_5_2[16] , \wRegInTop_5_2[15] , \wRegInTop_5_2[14] , 
        \wRegInTop_5_2[13] , \wRegInTop_5_2[12] , \wRegInTop_5_2[11] , 
        \wRegInTop_5_2[10] , \wRegInTop_5_2[9] , \wRegInTop_5_2[8] , 
        \wRegInTop_5_2[7] , \wRegInTop_5_2[6] , \wRegInTop_5_2[5] , 
        \wRegInTop_5_2[4] , \wRegInTop_5_2[3] , \wRegInTop_5_2[2] , 
        \wRegInTop_5_2[1] , \wRegInTop_5_2[0] }), .In2({\wRegInBot_5_2[31] , 
        \wRegInBot_5_2[30] , \wRegInBot_5_2[29] , \wRegInBot_5_2[28] , 
        \wRegInBot_5_2[27] , \wRegInBot_5_2[26] , \wRegInBot_5_2[25] , 
        \wRegInBot_5_2[24] , \wRegInBot_5_2[23] , \wRegInBot_5_2[22] , 
        \wRegInBot_5_2[21] , \wRegInBot_5_2[20] , \wRegInBot_5_2[19] , 
        \wRegInBot_5_2[18] , \wRegInBot_5_2[17] , \wRegInBot_5_2[16] , 
        \wRegInBot_5_2[15] , \wRegInBot_5_2[14] , \wRegInBot_5_2[13] , 
        \wRegInBot_5_2[12] , \wRegInBot_5_2[11] , \wRegInBot_5_2[10] , 
        \wRegInBot_5_2[9] , \wRegInBot_5_2[8] , \wRegInBot_5_2[7] , 
        \wRegInBot_5_2[6] , \wRegInBot_5_2[5] , \wRegInBot_5_2[4] , 
        \wRegInBot_5_2[3] , \wRegInBot_5_2[2] , \wRegInBot_5_2[1] , 
        \wRegInBot_5_2[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_17 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink49[31] , \ScanLink49[30] , \ScanLink49[29] , 
        \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , \ScanLink49[25] , 
        \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , \ScanLink49[21] , 
        \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , \ScanLink49[17] , 
        \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , \ScanLink49[13] , 
        \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , \ScanLink49[9] , 
        \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , \ScanLink49[5] , 
        \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , \ScanLink49[1] , 
        \ScanLink49[0] }), .ScanOut({\ScanLink48[31] , \ScanLink48[30] , 
        \ScanLink48[29] , \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , 
        \ScanLink48[25] , \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , 
        \ScanLink48[21] , \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , 
        \ScanLink48[17] , \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , 
        \ScanLink48[13] , \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , 
        \ScanLink48[9] , \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , 
        \ScanLink48[5] , \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , 
        \ScanLink48[1] , \ScanLink48[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_17[31] , \wRegOut_5_17[30] , 
        \wRegOut_5_17[29] , \wRegOut_5_17[28] , \wRegOut_5_17[27] , 
        \wRegOut_5_17[26] , \wRegOut_5_17[25] , \wRegOut_5_17[24] , 
        \wRegOut_5_17[23] , \wRegOut_5_17[22] , \wRegOut_5_17[21] , 
        \wRegOut_5_17[20] , \wRegOut_5_17[19] , \wRegOut_5_17[18] , 
        \wRegOut_5_17[17] , \wRegOut_5_17[16] , \wRegOut_5_17[15] , 
        \wRegOut_5_17[14] , \wRegOut_5_17[13] , \wRegOut_5_17[12] , 
        \wRegOut_5_17[11] , \wRegOut_5_17[10] , \wRegOut_5_17[9] , 
        \wRegOut_5_17[8] , \wRegOut_5_17[7] , \wRegOut_5_17[6] , 
        \wRegOut_5_17[5] , \wRegOut_5_17[4] , \wRegOut_5_17[3] , 
        \wRegOut_5_17[2] , \wRegOut_5_17[1] , \wRegOut_5_17[0] }), .Enable1(
        \wRegEnTop_5_17[0] ), .Enable2(\wRegEnBot_5_17[0] ), .In1({
        \wRegInTop_5_17[31] , \wRegInTop_5_17[30] , \wRegInTop_5_17[29] , 
        \wRegInTop_5_17[28] , \wRegInTop_5_17[27] , \wRegInTop_5_17[26] , 
        \wRegInTop_5_17[25] , \wRegInTop_5_17[24] , \wRegInTop_5_17[23] , 
        \wRegInTop_5_17[22] , \wRegInTop_5_17[21] , \wRegInTop_5_17[20] , 
        \wRegInTop_5_17[19] , \wRegInTop_5_17[18] , \wRegInTop_5_17[17] , 
        \wRegInTop_5_17[16] , \wRegInTop_5_17[15] , \wRegInTop_5_17[14] , 
        \wRegInTop_5_17[13] , \wRegInTop_5_17[12] , \wRegInTop_5_17[11] , 
        \wRegInTop_5_17[10] , \wRegInTop_5_17[9] , \wRegInTop_5_17[8] , 
        \wRegInTop_5_17[7] , \wRegInTop_5_17[6] , \wRegInTop_5_17[5] , 
        \wRegInTop_5_17[4] , \wRegInTop_5_17[3] , \wRegInTop_5_17[2] , 
        \wRegInTop_5_17[1] , \wRegInTop_5_17[0] }), .In2({\wRegInBot_5_17[31] , 
        \wRegInBot_5_17[30] , \wRegInBot_5_17[29] , \wRegInBot_5_17[28] , 
        \wRegInBot_5_17[27] , \wRegInBot_5_17[26] , \wRegInBot_5_17[25] , 
        \wRegInBot_5_17[24] , \wRegInBot_5_17[23] , \wRegInBot_5_17[22] , 
        \wRegInBot_5_17[21] , \wRegInBot_5_17[20] , \wRegInBot_5_17[19] , 
        \wRegInBot_5_17[18] , \wRegInBot_5_17[17] , \wRegInBot_5_17[16] , 
        \wRegInBot_5_17[15] , \wRegInBot_5_17[14] , \wRegInBot_5_17[13] , 
        \wRegInBot_5_17[12] , \wRegInBot_5_17[11] , \wRegInBot_5_17[10] , 
        \wRegInBot_5_17[9] , \wRegInBot_5_17[8] , \wRegInBot_5_17[7] , 
        \wRegInBot_5_17[6] , \wRegInBot_5_17[5] , \wRegInBot_5_17[4] , 
        \wRegInBot_5_17[3] , \wRegInBot_5_17[2] , \wRegInBot_5_17[1] , 
        \wRegInBot_5_17[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_30 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink62[31] , \ScanLink62[30] , \ScanLink62[29] , 
        \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , \ScanLink62[25] , 
        \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , \ScanLink62[21] , 
        \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , \ScanLink62[17] , 
        \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , \ScanLink62[13] , 
        \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , \ScanLink62[9] , 
        \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , \ScanLink62[5] , 
        \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , \ScanLink62[1] , 
        \ScanLink62[0] }), .ScanOut({\ScanLink61[31] , \ScanLink61[30] , 
        \ScanLink61[29] , \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , 
        \ScanLink61[25] , \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , 
        \ScanLink61[21] , \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , 
        \ScanLink61[17] , \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , 
        \ScanLink61[13] , \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , 
        \ScanLink61[9] , \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , 
        \ScanLink61[5] , \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , 
        \ScanLink61[1] , \ScanLink61[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_30[31] , \wRegOut_5_30[30] , 
        \wRegOut_5_30[29] , \wRegOut_5_30[28] , \wRegOut_5_30[27] , 
        \wRegOut_5_30[26] , \wRegOut_5_30[25] , \wRegOut_5_30[24] , 
        \wRegOut_5_30[23] , \wRegOut_5_30[22] , \wRegOut_5_30[21] , 
        \wRegOut_5_30[20] , \wRegOut_5_30[19] , \wRegOut_5_30[18] , 
        \wRegOut_5_30[17] , \wRegOut_5_30[16] , \wRegOut_5_30[15] , 
        \wRegOut_5_30[14] , \wRegOut_5_30[13] , \wRegOut_5_30[12] , 
        \wRegOut_5_30[11] , \wRegOut_5_30[10] , \wRegOut_5_30[9] , 
        \wRegOut_5_30[8] , \wRegOut_5_30[7] , \wRegOut_5_30[6] , 
        \wRegOut_5_30[5] , \wRegOut_5_30[4] , \wRegOut_5_30[3] , 
        \wRegOut_5_30[2] , \wRegOut_5_30[1] , \wRegOut_5_30[0] }), .Enable1(
        \wRegEnTop_5_30[0] ), .Enable2(\wRegEnBot_5_30[0] ), .In1({
        \wRegInTop_5_30[31] , \wRegInTop_5_30[30] , \wRegInTop_5_30[29] , 
        \wRegInTop_5_30[28] , \wRegInTop_5_30[27] , \wRegInTop_5_30[26] , 
        \wRegInTop_5_30[25] , \wRegInTop_5_30[24] , \wRegInTop_5_30[23] , 
        \wRegInTop_5_30[22] , \wRegInTop_5_30[21] , \wRegInTop_5_30[20] , 
        \wRegInTop_5_30[19] , \wRegInTop_5_30[18] , \wRegInTop_5_30[17] , 
        \wRegInTop_5_30[16] , \wRegInTop_5_30[15] , \wRegInTop_5_30[14] , 
        \wRegInTop_5_30[13] , \wRegInTop_5_30[12] , \wRegInTop_5_30[11] , 
        \wRegInTop_5_30[10] , \wRegInTop_5_30[9] , \wRegInTop_5_30[8] , 
        \wRegInTop_5_30[7] , \wRegInTop_5_30[6] , \wRegInTop_5_30[5] , 
        \wRegInTop_5_30[4] , \wRegInTop_5_30[3] , \wRegInTop_5_30[2] , 
        \wRegInTop_5_30[1] , \wRegInTop_5_30[0] }), .In2({\wRegInBot_5_30[31] , 
        \wRegInBot_5_30[30] , \wRegInBot_5_30[29] , \wRegInBot_5_30[28] , 
        \wRegInBot_5_30[27] , \wRegInBot_5_30[26] , \wRegInBot_5_30[25] , 
        \wRegInBot_5_30[24] , \wRegInBot_5_30[23] , \wRegInBot_5_30[22] , 
        \wRegInBot_5_30[21] , \wRegInBot_5_30[20] , \wRegInBot_5_30[19] , 
        \wRegInBot_5_30[18] , \wRegInBot_5_30[17] , \wRegInBot_5_30[16] , 
        \wRegInBot_5_30[15] , \wRegInBot_5_30[14] , \wRegInBot_5_30[13] , 
        \wRegInBot_5_30[12] , \wRegInBot_5_30[11] , \wRegInBot_5_30[10] , 
        \wRegInBot_5_30[9] , \wRegInBot_5_30[8] , \wRegInBot_5_30[7] , 
        \wRegInBot_5_30[6] , \wRegInBot_5_30[5] , \wRegInBot_5_30[4] , 
        \wRegInBot_5_30[3] , \wRegInBot_5_30[2] , \wRegInBot_5_30[1] , 
        \wRegInBot_5_30[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_74 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink202[31] , \ScanLink202[30] , \ScanLink202[29] , 
        \ScanLink202[28] , \ScanLink202[27] , \ScanLink202[26] , 
        \ScanLink202[25] , \ScanLink202[24] , \ScanLink202[23] , 
        \ScanLink202[22] , \ScanLink202[21] , \ScanLink202[20] , 
        \ScanLink202[19] , \ScanLink202[18] , \ScanLink202[17] , 
        \ScanLink202[16] , \ScanLink202[15] , \ScanLink202[14] , 
        \ScanLink202[13] , \ScanLink202[12] , \ScanLink202[11] , 
        \ScanLink202[10] , \ScanLink202[9] , \ScanLink202[8] , 
        \ScanLink202[7] , \ScanLink202[6] , \ScanLink202[5] , \ScanLink202[4] , 
        \ScanLink202[3] , \ScanLink202[2] , \ScanLink202[1] , \ScanLink202[0] 
        }), .ScanOut({\ScanLink201[31] , \ScanLink201[30] , \ScanLink201[29] , 
        \ScanLink201[28] , \ScanLink201[27] , \ScanLink201[26] , 
        \ScanLink201[25] , \ScanLink201[24] , \ScanLink201[23] , 
        \ScanLink201[22] , \ScanLink201[21] , \ScanLink201[20] , 
        \ScanLink201[19] , \ScanLink201[18] , \ScanLink201[17] , 
        \ScanLink201[16] , \ScanLink201[15] , \ScanLink201[14] , 
        \ScanLink201[13] , \ScanLink201[12] , \ScanLink201[11] , 
        \ScanLink201[10] , \ScanLink201[9] , \ScanLink201[8] , 
        \ScanLink201[7] , \ScanLink201[6] , \ScanLink201[5] , \ScanLink201[4] , 
        \ScanLink201[3] , \ScanLink201[2] , \ScanLink201[1] , \ScanLink201[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_74[31] , 
        \wRegOut_7_74[30] , \wRegOut_7_74[29] , \wRegOut_7_74[28] , 
        \wRegOut_7_74[27] , \wRegOut_7_74[26] , \wRegOut_7_74[25] , 
        \wRegOut_7_74[24] , \wRegOut_7_74[23] , \wRegOut_7_74[22] , 
        \wRegOut_7_74[21] , \wRegOut_7_74[20] , \wRegOut_7_74[19] , 
        \wRegOut_7_74[18] , \wRegOut_7_74[17] , \wRegOut_7_74[16] , 
        \wRegOut_7_74[15] , \wRegOut_7_74[14] , \wRegOut_7_74[13] , 
        \wRegOut_7_74[12] , \wRegOut_7_74[11] , \wRegOut_7_74[10] , 
        \wRegOut_7_74[9] , \wRegOut_7_74[8] , \wRegOut_7_74[7] , 
        \wRegOut_7_74[6] , \wRegOut_7_74[5] , \wRegOut_7_74[4] , 
        \wRegOut_7_74[3] , \wRegOut_7_74[2] , \wRegOut_7_74[1] , 
        \wRegOut_7_74[0] }), .Enable1(\wRegEnTop_7_74[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_74[31] , \wRegInTop_7_74[30] , \wRegInTop_7_74[29] , 
        \wRegInTop_7_74[28] , \wRegInTop_7_74[27] , \wRegInTop_7_74[26] , 
        \wRegInTop_7_74[25] , \wRegInTop_7_74[24] , \wRegInTop_7_74[23] , 
        \wRegInTop_7_74[22] , \wRegInTop_7_74[21] , \wRegInTop_7_74[20] , 
        \wRegInTop_7_74[19] , \wRegInTop_7_74[18] , \wRegInTop_7_74[17] , 
        \wRegInTop_7_74[16] , \wRegInTop_7_74[15] , \wRegInTop_7_74[14] , 
        \wRegInTop_7_74[13] , \wRegInTop_7_74[12] , \wRegInTop_7_74[11] , 
        \wRegInTop_7_74[10] , \wRegInTop_7_74[9] , \wRegInTop_7_74[8] , 
        \wRegInTop_7_74[7] , \wRegInTop_7_74[6] , \wRegInTop_7_74[5] , 
        \wRegInTop_7_74[4] , \wRegInTop_7_74[3] , \wRegInTop_7_74[2] , 
        \wRegInTop_7_74[1] , \wRegInTop_7_74[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_28[0] ), .P_In({\wRegOut_6_28[31] , 
        \wRegOut_6_28[30] , \wRegOut_6_28[29] , \wRegOut_6_28[28] , 
        \wRegOut_6_28[27] , \wRegOut_6_28[26] , \wRegOut_6_28[25] , 
        \wRegOut_6_28[24] , \wRegOut_6_28[23] , \wRegOut_6_28[22] , 
        \wRegOut_6_28[21] , \wRegOut_6_28[20] , \wRegOut_6_28[19] , 
        \wRegOut_6_28[18] , \wRegOut_6_28[17] , \wRegOut_6_28[16] , 
        \wRegOut_6_28[15] , \wRegOut_6_28[14] , \wRegOut_6_28[13] , 
        \wRegOut_6_28[12] , \wRegOut_6_28[11] , \wRegOut_6_28[10] , 
        \wRegOut_6_28[9] , \wRegOut_6_28[8] , \wRegOut_6_28[7] , 
        \wRegOut_6_28[6] , \wRegOut_6_28[5] , \wRegOut_6_28[4] , 
        \wRegOut_6_28[3] , \wRegOut_6_28[2] , \wRegOut_6_28[1] , 
        \wRegOut_6_28[0] }), .P_Out({\wRegInBot_6_28[31] , 
        \wRegInBot_6_28[30] , \wRegInBot_6_28[29] , \wRegInBot_6_28[28] , 
        \wRegInBot_6_28[27] , \wRegInBot_6_28[26] , \wRegInBot_6_28[25] , 
        \wRegInBot_6_28[24] , \wRegInBot_6_28[23] , \wRegInBot_6_28[22] , 
        \wRegInBot_6_28[21] , \wRegInBot_6_28[20] , \wRegInBot_6_28[19] , 
        \wRegInBot_6_28[18] , \wRegInBot_6_28[17] , \wRegInBot_6_28[16] , 
        \wRegInBot_6_28[15] , \wRegInBot_6_28[14] , \wRegInBot_6_28[13] , 
        \wRegInBot_6_28[12] , \wRegInBot_6_28[11] , \wRegInBot_6_28[10] , 
        \wRegInBot_6_28[9] , \wRegInBot_6_28[8] , \wRegInBot_6_28[7] , 
        \wRegInBot_6_28[6] , \wRegInBot_6_28[5] , \wRegInBot_6_28[4] , 
        \wRegInBot_6_28[3] , \wRegInBot_6_28[2] , \wRegInBot_6_28[1] , 
        \wRegInBot_6_28[0] }), .L_WR(\wRegEnTop_7_56[0] ), .L_In({
        \wRegOut_7_56[31] , \wRegOut_7_56[30] , \wRegOut_7_56[29] , 
        \wRegOut_7_56[28] , \wRegOut_7_56[27] , \wRegOut_7_56[26] , 
        \wRegOut_7_56[25] , \wRegOut_7_56[24] , \wRegOut_7_56[23] , 
        \wRegOut_7_56[22] , \wRegOut_7_56[21] , \wRegOut_7_56[20] , 
        \wRegOut_7_56[19] , \wRegOut_7_56[18] , \wRegOut_7_56[17] , 
        \wRegOut_7_56[16] , \wRegOut_7_56[15] , \wRegOut_7_56[14] , 
        \wRegOut_7_56[13] , \wRegOut_7_56[12] , \wRegOut_7_56[11] , 
        \wRegOut_7_56[10] , \wRegOut_7_56[9] , \wRegOut_7_56[8] , 
        \wRegOut_7_56[7] , \wRegOut_7_56[6] , \wRegOut_7_56[5] , 
        \wRegOut_7_56[4] , \wRegOut_7_56[3] , \wRegOut_7_56[2] , 
        \wRegOut_7_56[1] , \wRegOut_7_56[0] }), .L_Out({\wRegInTop_7_56[31] , 
        \wRegInTop_7_56[30] , \wRegInTop_7_56[29] , \wRegInTop_7_56[28] , 
        \wRegInTop_7_56[27] , \wRegInTop_7_56[26] , \wRegInTop_7_56[25] , 
        \wRegInTop_7_56[24] , \wRegInTop_7_56[23] , \wRegInTop_7_56[22] , 
        \wRegInTop_7_56[21] , \wRegInTop_7_56[20] , \wRegInTop_7_56[19] , 
        \wRegInTop_7_56[18] , \wRegInTop_7_56[17] , \wRegInTop_7_56[16] , 
        \wRegInTop_7_56[15] , \wRegInTop_7_56[14] , \wRegInTop_7_56[13] , 
        \wRegInTop_7_56[12] , \wRegInTop_7_56[11] , \wRegInTop_7_56[10] , 
        \wRegInTop_7_56[9] , \wRegInTop_7_56[8] , \wRegInTop_7_56[7] , 
        \wRegInTop_7_56[6] , \wRegInTop_7_56[5] , \wRegInTop_7_56[4] , 
        \wRegInTop_7_56[3] , \wRegInTop_7_56[2] , \wRegInTop_7_56[1] , 
        \wRegInTop_7_56[0] }), .R_WR(\wRegEnTop_7_57[0] ), .R_In({
        \wRegOut_7_57[31] , \wRegOut_7_57[30] , \wRegOut_7_57[29] , 
        \wRegOut_7_57[28] , \wRegOut_7_57[27] , \wRegOut_7_57[26] , 
        \wRegOut_7_57[25] , \wRegOut_7_57[24] , \wRegOut_7_57[23] , 
        \wRegOut_7_57[22] , \wRegOut_7_57[21] , \wRegOut_7_57[20] , 
        \wRegOut_7_57[19] , \wRegOut_7_57[18] , \wRegOut_7_57[17] , 
        \wRegOut_7_57[16] , \wRegOut_7_57[15] , \wRegOut_7_57[14] , 
        \wRegOut_7_57[13] , \wRegOut_7_57[12] , \wRegOut_7_57[11] , 
        \wRegOut_7_57[10] , \wRegOut_7_57[9] , \wRegOut_7_57[8] , 
        \wRegOut_7_57[7] , \wRegOut_7_57[6] , \wRegOut_7_57[5] , 
        \wRegOut_7_57[4] , \wRegOut_7_57[3] , \wRegOut_7_57[2] , 
        \wRegOut_7_57[1] , \wRegOut_7_57[0] }), .R_Out({\wRegInTop_7_57[31] , 
        \wRegInTop_7_57[30] , \wRegInTop_7_57[29] , \wRegInTop_7_57[28] , 
        \wRegInTop_7_57[27] , \wRegInTop_7_57[26] , \wRegInTop_7_57[25] , 
        \wRegInTop_7_57[24] , \wRegInTop_7_57[23] , \wRegInTop_7_57[22] , 
        \wRegInTop_7_57[21] , \wRegInTop_7_57[20] , \wRegInTop_7_57[19] , 
        \wRegInTop_7_57[18] , \wRegInTop_7_57[17] , \wRegInTop_7_57[16] , 
        \wRegInTop_7_57[15] , \wRegInTop_7_57[14] , \wRegInTop_7_57[13] , 
        \wRegInTop_7_57[12] , \wRegInTop_7_57[11] , \wRegInTop_7_57[10] , 
        \wRegInTop_7_57[9] , \wRegInTop_7_57[8] , \wRegInTop_7_57[7] , 
        \wRegInTop_7_57[6] , \wRegInTop_7_57[5] , \wRegInTop_7_57[4] , 
        \wRegInTop_7_57[3] , \wRegInTop_7_57[2] , \wRegInTop_7_57[1] , 
        \wRegInTop_7_57[0] }) );
    BHeap_Node_WIDTH32 BHN_5_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_18[0] ), .P_In({\wRegOut_5_18[31] , 
        \wRegOut_5_18[30] , \wRegOut_5_18[29] , \wRegOut_5_18[28] , 
        \wRegOut_5_18[27] , \wRegOut_5_18[26] , \wRegOut_5_18[25] , 
        \wRegOut_5_18[24] , \wRegOut_5_18[23] , \wRegOut_5_18[22] , 
        \wRegOut_5_18[21] , \wRegOut_5_18[20] , \wRegOut_5_18[19] , 
        \wRegOut_5_18[18] , \wRegOut_5_18[17] , \wRegOut_5_18[16] , 
        \wRegOut_5_18[15] , \wRegOut_5_18[14] , \wRegOut_5_18[13] , 
        \wRegOut_5_18[12] , \wRegOut_5_18[11] , \wRegOut_5_18[10] , 
        \wRegOut_5_18[9] , \wRegOut_5_18[8] , \wRegOut_5_18[7] , 
        \wRegOut_5_18[6] , \wRegOut_5_18[5] , \wRegOut_5_18[4] , 
        \wRegOut_5_18[3] , \wRegOut_5_18[2] , \wRegOut_5_18[1] , 
        \wRegOut_5_18[0] }), .P_Out({\wRegInBot_5_18[31] , 
        \wRegInBot_5_18[30] , \wRegInBot_5_18[29] , \wRegInBot_5_18[28] , 
        \wRegInBot_5_18[27] , \wRegInBot_5_18[26] , \wRegInBot_5_18[25] , 
        \wRegInBot_5_18[24] , \wRegInBot_5_18[23] , \wRegInBot_5_18[22] , 
        \wRegInBot_5_18[21] , \wRegInBot_5_18[20] , \wRegInBot_5_18[19] , 
        \wRegInBot_5_18[18] , \wRegInBot_5_18[17] , \wRegInBot_5_18[16] , 
        \wRegInBot_5_18[15] , \wRegInBot_5_18[14] , \wRegInBot_5_18[13] , 
        \wRegInBot_5_18[12] , \wRegInBot_5_18[11] , \wRegInBot_5_18[10] , 
        \wRegInBot_5_18[9] , \wRegInBot_5_18[8] , \wRegInBot_5_18[7] , 
        \wRegInBot_5_18[6] , \wRegInBot_5_18[5] , \wRegInBot_5_18[4] , 
        \wRegInBot_5_18[3] , \wRegInBot_5_18[2] , \wRegInBot_5_18[1] , 
        \wRegInBot_5_18[0] }), .L_WR(\wRegEnTop_6_36[0] ), .L_In({
        \wRegOut_6_36[31] , \wRegOut_6_36[30] , \wRegOut_6_36[29] , 
        \wRegOut_6_36[28] , \wRegOut_6_36[27] , \wRegOut_6_36[26] , 
        \wRegOut_6_36[25] , \wRegOut_6_36[24] , \wRegOut_6_36[23] , 
        \wRegOut_6_36[22] , \wRegOut_6_36[21] , \wRegOut_6_36[20] , 
        \wRegOut_6_36[19] , \wRegOut_6_36[18] , \wRegOut_6_36[17] , 
        \wRegOut_6_36[16] , \wRegOut_6_36[15] , \wRegOut_6_36[14] , 
        \wRegOut_6_36[13] , \wRegOut_6_36[12] , \wRegOut_6_36[11] , 
        \wRegOut_6_36[10] , \wRegOut_6_36[9] , \wRegOut_6_36[8] , 
        \wRegOut_6_36[7] , \wRegOut_6_36[6] , \wRegOut_6_36[5] , 
        \wRegOut_6_36[4] , \wRegOut_6_36[3] , \wRegOut_6_36[2] , 
        \wRegOut_6_36[1] , \wRegOut_6_36[0] }), .L_Out({\wRegInTop_6_36[31] , 
        \wRegInTop_6_36[30] , \wRegInTop_6_36[29] , \wRegInTop_6_36[28] , 
        \wRegInTop_6_36[27] , \wRegInTop_6_36[26] , \wRegInTop_6_36[25] , 
        \wRegInTop_6_36[24] , \wRegInTop_6_36[23] , \wRegInTop_6_36[22] , 
        \wRegInTop_6_36[21] , \wRegInTop_6_36[20] , \wRegInTop_6_36[19] , 
        \wRegInTop_6_36[18] , \wRegInTop_6_36[17] , \wRegInTop_6_36[16] , 
        \wRegInTop_6_36[15] , \wRegInTop_6_36[14] , \wRegInTop_6_36[13] , 
        \wRegInTop_6_36[12] , \wRegInTop_6_36[11] , \wRegInTop_6_36[10] , 
        \wRegInTop_6_36[9] , \wRegInTop_6_36[8] , \wRegInTop_6_36[7] , 
        \wRegInTop_6_36[6] , \wRegInTop_6_36[5] , \wRegInTop_6_36[4] , 
        \wRegInTop_6_36[3] , \wRegInTop_6_36[2] , \wRegInTop_6_36[1] , 
        \wRegInTop_6_36[0] }), .R_WR(\wRegEnTop_6_37[0] ), .R_In({
        \wRegOut_6_37[31] , \wRegOut_6_37[30] , \wRegOut_6_37[29] , 
        \wRegOut_6_37[28] , \wRegOut_6_37[27] , \wRegOut_6_37[26] , 
        \wRegOut_6_37[25] , \wRegOut_6_37[24] , \wRegOut_6_37[23] , 
        \wRegOut_6_37[22] , \wRegOut_6_37[21] , \wRegOut_6_37[20] , 
        \wRegOut_6_37[19] , \wRegOut_6_37[18] , \wRegOut_6_37[17] , 
        \wRegOut_6_37[16] , \wRegOut_6_37[15] , \wRegOut_6_37[14] , 
        \wRegOut_6_37[13] , \wRegOut_6_37[12] , \wRegOut_6_37[11] , 
        \wRegOut_6_37[10] , \wRegOut_6_37[9] , \wRegOut_6_37[8] , 
        \wRegOut_6_37[7] , \wRegOut_6_37[6] , \wRegOut_6_37[5] , 
        \wRegOut_6_37[4] , \wRegOut_6_37[3] , \wRegOut_6_37[2] , 
        \wRegOut_6_37[1] , \wRegOut_6_37[0] }), .R_Out({\wRegInTop_6_37[31] , 
        \wRegInTop_6_37[30] , \wRegInTop_6_37[29] , \wRegInTop_6_37[28] , 
        \wRegInTop_6_37[27] , \wRegInTop_6_37[26] , \wRegInTop_6_37[25] , 
        \wRegInTop_6_37[24] , \wRegInTop_6_37[23] , \wRegInTop_6_37[22] , 
        \wRegInTop_6_37[21] , \wRegInTop_6_37[20] , \wRegInTop_6_37[19] , 
        \wRegInTop_6_37[18] , \wRegInTop_6_37[17] , \wRegInTop_6_37[16] , 
        \wRegInTop_6_37[15] , \wRegInTop_6_37[14] , \wRegInTop_6_37[13] , 
        \wRegInTop_6_37[12] , \wRegInTop_6_37[11] , \wRegInTop_6_37[10] , 
        \wRegInTop_6_37[9] , \wRegInTop_6_37[8] , \wRegInTop_6_37[7] , 
        \wRegInTop_6_37[6] , \wRegInTop_6_37[5] , \wRegInTop_6_37[4] , 
        \wRegInTop_6_37[3] , \wRegInTop_6_37[2] , \wRegInTop_6_37[1] , 
        \wRegInTop_6_37[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_27 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink91[31] , \ScanLink91[30] , \ScanLink91[29] , 
        \ScanLink91[28] , \ScanLink91[27] , \ScanLink91[26] , \ScanLink91[25] , 
        \ScanLink91[24] , \ScanLink91[23] , \ScanLink91[22] , \ScanLink91[21] , 
        \ScanLink91[20] , \ScanLink91[19] , \ScanLink91[18] , \ScanLink91[17] , 
        \ScanLink91[16] , \ScanLink91[15] , \ScanLink91[14] , \ScanLink91[13] , 
        \ScanLink91[12] , \ScanLink91[11] , \ScanLink91[10] , \ScanLink91[9] , 
        \ScanLink91[8] , \ScanLink91[7] , \ScanLink91[6] , \ScanLink91[5] , 
        \ScanLink91[4] , \ScanLink91[3] , \ScanLink91[2] , \ScanLink91[1] , 
        \ScanLink91[0] }), .ScanOut({\ScanLink90[31] , \ScanLink90[30] , 
        \ScanLink90[29] , \ScanLink90[28] , \ScanLink90[27] , \ScanLink90[26] , 
        \ScanLink90[25] , \ScanLink90[24] , \ScanLink90[23] , \ScanLink90[22] , 
        \ScanLink90[21] , \ScanLink90[20] , \ScanLink90[19] , \ScanLink90[18] , 
        \ScanLink90[17] , \ScanLink90[16] , \ScanLink90[15] , \ScanLink90[14] , 
        \ScanLink90[13] , \ScanLink90[12] , \ScanLink90[11] , \ScanLink90[10] , 
        \ScanLink90[9] , \ScanLink90[8] , \ScanLink90[7] , \ScanLink90[6] , 
        \ScanLink90[5] , \ScanLink90[4] , \ScanLink90[3] , \ScanLink90[2] , 
        \ScanLink90[1] , \ScanLink90[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_27[31] , \wRegOut_6_27[30] , 
        \wRegOut_6_27[29] , \wRegOut_6_27[28] , \wRegOut_6_27[27] , 
        \wRegOut_6_27[26] , \wRegOut_6_27[25] , \wRegOut_6_27[24] , 
        \wRegOut_6_27[23] , \wRegOut_6_27[22] , \wRegOut_6_27[21] , 
        \wRegOut_6_27[20] , \wRegOut_6_27[19] , \wRegOut_6_27[18] , 
        \wRegOut_6_27[17] , \wRegOut_6_27[16] , \wRegOut_6_27[15] , 
        \wRegOut_6_27[14] , \wRegOut_6_27[13] , \wRegOut_6_27[12] , 
        \wRegOut_6_27[11] , \wRegOut_6_27[10] , \wRegOut_6_27[9] , 
        \wRegOut_6_27[8] , \wRegOut_6_27[7] , \wRegOut_6_27[6] , 
        \wRegOut_6_27[5] , \wRegOut_6_27[4] , \wRegOut_6_27[3] , 
        \wRegOut_6_27[2] , \wRegOut_6_27[1] , \wRegOut_6_27[0] }), .Enable1(
        \wRegEnTop_6_27[0] ), .Enable2(\wRegEnBot_6_27[0] ), .In1({
        \wRegInTop_6_27[31] , \wRegInTop_6_27[30] , \wRegInTop_6_27[29] , 
        \wRegInTop_6_27[28] , \wRegInTop_6_27[27] , \wRegInTop_6_27[26] , 
        \wRegInTop_6_27[25] , \wRegInTop_6_27[24] , \wRegInTop_6_27[23] , 
        \wRegInTop_6_27[22] , \wRegInTop_6_27[21] , \wRegInTop_6_27[20] , 
        \wRegInTop_6_27[19] , \wRegInTop_6_27[18] , \wRegInTop_6_27[17] , 
        \wRegInTop_6_27[16] , \wRegInTop_6_27[15] , \wRegInTop_6_27[14] , 
        \wRegInTop_6_27[13] , \wRegInTop_6_27[12] , \wRegInTop_6_27[11] , 
        \wRegInTop_6_27[10] , \wRegInTop_6_27[9] , \wRegInTop_6_27[8] , 
        \wRegInTop_6_27[7] , \wRegInTop_6_27[6] , \wRegInTop_6_27[5] , 
        \wRegInTop_6_27[4] , \wRegInTop_6_27[3] , \wRegInTop_6_27[2] , 
        \wRegInTop_6_27[1] , \wRegInTop_6_27[0] }), .In2({\wRegInBot_6_27[31] , 
        \wRegInBot_6_27[30] , \wRegInBot_6_27[29] , \wRegInBot_6_27[28] , 
        \wRegInBot_6_27[27] , \wRegInBot_6_27[26] , \wRegInBot_6_27[25] , 
        \wRegInBot_6_27[24] , \wRegInBot_6_27[23] , \wRegInBot_6_27[22] , 
        \wRegInBot_6_27[21] , \wRegInBot_6_27[20] , \wRegInBot_6_27[19] , 
        \wRegInBot_6_27[18] , \wRegInBot_6_27[17] , \wRegInBot_6_27[16] , 
        \wRegInBot_6_27[15] , \wRegInBot_6_27[14] , \wRegInBot_6_27[13] , 
        \wRegInBot_6_27[12] , \wRegInBot_6_27[11] , \wRegInBot_6_27[10] , 
        \wRegInBot_6_27[9] , \wRegInBot_6_27[8] , \wRegInBot_6_27[7] , 
        \wRegInBot_6_27[6] , \wRegInBot_6_27[5] , \wRegInBot_6_27[4] , 
        \wRegInBot_6_27[3] , \wRegInBot_6_27[2] , \wRegInBot_6_27[1] , 
        \wRegInBot_6_27[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_53 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink181[31] , \ScanLink181[30] , \ScanLink181[29] , 
        \ScanLink181[28] , \ScanLink181[27] , \ScanLink181[26] , 
        \ScanLink181[25] , \ScanLink181[24] , \ScanLink181[23] , 
        \ScanLink181[22] , \ScanLink181[21] , \ScanLink181[20] , 
        \ScanLink181[19] , \ScanLink181[18] , \ScanLink181[17] , 
        \ScanLink181[16] , \ScanLink181[15] , \ScanLink181[14] , 
        \ScanLink181[13] , \ScanLink181[12] , \ScanLink181[11] , 
        \ScanLink181[10] , \ScanLink181[9] , \ScanLink181[8] , 
        \ScanLink181[7] , \ScanLink181[6] , \ScanLink181[5] , \ScanLink181[4] , 
        \ScanLink181[3] , \ScanLink181[2] , \ScanLink181[1] , \ScanLink181[0] 
        }), .ScanOut({\ScanLink180[31] , \ScanLink180[30] , \ScanLink180[29] , 
        \ScanLink180[28] , \ScanLink180[27] , \ScanLink180[26] , 
        \ScanLink180[25] , \ScanLink180[24] , \ScanLink180[23] , 
        \ScanLink180[22] , \ScanLink180[21] , \ScanLink180[20] , 
        \ScanLink180[19] , \ScanLink180[18] , \ScanLink180[17] , 
        \ScanLink180[16] , \ScanLink180[15] , \ScanLink180[14] , 
        \ScanLink180[13] , \ScanLink180[12] , \ScanLink180[11] , 
        \ScanLink180[10] , \ScanLink180[9] , \ScanLink180[8] , 
        \ScanLink180[7] , \ScanLink180[6] , \ScanLink180[5] , \ScanLink180[4] , 
        \ScanLink180[3] , \ScanLink180[2] , \ScanLink180[1] , \ScanLink180[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_53[31] , 
        \wRegOut_7_53[30] , \wRegOut_7_53[29] , \wRegOut_7_53[28] , 
        \wRegOut_7_53[27] , \wRegOut_7_53[26] , \wRegOut_7_53[25] , 
        \wRegOut_7_53[24] , \wRegOut_7_53[23] , \wRegOut_7_53[22] , 
        \wRegOut_7_53[21] , \wRegOut_7_53[20] , \wRegOut_7_53[19] , 
        \wRegOut_7_53[18] , \wRegOut_7_53[17] , \wRegOut_7_53[16] , 
        \wRegOut_7_53[15] , \wRegOut_7_53[14] , \wRegOut_7_53[13] , 
        \wRegOut_7_53[12] , \wRegOut_7_53[11] , \wRegOut_7_53[10] , 
        \wRegOut_7_53[9] , \wRegOut_7_53[8] , \wRegOut_7_53[7] , 
        \wRegOut_7_53[6] , \wRegOut_7_53[5] , \wRegOut_7_53[4] , 
        \wRegOut_7_53[3] , \wRegOut_7_53[2] , \wRegOut_7_53[1] , 
        \wRegOut_7_53[0] }), .Enable1(\wRegEnTop_7_53[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_53[31] , \wRegInTop_7_53[30] , \wRegInTop_7_53[29] , 
        \wRegInTop_7_53[28] , \wRegInTop_7_53[27] , \wRegInTop_7_53[26] , 
        \wRegInTop_7_53[25] , \wRegInTop_7_53[24] , \wRegInTop_7_53[23] , 
        \wRegInTop_7_53[22] , \wRegInTop_7_53[21] , \wRegInTop_7_53[20] , 
        \wRegInTop_7_53[19] , \wRegInTop_7_53[18] , \wRegInTop_7_53[17] , 
        \wRegInTop_7_53[16] , \wRegInTop_7_53[15] , \wRegInTop_7_53[14] , 
        \wRegInTop_7_53[13] , \wRegInTop_7_53[12] , \wRegInTop_7_53[11] , 
        \wRegInTop_7_53[10] , \wRegInTop_7_53[9] , \wRegInTop_7_53[8] , 
        \wRegInTop_7_53[7] , \wRegInTop_7_53[6] , \wRegInTop_7_53[5] , 
        \wRegInTop_7_53[4] , \wRegInTop_7_53[3] , \wRegInTop_7_53[2] , 
        \wRegInTop_7_53[1] , \wRegInTop_7_53[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_49 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink113[31] , \ScanLink113[30] , \ScanLink113[29] , 
        \ScanLink113[28] , \ScanLink113[27] , \ScanLink113[26] , 
        \ScanLink113[25] , \ScanLink113[24] , \ScanLink113[23] , 
        \ScanLink113[22] , \ScanLink113[21] , \ScanLink113[20] , 
        \ScanLink113[19] , \ScanLink113[18] , \ScanLink113[17] , 
        \ScanLink113[16] , \ScanLink113[15] , \ScanLink113[14] , 
        \ScanLink113[13] , \ScanLink113[12] , \ScanLink113[11] , 
        \ScanLink113[10] , \ScanLink113[9] , \ScanLink113[8] , 
        \ScanLink113[7] , \ScanLink113[6] , \ScanLink113[5] , \ScanLink113[4] , 
        \ScanLink113[3] , \ScanLink113[2] , \ScanLink113[1] , \ScanLink113[0] 
        }), .ScanOut({\ScanLink112[31] , \ScanLink112[30] , \ScanLink112[29] , 
        \ScanLink112[28] , \ScanLink112[27] , \ScanLink112[26] , 
        \ScanLink112[25] , \ScanLink112[24] , \ScanLink112[23] , 
        \ScanLink112[22] , \ScanLink112[21] , \ScanLink112[20] , 
        \ScanLink112[19] , \ScanLink112[18] , \ScanLink112[17] , 
        \ScanLink112[16] , \ScanLink112[15] , \ScanLink112[14] , 
        \ScanLink112[13] , \ScanLink112[12] , \ScanLink112[11] , 
        \ScanLink112[10] , \ScanLink112[9] , \ScanLink112[8] , 
        \ScanLink112[7] , \ScanLink112[6] , \ScanLink112[5] , \ScanLink112[4] , 
        \ScanLink112[3] , \ScanLink112[2] , \ScanLink112[1] , \ScanLink112[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_49[31] , 
        \wRegOut_6_49[30] , \wRegOut_6_49[29] , \wRegOut_6_49[28] , 
        \wRegOut_6_49[27] , \wRegOut_6_49[26] , \wRegOut_6_49[25] , 
        \wRegOut_6_49[24] , \wRegOut_6_49[23] , \wRegOut_6_49[22] , 
        \wRegOut_6_49[21] , \wRegOut_6_49[20] , \wRegOut_6_49[19] , 
        \wRegOut_6_49[18] , \wRegOut_6_49[17] , \wRegOut_6_49[16] , 
        \wRegOut_6_49[15] , \wRegOut_6_49[14] , \wRegOut_6_49[13] , 
        \wRegOut_6_49[12] , \wRegOut_6_49[11] , \wRegOut_6_49[10] , 
        \wRegOut_6_49[9] , \wRegOut_6_49[8] , \wRegOut_6_49[7] , 
        \wRegOut_6_49[6] , \wRegOut_6_49[5] , \wRegOut_6_49[4] , 
        \wRegOut_6_49[3] , \wRegOut_6_49[2] , \wRegOut_6_49[1] , 
        \wRegOut_6_49[0] }), .Enable1(\wRegEnTop_6_49[0] ), .Enable2(
        \wRegEnBot_6_49[0] ), .In1({\wRegInTop_6_49[31] , \wRegInTop_6_49[30] , 
        \wRegInTop_6_49[29] , \wRegInTop_6_49[28] , \wRegInTop_6_49[27] , 
        \wRegInTop_6_49[26] , \wRegInTop_6_49[25] , \wRegInTop_6_49[24] , 
        \wRegInTop_6_49[23] , \wRegInTop_6_49[22] , \wRegInTop_6_49[21] , 
        \wRegInTop_6_49[20] , \wRegInTop_6_49[19] , \wRegInTop_6_49[18] , 
        \wRegInTop_6_49[17] , \wRegInTop_6_49[16] , \wRegInTop_6_49[15] , 
        \wRegInTop_6_49[14] , \wRegInTop_6_49[13] , \wRegInTop_6_49[12] , 
        \wRegInTop_6_49[11] , \wRegInTop_6_49[10] , \wRegInTop_6_49[9] , 
        \wRegInTop_6_49[8] , \wRegInTop_6_49[7] , \wRegInTop_6_49[6] , 
        \wRegInTop_6_49[5] , \wRegInTop_6_49[4] , \wRegInTop_6_49[3] , 
        \wRegInTop_6_49[2] , \wRegInTop_6_49[1] , \wRegInTop_6_49[0] }), .In2(
        {\wRegInBot_6_49[31] , \wRegInBot_6_49[30] , \wRegInBot_6_49[29] , 
        \wRegInBot_6_49[28] , \wRegInBot_6_49[27] , \wRegInBot_6_49[26] , 
        \wRegInBot_6_49[25] , \wRegInBot_6_49[24] , \wRegInBot_6_49[23] , 
        \wRegInBot_6_49[22] , \wRegInBot_6_49[21] , \wRegInBot_6_49[20] , 
        \wRegInBot_6_49[19] , \wRegInBot_6_49[18] , \wRegInBot_6_49[17] , 
        \wRegInBot_6_49[16] , \wRegInBot_6_49[15] , \wRegInBot_6_49[14] , 
        \wRegInBot_6_49[13] , \wRegInBot_6_49[12] , \wRegInBot_6_49[11] , 
        \wRegInBot_6_49[10] , \wRegInBot_6_49[9] , \wRegInBot_6_49[8] , 
        \wRegInBot_6_49[7] , \wRegInBot_6_49[6] , \wRegInBot_6_49[5] , 
        \wRegInBot_6_49[4] , \wRegInBot_6_49[3] , \wRegInBot_6_49[2] , 
        \wRegInBot_6_49[1] , \wRegInBot_6_49[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_91 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink219[31] , \ScanLink219[30] , \ScanLink219[29] , 
        \ScanLink219[28] , \ScanLink219[27] , \ScanLink219[26] , 
        \ScanLink219[25] , \ScanLink219[24] , \ScanLink219[23] , 
        \ScanLink219[22] , \ScanLink219[21] , \ScanLink219[20] , 
        \ScanLink219[19] , \ScanLink219[18] , \ScanLink219[17] , 
        \ScanLink219[16] , \ScanLink219[15] , \ScanLink219[14] , 
        \ScanLink219[13] , \ScanLink219[12] , \ScanLink219[11] , 
        \ScanLink219[10] , \ScanLink219[9] , \ScanLink219[8] , 
        \ScanLink219[7] , \ScanLink219[6] , \ScanLink219[5] , \ScanLink219[4] , 
        \ScanLink219[3] , \ScanLink219[2] , \ScanLink219[1] , \ScanLink219[0] 
        }), .ScanOut({\ScanLink218[31] , \ScanLink218[30] , \ScanLink218[29] , 
        \ScanLink218[28] , \ScanLink218[27] , \ScanLink218[26] , 
        \ScanLink218[25] , \ScanLink218[24] , \ScanLink218[23] , 
        \ScanLink218[22] , \ScanLink218[21] , \ScanLink218[20] , 
        \ScanLink218[19] , \ScanLink218[18] , \ScanLink218[17] , 
        \ScanLink218[16] , \ScanLink218[15] , \ScanLink218[14] , 
        \ScanLink218[13] , \ScanLink218[12] , \ScanLink218[11] , 
        \ScanLink218[10] , \ScanLink218[9] , \ScanLink218[8] , 
        \ScanLink218[7] , \ScanLink218[6] , \ScanLink218[5] , \ScanLink218[4] , 
        \ScanLink218[3] , \ScanLink218[2] , \ScanLink218[1] , \ScanLink218[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_91[31] , 
        \wRegOut_7_91[30] , \wRegOut_7_91[29] , \wRegOut_7_91[28] , 
        \wRegOut_7_91[27] , \wRegOut_7_91[26] , \wRegOut_7_91[25] , 
        \wRegOut_7_91[24] , \wRegOut_7_91[23] , \wRegOut_7_91[22] , 
        \wRegOut_7_91[21] , \wRegOut_7_91[20] , \wRegOut_7_91[19] , 
        \wRegOut_7_91[18] , \wRegOut_7_91[17] , \wRegOut_7_91[16] , 
        \wRegOut_7_91[15] , \wRegOut_7_91[14] , \wRegOut_7_91[13] , 
        \wRegOut_7_91[12] , \wRegOut_7_91[11] , \wRegOut_7_91[10] , 
        \wRegOut_7_91[9] , \wRegOut_7_91[8] , \wRegOut_7_91[7] , 
        \wRegOut_7_91[6] , \wRegOut_7_91[5] , \wRegOut_7_91[4] , 
        \wRegOut_7_91[3] , \wRegOut_7_91[2] , \wRegOut_7_91[1] , 
        \wRegOut_7_91[0] }), .Enable1(\wRegEnTop_7_91[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_91[31] , \wRegInTop_7_91[30] , \wRegInTop_7_91[29] , 
        \wRegInTop_7_91[28] , \wRegInTop_7_91[27] , \wRegInTop_7_91[26] , 
        \wRegInTop_7_91[25] , \wRegInTop_7_91[24] , \wRegInTop_7_91[23] , 
        \wRegInTop_7_91[22] , \wRegInTop_7_91[21] , \wRegInTop_7_91[20] , 
        \wRegInTop_7_91[19] , \wRegInTop_7_91[18] , \wRegInTop_7_91[17] , 
        \wRegInTop_7_91[16] , \wRegInTop_7_91[15] , \wRegInTop_7_91[14] , 
        \wRegInTop_7_91[13] , \wRegInTop_7_91[12] , \wRegInTop_7_91[11] , 
        \wRegInTop_7_91[10] , \wRegInTop_7_91[9] , \wRegInTop_7_91[8] , 
        \wRegInTop_7_91[7] , \wRegInTop_7_91[6] , \wRegInTop_7_91[5] , 
        \wRegInTop_7_91[4] , \wRegInTop_7_91[3] , \wRegInTop_7_91[2] , 
        \wRegInTop_7_91[1] , \wRegInTop_7_91[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_0[0] ), .P_In({\wRegOut_5_0[31] , 
        \wRegOut_5_0[30] , \wRegOut_5_0[29] , \wRegOut_5_0[28] , 
        \wRegOut_5_0[27] , \wRegOut_5_0[26] , \wRegOut_5_0[25] , 
        \wRegOut_5_0[24] , \wRegOut_5_0[23] , \wRegOut_5_0[22] , 
        \wRegOut_5_0[21] , \wRegOut_5_0[20] , \wRegOut_5_0[19] , 
        \wRegOut_5_0[18] , \wRegOut_5_0[17] , \wRegOut_5_0[16] , 
        \wRegOut_5_0[15] , \wRegOut_5_0[14] , \wRegOut_5_0[13] , 
        \wRegOut_5_0[12] , \wRegOut_5_0[11] , \wRegOut_5_0[10] , 
        \wRegOut_5_0[9] , \wRegOut_5_0[8] , \wRegOut_5_0[7] , \wRegOut_5_0[6] , 
        \wRegOut_5_0[5] , \wRegOut_5_0[4] , \wRegOut_5_0[3] , \wRegOut_5_0[2] , 
        \wRegOut_5_0[1] , \wRegOut_5_0[0] }), .P_Out({\wRegInBot_5_0[31] , 
        \wRegInBot_5_0[30] , \wRegInBot_5_0[29] , \wRegInBot_5_0[28] , 
        \wRegInBot_5_0[27] , \wRegInBot_5_0[26] , \wRegInBot_5_0[25] , 
        \wRegInBot_5_0[24] , \wRegInBot_5_0[23] , \wRegInBot_5_0[22] , 
        \wRegInBot_5_0[21] , \wRegInBot_5_0[20] , \wRegInBot_5_0[19] , 
        \wRegInBot_5_0[18] , \wRegInBot_5_0[17] , \wRegInBot_5_0[16] , 
        \wRegInBot_5_0[15] , \wRegInBot_5_0[14] , \wRegInBot_5_0[13] , 
        \wRegInBot_5_0[12] , \wRegInBot_5_0[11] , \wRegInBot_5_0[10] , 
        \wRegInBot_5_0[9] , \wRegInBot_5_0[8] , \wRegInBot_5_0[7] , 
        \wRegInBot_5_0[6] , \wRegInBot_5_0[5] , \wRegInBot_5_0[4] , 
        \wRegInBot_5_0[3] , \wRegInBot_5_0[2] , \wRegInBot_5_0[1] , 
        \wRegInBot_5_0[0] }), .L_WR(\wRegEnTop_6_0[0] ), .L_In({
        \wRegOut_6_0[31] , \wRegOut_6_0[30] , \wRegOut_6_0[29] , 
        \wRegOut_6_0[28] , \wRegOut_6_0[27] , \wRegOut_6_0[26] , 
        \wRegOut_6_0[25] , \wRegOut_6_0[24] , \wRegOut_6_0[23] , 
        \wRegOut_6_0[22] , \wRegOut_6_0[21] , \wRegOut_6_0[20] , 
        \wRegOut_6_0[19] , \wRegOut_6_0[18] , \wRegOut_6_0[17] , 
        \wRegOut_6_0[16] , \wRegOut_6_0[15] , \wRegOut_6_0[14] , 
        \wRegOut_6_0[13] , \wRegOut_6_0[12] , \wRegOut_6_0[11] , 
        \wRegOut_6_0[10] , \wRegOut_6_0[9] , \wRegOut_6_0[8] , 
        \wRegOut_6_0[7] , \wRegOut_6_0[6] , \wRegOut_6_0[5] , \wRegOut_6_0[4] , 
        \wRegOut_6_0[3] , \wRegOut_6_0[2] , \wRegOut_6_0[1] , \wRegOut_6_0[0] 
        }), .L_Out({\wRegInTop_6_0[31] , \wRegInTop_6_0[30] , 
        \wRegInTop_6_0[29] , \wRegInTop_6_0[28] , \wRegInTop_6_0[27] , 
        \wRegInTop_6_0[26] , \wRegInTop_6_0[25] , \wRegInTop_6_0[24] , 
        \wRegInTop_6_0[23] , \wRegInTop_6_0[22] , \wRegInTop_6_0[21] , 
        \wRegInTop_6_0[20] , \wRegInTop_6_0[19] , \wRegInTop_6_0[18] , 
        \wRegInTop_6_0[17] , \wRegInTop_6_0[16] , \wRegInTop_6_0[15] , 
        \wRegInTop_6_0[14] , \wRegInTop_6_0[13] , \wRegInTop_6_0[12] , 
        \wRegInTop_6_0[11] , \wRegInTop_6_0[10] , \wRegInTop_6_0[9] , 
        \wRegInTop_6_0[8] , \wRegInTop_6_0[7] , \wRegInTop_6_0[6] , 
        \wRegInTop_6_0[5] , \wRegInTop_6_0[4] , \wRegInTop_6_0[3] , 
        \wRegInTop_6_0[2] , \wRegInTop_6_0[1] , \wRegInTop_6_0[0] }), .R_WR(
        \wRegEnTop_6_1[0] ), .R_In({\wRegOut_6_1[31] , \wRegOut_6_1[30] , 
        \wRegOut_6_1[29] , \wRegOut_6_1[28] , \wRegOut_6_1[27] , 
        \wRegOut_6_1[26] , \wRegOut_6_1[25] , \wRegOut_6_1[24] , 
        \wRegOut_6_1[23] , \wRegOut_6_1[22] , \wRegOut_6_1[21] , 
        \wRegOut_6_1[20] , \wRegOut_6_1[19] , \wRegOut_6_1[18] , 
        \wRegOut_6_1[17] , \wRegOut_6_1[16] , \wRegOut_6_1[15] , 
        \wRegOut_6_1[14] , \wRegOut_6_1[13] , \wRegOut_6_1[12] , 
        \wRegOut_6_1[11] , \wRegOut_6_1[10] , \wRegOut_6_1[9] , 
        \wRegOut_6_1[8] , \wRegOut_6_1[7] , \wRegOut_6_1[6] , \wRegOut_6_1[5] , 
        \wRegOut_6_1[4] , \wRegOut_6_1[3] , \wRegOut_6_1[2] , \wRegOut_6_1[1] , 
        \wRegOut_6_1[0] }), .R_Out({\wRegInTop_6_1[31] , \wRegInTop_6_1[30] , 
        \wRegInTop_6_1[29] , \wRegInTop_6_1[28] , \wRegInTop_6_1[27] , 
        \wRegInTop_6_1[26] , \wRegInTop_6_1[25] , \wRegInTop_6_1[24] , 
        \wRegInTop_6_1[23] , \wRegInTop_6_1[22] , \wRegInTop_6_1[21] , 
        \wRegInTop_6_1[20] , \wRegInTop_6_1[19] , \wRegInTop_6_1[18] , 
        \wRegInTop_6_1[17] , \wRegInTop_6_1[16] , \wRegInTop_6_1[15] , 
        \wRegInTop_6_1[14] , \wRegInTop_6_1[13] , \wRegInTop_6_1[12] , 
        \wRegInTop_6_1[11] , \wRegInTop_6_1[10] , \wRegInTop_6_1[9] , 
        \wRegInTop_6_1[8] , \wRegInTop_6_1[7] , \wRegInTop_6_1[6] , 
        \wRegInTop_6_1[5] , \wRegInTop_6_1[4] , \wRegInTop_6_1[3] , 
        \wRegInTop_6_1[2] , \wRegInTop_6_1[1] , \wRegInTop_6_1[0] }) );
    BHeap_Node_WIDTH32 BHN_6_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_61[0] ), .P_In({\wRegOut_6_61[31] , 
        \wRegOut_6_61[30] , \wRegOut_6_61[29] , \wRegOut_6_61[28] , 
        \wRegOut_6_61[27] , \wRegOut_6_61[26] , \wRegOut_6_61[25] , 
        \wRegOut_6_61[24] , \wRegOut_6_61[23] , \wRegOut_6_61[22] , 
        \wRegOut_6_61[21] , \wRegOut_6_61[20] , \wRegOut_6_61[19] , 
        \wRegOut_6_61[18] , \wRegOut_6_61[17] , \wRegOut_6_61[16] , 
        \wRegOut_6_61[15] , \wRegOut_6_61[14] , \wRegOut_6_61[13] , 
        \wRegOut_6_61[12] , \wRegOut_6_61[11] , \wRegOut_6_61[10] , 
        \wRegOut_6_61[9] , \wRegOut_6_61[8] , \wRegOut_6_61[7] , 
        \wRegOut_6_61[6] , \wRegOut_6_61[5] , \wRegOut_6_61[4] , 
        \wRegOut_6_61[3] , \wRegOut_6_61[2] , \wRegOut_6_61[1] , 
        \wRegOut_6_61[0] }), .P_Out({\wRegInBot_6_61[31] , 
        \wRegInBot_6_61[30] , \wRegInBot_6_61[29] , \wRegInBot_6_61[28] , 
        \wRegInBot_6_61[27] , \wRegInBot_6_61[26] , \wRegInBot_6_61[25] , 
        \wRegInBot_6_61[24] , \wRegInBot_6_61[23] , \wRegInBot_6_61[22] , 
        \wRegInBot_6_61[21] , \wRegInBot_6_61[20] , \wRegInBot_6_61[19] , 
        \wRegInBot_6_61[18] , \wRegInBot_6_61[17] , \wRegInBot_6_61[16] , 
        \wRegInBot_6_61[15] , \wRegInBot_6_61[14] , \wRegInBot_6_61[13] , 
        \wRegInBot_6_61[12] , \wRegInBot_6_61[11] , \wRegInBot_6_61[10] , 
        \wRegInBot_6_61[9] , \wRegInBot_6_61[8] , \wRegInBot_6_61[7] , 
        \wRegInBot_6_61[6] , \wRegInBot_6_61[5] , \wRegInBot_6_61[4] , 
        \wRegInBot_6_61[3] , \wRegInBot_6_61[2] , \wRegInBot_6_61[1] , 
        \wRegInBot_6_61[0] }), .L_WR(\wRegEnTop_7_122[0] ), .L_In({
        \wRegOut_7_122[31] , \wRegOut_7_122[30] , \wRegOut_7_122[29] , 
        \wRegOut_7_122[28] , \wRegOut_7_122[27] , \wRegOut_7_122[26] , 
        \wRegOut_7_122[25] , \wRegOut_7_122[24] , \wRegOut_7_122[23] , 
        \wRegOut_7_122[22] , \wRegOut_7_122[21] , \wRegOut_7_122[20] , 
        \wRegOut_7_122[19] , \wRegOut_7_122[18] , \wRegOut_7_122[17] , 
        \wRegOut_7_122[16] , \wRegOut_7_122[15] , \wRegOut_7_122[14] , 
        \wRegOut_7_122[13] , \wRegOut_7_122[12] , \wRegOut_7_122[11] , 
        \wRegOut_7_122[10] , \wRegOut_7_122[9] , \wRegOut_7_122[8] , 
        \wRegOut_7_122[7] , \wRegOut_7_122[6] , \wRegOut_7_122[5] , 
        \wRegOut_7_122[4] , \wRegOut_7_122[3] , \wRegOut_7_122[2] , 
        \wRegOut_7_122[1] , \wRegOut_7_122[0] }), .L_Out({
        \wRegInTop_7_122[31] , \wRegInTop_7_122[30] , \wRegInTop_7_122[29] , 
        \wRegInTop_7_122[28] , \wRegInTop_7_122[27] , \wRegInTop_7_122[26] , 
        \wRegInTop_7_122[25] , \wRegInTop_7_122[24] , \wRegInTop_7_122[23] , 
        \wRegInTop_7_122[22] , \wRegInTop_7_122[21] , \wRegInTop_7_122[20] , 
        \wRegInTop_7_122[19] , \wRegInTop_7_122[18] , \wRegInTop_7_122[17] , 
        \wRegInTop_7_122[16] , \wRegInTop_7_122[15] , \wRegInTop_7_122[14] , 
        \wRegInTop_7_122[13] , \wRegInTop_7_122[12] , \wRegInTop_7_122[11] , 
        \wRegInTop_7_122[10] , \wRegInTop_7_122[9] , \wRegInTop_7_122[8] , 
        \wRegInTop_7_122[7] , \wRegInTop_7_122[6] , \wRegInTop_7_122[5] , 
        \wRegInTop_7_122[4] , \wRegInTop_7_122[3] , \wRegInTop_7_122[2] , 
        \wRegInTop_7_122[1] , \wRegInTop_7_122[0] }), .R_WR(
        \wRegEnTop_7_123[0] ), .R_In({\wRegOut_7_123[31] , \wRegOut_7_123[30] , 
        \wRegOut_7_123[29] , \wRegOut_7_123[28] , \wRegOut_7_123[27] , 
        \wRegOut_7_123[26] , \wRegOut_7_123[25] , \wRegOut_7_123[24] , 
        \wRegOut_7_123[23] , \wRegOut_7_123[22] , \wRegOut_7_123[21] , 
        \wRegOut_7_123[20] , \wRegOut_7_123[19] , \wRegOut_7_123[18] , 
        \wRegOut_7_123[17] , \wRegOut_7_123[16] , \wRegOut_7_123[15] , 
        \wRegOut_7_123[14] , \wRegOut_7_123[13] , \wRegOut_7_123[12] , 
        \wRegOut_7_123[11] , \wRegOut_7_123[10] , \wRegOut_7_123[9] , 
        \wRegOut_7_123[8] , \wRegOut_7_123[7] , \wRegOut_7_123[6] , 
        \wRegOut_7_123[5] , \wRegOut_7_123[4] , \wRegOut_7_123[3] , 
        \wRegOut_7_123[2] , \wRegOut_7_123[1] , \wRegOut_7_123[0] }), .R_Out({
        \wRegInTop_7_123[31] , \wRegInTop_7_123[30] , \wRegInTop_7_123[29] , 
        \wRegInTop_7_123[28] , \wRegInTop_7_123[27] , \wRegInTop_7_123[26] , 
        \wRegInTop_7_123[25] , \wRegInTop_7_123[24] , \wRegInTop_7_123[23] , 
        \wRegInTop_7_123[22] , \wRegInTop_7_123[21] , \wRegInTop_7_123[20] , 
        \wRegInTop_7_123[19] , \wRegInTop_7_123[18] , \wRegInTop_7_123[17] , 
        \wRegInTop_7_123[16] , \wRegInTop_7_123[15] , \wRegInTop_7_123[14] , 
        \wRegInTop_7_123[13] , \wRegInTop_7_123[12] , \wRegInTop_7_123[11] , 
        \wRegInTop_7_123[10] , \wRegInTop_7_123[9] , \wRegInTop_7_123[8] , 
        \wRegInTop_7_123[7] , \wRegInTop_7_123[6] , \wRegInTop_7_123[5] , 
        \wRegInTop_7_123[4] , \wRegInTop_7_123[3] , \wRegInTop_7_123[2] , 
        \wRegInTop_7_123[1] , \wRegInTop_7_123[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_52 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink116[31] , \ScanLink116[30] , \ScanLink116[29] , 
        \ScanLink116[28] , \ScanLink116[27] , \ScanLink116[26] , 
        \ScanLink116[25] , \ScanLink116[24] , \ScanLink116[23] , 
        \ScanLink116[22] , \ScanLink116[21] , \ScanLink116[20] , 
        \ScanLink116[19] , \ScanLink116[18] , \ScanLink116[17] , 
        \ScanLink116[16] , \ScanLink116[15] , \ScanLink116[14] , 
        \ScanLink116[13] , \ScanLink116[12] , \ScanLink116[11] , 
        \ScanLink116[10] , \ScanLink116[9] , \ScanLink116[8] , 
        \ScanLink116[7] , \ScanLink116[6] , \ScanLink116[5] , \ScanLink116[4] , 
        \ScanLink116[3] , \ScanLink116[2] , \ScanLink116[1] , \ScanLink116[0] 
        }), .ScanOut({\ScanLink115[31] , \ScanLink115[30] , \ScanLink115[29] , 
        \ScanLink115[28] , \ScanLink115[27] , \ScanLink115[26] , 
        \ScanLink115[25] , \ScanLink115[24] , \ScanLink115[23] , 
        \ScanLink115[22] , \ScanLink115[21] , \ScanLink115[20] , 
        \ScanLink115[19] , \ScanLink115[18] , \ScanLink115[17] , 
        \ScanLink115[16] , \ScanLink115[15] , \ScanLink115[14] , 
        \ScanLink115[13] , \ScanLink115[12] , \ScanLink115[11] , 
        \ScanLink115[10] , \ScanLink115[9] , \ScanLink115[8] , 
        \ScanLink115[7] , \ScanLink115[6] , \ScanLink115[5] , \ScanLink115[4] , 
        \ScanLink115[3] , \ScanLink115[2] , \ScanLink115[1] , \ScanLink115[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_52[31] , 
        \wRegOut_6_52[30] , \wRegOut_6_52[29] , \wRegOut_6_52[28] , 
        \wRegOut_6_52[27] , \wRegOut_6_52[26] , \wRegOut_6_52[25] , 
        \wRegOut_6_52[24] , \wRegOut_6_52[23] , \wRegOut_6_52[22] , 
        \wRegOut_6_52[21] , \wRegOut_6_52[20] , \wRegOut_6_52[19] , 
        \wRegOut_6_52[18] , \wRegOut_6_52[17] , \wRegOut_6_52[16] , 
        \wRegOut_6_52[15] , \wRegOut_6_52[14] , \wRegOut_6_52[13] , 
        \wRegOut_6_52[12] , \wRegOut_6_52[11] , \wRegOut_6_52[10] , 
        \wRegOut_6_52[9] , \wRegOut_6_52[8] , \wRegOut_6_52[7] , 
        \wRegOut_6_52[6] , \wRegOut_6_52[5] , \wRegOut_6_52[4] , 
        \wRegOut_6_52[3] , \wRegOut_6_52[2] , \wRegOut_6_52[1] , 
        \wRegOut_6_52[0] }), .Enable1(\wRegEnTop_6_52[0] ), .Enable2(
        \wRegEnBot_6_52[0] ), .In1({\wRegInTop_6_52[31] , \wRegInTop_6_52[30] , 
        \wRegInTop_6_52[29] , \wRegInTop_6_52[28] , \wRegInTop_6_52[27] , 
        \wRegInTop_6_52[26] , \wRegInTop_6_52[25] , \wRegInTop_6_52[24] , 
        \wRegInTop_6_52[23] , \wRegInTop_6_52[22] , \wRegInTop_6_52[21] , 
        \wRegInTop_6_52[20] , \wRegInTop_6_52[19] , \wRegInTop_6_52[18] , 
        \wRegInTop_6_52[17] , \wRegInTop_6_52[16] , \wRegInTop_6_52[15] , 
        \wRegInTop_6_52[14] , \wRegInTop_6_52[13] , \wRegInTop_6_52[12] , 
        \wRegInTop_6_52[11] , \wRegInTop_6_52[10] , \wRegInTop_6_52[9] , 
        \wRegInTop_6_52[8] , \wRegInTop_6_52[7] , \wRegInTop_6_52[6] , 
        \wRegInTop_6_52[5] , \wRegInTop_6_52[4] , \wRegInTop_6_52[3] , 
        \wRegInTop_6_52[2] , \wRegInTop_6_52[1] , \wRegInTop_6_52[0] }), .In2(
        {\wRegInBot_6_52[31] , \wRegInBot_6_52[30] , \wRegInBot_6_52[29] , 
        \wRegInBot_6_52[28] , \wRegInBot_6_52[27] , \wRegInBot_6_52[26] , 
        \wRegInBot_6_52[25] , \wRegInBot_6_52[24] , \wRegInBot_6_52[23] , 
        \wRegInBot_6_52[22] , \wRegInBot_6_52[21] , \wRegInBot_6_52[20] , 
        \wRegInBot_6_52[19] , \wRegInBot_6_52[18] , \wRegInBot_6_52[17] , 
        \wRegInBot_6_52[16] , \wRegInBot_6_52[15] , \wRegInBot_6_52[14] , 
        \wRegInBot_6_52[13] , \wRegInBot_6_52[12] , \wRegInBot_6_52[11] , 
        \wRegInBot_6_52[10] , \wRegInBot_6_52[9] , \wRegInBot_6_52[8] , 
        \wRegInBot_6_52[7] , \wRegInBot_6_52[6] , \wRegInBot_6_52[5] , 
        \wRegInBot_6_52[4] , \wRegInBot_6_52[3] , \wRegInBot_6_52[2] , 
        \wRegInBot_6_52[1] , \wRegInBot_6_52[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_115 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink243[31] , \ScanLink243[30] , \ScanLink243[29] , 
        \ScanLink243[28] , \ScanLink243[27] , \ScanLink243[26] , 
        \ScanLink243[25] , \ScanLink243[24] , \ScanLink243[23] , 
        \ScanLink243[22] , \ScanLink243[21] , \ScanLink243[20] , 
        \ScanLink243[19] , \ScanLink243[18] , \ScanLink243[17] , 
        \ScanLink243[16] , \ScanLink243[15] , \ScanLink243[14] , 
        \ScanLink243[13] , \ScanLink243[12] , \ScanLink243[11] , 
        \ScanLink243[10] , \ScanLink243[9] , \ScanLink243[8] , 
        \ScanLink243[7] , \ScanLink243[6] , \ScanLink243[5] , \ScanLink243[4] , 
        \ScanLink243[3] , \ScanLink243[2] , \ScanLink243[1] , \ScanLink243[0] 
        }), .ScanOut({\ScanLink242[31] , \ScanLink242[30] , \ScanLink242[29] , 
        \ScanLink242[28] , \ScanLink242[27] , \ScanLink242[26] , 
        \ScanLink242[25] , \ScanLink242[24] , \ScanLink242[23] , 
        \ScanLink242[22] , \ScanLink242[21] , \ScanLink242[20] , 
        \ScanLink242[19] , \ScanLink242[18] , \ScanLink242[17] , 
        \ScanLink242[16] , \ScanLink242[15] , \ScanLink242[14] , 
        \ScanLink242[13] , \ScanLink242[12] , \ScanLink242[11] , 
        \ScanLink242[10] , \ScanLink242[9] , \ScanLink242[8] , 
        \ScanLink242[7] , \ScanLink242[6] , \ScanLink242[5] , \ScanLink242[4] , 
        \ScanLink242[3] , \ScanLink242[2] , \ScanLink242[1] , \ScanLink242[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_115[31] , 
        \wRegOut_7_115[30] , \wRegOut_7_115[29] , \wRegOut_7_115[28] , 
        \wRegOut_7_115[27] , \wRegOut_7_115[26] , \wRegOut_7_115[25] , 
        \wRegOut_7_115[24] , \wRegOut_7_115[23] , \wRegOut_7_115[22] , 
        \wRegOut_7_115[21] , \wRegOut_7_115[20] , \wRegOut_7_115[19] , 
        \wRegOut_7_115[18] , \wRegOut_7_115[17] , \wRegOut_7_115[16] , 
        \wRegOut_7_115[15] , \wRegOut_7_115[14] , \wRegOut_7_115[13] , 
        \wRegOut_7_115[12] , \wRegOut_7_115[11] , \wRegOut_7_115[10] , 
        \wRegOut_7_115[9] , \wRegOut_7_115[8] , \wRegOut_7_115[7] , 
        \wRegOut_7_115[6] , \wRegOut_7_115[5] , \wRegOut_7_115[4] , 
        \wRegOut_7_115[3] , \wRegOut_7_115[2] , \wRegOut_7_115[1] , 
        \wRegOut_7_115[0] }), .Enable1(\wRegEnTop_7_115[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_115[31] , \wRegInTop_7_115[30] , 
        \wRegInTop_7_115[29] , \wRegInTop_7_115[28] , \wRegInTop_7_115[27] , 
        \wRegInTop_7_115[26] , \wRegInTop_7_115[25] , \wRegInTop_7_115[24] , 
        \wRegInTop_7_115[23] , \wRegInTop_7_115[22] , \wRegInTop_7_115[21] , 
        \wRegInTop_7_115[20] , \wRegInTop_7_115[19] , \wRegInTop_7_115[18] , 
        \wRegInTop_7_115[17] , \wRegInTop_7_115[16] , \wRegInTop_7_115[15] , 
        \wRegInTop_7_115[14] , \wRegInTop_7_115[13] , \wRegInTop_7_115[12] , 
        \wRegInTop_7_115[11] , \wRegInTop_7_115[10] , \wRegInTop_7_115[9] , 
        \wRegInTop_7_115[8] , \wRegInTop_7_115[7] , \wRegInTop_7_115[6] , 
        \wRegInTop_7_115[5] , \wRegInTop_7_115[4] , \wRegInTop_7_115[3] , 
        \wRegInTop_7_115[2] , \wRegInTop_7_115[1] , \wRegInTop_7_115[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_46[0] ), .P_In({\wRegOut_6_46[31] , 
        \wRegOut_6_46[30] , \wRegOut_6_46[29] , \wRegOut_6_46[28] , 
        \wRegOut_6_46[27] , \wRegOut_6_46[26] , \wRegOut_6_46[25] , 
        \wRegOut_6_46[24] , \wRegOut_6_46[23] , \wRegOut_6_46[22] , 
        \wRegOut_6_46[21] , \wRegOut_6_46[20] , \wRegOut_6_46[19] , 
        \wRegOut_6_46[18] , \wRegOut_6_46[17] , \wRegOut_6_46[16] , 
        \wRegOut_6_46[15] , \wRegOut_6_46[14] , \wRegOut_6_46[13] , 
        \wRegOut_6_46[12] , \wRegOut_6_46[11] , \wRegOut_6_46[10] , 
        \wRegOut_6_46[9] , \wRegOut_6_46[8] , \wRegOut_6_46[7] , 
        \wRegOut_6_46[6] , \wRegOut_6_46[5] , \wRegOut_6_46[4] , 
        \wRegOut_6_46[3] , \wRegOut_6_46[2] , \wRegOut_6_46[1] , 
        \wRegOut_6_46[0] }), .P_Out({\wRegInBot_6_46[31] , 
        \wRegInBot_6_46[30] , \wRegInBot_6_46[29] , \wRegInBot_6_46[28] , 
        \wRegInBot_6_46[27] , \wRegInBot_6_46[26] , \wRegInBot_6_46[25] , 
        \wRegInBot_6_46[24] , \wRegInBot_6_46[23] , \wRegInBot_6_46[22] , 
        \wRegInBot_6_46[21] , \wRegInBot_6_46[20] , \wRegInBot_6_46[19] , 
        \wRegInBot_6_46[18] , \wRegInBot_6_46[17] , \wRegInBot_6_46[16] , 
        \wRegInBot_6_46[15] , \wRegInBot_6_46[14] , \wRegInBot_6_46[13] , 
        \wRegInBot_6_46[12] , \wRegInBot_6_46[11] , \wRegInBot_6_46[10] , 
        \wRegInBot_6_46[9] , \wRegInBot_6_46[8] , \wRegInBot_6_46[7] , 
        \wRegInBot_6_46[6] , \wRegInBot_6_46[5] , \wRegInBot_6_46[4] , 
        \wRegInBot_6_46[3] , \wRegInBot_6_46[2] , \wRegInBot_6_46[1] , 
        \wRegInBot_6_46[0] }), .L_WR(\wRegEnTop_7_92[0] ), .L_In({
        \wRegOut_7_92[31] , \wRegOut_7_92[30] , \wRegOut_7_92[29] , 
        \wRegOut_7_92[28] , \wRegOut_7_92[27] , \wRegOut_7_92[26] , 
        \wRegOut_7_92[25] , \wRegOut_7_92[24] , \wRegOut_7_92[23] , 
        \wRegOut_7_92[22] , \wRegOut_7_92[21] , \wRegOut_7_92[20] , 
        \wRegOut_7_92[19] , \wRegOut_7_92[18] , \wRegOut_7_92[17] , 
        \wRegOut_7_92[16] , \wRegOut_7_92[15] , \wRegOut_7_92[14] , 
        \wRegOut_7_92[13] , \wRegOut_7_92[12] , \wRegOut_7_92[11] , 
        \wRegOut_7_92[10] , \wRegOut_7_92[9] , \wRegOut_7_92[8] , 
        \wRegOut_7_92[7] , \wRegOut_7_92[6] , \wRegOut_7_92[5] , 
        \wRegOut_7_92[4] , \wRegOut_7_92[3] , \wRegOut_7_92[2] , 
        \wRegOut_7_92[1] , \wRegOut_7_92[0] }), .L_Out({\wRegInTop_7_92[31] , 
        \wRegInTop_7_92[30] , \wRegInTop_7_92[29] , \wRegInTop_7_92[28] , 
        \wRegInTop_7_92[27] , \wRegInTop_7_92[26] , \wRegInTop_7_92[25] , 
        \wRegInTop_7_92[24] , \wRegInTop_7_92[23] , \wRegInTop_7_92[22] , 
        \wRegInTop_7_92[21] , \wRegInTop_7_92[20] , \wRegInTop_7_92[19] , 
        \wRegInTop_7_92[18] , \wRegInTop_7_92[17] , \wRegInTop_7_92[16] , 
        \wRegInTop_7_92[15] , \wRegInTop_7_92[14] , \wRegInTop_7_92[13] , 
        \wRegInTop_7_92[12] , \wRegInTop_7_92[11] , \wRegInTop_7_92[10] , 
        \wRegInTop_7_92[9] , \wRegInTop_7_92[8] , \wRegInTop_7_92[7] , 
        \wRegInTop_7_92[6] , \wRegInTop_7_92[5] , \wRegInTop_7_92[4] , 
        \wRegInTop_7_92[3] , \wRegInTop_7_92[2] , \wRegInTop_7_92[1] , 
        \wRegInTop_7_92[0] }), .R_WR(\wRegEnTop_7_93[0] ), .R_In({
        \wRegOut_7_93[31] , \wRegOut_7_93[30] , \wRegOut_7_93[29] , 
        \wRegOut_7_93[28] , \wRegOut_7_93[27] , \wRegOut_7_93[26] , 
        \wRegOut_7_93[25] , \wRegOut_7_93[24] , \wRegOut_7_93[23] , 
        \wRegOut_7_93[22] , \wRegOut_7_93[21] , \wRegOut_7_93[20] , 
        \wRegOut_7_93[19] , \wRegOut_7_93[18] , \wRegOut_7_93[17] , 
        \wRegOut_7_93[16] , \wRegOut_7_93[15] , \wRegOut_7_93[14] , 
        \wRegOut_7_93[13] , \wRegOut_7_93[12] , \wRegOut_7_93[11] , 
        \wRegOut_7_93[10] , \wRegOut_7_93[9] , \wRegOut_7_93[8] , 
        \wRegOut_7_93[7] , \wRegOut_7_93[6] , \wRegOut_7_93[5] , 
        \wRegOut_7_93[4] , \wRegOut_7_93[3] , \wRegOut_7_93[2] , 
        \wRegOut_7_93[1] , \wRegOut_7_93[0] }), .R_Out({\wRegInTop_7_93[31] , 
        \wRegInTop_7_93[30] , \wRegInTop_7_93[29] , \wRegInTop_7_93[28] , 
        \wRegInTop_7_93[27] , \wRegInTop_7_93[26] , \wRegInTop_7_93[25] , 
        \wRegInTop_7_93[24] , \wRegInTop_7_93[23] , \wRegInTop_7_93[22] , 
        \wRegInTop_7_93[21] , \wRegInTop_7_93[20] , \wRegInTop_7_93[19] , 
        \wRegInTop_7_93[18] , \wRegInTop_7_93[17] , \wRegInTop_7_93[16] , 
        \wRegInTop_7_93[15] , \wRegInTop_7_93[14] , \wRegInTop_7_93[13] , 
        \wRegInTop_7_93[12] , \wRegInTop_7_93[11] , \wRegInTop_7_93[10] , 
        \wRegInTop_7_93[9] , \wRegInTop_7_93[8] , \wRegInTop_7_93[7] , 
        \wRegInTop_7_93[6] , \wRegInTop_7_93[5] , \wRegInTop_7_93[4] , 
        \wRegInTop_7_93[3] , \wRegInTop_7_93[2] , \wRegInTop_7_93[1] , 
        \wRegInTop_7_93[0] }) );
    BHeap_Node_WIDTH32 BHN_4_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_0[0] ), .P_In({\wRegOut_4_0[31] , 
        \wRegOut_4_0[30] , \wRegOut_4_0[29] , \wRegOut_4_0[28] , 
        \wRegOut_4_0[27] , \wRegOut_4_0[26] , \wRegOut_4_0[25] , 
        \wRegOut_4_0[24] , \wRegOut_4_0[23] , \wRegOut_4_0[22] , 
        \wRegOut_4_0[21] , \wRegOut_4_0[20] , \wRegOut_4_0[19] , 
        \wRegOut_4_0[18] , \wRegOut_4_0[17] , \wRegOut_4_0[16] , 
        \wRegOut_4_0[15] , \wRegOut_4_0[14] , \wRegOut_4_0[13] , 
        \wRegOut_4_0[12] , \wRegOut_4_0[11] , \wRegOut_4_0[10] , 
        \wRegOut_4_0[9] , \wRegOut_4_0[8] , \wRegOut_4_0[7] , \wRegOut_4_0[6] , 
        \wRegOut_4_0[5] , \wRegOut_4_0[4] , \wRegOut_4_0[3] , \wRegOut_4_0[2] , 
        \wRegOut_4_0[1] , \wRegOut_4_0[0] }), .P_Out({\wRegInBot_4_0[31] , 
        \wRegInBot_4_0[30] , \wRegInBot_4_0[29] , \wRegInBot_4_0[28] , 
        \wRegInBot_4_0[27] , \wRegInBot_4_0[26] , \wRegInBot_4_0[25] , 
        \wRegInBot_4_0[24] , \wRegInBot_4_0[23] , \wRegInBot_4_0[22] , 
        \wRegInBot_4_0[21] , \wRegInBot_4_0[20] , \wRegInBot_4_0[19] , 
        \wRegInBot_4_0[18] , \wRegInBot_4_0[17] , \wRegInBot_4_0[16] , 
        \wRegInBot_4_0[15] , \wRegInBot_4_0[14] , \wRegInBot_4_0[13] , 
        \wRegInBot_4_0[12] , \wRegInBot_4_0[11] , \wRegInBot_4_0[10] , 
        \wRegInBot_4_0[9] , \wRegInBot_4_0[8] , \wRegInBot_4_0[7] , 
        \wRegInBot_4_0[6] , \wRegInBot_4_0[5] , \wRegInBot_4_0[4] , 
        \wRegInBot_4_0[3] , \wRegInBot_4_0[2] , \wRegInBot_4_0[1] , 
        \wRegInBot_4_0[0] }), .L_WR(\wRegEnTop_5_0[0] ), .L_In({
        \wRegOut_5_0[31] , \wRegOut_5_0[30] , \wRegOut_5_0[29] , 
        \wRegOut_5_0[28] , \wRegOut_5_0[27] , \wRegOut_5_0[26] , 
        \wRegOut_5_0[25] , \wRegOut_5_0[24] , \wRegOut_5_0[23] , 
        \wRegOut_5_0[22] , \wRegOut_5_0[21] , \wRegOut_5_0[20] , 
        \wRegOut_5_0[19] , \wRegOut_5_0[18] , \wRegOut_5_0[17] , 
        \wRegOut_5_0[16] , \wRegOut_5_0[15] , \wRegOut_5_0[14] , 
        \wRegOut_5_0[13] , \wRegOut_5_0[12] , \wRegOut_5_0[11] , 
        \wRegOut_5_0[10] , \wRegOut_5_0[9] , \wRegOut_5_0[8] , 
        \wRegOut_5_0[7] , \wRegOut_5_0[6] , \wRegOut_5_0[5] , \wRegOut_5_0[4] , 
        \wRegOut_5_0[3] , \wRegOut_5_0[2] , \wRegOut_5_0[1] , \wRegOut_5_0[0] 
        }), .L_Out({\wRegInTop_5_0[31] , \wRegInTop_5_0[30] , 
        \wRegInTop_5_0[29] , \wRegInTop_5_0[28] , \wRegInTop_5_0[27] , 
        \wRegInTop_5_0[26] , \wRegInTop_5_0[25] , \wRegInTop_5_0[24] , 
        \wRegInTop_5_0[23] , \wRegInTop_5_0[22] , \wRegInTop_5_0[21] , 
        \wRegInTop_5_0[20] , \wRegInTop_5_0[19] , \wRegInTop_5_0[18] , 
        \wRegInTop_5_0[17] , \wRegInTop_5_0[16] , \wRegInTop_5_0[15] , 
        \wRegInTop_5_0[14] , \wRegInTop_5_0[13] , \wRegInTop_5_0[12] , 
        \wRegInTop_5_0[11] , \wRegInTop_5_0[10] , \wRegInTop_5_0[9] , 
        \wRegInTop_5_0[8] , \wRegInTop_5_0[7] , \wRegInTop_5_0[6] , 
        \wRegInTop_5_0[5] , \wRegInTop_5_0[4] , \wRegInTop_5_0[3] , 
        \wRegInTop_5_0[2] , \wRegInTop_5_0[1] , \wRegInTop_5_0[0] }), .R_WR(
        \wRegEnTop_5_1[0] ), .R_In({\wRegOut_5_1[31] , \wRegOut_5_1[30] , 
        \wRegOut_5_1[29] , \wRegOut_5_1[28] , \wRegOut_5_1[27] , 
        \wRegOut_5_1[26] , \wRegOut_5_1[25] , \wRegOut_5_1[24] , 
        \wRegOut_5_1[23] , \wRegOut_5_1[22] , \wRegOut_5_1[21] , 
        \wRegOut_5_1[20] , \wRegOut_5_1[19] , \wRegOut_5_1[18] , 
        \wRegOut_5_1[17] , \wRegOut_5_1[16] , \wRegOut_5_1[15] , 
        \wRegOut_5_1[14] , \wRegOut_5_1[13] , \wRegOut_5_1[12] , 
        \wRegOut_5_1[11] , \wRegOut_5_1[10] , \wRegOut_5_1[9] , 
        \wRegOut_5_1[8] , \wRegOut_5_1[7] , \wRegOut_5_1[6] , \wRegOut_5_1[5] , 
        \wRegOut_5_1[4] , \wRegOut_5_1[3] , \wRegOut_5_1[2] , \wRegOut_5_1[1] , 
        \wRegOut_5_1[0] }), .R_Out({\wRegInTop_5_1[31] , \wRegInTop_5_1[30] , 
        \wRegInTop_5_1[29] , \wRegInTop_5_1[28] , \wRegInTop_5_1[27] , 
        \wRegInTop_5_1[26] , \wRegInTop_5_1[25] , \wRegInTop_5_1[24] , 
        \wRegInTop_5_1[23] , \wRegInTop_5_1[22] , \wRegInTop_5_1[21] , 
        \wRegInTop_5_1[20] , \wRegInTop_5_1[19] , \wRegInTop_5_1[18] , 
        \wRegInTop_5_1[17] , \wRegInTop_5_1[16] , \wRegInTop_5_1[15] , 
        \wRegInTop_5_1[14] , \wRegInTop_5_1[13] , \wRegInTop_5_1[12] , 
        \wRegInTop_5_1[11] , \wRegInTop_5_1[10] , \wRegInTop_5_1[9] , 
        \wRegInTop_5_1[8] , \wRegInTop_5_1[7] , \wRegInTop_5_1[6] , 
        \wRegInTop_5_1[5] , \wRegInTop_5_1[4] , \wRegInTop_5_1[3] , 
        \wRegInTop_5_1[2] , \wRegInTop_5_1[1] , \wRegInTop_5_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_26 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink154[31] , \ScanLink154[30] , \ScanLink154[29] , 
        \ScanLink154[28] , \ScanLink154[27] , \ScanLink154[26] , 
        \ScanLink154[25] , \ScanLink154[24] , \ScanLink154[23] , 
        \ScanLink154[22] , \ScanLink154[21] , \ScanLink154[20] , 
        \ScanLink154[19] , \ScanLink154[18] , \ScanLink154[17] , 
        \ScanLink154[16] , \ScanLink154[15] , \ScanLink154[14] , 
        \ScanLink154[13] , \ScanLink154[12] , \ScanLink154[11] , 
        \ScanLink154[10] , \ScanLink154[9] , \ScanLink154[8] , 
        \ScanLink154[7] , \ScanLink154[6] , \ScanLink154[5] , \ScanLink154[4] , 
        \ScanLink154[3] , \ScanLink154[2] , \ScanLink154[1] , \ScanLink154[0] 
        }), .ScanOut({\ScanLink153[31] , \ScanLink153[30] , \ScanLink153[29] , 
        \ScanLink153[28] , \ScanLink153[27] , \ScanLink153[26] , 
        \ScanLink153[25] , \ScanLink153[24] , \ScanLink153[23] , 
        \ScanLink153[22] , \ScanLink153[21] , \ScanLink153[20] , 
        \ScanLink153[19] , \ScanLink153[18] , \ScanLink153[17] , 
        \ScanLink153[16] , \ScanLink153[15] , \ScanLink153[14] , 
        \ScanLink153[13] , \ScanLink153[12] , \ScanLink153[11] , 
        \ScanLink153[10] , \ScanLink153[9] , \ScanLink153[8] , 
        \ScanLink153[7] , \ScanLink153[6] , \ScanLink153[5] , \ScanLink153[4] , 
        \ScanLink153[3] , \ScanLink153[2] , \ScanLink153[1] , \ScanLink153[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_26[31] , 
        \wRegOut_7_26[30] , \wRegOut_7_26[29] , \wRegOut_7_26[28] , 
        \wRegOut_7_26[27] , \wRegOut_7_26[26] , \wRegOut_7_26[25] , 
        \wRegOut_7_26[24] , \wRegOut_7_26[23] , \wRegOut_7_26[22] , 
        \wRegOut_7_26[21] , \wRegOut_7_26[20] , \wRegOut_7_26[19] , 
        \wRegOut_7_26[18] , \wRegOut_7_26[17] , \wRegOut_7_26[16] , 
        \wRegOut_7_26[15] , \wRegOut_7_26[14] , \wRegOut_7_26[13] , 
        \wRegOut_7_26[12] , \wRegOut_7_26[11] , \wRegOut_7_26[10] , 
        \wRegOut_7_26[9] , \wRegOut_7_26[8] , \wRegOut_7_26[7] , 
        \wRegOut_7_26[6] , \wRegOut_7_26[5] , \wRegOut_7_26[4] , 
        \wRegOut_7_26[3] , \wRegOut_7_26[2] , \wRegOut_7_26[1] , 
        \wRegOut_7_26[0] }), .Enable1(\wRegEnTop_7_26[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_26[31] , \wRegInTop_7_26[30] , \wRegInTop_7_26[29] , 
        \wRegInTop_7_26[28] , \wRegInTop_7_26[27] , \wRegInTop_7_26[26] , 
        \wRegInTop_7_26[25] , \wRegInTop_7_26[24] , \wRegInTop_7_26[23] , 
        \wRegInTop_7_26[22] , \wRegInTop_7_26[21] , \wRegInTop_7_26[20] , 
        \wRegInTop_7_26[19] , \wRegInTop_7_26[18] , \wRegInTop_7_26[17] , 
        \wRegInTop_7_26[16] , \wRegInTop_7_26[15] , \wRegInTop_7_26[14] , 
        \wRegInTop_7_26[13] , \wRegInTop_7_26[12] , \wRegInTop_7_26[11] , 
        \wRegInTop_7_26[10] , \wRegInTop_7_26[9] , \wRegInTop_7_26[8] , 
        \wRegInTop_7_26[7] , \wRegInTop_7_26[6] , \wRegInTop_7_26[5] , 
        \wRegInTop_7_26[4] , \wRegInTop_7_26[3] , \wRegInTop_7_26[2] , 
        \wRegInTop_7_26[1] , \wRegInTop_7_26[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink71[31] , \ScanLink71[30] , \ScanLink71[29] , 
        \ScanLink71[28] , \ScanLink71[27] , \ScanLink71[26] , \ScanLink71[25] , 
        \ScanLink71[24] , \ScanLink71[23] , \ScanLink71[22] , \ScanLink71[21] , 
        \ScanLink71[20] , \ScanLink71[19] , \ScanLink71[18] , \ScanLink71[17] , 
        \ScanLink71[16] , \ScanLink71[15] , \ScanLink71[14] , \ScanLink71[13] , 
        \ScanLink71[12] , \ScanLink71[11] , \ScanLink71[10] , \ScanLink71[9] , 
        \ScanLink71[8] , \ScanLink71[7] , \ScanLink71[6] , \ScanLink71[5] , 
        \ScanLink71[4] , \ScanLink71[3] , \ScanLink71[2] , \ScanLink71[1] , 
        \ScanLink71[0] }), .ScanOut({\ScanLink70[31] , \ScanLink70[30] , 
        \ScanLink70[29] , \ScanLink70[28] , \ScanLink70[27] , \ScanLink70[26] , 
        \ScanLink70[25] , \ScanLink70[24] , \ScanLink70[23] , \ScanLink70[22] , 
        \ScanLink70[21] , \ScanLink70[20] , \ScanLink70[19] , \ScanLink70[18] , 
        \ScanLink70[17] , \ScanLink70[16] , \ScanLink70[15] , \ScanLink70[14] , 
        \ScanLink70[13] , \ScanLink70[12] , \ScanLink70[11] , \ScanLink70[10] , 
        \ScanLink70[9] , \ScanLink70[8] , \ScanLink70[7] , \ScanLink70[6] , 
        \ScanLink70[5] , \ScanLink70[4] , \ScanLink70[3] , \ScanLink70[2] , 
        \ScanLink70[1] , \ScanLink70[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_7[31] , \wRegOut_6_7[30] , \wRegOut_6_7[29] , 
        \wRegOut_6_7[28] , \wRegOut_6_7[27] , \wRegOut_6_7[26] , 
        \wRegOut_6_7[25] , \wRegOut_6_7[24] , \wRegOut_6_7[23] , 
        \wRegOut_6_7[22] , \wRegOut_6_7[21] , \wRegOut_6_7[20] , 
        \wRegOut_6_7[19] , \wRegOut_6_7[18] , \wRegOut_6_7[17] , 
        \wRegOut_6_7[16] , \wRegOut_6_7[15] , \wRegOut_6_7[14] , 
        \wRegOut_6_7[13] , \wRegOut_6_7[12] , \wRegOut_6_7[11] , 
        \wRegOut_6_7[10] , \wRegOut_6_7[9] , \wRegOut_6_7[8] , 
        \wRegOut_6_7[7] , \wRegOut_6_7[6] , \wRegOut_6_7[5] , \wRegOut_6_7[4] , 
        \wRegOut_6_7[3] , \wRegOut_6_7[2] , \wRegOut_6_7[1] , \wRegOut_6_7[0] 
        }), .Enable1(\wRegEnTop_6_7[0] ), .Enable2(\wRegEnBot_6_7[0] ), .In1({
        \wRegInTop_6_7[31] , \wRegInTop_6_7[30] , \wRegInTop_6_7[29] , 
        \wRegInTop_6_7[28] , \wRegInTop_6_7[27] , \wRegInTop_6_7[26] , 
        \wRegInTop_6_7[25] , \wRegInTop_6_7[24] , \wRegInTop_6_7[23] , 
        \wRegInTop_6_7[22] , \wRegInTop_6_7[21] , \wRegInTop_6_7[20] , 
        \wRegInTop_6_7[19] , \wRegInTop_6_7[18] , \wRegInTop_6_7[17] , 
        \wRegInTop_6_7[16] , \wRegInTop_6_7[15] , \wRegInTop_6_7[14] , 
        \wRegInTop_6_7[13] , \wRegInTop_6_7[12] , \wRegInTop_6_7[11] , 
        \wRegInTop_6_7[10] , \wRegInTop_6_7[9] , \wRegInTop_6_7[8] , 
        \wRegInTop_6_7[7] , \wRegInTop_6_7[6] , \wRegInTop_6_7[5] , 
        \wRegInTop_6_7[4] , \wRegInTop_6_7[3] , \wRegInTop_6_7[2] , 
        \wRegInTop_6_7[1] , \wRegInTop_6_7[0] }), .In2({\wRegInBot_6_7[31] , 
        \wRegInBot_6_7[30] , \wRegInBot_6_7[29] , \wRegInBot_6_7[28] , 
        \wRegInBot_6_7[27] , \wRegInBot_6_7[26] , \wRegInBot_6_7[25] , 
        \wRegInBot_6_7[24] , \wRegInBot_6_7[23] , \wRegInBot_6_7[22] , 
        \wRegInBot_6_7[21] , \wRegInBot_6_7[20] , \wRegInBot_6_7[19] , 
        \wRegInBot_6_7[18] , \wRegInBot_6_7[17] , \wRegInBot_6_7[16] , 
        \wRegInBot_6_7[15] , \wRegInBot_6_7[14] , \wRegInBot_6_7[13] , 
        \wRegInBot_6_7[12] , \wRegInBot_6_7[11] , \wRegInBot_6_7[10] , 
        \wRegInBot_6_7[9] , \wRegInBot_6_7[8] , \wRegInBot_6_7[7] , 
        \wRegInBot_6_7[6] , \wRegInBot_6_7[5] , \wRegInBot_6_7[4] , 
        \wRegInBot_6_7[3] , \wRegInBot_6_7[2] , \wRegInBot_6_7[1] , 
        \wRegInBot_6_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_48 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink176[31] , \ScanLink176[30] , \ScanLink176[29] , 
        \ScanLink176[28] , \ScanLink176[27] , \ScanLink176[26] , 
        \ScanLink176[25] , \ScanLink176[24] , \ScanLink176[23] , 
        \ScanLink176[22] , \ScanLink176[21] , \ScanLink176[20] , 
        \ScanLink176[19] , \ScanLink176[18] , \ScanLink176[17] , 
        \ScanLink176[16] , \ScanLink176[15] , \ScanLink176[14] , 
        \ScanLink176[13] , \ScanLink176[12] , \ScanLink176[11] , 
        \ScanLink176[10] , \ScanLink176[9] , \ScanLink176[8] , 
        \ScanLink176[7] , \ScanLink176[6] , \ScanLink176[5] , \ScanLink176[4] , 
        \ScanLink176[3] , \ScanLink176[2] , \ScanLink176[1] , \ScanLink176[0] 
        }), .ScanOut({\ScanLink175[31] , \ScanLink175[30] , \ScanLink175[29] , 
        \ScanLink175[28] , \ScanLink175[27] , \ScanLink175[26] , 
        \ScanLink175[25] , \ScanLink175[24] , \ScanLink175[23] , 
        \ScanLink175[22] , \ScanLink175[21] , \ScanLink175[20] , 
        \ScanLink175[19] , \ScanLink175[18] , \ScanLink175[17] , 
        \ScanLink175[16] , \ScanLink175[15] , \ScanLink175[14] , 
        \ScanLink175[13] , \ScanLink175[12] , \ScanLink175[11] , 
        \ScanLink175[10] , \ScanLink175[9] , \ScanLink175[8] , 
        \ScanLink175[7] , \ScanLink175[6] , \ScanLink175[5] , \ScanLink175[4] , 
        \ScanLink175[3] , \ScanLink175[2] , \ScanLink175[1] , \ScanLink175[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_48[31] , 
        \wRegOut_7_48[30] , \wRegOut_7_48[29] , \wRegOut_7_48[28] , 
        \wRegOut_7_48[27] , \wRegOut_7_48[26] , \wRegOut_7_48[25] , 
        \wRegOut_7_48[24] , \wRegOut_7_48[23] , \wRegOut_7_48[22] , 
        \wRegOut_7_48[21] , \wRegOut_7_48[20] , \wRegOut_7_48[19] , 
        \wRegOut_7_48[18] , \wRegOut_7_48[17] , \wRegOut_7_48[16] , 
        \wRegOut_7_48[15] , \wRegOut_7_48[14] , \wRegOut_7_48[13] , 
        \wRegOut_7_48[12] , \wRegOut_7_48[11] , \wRegOut_7_48[10] , 
        \wRegOut_7_48[9] , \wRegOut_7_48[8] , \wRegOut_7_48[7] , 
        \wRegOut_7_48[6] , \wRegOut_7_48[5] , \wRegOut_7_48[4] , 
        \wRegOut_7_48[3] , \wRegOut_7_48[2] , \wRegOut_7_48[1] , 
        \wRegOut_7_48[0] }), .Enable1(\wRegEnTop_7_48[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_48[31] , \wRegInTop_7_48[30] , \wRegInTop_7_48[29] , 
        \wRegInTop_7_48[28] , \wRegInTop_7_48[27] , \wRegInTop_7_48[26] , 
        \wRegInTop_7_48[25] , \wRegInTop_7_48[24] , \wRegInTop_7_48[23] , 
        \wRegInTop_7_48[22] , \wRegInTop_7_48[21] , \wRegInTop_7_48[20] , 
        \wRegInTop_7_48[19] , \wRegInTop_7_48[18] , \wRegInTop_7_48[17] , 
        \wRegInTop_7_48[16] , \wRegInTop_7_48[15] , \wRegInTop_7_48[14] , 
        \wRegInTop_7_48[13] , \wRegInTop_7_48[12] , \wRegInTop_7_48[11] , 
        \wRegInTop_7_48[10] , \wRegInTop_7_48[9] , \wRegInTop_7_48[8] , 
        \wRegInTop_7_48[7] , \wRegInTop_7_48[6] , \wRegInTop_7_48[5] , 
        \wRegInTop_7_48[4] , \wRegInTop_7_48[3] , \wRegInTop_7_48[2] , 
        \wRegInTop_7_48[1] , \wRegInTop_7_48[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_24[0] ), .P_In({\wRegOut_5_24[31] , 
        \wRegOut_5_24[30] , \wRegOut_5_24[29] , \wRegOut_5_24[28] , 
        \wRegOut_5_24[27] , \wRegOut_5_24[26] , \wRegOut_5_24[25] , 
        \wRegOut_5_24[24] , \wRegOut_5_24[23] , \wRegOut_5_24[22] , 
        \wRegOut_5_24[21] , \wRegOut_5_24[20] , \wRegOut_5_24[19] , 
        \wRegOut_5_24[18] , \wRegOut_5_24[17] , \wRegOut_5_24[16] , 
        \wRegOut_5_24[15] , \wRegOut_5_24[14] , \wRegOut_5_24[13] , 
        \wRegOut_5_24[12] , \wRegOut_5_24[11] , \wRegOut_5_24[10] , 
        \wRegOut_5_24[9] , \wRegOut_5_24[8] , \wRegOut_5_24[7] , 
        \wRegOut_5_24[6] , \wRegOut_5_24[5] , \wRegOut_5_24[4] , 
        \wRegOut_5_24[3] , \wRegOut_5_24[2] , \wRegOut_5_24[1] , 
        \wRegOut_5_24[0] }), .P_Out({\wRegInBot_5_24[31] , 
        \wRegInBot_5_24[30] , \wRegInBot_5_24[29] , \wRegInBot_5_24[28] , 
        \wRegInBot_5_24[27] , \wRegInBot_5_24[26] , \wRegInBot_5_24[25] , 
        \wRegInBot_5_24[24] , \wRegInBot_5_24[23] , \wRegInBot_5_24[22] , 
        \wRegInBot_5_24[21] , \wRegInBot_5_24[20] , \wRegInBot_5_24[19] , 
        \wRegInBot_5_24[18] , \wRegInBot_5_24[17] , \wRegInBot_5_24[16] , 
        \wRegInBot_5_24[15] , \wRegInBot_5_24[14] , \wRegInBot_5_24[13] , 
        \wRegInBot_5_24[12] , \wRegInBot_5_24[11] , \wRegInBot_5_24[10] , 
        \wRegInBot_5_24[9] , \wRegInBot_5_24[8] , \wRegInBot_5_24[7] , 
        \wRegInBot_5_24[6] , \wRegInBot_5_24[5] , \wRegInBot_5_24[4] , 
        \wRegInBot_5_24[3] , \wRegInBot_5_24[2] , \wRegInBot_5_24[1] , 
        \wRegInBot_5_24[0] }), .L_WR(\wRegEnTop_6_48[0] ), .L_In({
        \wRegOut_6_48[31] , \wRegOut_6_48[30] , \wRegOut_6_48[29] , 
        \wRegOut_6_48[28] , \wRegOut_6_48[27] , \wRegOut_6_48[26] , 
        \wRegOut_6_48[25] , \wRegOut_6_48[24] , \wRegOut_6_48[23] , 
        \wRegOut_6_48[22] , \wRegOut_6_48[21] , \wRegOut_6_48[20] , 
        \wRegOut_6_48[19] , \wRegOut_6_48[18] , \wRegOut_6_48[17] , 
        \wRegOut_6_48[16] , \wRegOut_6_48[15] , \wRegOut_6_48[14] , 
        \wRegOut_6_48[13] , \wRegOut_6_48[12] , \wRegOut_6_48[11] , 
        \wRegOut_6_48[10] , \wRegOut_6_48[9] , \wRegOut_6_48[8] , 
        \wRegOut_6_48[7] , \wRegOut_6_48[6] , \wRegOut_6_48[5] , 
        \wRegOut_6_48[4] , \wRegOut_6_48[3] , \wRegOut_6_48[2] , 
        \wRegOut_6_48[1] , \wRegOut_6_48[0] }), .L_Out({\wRegInTop_6_48[31] , 
        \wRegInTop_6_48[30] , \wRegInTop_6_48[29] , \wRegInTop_6_48[28] , 
        \wRegInTop_6_48[27] , \wRegInTop_6_48[26] , \wRegInTop_6_48[25] , 
        \wRegInTop_6_48[24] , \wRegInTop_6_48[23] , \wRegInTop_6_48[22] , 
        \wRegInTop_6_48[21] , \wRegInTop_6_48[20] , \wRegInTop_6_48[19] , 
        \wRegInTop_6_48[18] , \wRegInTop_6_48[17] , \wRegInTop_6_48[16] , 
        \wRegInTop_6_48[15] , \wRegInTop_6_48[14] , \wRegInTop_6_48[13] , 
        \wRegInTop_6_48[12] , \wRegInTop_6_48[11] , \wRegInTop_6_48[10] , 
        \wRegInTop_6_48[9] , \wRegInTop_6_48[8] , \wRegInTop_6_48[7] , 
        \wRegInTop_6_48[6] , \wRegInTop_6_48[5] , \wRegInTop_6_48[4] , 
        \wRegInTop_6_48[3] , \wRegInTop_6_48[2] , \wRegInTop_6_48[1] , 
        \wRegInTop_6_48[0] }), .R_WR(\wRegEnTop_6_49[0] ), .R_In({
        \wRegOut_6_49[31] , \wRegOut_6_49[30] , \wRegOut_6_49[29] , 
        \wRegOut_6_49[28] , \wRegOut_6_49[27] , \wRegOut_6_49[26] , 
        \wRegOut_6_49[25] , \wRegOut_6_49[24] , \wRegOut_6_49[23] , 
        \wRegOut_6_49[22] , \wRegOut_6_49[21] , \wRegOut_6_49[20] , 
        \wRegOut_6_49[19] , \wRegOut_6_49[18] , \wRegOut_6_49[17] , 
        \wRegOut_6_49[16] , \wRegOut_6_49[15] , \wRegOut_6_49[14] , 
        \wRegOut_6_49[13] , \wRegOut_6_49[12] , \wRegOut_6_49[11] , 
        \wRegOut_6_49[10] , \wRegOut_6_49[9] , \wRegOut_6_49[8] , 
        \wRegOut_6_49[7] , \wRegOut_6_49[6] , \wRegOut_6_49[5] , 
        \wRegOut_6_49[4] , \wRegOut_6_49[3] , \wRegOut_6_49[2] , 
        \wRegOut_6_49[1] , \wRegOut_6_49[0] }), .R_Out({\wRegInTop_6_49[31] , 
        \wRegInTop_6_49[30] , \wRegInTop_6_49[29] , \wRegInTop_6_49[28] , 
        \wRegInTop_6_49[27] , \wRegInTop_6_49[26] , \wRegInTop_6_49[25] , 
        \wRegInTop_6_49[24] , \wRegInTop_6_49[23] , \wRegInTop_6_49[22] , 
        \wRegInTop_6_49[21] , \wRegInTop_6_49[20] , \wRegInTop_6_49[19] , 
        \wRegInTop_6_49[18] , \wRegInTop_6_49[17] , \wRegInTop_6_49[16] , 
        \wRegInTop_6_49[15] , \wRegInTop_6_49[14] , \wRegInTop_6_49[13] , 
        \wRegInTop_6_49[12] , \wRegInTop_6_49[11] , \wRegInTop_6_49[10] , 
        \wRegInTop_6_49[9] , \wRegInTop_6_49[8] , \wRegInTop_6_49[7] , 
        \wRegInTop_6_49[6] , \wRegInTop_6_49[5] , \wRegInTop_6_49[4] , 
        \wRegInTop_6_49[3] , \wRegInTop_6_49[2] , \wRegInTop_6_49[1] , 
        \wRegInTop_6_49[0] }) );
    BHeap_Node_WIDTH32 BHN_5_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_11[0] ), .P_In({\wRegOut_5_11[31] , 
        \wRegOut_5_11[30] , \wRegOut_5_11[29] , \wRegOut_5_11[28] , 
        \wRegOut_5_11[27] , \wRegOut_5_11[26] , \wRegOut_5_11[25] , 
        \wRegOut_5_11[24] , \wRegOut_5_11[23] , \wRegOut_5_11[22] , 
        \wRegOut_5_11[21] , \wRegOut_5_11[20] , \wRegOut_5_11[19] , 
        \wRegOut_5_11[18] , \wRegOut_5_11[17] , \wRegOut_5_11[16] , 
        \wRegOut_5_11[15] , \wRegOut_5_11[14] , \wRegOut_5_11[13] , 
        \wRegOut_5_11[12] , \wRegOut_5_11[11] , \wRegOut_5_11[10] , 
        \wRegOut_5_11[9] , \wRegOut_5_11[8] , \wRegOut_5_11[7] , 
        \wRegOut_5_11[6] , \wRegOut_5_11[5] , \wRegOut_5_11[4] , 
        \wRegOut_5_11[3] , \wRegOut_5_11[2] , \wRegOut_5_11[1] , 
        \wRegOut_5_11[0] }), .P_Out({\wRegInBot_5_11[31] , 
        \wRegInBot_5_11[30] , \wRegInBot_5_11[29] , \wRegInBot_5_11[28] , 
        \wRegInBot_5_11[27] , \wRegInBot_5_11[26] , \wRegInBot_5_11[25] , 
        \wRegInBot_5_11[24] , \wRegInBot_5_11[23] , \wRegInBot_5_11[22] , 
        \wRegInBot_5_11[21] , \wRegInBot_5_11[20] , \wRegInBot_5_11[19] , 
        \wRegInBot_5_11[18] , \wRegInBot_5_11[17] , \wRegInBot_5_11[16] , 
        \wRegInBot_5_11[15] , \wRegInBot_5_11[14] , \wRegInBot_5_11[13] , 
        \wRegInBot_5_11[12] , \wRegInBot_5_11[11] , \wRegInBot_5_11[10] , 
        \wRegInBot_5_11[9] , \wRegInBot_5_11[8] , \wRegInBot_5_11[7] , 
        \wRegInBot_5_11[6] , \wRegInBot_5_11[5] , \wRegInBot_5_11[4] , 
        \wRegInBot_5_11[3] , \wRegInBot_5_11[2] , \wRegInBot_5_11[1] , 
        \wRegInBot_5_11[0] }), .L_WR(\wRegEnTop_6_22[0] ), .L_In({
        \wRegOut_6_22[31] , \wRegOut_6_22[30] , \wRegOut_6_22[29] , 
        \wRegOut_6_22[28] , \wRegOut_6_22[27] , \wRegOut_6_22[26] , 
        \wRegOut_6_22[25] , \wRegOut_6_22[24] , \wRegOut_6_22[23] , 
        \wRegOut_6_22[22] , \wRegOut_6_22[21] , \wRegOut_6_22[20] , 
        \wRegOut_6_22[19] , \wRegOut_6_22[18] , \wRegOut_6_22[17] , 
        \wRegOut_6_22[16] , \wRegOut_6_22[15] , \wRegOut_6_22[14] , 
        \wRegOut_6_22[13] , \wRegOut_6_22[12] , \wRegOut_6_22[11] , 
        \wRegOut_6_22[10] , \wRegOut_6_22[9] , \wRegOut_6_22[8] , 
        \wRegOut_6_22[7] , \wRegOut_6_22[6] , \wRegOut_6_22[5] , 
        \wRegOut_6_22[4] , \wRegOut_6_22[3] , \wRegOut_6_22[2] , 
        \wRegOut_6_22[1] , \wRegOut_6_22[0] }), .L_Out({\wRegInTop_6_22[31] , 
        \wRegInTop_6_22[30] , \wRegInTop_6_22[29] , \wRegInTop_6_22[28] , 
        \wRegInTop_6_22[27] , \wRegInTop_6_22[26] , \wRegInTop_6_22[25] , 
        \wRegInTop_6_22[24] , \wRegInTop_6_22[23] , \wRegInTop_6_22[22] , 
        \wRegInTop_6_22[21] , \wRegInTop_6_22[20] , \wRegInTop_6_22[19] , 
        \wRegInTop_6_22[18] , \wRegInTop_6_22[17] , \wRegInTop_6_22[16] , 
        \wRegInTop_6_22[15] , \wRegInTop_6_22[14] , \wRegInTop_6_22[13] , 
        \wRegInTop_6_22[12] , \wRegInTop_6_22[11] , \wRegInTop_6_22[10] , 
        \wRegInTop_6_22[9] , \wRegInTop_6_22[8] , \wRegInTop_6_22[7] , 
        \wRegInTop_6_22[6] , \wRegInTop_6_22[5] , \wRegInTop_6_22[4] , 
        \wRegInTop_6_22[3] , \wRegInTop_6_22[2] , \wRegInTop_6_22[1] , 
        \wRegInTop_6_22[0] }), .R_WR(\wRegEnTop_6_23[0] ), .R_In({
        \wRegOut_6_23[31] , \wRegOut_6_23[30] , \wRegOut_6_23[29] , 
        \wRegOut_6_23[28] , \wRegOut_6_23[27] , \wRegOut_6_23[26] , 
        \wRegOut_6_23[25] , \wRegOut_6_23[24] , \wRegOut_6_23[23] , 
        \wRegOut_6_23[22] , \wRegOut_6_23[21] , \wRegOut_6_23[20] , 
        \wRegOut_6_23[19] , \wRegOut_6_23[18] , \wRegOut_6_23[17] , 
        \wRegOut_6_23[16] , \wRegOut_6_23[15] , \wRegOut_6_23[14] , 
        \wRegOut_6_23[13] , \wRegOut_6_23[12] , \wRegOut_6_23[11] , 
        \wRegOut_6_23[10] , \wRegOut_6_23[9] , \wRegOut_6_23[8] , 
        \wRegOut_6_23[7] , \wRegOut_6_23[6] , \wRegOut_6_23[5] , 
        \wRegOut_6_23[4] , \wRegOut_6_23[3] , \wRegOut_6_23[2] , 
        \wRegOut_6_23[1] , \wRegOut_6_23[0] }), .R_Out({\wRegInTop_6_23[31] , 
        \wRegInTop_6_23[30] , \wRegInTop_6_23[29] , \wRegInTop_6_23[28] , 
        \wRegInTop_6_23[27] , \wRegInTop_6_23[26] , \wRegInTop_6_23[25] , 
        \wRegInTop_6_23[24] , \wRegInTop_6_23[23] , \wRegInTop_6_23[22] , 
        \wRegInTop_6_23[21] , \wRegInTop_6_23[20] , \wRegInTop_6_23[19] , 
        \wRegInTop_6_23[18] , \wRegInTop_6_23[17] , \wRegInTop_6_23[16] , 
        \wRegInTop_6_23[15] , \wRegInTop_6_23[14] , \wRegInTop_6_23[13] , 
        \wRegInTop_6_23[12] , \wRegInTop_6_23[11] , \wRegInTop_6_23[10] , 
        \wRegInTop_6_23[9] , \wRegInTop_6_23[8] , \wRegInTop_6_23[7] , 
        \wRegInTop_6_23[6] , \wRegInTop_6_23[5] , \wRegInTop_6_23[4] , 
        \wRegInTop_6_23[3] , \wRegInTop_6_23[2] , \wRegInTop_6_23[1] , 
        \wRegInTop_6_23[0] }) );
    BHeap_Node_WIDTH32 BHN_6_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_14[0] ), .P_In({\wRegOut_6_14[31] , 
        \wRegOut_6_14[30] , \wRegOut_6_14[29] , \wRegOut_6_14[28] , 
        \wRegOut_6_14[27] , \wRegOut_6_14[26] , \wRegOut_6_14[25] , 
        \wRegOut_6_14[24] , \wRegOut_6_14[23] , \wRegOut_6_14[22] , 
        \wRegOut_6_14[21] , \wRegOut_6_14[20] , \wRegOut_6_14[19] , 
        \wRegOut_6_14[18] , \wRegOut_6_14[17] , \wRegOut_6_14[16] , 
        \wRegOut_6_14[15] , \wRegOut_6_14[14] , \wRegOut_6_14[13] , 
        \wRegOut_6_14[12] , \wRegOut_6_14[11] , \wRegOut_6_14[10] , 
        \wRegOut_6_14[9] , \wRegOut_6_14[8] , \wRegOut_6_14[7] , 
        \wRegOut_6_14[6] , \wRegOut_6_14[5] , \wRegOut_6_14[4] , 
        \wRegOut_6_14[3] , \wRegOut_6_14[2] , \wRegOut_6_14[1] , 
        \wRegOut_6_14[0] }), .P_Out({\wRegInBot_6_14[31] , 
        \wRegInBot_6_14[30] , \wRegInBot_6_14[29] , \wRegInBot_6_14[28] , 
        \wRegInBot_6_14[27] , \wRegInBot_6_14[26] , \wRegInBot_6_14[25] , 
        \wRegInBot_6_14[24] , \wRegInBot_6_14[23] , \wRegInBot_6_14[22] , 
        \wRegInBot_6_14[21] , \wRegInBot_6_14[20] , \wRegInBot_6_14[19] , 
        \wRegInBot_6_14[18] , \wRegInBot_6_14[17] , \wRegInBot_6_14[16] , 
        \wRegInBot_6_14[15] , \wRegInBot_6_14[14] , \wRegInBot_6_14[13] , 
        \wRegInBot_6_14[12] , \wRegInBot_6_14[11] , \wRegInBot_6_14[10] , 
        \wRegInBot_6_14[9] , \wRegInBot_6_14[8] , \wRegInBot_6_14[7] , 
        \wRegInBot_6_14[6] , \wRegInBot_6_14[5] , \wRegInBot_6_14[4] , 
        \wRegInBot_6_14[3] , \wRegInBot_6_14[2] , \wRegInBot_6_14[1] , 
        \wRegInBot_6_14[0] }), .L_WR(\wRegEnTop_7_28[0] ), .L_In({
        \wRegOut_7_28[31] , \wRegOut_7_28[30] , \wRegOut_7_28[29] , 
        \wRegOut_7_28[28] , \wRegOut_7_28[27] , \wRegOut_7_28[26] , 
        \wRegOut_7_28[25] , \wRegOut_7_28[24] , \wRegOut_7_28[23] , 
        \wRegOut_7_28[22] , \wRegOut_7_28[21] , \wRegOut_7_28[20] , 
        \wRegOut_7_28[19] , \wRegOut_7_28[18] , \wRegOut_7_28[17] , 
        \wRegOut_7_28[16] , \wRegOut_7_28[15] , \wRegOut_7_28[14] , 
        \wRegOut_7_28[13] , \wRegOut_7_28[12] , \wRegOut_7_28[11] , 
        \wRegOut_7_28[10] , \wRegOut_7_28[9] , \wRegOut_7_28[8] , 
        \wRegOut_7_28[7] , \wRegOut_7_28[6] , \wRegOut_7_28[5] , 
        \wRegOut_7_28[4] , \wRegOut_7_28[3] , \wRegOut_7_28[2] , 
        \wRegOut_7_28[1] , \wRegOut_7_28[0] }), .L_Out({\wRegInTop_7_28[31] , 
        \wRegInTop_7_28[30] , \wRegInTop_7_28[29] , \wRegInTop_7_28[28] , 
        \wRegInTop_7_28[27] , \wRegInTop_7_28[26] , \wRegInTop_7_28[25] , 
        \wRegInTop_7_28[24] , \wRegInTop_7_28[23] , \wRegInTop_7_28[22] , 
        \wRegInTop_7_28[21] , \wRegInTop_7_28[20] , \wRegInTop_7_28[19] , 
        \wRegInTop_7_28[18] , \wRegInTop_7_28[17] , \wRegInTop_7_28[16] , 
        \wRegInTop_7_28[15] , \wRegInTop_7_28[14] , \wRegInTop_7_28[13] , 
        \wRegInTop_7_28[12] , \wRegInTop_7_28[11] , \wRegInTop_7_28[10] , 
        \wRegInTop_7_28[9] , \wRegInTop_7_28[8] , \wRegInTop_7_28[7] , 
        \wRegInTop_7_28[6] , \wRegInTop_7_28[5] , \wRegInTop_7_28[4] , 
        \wRegInTop_7_28[3] , \wRegInTop_7_28[2] , \wRegInTop_7_28[1] , 
        \wRegInTop_7_28[0] }), .R_WR(\wRegEnTop_7_29[0] ), .R_In({
        \wRegOut_7_29[31] , \wRegOut_7_29[30] , \wRegOut_7_29[29] , 
        \wRegOut_7_29[28] , \wRegOut_7_29[27] , \wRegOut_7_29[26] , 
        \wRegOut_7_29[25] , \wRegOut_7_29[24] , \wRegOut_7_29[23] , 
        \wRegOut_7_29[22] , \wRegOut_7_29[21] , \wRegOut_7_29[20] , 
        \wRegOut_7_29[19] , \wRegOut_7_29[18] , \wRegOut_7_29[17] , 
        \wRegOut_7_29[16] , \wRegOut_7_29[15] , \wRegOut_7_29[14] , 
        \wRegOut_7_29[13] , \wRegOut_7_29[12] , \wRegOut_7_29[11] , 
        \wRegOut_7_29[10] , \wRegOut_7_29[9] , \wRegOut_7_29[8] , 
        \wRegOut_7_29[7] , \wRegOut_7_29[6] , \wRegOut_7_29[5] , 
        \wRegOut_7_29[4] , \wRegOut_7_29[3] , \wRegOut_7_29[2] , 
        \wRegOut_7_29[1] , \wRegOut_7_29[0] }), .R_Out({\wRegInTop_7_29[31] , 
        \wRegInTop_7_29[30] , \wRegInTop_7_29[29] , \wRegInTop_7_29[28] , 
        \wRegInTop_7_29[27] , \wRegInTop_7_29[26] , \wRegInTop_7_29[25] , 
        \wRegInTop_7_29[24] , \wRegInTop_7_29[23] , \wRegInTop_7_29[22] , 
        \wRegInTop_7_29[21] , \wRegInTop_7_29[20] , \wRegInTop_7_29[19] , 
        \wRegInTop_7_29[18] , \wRegInTop_7_29[17] , \wRegInTop_7_29[16] , 
        \wRegInTop_7_29[15] , \wRegInTop_7_29[14] , \wRegInTop_7_29[13] , 
        \wRegInTop_7_29[12] , \wRegInTop_7_29[11] , \wRegInTop_7_29[10] , 
        \wRegInTop_7_29[9] , \wRegInTop_7_29[8] , \wRegInTop_7_29[7] , 
        \wRegInTop_7_29[6] , \wRegInTop_7_29[5] , \wRegInTop_7_29[4] , 
        \wRegInTop_7_29[3] , \wRegInTop_7_29[2] , \wRegInTop_7_29[1] , 
        \wRegInTop_7_29[0] }) );
    BHeap_Node_WIDTH32 BHN_6_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_33[0] ), .P_In({\wRegOut_6_33[31] , 
        \wRegOut_6_33[30] , \wRegOut_6_33[29] , \wRegOut_6_33[28] , 
        \wRegOut_6_33[27] , \wRegOut_6_33[26] , \wRegOut_6_33[25] , 
        \wRegOut_6_33[24] , \wRegOut_6_33[23] , \wRegOut_6_33[22] , 
        \wRegOut_6_33[21] , \wRegOut_6_33[20] , \wRegOut_6_33[19] , 
        \wRegOut_6_33[18] , \wRegOut_6_33[17] , \wRegOut_6_33[16] , 
        \wRegOut_6_33[15] , \wRegOut_6_33[14] , \wRegOut_6_33[13] , 
        \wRegOut_6_33[12] , \wRegOut_6_33[11] , \wRegOut_6_33[10] , 
        \wRegOut_6_33[9] , \wRegOut_6_33[8] , \wRegOut_6_33[7] , 
        \wRegOut_6_33[6] , \wRegOut_6_33[5] , \wRegOut_6_33[4] , 
        \wRegOut_6_33[3] , \wRegOut_6_33[2] , \wRegOut_6_33[1] , 
        \wRegOut_6_33[0] }), .P_Out({\wRegInBot_6_33[31] , 
        \wRegInBot_6_33[30] , \wRegInBot_6_33[29] , \wRegInBot_6_33[28] , 
        \wRegInBot_6_33[27] , \wRegInBot_6_33[26] , \wRegInBot_6_33[25] , 
        \wRegInBot_6_33[24] , \wRegInBot_6_33[23] , \wRegInBot_6_33[22] , 
        \wRegInBot_6_33[21] , \wRegInBot_6_33[20] , \wRegInBot_6_33[19] , 
        \wRegInBot_6_33[18] , \wRegInBot_6_33[17] , \wRegInBot_6_33[16] , 
        \wRegInBot_6_33[15] , \wRegInBot_6_33[14] , \wRegInBot_6_33[13] , 
        \wRegInBot_6_33[12] , \wRegInBot_6_33[11] , \wRegInBot_6_33[10] , 
        \wRegInBot_6_33[9] , \wRegInBot_6_33[8] , \wRegInBot_6_33[7] , 
        \wRegInBot_6_33[6] , \wRegInBot_6_33[5] , \wRegInBot_6_33[4] , 
        \wRegInBot_6_33[3] , \wRegInBot_6_33[2] , \wRegInBot_6_33[1] , 
        \wRegInBot_6_33[0] }), .L_WR(\wRegEnTop_7_66[0] ), .L_In({
        \wRegOut_7_66[31] , \wRegOut_7_66[30] , \wRegOut_7_66[29] , 
        \wRegOut_7_66[28] , \wRegOut_7_66[27] , \wRegOut_7_66[26] , 
        \wRegOut_7_66[25] , \wRegOut_7_66[24] , \wRegOut_7_66[23] , 
        \wRegOut_7_66[22] , \wRegOut_7_66[21] , \wRegOut_7_66[20] , 
        \wRegOut_7_66[19] , \wRegOut_7_66[18] , \wRegOut_7_66[17] , 
        \wRegOut_7_66[16] , \wRegOut_7_66[15] , \wRegOut_7_66[14] , 
        \wRegOut_7_66[13] , \wRegOut_7_66[12] , \wRegOut_7_66[11] , 
        \wRegOut_7_66[10] , \wRegOut_7_66[9] , \wRegOut_7_66[8] , 
        \wRegOut_7_66[7] , \wRegOut_7_66[6] , \wRegOut_7_66[5] , 
        \wRegOut_7_66[4] , \wRegOut_7_66[3] , \wRegOut_7_66[2] , 
        \wRegOut_7_66[1] , \wRegOut_7_66[0] }), .L_Out({\wRegInTop_7_66[31] , 
        \wRegInTop_7_66[30] , \wRegInTop_7_66[29] , \wRegInTop_7_66[28] , 
        \wRegInTop_7_66[27] , \wRegInTop_7_66[26] , \wRegInTop_7_66[25] , 
        \wRegInTop_7_66[24] , \wRegInTop_7_66[23] , \wRegInTop_7_66[22] , 
        \wRegInTop_7_66[21] , \wRegInTop_7_66[20] , \wRegInTop_7_66[19] , 
        \wRegInTop_7_66[18] , \wRegInTop_7_66[17] , \wRegInTop_7_66[16] , 
        \wRegInTop_7_66[15] , \wRegInTop_7_66[14] , \wRegInTop_7_66[13] , 
        \wRegInTop_7_66[12] , \wRegInTop_7_66[11] , \wRegInTop_7_66[10] , 
        \wRegInTop_7_66[9] , \wRegInTop_7_66[8] , \wRegInTop_7_66[7] , 
        \wRegInTop_7_66[6] , \wRegInTop_7_66[5] , \wRegInTop_7_66[4] , 
        \wRegInTop_7_66[3] , \wRegInTop_7_66[2] , \wRegInTop_7_66[1] , 
        \wRegInTop_7_66[0] }), .R_WR(\wRegEnTop_7_67[0] ), .R_In({
        \wRegOut_7_67[31] , \wRegOut_7_67[30] , \wRegOut_7_67[29] , 
        \wRegOut_7_67[28] , \wRegOut_7_67[27] , \wRegOut_7_67[26] , 
        \wRegOut_7_67[25] , \wRegOut_7_67[24] , \wRegOut_7_67[23] , 
        \wRegOut_7_67[22] , \wRegOut_7_67[21] , \wRegOut_7_67[20] , 
        \wRegOut_7_67[19] , \wRegOut_7_67[18] , \wRegOut_7_67[17] , 
        \wRegOut_7_67[16] , \wRegOut_7_67[15] , \wRegOut_7_67[14] , 
        \wRegOut_7_67[13] , \wRegOut_7_67[12] , \wRegOut_7_67[11] , 
        \wRegOut_7_67[10] , \wRegOut_7_67[9] , \wRegOut_7_67[8] , 
        \wRegOut_7_67[7] , \wRegOut_7_67[6] , \wRegOut_7_67[5] , 
        \wRegOut_7_67[4] , \wRegOut_7_67[3] , \wRegOut_7_67[2] , 
        \wRegOut_7_67[1] , \wRegOut_7_67[0] }), .R_Out({\wRegInTop_7_67[31] , 
        \wRegInTop_7_67[30] , \wRegInTop_7_67[29] , \wRegInTop_7_67[28] , 
        \wRegInTop_7_67[27] , \wRegInTop_7_67[26] , \wRegInTop_7_67[25] , 
        \wRegInTop_7_67[24] , \wRegInTop_7_67[23] , \wRegInTop_7_67[22] , 
        \wRegInTop_7_67[21] , \wRegInTop_7_67[20] , \wRegInTop_7_67[19] , 
        \wRegInTop_7_67[18] , \wRegInTop_7_67[17] , \wRegInTop_7_67[16] , 
        \wRegInTop_7_67[15] , \wRegInTop_7_67[14] , \wRegInTop_7_67[13] , 
        \wRegInTop_7_67[12] , \wRegInTop_7_67[11] , \wRegInTop_7_67[10] , 
        \wRegInTop_7_67[9] , \wRegInTop_7_67[8] , \wRegInTop_7_67[7] , 
        \wRegInTop_7_67[6] , \wRegInTop_7_67[5] , \wRegInTop_7_67[4] , 
        \wRegInTop_7_67[3] , \wRegInTop_7_67[2] , \wRegInTop_7_67[1] , 
        \wRegInTop_7_67[0] }) );
    BHeap_Node_WIDTH32 BHN_6_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_21[0] ), .P_In({\wRegOut_6_21[31] , 
        \wRegOut_6_21[30] , \wRegOut_6_21[29] , \wRegOut_6_21[28] , 
        \wRegOut_6_21[27] , \wRegOut_6_21[26] , \wRegOut_6_21[25] , 
        \wRegOut_6_21[24] , \wRegOut_6_21[23] , \wRegOut_6_21[22] , 
        \wRegOut_6_21[21] , \wRegOut_6_21[20] , \wRegOut_6_21[19] , 
        \wRegOut_6_21[18] , \wRegOut_6_21[17] , \wRegOut_6_21[16] , 
        \wRegOut_6_21[15] , \wRegOut_6_21[14] , \wRegOut_6_21[13] , 
        \wRegOut_6_21[12] , \wRegOut_6_21[11] , \wRegOut_6_21[10] , 
        \wRegOut_6_21[9] , \wRegOut_6_21[8] , \wRegOut_6_21[7] , 
        \wRegOut_6_21[6] , \wRegOut_6_21[5] , \wRegOut_6_21[4] , 
        \wRegOut_6_21[3] , \wRegOut_6_21[2] , \wRegOut_6_21[1] , 
        \wRegOut_6_21[0] }), .P_Out({\wRegInBot_6_21[31] , 
        \wRegInBot_6_21[30] , \wRegInBot_6_21[29] , \wRegInBot_6_21[28] , 
        \wRegInBot_6_21[27] , \wRegInBot_6_21[26] , \wRegInBot_6_21[25] , 
        \wRegInBot_6_21[24] , \wRegInBot_6_21[23] , \wRegInBot_6_21[22] , 
        \wRegInBot_6_21[21] , \wRegInBot_6_21[20] , \wRegInBot_6_21[19] , 
        \wRegInBot_6_21[18] , \wRegInBot_6_21[17] , \wRegInBot_6_21[16] , 
        \wRegInBot_6_21[15] , \wRegInBot_6_21[14] , \wRegInBot_6_21[13] , 
        \wRegInBot_6_21[12] , \wRegInBot_6_21[11] , \wRegInBot_6_21[10] , 
        \wRegInBot_6_21[9] , \wRegInBot_6_21[8] , \wRegInBot_6_21[7] , 
        \wRegInBot_6_21[6] , \wRegInBot_6_21[5] , \wRegInBot_6_21[4] , 
        \wRegInBot_6_21[3] , \wRegInBot_6_21[2] , \wRegInBot_6_21[1] , 
        \wRegInBot_6_21[0] }), .L_WR(\wRegEnTop_7_42[0] ), .L_In({
        \wRegOut_7_42[31] , \wRegOut_7_42[30] , \wRegOut_7_42[29] , 
        \wRegOut_7_42[28] , \wRegOut_7_42[27] , \wRegOut_7_42[26] , 
        \wRegOut_7_42[25] , \wRegOut_7_42[24] , \wRegOut_7_42[23] , 
        \wRegOut_7_42[22] , \wRegOut_7_42[21] , \wRegOut_7_42[20] , 
        \wRegOut_7_42[19] , \wRegOut_7_42[18] , \wRegOut_7_42[17] , 
        \wRegOut_7_42[16] , \wRegOut_7_42[15] , \wRegOut_7_42[14] , 
        \wRegOut_7_42[13] , \wRegOut_7_42[12] , \wRegOut_7_42[11] , 
        \wRegOut_7_42[10] , \wRegOut_7_42[9] , \wRegOut_7_42[8] , 
        \wRegOut_7_42[7] , \wRegOut_7_42[6] , \wRegOut_7_42[5] , 
        \wRegOut_7_42[4] , \wRegOut_7_42[3] , \wRegOut_7_42[2] , 
        \wRegOut_7_42[1] , \wRegOut_7_42[0] }), .L_Out({\wRegInTop_7_42[31] , 
        \wRegInTop_7_42[30] , \wRegInTop_7_42[29] , \wRegInTop_7_42[28] , 
        \wRegInTop_7_42[27] , \wRegInTop_7_42[26] , \wRegInTop_7_42[25] , 
        \wRegInTop_7_42[24] , \wRegInTop_7_42[23] , \wRegInTop_7_42[22] , 
        \wRegInTop_7_42[21] , \wRegInTop_7_42[20] , \wRegInTop_7_42[19] , 
        \wRegInTop_7_42[18] , \wRegInTop_7_42[17] , \wRegInTop_7_42[16] , 
        \wRegInTop_7_42[15] , \wRegInTop_7_42[14] , \wRegInTop_7_42[13] , 
        \wRegInTop_7_42[12] , \wRegInTop_7_42[11] , \wRegInTop_7_42[10] , 
        \wRegInTop_7_42[9] , \wRegInTop_7_42[8] , \wRegInTop_7_42[7] , 
        \wRegInTop_7_42[6] , \wRegInTop_7_42[5] , \wRegInTop_7_42[4] , 
        \wRegInTop_7_42[3] , \wRegInTop_7_42[2] , \wRegInTop_7_42[1] , 
        \wRegInTop_7_42[0] }), .R_WR(\wRegEnTop_7_43[0] ), .R_In({
        \wRegOut_7_43[31] , \wRegOut_7_43[30] , \wRegOut_7_43[29] , 
        \wRegOut_7_43[28] , \wRegOut_7_43[27] , \wRegOut_7_43[26] , 
        \wRegOut_7_43[25] , \wRegOut_7_43[24] , \wRegOut_7_43[23] , 
        \wRegOut_7_43[22] , \wRegOut_7_43[21] , \wRegOut_7_43[20] , 
        \wRegOut_7_43[19] , \wRegOut_7_43[18] , \wRegOut_7_43[17] , 
        \wRegOut_7_43[16] , \wRegOut_7_43[15] , \wRegOut_7_43[14] , 
        \wRegOut_7_43[13] , \wRegOut_7_43[12] , \wRegOut_7_43[11] , 
        \wRegOut_7_43[10] , \wRegOut_7_43[9] , \wRegOut_7_43[8] , 
        \wRegOut_7_43[7] , \wRegOut_7_43[6] , \wRegOut_7_43[5] , 
        \wRegOut_7_43[4] , \wRegOut_7_43[3] , \wRegOut_7_43[2] , 
        \wRegOut_7_43[1] , \wRegOut_7_43[0] }), .R_Out({\wRegInTop_7_43[31] , 
        \wRegInTop_7_43[30] , \wRegInTop_7_43[29] , \wRegInTop_7_43[28] , 
        \wRegInTop_7_43[27] , \wRegInTop_7_43[26] , \wRegInTop_7_43[25] , 
        \wRegInTop_7_43[24] , \wRegInTop_7_43[23] , \wRegInTop_7_43[22] , 
        \wRegInTop_7_43[21] , \wRegInTop_7_43[20] , \wRegInTop_7_43[19] , 
        \wRegInTop_7_43[18] , \wRegInTop_7_43[17] , \wRegInTop_7_43[16] , 
        \wRegInTop_7_43[15] , \wRegInTop_7_43[14] , \wRegInTop_7_43[13] , 
        \wRegInTop_7_43[12] , \wRegInTop_7_43[11] , \wRegInTop_7_43[10] , 
        \wRegInTop_7_43[9] , \wRegInTop_7_43[8] , \wRegInTop_7_43[7] , 
        \wRegInTop_7_43[6] , \wRegInTop_7_43[5] , \wRegInTop_7_43[4] , 
        \wRegInTop_7_43[3] , \wRegInTop_7_43[2] , \wRegInTop_7_43[1] , 
        \wRegInTop_7_43[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_40 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink104[31] , \ScanLink104[30] , \ScanLink104[29] , 
        \ScanLink104[28] , \ScanLink104[27] , \ScanLink104[26] , 
        \ScanLink104[25] , \ScanLink104[24] , \ScanLink104[23] , 
        \ScanLink104[22] , \ScanLink104[21] , \ScanLink104[20] , 
        \ScanLink104[19] , \ScanLink104[18] , \ScanLink104[17] , 
        \ScanLink104[16] , \ScanLink104[15] , \ScanLink104[14] , 
        \ScanLink104[13] , \ScanLink104[12] , \ScanLink104[11] , 
        \ScanLink104[10] , \ScanLink104[9] , \ScanLink104[8] , 
        \ScanLink104[7] , \ScanLink104[6] , \ScanLink104[5] , \ScanLink104[4] , 
        \ScanLink104[3] , \ScanLink104[2] , \ScanLink104[1] , \ScanLink104[0] 
        }), .ScanOut({\ScanLink103[31] , \ScanLink103[30] , \ScanLink103[29] , 
        \ScanLink103[28] , \ScanLink103[27] , \ScanLink103[26] , 
        \ScanLink103[25] , \ScanLink103[24] , \ScanLink103[23] , 
        \ScanLink103[22] , \ScanLink103[21] , \ScanLink103[20] , 
        \ScanLink103[19] , \ScanLink103[18] , \ScanLink103[17] , 
        \ScanLink103[16] , \ScanLink103[15] , \ScanLink103[14] , 
        \ScanLink103[13] , \ScanLink103[12] , \ScanLink103[11] , 
        \ScanLink103[10] , \ScanLink103[9] , \ScanLink103[8] , 
        \ScanLink103[7] , \ScanLink103[6] , \ScanLink103[5] , \ScanLink103[4] , 
        \ScanLink103[3] , \ScanLink103[2] , \ScanLink103[1] , \ScanLink103[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_40[31] , 
        \wRegOut_6_40[30] , \wRegOut_6_40[29] , \wRegOut_6_40[28] , 
        \wRegOut_6_40[27] , \wRegOut_6_40[26] , \wRegOut_6_40[25] , 
        \wRegOut_6_40[24] , \wRegOut_6_40[23] , \wRegOut_6_40[22] , 
        \wRegOut_6_40[21] , \wRegOut_6_40[20] , \wRegOut_6_40[19] , 
        \wRegOut_6_40[18] , \wRegOut_6_40[17] , \wRegOut_6_40[16] , 
        \wRegOut_6_40[15] , \wRegOut_6_40[14] , \wRegOut_6_40[13] , 
        \wRegOut_6_40[12] , \wRegOut_6_40[11] , \wRegOut_6_40[10] , 
        \wRegOut_6_40[9] , \wRegOut_6_40[8] , \wRegOut_6_40[7] , 
        \wRegOut_6_40[6] , \wRegOut_6_40[5] , \wRegOut_6_40[4] , 
        \wRegOut_6_40[3] , \wRegOut_6_40[2] , \wRegOut_6_40[1] , 
        \wRegOut_6_40[0] }), .Enable1(\wRegEnTop_6_40[0] ), .Enable2(
        \wRegEnBot_6_40[0] ), .In1({\wRegInTop_6_40[31] , \wRegInTop_6_40[30] , 
        \wRegInTop_6_40[29] , \wRegInTop_6_40[28] , \wRegInTop_6_40[27] , 
        \wRegInTop_6_40[26] , \wRegInTop_6_40[25] , \wRegInTop_6_40[24] , 
        \wRegInTop_6_40[23] , \wRegInTop_6_40[22] , \wRegInTop_6_40[21] , 
        \wRegInTop_6_40[20] , \wRegInTop_6_40[19] , \wRegInTop_6_40[18] , 
        \wRegInTop_6_40[17] , \wRegInTop_6_40[16] , \wRegInTop_6_40[15] , 
        \wRegInTop_6_40[14] , \wRegInTop_6_40[13] , \wRegInTop_6_40[12] , 
        \wRegInTop_6_40[11] , \wRegInTop_6_40[10] , \wRegInTop_6_40[9] , 
        \wRegInTop_6_40[8] , \wRegInTop_6_40[7] , \wRegInTop_6_40[6] , 
        \wRegInTop_6_40[5] , \wRegInTop_6_40[4] , \wRegInTop_6_40[3] , 
        \wRegInTop_6_40[2] , \wRegInTop_6_40[1] , \wRegInTop_6_40[0] }), .In2(
        {\wRegInBot_6_40[31] , \wRegInBot_6_40[30] , \wRegInBot_6_40[29] , 
        \wRegInBot_6_40[28] , \wRegInBot_6_40[27] , \wRegInBot_6_40[26] , 
        \wRegInBot_6_40[25] , \wRegInBot_6_40[24] , \wRegInBot_6_40[23] , 
        \wRegInBot_6_40[22] , \wRegInBot_6_40[21] , \wRegInBot_6_40[20] , 
        \wRegInBot_6_40[19] , \wRegInBot_6_40[18] , \wRegInBot_6_40[17] , 
        \wRegInBot_6_40[16] , \wRegInBot_6_40[15] , \wRegInBot_6_40[14] , 
        \wRegInBot_6_40[13] , \wRegInBot_6_40[12] , \wRegInBot_6_40[11] , 
        \wRegInBot_6_40[10] , \wRegInBot_6_40[9] , \wRegInBot_6_40[8] , 
        \wRegInBot_6_40[7] , \wRegInBot_6_40[6] , \wRegInBot_6_40[5] , 
        \wRegInBot_6_40[4] , \wRegInBot_6_40[3] , \wRegInBot_6_40[2] , 
        \wRegInBot_6_40[1] , \wRegInBot_6_40[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink141[31] , \ScanLink141[30] , \ScanLink141[29] , 
        \ScanLink141[28] , \ScanLink141[27] , \ScanLink141[26] , 
        \ScanLink141[25] , \ScanLink141[24] , \ScanLink141[23] , 
        \ScanLink141[22] , \ScanLink141[21] , \ScanLink141[20] , 
        \ScanLink141[19] , \ScanLink141[18] , \ScanLink141[17] , 
        \ScanLink141[16] , \ScanLink141[15] , \ScanLink141[14] , 
        \ScanLink141[13] , \ScanLink141[12] , \ScanLink141[11] , 
        \ScanLink141[10] , \ScanLink141[9] , \ScanLink141[8] , 
        \ScanLink141[7] , \ScanLink141[6] , \ScanLink141[5] , \ScanLink141[4] , 
        \ScanLink141[3] , \ScanLink141[2] , \ScanLink141[1] , \ScanLink141[0] 
        }), .ScanOut({\ScanLink140[31] , \ScanLink140[30] , \ScanLink140[29] , 
        \ScanLink140[28] , \ScanLink140[27] , \ScanLink140[26] , 
        \ScanLink140[25] , \ScanLink140[24] , \ScanLink140[23] , 
        \ScanLink140[22] , \ScanLink140[21] , \ScanLink140[20] , 
        \ScanLink140[19] , \ScanLink140[18] , \ScanLink140[17] , 
        \ScanLink140[16] , \ScanLink140[15] , \ScanLink140[14] , 
        \ScanLink140[13] , \ScanLink140[12] , \ScanLink140[11] , 
        \ScanLink140[10] , \ScanLink140[9] , \ScanLink140[8] , 
        \ScanLink140[7] , \ScanLink140[6] , \ScanLink140[5] , \ScanLink140[4] , 
        \ScanLink140[3] , \ScanLink140[2] , \ScanLink140[1] , \ScanLink140[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_13[31] , 
        \wRegOut_7_13[30] , \wRegOut_7_13[29] , \wRegOut_7_13[28] , 
        \wRegOut_7_13[27] , \wRegOut_7_13[26] , \wRegOut_7_13[25] , 
        \wRegOut_7_13[24] , \wRegOut_7_13[23] , \wRegOut_7_13[22] , 
        \wRegOut_7_13[21] , \wRegOut_7_13[20] , \wRegOut_7_13[19] , 
        \wRegOut_7_13[18] , \wRegOut_7_13[17] , \wRegOut_7_13[16] , 
        \wRegOut_7_13[15] , \wRegOut_7_13[14] , \wRegOut_7_13[13] , 
        \wRegOut_7_13[12] , \wRegOut_7_13[11] , \wRegOut_7_13[10] , 
        \wRegOut_7_13[9] , \wRegOut_7_13[8] , \wRegOut_7_13[7] , 
        \wRegOut_7_13[6] , \wRegOut_7_13[5] , \wRegOut_7_13[4] , 
        \wRegOut_7_13[3] , \wRegOut_7_13[2] , \wRegOut_7_13[1] , 
        \wRegOut_7_13[0] }), .Enable1(\wRegEnTop_7_13[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_13[31] , \wRegInTop_7_13[30] , \wRegInTop_7_13[29] , 
        \wRegInTop_7_13[28] , \wRegInTop_7_13[27] , \wRegInTop_7_13[26] , 
        \wRegInTop_7_13[25] , \wRegInTop_7_13[24] , \wRegInTop_7_13[23] , 
        \wRegInTop_7_13[22] , \wRegInTop_7_13[21] , \wRegInTop_7_13[20] , 
        \wRegInTop_7_13[19] , \wRegInTop_7_13[18] , \wRegInTop_7_13[17] , 
        \wRegInTop_7_13[16] , \wRegInTop_7_13[15] , \wRegInTop_7_13[14] , 
        \wRegInTop_7_13[13] , \wRegInTop_7_13[12] , \wRegInTop_7_13[11] , 
        \wRegInTop_7_13[10] , \wRegInTop_7_13[9] , \wRegInTop_7_13[8] , 
        \wRegInTop_7_13[7] , \wRegInTop_7_13[6] , \wRegInTop_7_13[5] , 
        \wRegInTop_7_13[4] , \wRegInTop_7_13[3] , \wRegInTop_7_13[2] , 
        \wRegInTop_7_13[1] , \wRegInTop_7_13[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_98 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink226[31] , \ScanLink226[30] , \ScanLink226[29] , 
        \ScanLink226[28] , \ScanLink226[27] , \ScanLink226[26] , 
        \ScanLink226[25] , \ScanLink226[24] , \ScanLink226[23] , 
        \ScanLink226[22] , \ScanLink226[21] , \ScanLink226[20] , 
        \ScanLink226[19] , \ScanLink226[18] , \ScanLink226[17] , 
        \ScanLink226[16] , \ScanLink226[15] , \ScanLink226[14] , 
        \ScanLink226[13] , \ScanLink226[12] , \ScanLink226[11] , 
        \ScanLink226[10] , \ScanLink226[9] , \ScanLink226[8] , 
        \ScanLink226[7] , \ScanLink226[6] , \ScanLink226[5] , \ScanLink226[4] , 
        \ScanLink226[3] , \ScanLink226[2] , \ScanLink226[1] , \ScanLink226[0] 
        }), .ScanOut({\ScanLink225[31] , \ScanLink225[30] , \ScanLink225[29] , 
        \ScanLink225[28] , \ScanLink225[27] , \ScanLink225[26] , 
        \ScanLink225[25] , \ScanLink225[24] , \ScanLink225[23] , 
        \ScanLink225[22] , \ScanLink225[21] , \ScanLink225[20] , 
        \ScanLink225[19] , \ScanLink225[18] , \ScanLink225[17] , 
        \ScanLink225[16] , \ScanLink225[15] , \ScanLink225[14] , 
        \ScanLink225[13] , \ScanLink225[12] , \ScanLink225[11] , 
        \ScanLink225[10] , \ScanLink225[9] , \ScanLink225[8] , 
        \ScanLink225[7] , \ScanLink225[6] , \ScanLink225[5] , \ScanLink225[4] , 
        \ScanLink225[3] , \ScanLink225[2] , \ScanLink225[1] , \ScanLink225[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_98[31] , 
        \wRegOut_7_98[30] , \wRegOut_7_98[29] , \wRegOut_7_98[28] , 
        \wRegOut_7_98[27] , \wRegOut_7_98[26] , \wRegOut_7_98[25] , 
        \wRegOut_7_98[24] , \wRegOut_7_98[23] , \wRegOut_7_98[22] , 
        \wRegOut_7_98[21] , \wRegOut_7_98[20] , \wRegOut_7_98[19] , 
        \wRegOut_7_98[18] , \wRegOut_7_98[17] , \wRegOut_7_98[16] , 
        \wRegOut_7_98[15] , \wRegOut_7_98[14] , \wRegOut_7_98[13] , 
        \wRegOut_7_98[12] , \wRegOut_7_98[11] , \wRegOut_7_98[10] , 
        \wRegOut_7_98[9] , \wRegOut_7_98[8] , \wRegOut_7_98[7] , 
        \wRegOut_7_98[6] , \wRegOut_7_98[5] , \wRegOut_7_98[4] , 
        \wRegOut_7_98[3] , \wRegOut_7_98[2] , \wRegOut_7_98[1] , 
        \wRegOut_7_98[0] }), .Enable1(\wRegEnTop_7_98[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_98[31] , \wRegInTop_7_98[30] , \wRegInTop_7_98[29] , 
        \wRegInTop_7_98[28] , \wRegInTop_7_98[27] , \wRegInTop_7_98[26] , 
        \wRegInTop_7_98[25] , \wRegInTop_7_98[24] , \wRegInTop_7_98[23] , 
        \wRegInTop_7_98[22] , \wRegInTop_7_98[21] , \wRegInTop_7_98[20] , 
        \wRegInTop_7_98[19] , \wRegInTop_7_98[18] , \wRegInTop_7_98[17] , 
        \wRegInTop_7_98[16] , \wRegInTop_7_98[15] , \wRegInTop_7_98[14] , 
        \wRegInTop_7_98[13] , \wRegInTop_7_98[12] , \wRegInTop_7_98[11] , 
        \wRegInTop_7_98[10] , \wRegInTop_7_98[9] , \wRegInTop_7_98[8] , 
        \wRegInTop_7_98[7] , \wRegInTop_7_98[6] , \wRegInTop_7_98[5] , 
        \wRegInTop_7_98[4] , \wRegInTop_7_98[3] , \wRegInTop_7_98[2] , 
        \wRegInTop_7_98[1] , \wRegInTop_7_98[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_107 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink235[31] , \ScanLink235[30] , \ScanLink235[29] , 
        \ScanLink235[28] , \ScanLink235[27] , \ScanLink235[26] , 
        \ScanLink235[25] , \ScanLink235[24] , \ScanLink235[23] , 
        \ScanLink235[22] , \ScanLink235[21] , \ScanLink235[20] , 
        \ScanLink235[19] , \ScanLink235[18] , \ScanLink235[17] , 
        \ScanLink235[16] , \ScanLink235[15] , \ScanLink235[14] , 
        \ScanLink235[13] , \ScanLink235[12] , \ScanLink235[11] , 
        \ScanLink235[10] , \ScanLink235[9] , \ScanLink235[8] , 
        \ScanLink235[7] , \ScanLink235[6] , \ScanLink235[5] , \ScanLink235[4] , 
        \ScanLink235[3] , \ScanLink235[2] , \ScanLink235[1] , \ScanLink235[0] 
        }), .ScanOut({\ScanLink234[31] , \ScanLink234[30] , \ScanLink234[29] , 
        \ScanLink234[28] , \ScanLink234[27] , \ScanLink234[26] , 
        \ScanLink234[25] , \ScanLink234[24] , \ScanLink234[23] , 
        \ScanLink234[22] , \ScanLink234[21] , \ScanLink234[20] , 
        \ScanLink234[19] , \ScanLink234[18] , \ScanLink234[17] , 
        \ScanLink234[16] , \ScanLink234[15] , \ScanLink234[14] , 
        \ScanLink234[13] , \ScanLink234[12] , \ScanLink234[11] , 
        \ScanLink234[10] , \ScanLink234[9] , \ScanLink234[8] , 
        \ScanLink234[7] , \ScanLink234[6] , \ScanLink234[5] , \ScanLink234[4] , 
        \ScanLink234[3] , \ScanLink234[2] , \ScanLink234[1] , \ScanLink234[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_107[31] , 
        \wRegOut_7_107[30] , \wRegOut_7_107[29] , \wRegOut_7_107[28] , 
        \wRegOut_7_107[27] , \wRegOut_7_107[26] , \wRegOut_7_107[25] , 
        \wRegOut_7_107[24] , \wRegOut_7_107[23] , \wRegOut_7_107[22] , 
        \wRegOut_7_107[21] , \wRegOut_7_107[20] , \wRegOut_7_107[19] , 
        \wRegOut_7_107[18] , \wRegOut_7_107[17] , \wRegOut_7_107[16] , 
        \wRegOut_7_107[15] , \wRegOut_7_107[14] , \wRegOut_7_107[13] , 
        \wRegOut_7_107[12] , \wRegOut_7_107[11] , \wRegOut_7_107[10] , 
        \wRegOut_7_107[9] , \wRegOut_7_107[8] , \wRegOut_7_107[7] , 
        \wRegOut_7_107[6] , \wRegOut_7_107[5] , \wRegOut_7_107[4] , 
        \wRegOut_7_107[3] , \wRegOut_7_107[2] , \wRegOut_7_107[1] , 
        \wRegOut_7_107[0] }), .Enable1(\wRegEnTop_7_107[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_107[31] , \wRegInTop_7_107[30] , 
        \wRegInTop_7_107[29] , \wRegInTop_7_107[28] , \wRegInTop_7_107[27] , 
        \wRegInTop_7_107[26] , \wRegInTop_7_107[25] , \wRegInTop_7_107[24] , 
        \wRegInTop_7_107[23] , \wRegInTop_7_107[22] , \wRegInTop_7_107[21] , 
        \wRegInTop_7_107[20] , \wRegInTop_7_107[19] , \wRegInTop_7_107[18] , 
        \wRegInTop_7_107[17] , \wRegInTop_7_107[16] , \wRegInTop_7_107[15] , 
        \wRegInTop_7_107[14] , \wRegInTop_7_107[13] , \wRegInTop_7_107[12] , 
        \wRegInTop_7_107[11] , \wRegInTop_7_107[10] , \wRegInTop_7_107[9] , 
        \wRegInTop_7_107[8] , \wRegInTop_7_107[7] , \wRegInTop_7_107[6] , 
        \wRegInTop_7_107[5] , \wRegInTop_7_107[4] , \wRegInTop_7_107[3] , 
        \wRegInTop_7_107[2] , \wRegInTop_7_107[1] , \wRegInTop_7_107[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_9[0] ), .P_In({\wRegOut_5_9[31] , 
        \wRegOut_5_9[30] , \wRegOut_5_9[29] , \wRegOut_5_9[28] , 
        \wRegOut_5_9[27] , \wRegOut_5_9[26] , \wRegOut_5_9[25] , 
        \wRegOut_5_9[24] , \wRegOut_5_9[23] , \wRegOut_5_9[22] , 
        \wRegOut_5_9[21] , \wRegOut_5_9[20] , \wRegOut_5_9[19] , 
        \wRegOut_5_9[18] , \wRegOut_5_9[17] , \wRegOut_5_9[16] , 
        \wRegOut_5_9[15] , \wRegOut_5_9[14] , \wRegOut_5_9[13] , 
        \wRegOut_5_9[12] , \wRegOut_5_9[11] , \wRegOut_5_9[10] , 
        \wRegOut_5_9[9] , \wRegOut_5_9[8] , \wRegOut_5_9[7] , \wRegOut_5_9[6] , 
        \wRegOut_5_9[5] , \wRegOut_5_9[4] , \wRegOut_5_9[3] , \wRegOut_5_9[2] , 
        \wRegOut_5_9[1] , \wRegOut_5_9[0] }), .P_Out({\wRegInBot_5_9[31] , 
        \wRegInBot_5_9[30] , \wRegInBot_5_9[29] , \wRegInBot_5_9[28] , 
        \wRegInBot_5_9[27] , \wRegInBot_5_9[26] , \wRegInBot_5_9[25] , 
        \wRegInBot_5_9[24] , \wRegInBot_5_9[23] , \wRegInBot_5_9[22] , 
        \wRegInBot_5_9[21] , \wRegInBot_5_9[20] , \wRegInBot_5_9[19] , 
        \wRegInBot_5_9[18] , \wRegInBot_5_9[17] , \wRegInBot_5_9[16] , 
        \wRegInBot_5_9[15] , \wRegInBot_5_9[14] , \wRegInBot_5_9[13] , 
        \wRegInBot_5_9[12] , \wRegInBot_5_9[11] , \wRegInBot_5_9[10] , 
        \wRegInBot_5_9[9] , \wRegInBot_5_9[8] , \wRegInBot_5_9[7] , 
        \wRegInBot_5_9[6] , \wRegInBot_5_9[5] , \wRegInBot_5_9[4] , 
        \wRegInBot_5_9[3] , \wRegInBot_5_9[2] , \wRegInBot_5_9[1] , 
        \wRegInBot_5_9[0] }), .L_WR(\wRegEnTop_6_18[0] ), .L_In({
        \wRegOut_6_18[31] , \wRegOut_6_18[30] , \wRegOut_6_18[29] , 
        \wRegOut_6_18[28] , \wRegOut_6_18[27] , \wRegOut_6_18[26] , 
        \wRegOut_6_18[25] , \wRegOut_6_18[24] , \wRegOut_6_18[23] , 
        \wRegOut_6_18[22] , \wRegOut_6_18[21] , \wRegOut_6_18[20] , 
        \wRegOut_6_18[19] , \wRegOut_6_18[18] , \wRegOut_6_18[17] , 
        \wRegOut_6_18[16] , \wRegOut_6_18[15] , \wRegOut_6_18[14] , 
        \wRegOut_6_18[13] , \wRegOut_6_18[12] , \wRegOut_6_18[11] , 
        \wRegOut_6_18[10] , \wRegOut_6_18[9] , \wRegOut_6_18[8] , 
        \wRegOut_6_18[7] , \wRegOut_6_18[6] , \wRegOut_6_18[5] , 
        \wRegOut_6_18[4] , \wRegOut_6_18[3] , \wRegOut_6_18[2] , 
        \wRegOut_6_18[1] , \wRegOut_6_18[0] }), .L_Out({\wRegInTop_6_18[31] , 
        \wRegInTop_6_18[30] , \wRegInTop_6_18[29] , \wRegInTop_6_18[28] , 
        \wRegInTop_6_18[27] , \wRegInTop_6_18[26] , \wRegInTop_6_18[25] , 
        \wRegInTop_6_18[24] , \wRegInTop_6_18[23] , \wRegInTop_6_18[22] , 
        \wRegInTop_6_18[21] , \wRegInTop_6_18[20] , \wRegInTop_6_18[19] , 
        \wRegInTop_6_18[18] , \wRegInTop_6_18[17] , \wRegInTop_6_18[16] , 
        \wRegInTop_6_18[15] , \wRegInTop_6_18[14] , \wRegInTop_6_18[13] , 
        \wRegInTop_6_18[12] , \wRegInTop_6_18[11] , \wRegInTop_6_18[10] , 
        \wRegInTop_6_18[9] , \wRegInTop_6_18[8] , \wRegInTop_6_18[7] , 
        \wRegInTop_6_18[6] , \wRegInTop_6_18[5] , \wRegInTop_6_18[4] , 
        \wRegInTop_6_18[3] , \wRegInTop_6_18[2] , \wRegInTop_6_18[1] , 
        \wRegInTop_6_18[0] }), .R_WR(\wRegEnTop_6_19[0] ), .R_In({
        \wRegOut_6_19[31] , \wRegOut_6_19[30] , \wRegOut_6_19[29] , 
        \wRegOut_6_19[28] , \wRegOut_6_19[27] , \wRegOut_6_19[26] , 
        \wRegOut_6_19[25] , \wRegOut_6_19[24] , \wRegOut_6_19[23] , 
        \wRegOut_6_19[22] , \wRegOut_6_19[21] , \wRegOut_6_19[20] , 
        \wRegOut_6_19[19] , \wRegOut_6_19[18] , \wRegOut_6_19[17] , 
        \wRegOut_6_19[16] , \wRegOut_6_19[15] , \wRegOut_6_19[14] , 
        \wRegOut_6_19[13] , \wRegOut_6_19[12] , \wRegOut_6_19[11] , 
        \wRegOut_6_19[10] , \wRegOut_6_19[9] , \wRegOut_6_19[8] , 
        \wRegOut_6_19[7] , \wRegOut_6_19[6] , \wRegOut_6_19[5] , 
        \wRegOut_6_19[4] , \wRegOut_6_19[3] , \wRegOut_6_19[2] , 
        \wRegOut_6_19[1] , \wRegOut_6_19[0] }), .R_Out({\wRegInTop_6_19[31] , 
        \wRegInTop_6_19[30] , \wRegInTop_6_19[29] , \wRegInTop_6_19[28] , 
        \wRegInTop_6_19[27] , \wRegInTop_6_19[26] , \wRegInTop_6_19[25] , 
        \wRegInTop_6_19[24] , \wRegInTop_6_19[23] , \wRegInTop_6_19[22] , 
        \wRegInTop_6_19[21] , \wRegInTop_6_19[20] , \wRegInTop_6_19[19] , 
        \wRegInTop_6_19[18] , \wRegInTop_6_19[17] , \wRegInTop_6_19[16] , 
        \wRegInTop_6_19[15] , \wRegInTop_6_19[14] , \wRegInTop_6_19[13] , 
        \wRegInTop_6_19[12] , \wRegInTop_6_19[11] , \wRegInTop_6_19[10] , 
        \wRegInTop_6_19[9] , \wRegInTop_6_19[8] , \wRegInTop_6_19[7] , 
        \wRegInTop_6_19[6] , \wRegInTop_6_19[5] , \wRegInTop_6_19[4] , 
        \wRegInTop_6_19[3] , \wRegInTop_6_19[2] , \wRegInTop_6_19[1] , 
        \wRegInTop_6_19[0] }) );
    BHeap_Node_WIDTH32 BHN_2_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_2[0] ), .P_WR(\wRegEnBot_2_3[0] ), .P_In({\wRegOut_2_3[31] , 
        \wRegOut_2_3[30] , \wRegOut_2_3[29] , \wRegOut_2_3[28] , 
        \wRegOut_2_3[27] , \wRegOut_2_3[26] , \wRegOut_2_3[25] , 
        \wRegOut_2_3[24] , \wRegOut_2_3[23] , \wRegOut_2_3[22] , 
        \wRegOut_2_3[21] , \wRegOut_2_3[20] , \wRegOut_2_3[19] , 
        \wRegOut_2_3[18] , \wRegOut_2_3[17] , \wRegOut_2_3[16] , 
        \wRegOut_2_3[15] , \wRegOut_2_3[14] , \wRegOut_2_3[13] , 
        \wRegOut_2_3[12] , \wRegOut_2_3[11] , \wRegOut_2_3[10] , 
        \wRegOut_2_3[9] , \wRegOut_2_3[8] , \wRegOut_2_3[7] , \wRegOut_2_3[6] , 
        \wRegOut_2_3[5] , \wRegOut_2_3[4] , \wRegOut_2_3[3] , \wRegOut_2_3[2] , 
        \wRegOut_2_3[1] , \wRegOut_2_3[0] }), .P_Out({\wRegInBot_2_3[31] , 
        \wRegInBot_2_3[30] , \wRegInBot_2_3[29] , \wRegInBot_2_3[28] , 
        \wRegInBot_2_3[27] , \wRegInBot_2_3[26] , \wRegInBot_2_3[25] , 
        \wRegInBot_2_3[24] , \wRegInBot_2_3[23] , \wRegInBot_2_3[22] , 
        \wRegInBot_2_3[21] , \wRegInBot_2_3[20] , \wRegInBot_2_3[19] , 
        \wRegInBot_2_3[18] , \wRegInBot_2_3[17] , \wRegInBot_2_3[16] , 
        \wRegInBot_2_3[15] , \wRegInBot_2_3[14] , \wRegInBot_2_3[13] , 
        \wRegInBot_2_3[12] , \wRegInBot_2_3[11] , \wRegInBot_2_3[10] , 
        \wRegInBot_2_3[9] , \wRegInBot_2_3[8] , \wRegInBot_2_3[7] , 
        \wRegInBot_2_3[6] , \wRegInBot_2_3[5] , \wRegInBot_2_3[4] , 
        \wRegInBot_2_3[3] , \wRegInBot_2_3[2] , \wRegInBot_2_3[1] , 
        \wRegInBot_2_3[0] }), .L_WR(\wRegEnTop_3_6[0] ), .L_In({
        \wRegOut_3_6[31] , \wRegOut_3_6[30] , \wRegOut_3_6[29] , 
        \wRegOut_3_6[28] , \wRegOut_3_6[27] , \wRegOut_3_6[26] , 
        \wRegOut_3_6[25] , \wRegOut_3_6[24] , \wRegOut_3_6[23] , 
        \wRegOut_3_6[22] , \wRegOut_3_6[21] , \wRegOut_3_6[20] , 
        \wRegOut_3_6[19] , \wRegOut_3_6[18] , \wRegOut_3_6[17] , 
        \wRegOut_3_6[16] , \wRegOut_3_6[15] , \wRegOut_3_6[14] , 
        \wRegOut_3_6[13] , \wRegOut_3_6[12] , \wRegOut_3_6[11] , 
        \wRegOut_3_6[10] , \wRegOut_3_6[9] , \wRegOut_3_6[8] , 
        \wRegOut_3_6[7] , \wRegOut_3_6[6] , \wRegOut_3_6[5] , \wRegOut_3_6[4] , 
        \wRegOut_3_6[3] , \wRegOut_3_6[2] , \wRegOut_3_6[1] , \wRegOut_3_6[0] 
        }), .L_Out({\wRegInTop_3_6[31] , \wRegInTop_3_6[30] , 
        \wRegInTop_3_6[29] , \wRegInTop_3_6[28] , \wRegInTop_3_6[27] , 
        \wRegInTop_3_6[26] , \wRegInTop_3_6[25] , \wRegInTop_3_6[24] , 
        \wRegInTop_3_6[23] , \wRegInTop_3_6[22] , \wRegInTop_3_6[21] , 
        \wRegInTop_3_6[20] , \wRegInTop_3_6[19] , \wRegInTop_3_6[18] , 
        \wRegInTop_3_6[17] , \wRegInTop_3_6[16] , \wRegInTop_3_6[15] , 
        \wRegInTop_3_6[14] , \wRegInTop_3_6[13] , \wRegInTop_3_6[12] , 
        \wRegInTop_3_6[11] , \wRegInTop_3_6[10] , \wRegInTop_3_6[9] , 
        \wRegInTop_3_6[8] , \wRegInTop_3_6[7] , \wRegInTop_3_6[6] , 
        \wRegInTop_3_6[5] , \wRegInTop_3_6[4] , \wRegInTop_3_6[3] , 
        \wRegInTop_3_6[2] , \wRegInTop_3_6[1] , \wRegInTop_3_6[0] }), .R_WR(
        \wRegEnTop_3_7[0] ), .R_In({\wRegOut_3_7[31] , \wRegOut_3_7[30] , 
        \wRegOut_3_7[29] , \wRegOut_3_7[28] , \wRegOut_3_7[27] , 
        \wRegOut_3_7[26] , \wRegOut_3_7[25] , \wRegOut_3_7[24] , 
        \wRegOut_3_7[23] , \wRegOut_3_7[22] , \wRegOut_3_7[21] , 
        \wRegOut_3_7[20] , \wRegOut_3_7[19] , \wRegOut_3_7[18] , 
        \wRegOut_3_7[17] , \wRegOut_3_7[16] , \wRegOut_3_7[15] , 
        \wRegOut_3_7[14] , \wRegOut_3_7[13] , \wRegOut_3_7[12] , 
        \wRegOut_3_7[11] , \wRegOut_3_7[10] , \wRegOut_3_7[9] , 
        \wRegOut_3_7[8] , \wRegOut_3_7[7] , \wRegOut_3_7[6] , \wRegOut_3_7[5] , 
        \wRegOut_3_7[4] , \wRegOut_3_7[3] , \wRegOut_3_7[2] , \wRegOut_3_7[1] , 
        \wRegOut_3_7[0] }), .R_Out({\wRegInTop_3_7[31] , \wRegInTop_3_7[30] , 
        \wRegInTop_3_7[29] , \wRegInTop_3_7[28] , \wRegInTop_3_7[27] , 
        \wRegInTop_3_7[26] , \wRegInTop_3_7[25] , \wRegInTop_3_7[24] , 
        \wRegInTop_3_7[23] , \wRegInTop_3_7[22] , \wRegInTop_3_7[21] , 
        \wRegInTop_3_7[20] , \wRegInTop_3_7[19] , \wRegInTop_3_7[18] , 
        \wRegInTop_3_7[17] , \wRegInTop_3_7[16] , \wRegInTop_3_7[15] , 
        \wRegInTop_3_7[14] , \wRegInTop_3_7[13] , \wRegInTop_3_7[12] , 
        \wRegInTop_3_7[11] , \wRegInTop_3_7[10] , \wRegInTop_3_7[9] , 
        \wRegInTop_3_7[8] , \wRegInTop_3_7[7] , \wRegInTop_3_7[6] , 
        \wRegInTop_3_7[5] , \wRegInTop_3_7[4] , \wRegInTop_3_7[3] , 
        \wRegInTop_3_7[2] , \wRegInTop_3_7[1] , \wRegInTop_3_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_34 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink162[31] , \ScanLink162[30] , \ScanLink162[29] , 
        \ScanLink162[28] , \ScanLink162[27] , \ScanLink162[26] , 
        \ScanLink162[25] , \ScanLink162[24] , \ScanLink162[23] , 
        \ScanLink162[22] , \ScanLink162[21] , \ScanLink162[20] , 
        \ScanLink162[19] , \ScanLink162[18] , \ScanLink162[17] , 
        \ScanLink162[16] , \ScanLink162[15] , \ScanLink162[14] , 
        \ScanLink162[13] , \ScanLink162[12] , \ScanLink162[11] , 
        \ScanLink162[10] , \ScanLink162[9] , \ScanLink162[8] , 
        \ScanLink162[7] , \ScanLink162[6] , \ScanLink162[5] , \ScanLink162[4] , 
        \ScanLink162[3] , \ScanLink162[2] , \ScanLink162[1] , \ScanLink162[0] 
        }), .ScanOut({\ScanLink161[31] , \ScanLink161[30] , \ScanLink161[29] , 
        \ScanLink161[28] , \ScanLink161[27] , \ScanLink161[26] , 
        \ScanLink161[25] , \ScanLink161[24] , \ScanLink161[23] , 
        \ScanLink161[22] , \ScanLink161[21] , \ScanLink161[20] , 
        \ScanLink161[19] , \ScanLink161[18] , \ScanLink161[17] , 
        \ScanLink161[16] , \ScanLink161[15] , \ScanLink161[14] , 
        \ScanLink161[13] , \ScanLink161[12] , \ScanLink161[11] , 
        \ScanLink161[10] , \ScanLink161[9] , \ScanLink161[8] , 
        \ScanLink161[7] , \ScanLink161[6] , \ScanLink161[5] , \ScanLink161[4] , 
        \ScanLink161[3] , \ScanLink161[2] , \ScanLink161[1] , \ScanLink161[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_34[31] , 
        \wRegOut_7_34[30] , \wRegOut_7_34[29] , \wRegOut_7_34[28] , 
        \wRegOut_7_34[27] , \wRegOut_7_34[26] , \wRegOut_7_34[25] , 
        \wRegOut_7_34[24] , \wRegOut_7_34[23] , \wRegOut_7_34[22] , 
        \wRegOut_7_34[21] , \wRegOut_7_34[20] , \wRegOut_7_34[19] , 
        \wRegOut_7_34[18] , \wRegOut_7_34[17] , \wRegOut_7_34[16] , 
        \wRegOut_7_34[15] , \wRegOut_7_34[14] , \wRegOut_7_34[13] , 
        \wRegOut_7_34[12] , \wRegOut_7_34[11] , \wRegOut_7_34[10] , 
        \wRegOut_7_34[9] , \wRegOut_7_34[8] , \wRegOut_7_34[7] , 
        \wRegOut_7_34[6] , \wRegOut_7_34[5] , \wRegOut_7_34[4] , 
        \wRegOut_7_34[3] , \wRegOut_7_34[2] , \wRegOut_7_34[1] , 
        \wRegOut_7_34[0] }), .Enable1(\wRegEnTop_7_34[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_34[31] , \wRegInTop_7_34[30] , \wRegInTop_7_34[29] , 
        \wRegInTop_7_34[28] , \wRegInTop_7_34[27] , \wRegInTop_7_34[26] , 
        \wRegInTop_7_34[25] , \wRegInTop_7_34[24] , \wRegInTop_7_34[23] , 
        \wRegInTop_7_34[22] , \wRegInTop_7_34[21] , \wRegInTop_7_34[20] , 
        \wRegInTop_7_34[19] , \wRegInTop_7_34[18] , \wRegInTop_7_34[17] , 
        \wRegInTop_7_34[16] , \wRegInTop_7_34[15] , \wRegInTop_7_34[14] , 
        \wRegInTop_7_34[13] , \wRegInTop_7_34[12] , \wRegInTop_7_34[11] , 
        \wRegInTop_7_34[10] , \wRegInTop_7_34[9] , \wRegInTop_7_34[8] , 
        \wRegInTop_7_34[7] , \wRegInTop_7_34[6] , \wRegInTop_7_34[5] , 
        \wRegInTop_7_34[4] , \wRegInTop_7_34[3] , \wRegInTop_7_34[2] , 
        \wRegInTop_7_34[1] , \wRegInTop_7_34[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_120 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink248[31] , \ScanLink248[30] , \ScanLink248[29] , 
        \ScanLink248[28] , \ScanLink248[27] , \ScanLink248[26] , 
        \ScanLink248[25] , \ScanLink248[24] , \ScanLink248[23] , 
        \ScanLink248[22] , \ScanLink248[21] , \ScanLink248[20] , 
        \ScanLink248[19] , \ScanLink248[18] , \ScanLink248[17] , 
        \ScanLink248[16] , \ScanLink248[15] , \ScanLink248[14] , 
        \ScanLink248[13] , \ScanLink248[12] , \ScanLink248[11] , 
        \ScanLink248[10] , \ScanLink248[9] , \ScanLink248[8] , 
        \ScanLink248[7] , \ScanLink248[6] , \ScanLink248[5] , \ScanLink248[4] , 
        \ScanLink248[3] , \ScanLink248[2] , \ScanLink248[1] , \ScanLink248[0] 
        }), .ScanOut({\ScanLink247[31] , \ScanLink247[30] , \ScanLink247[29] , 
        \ScanLink247[28] , \ScanLink247[27] , \ScanLink247[26] , 
        \ScanLink247[25] , \ScanLink247[24] , \ScanLink247[23] , 
        \ScanLink247[22] , \ScanLink247[21] , \ScanLink247[20] , 
        \ScanLink247[19] , \ScanLink247[18] , \ScanLink247[17] , 
        \ScanLink247[16] , \ScanLink247[15] , \ScanLink247[14] , 
        \ScanLink247[13] , \ScanLink247[12] , \ScanLink247[11] , 
        \ScanLink247[10] , \ScanLink247[9] , \ScanLink247[8] , 
        \ScanLink247[7] , \ScanLink247[6] , \ScanLink247[5] , \ScanLink247[4] , 
        \ScanLink247[3] , \ScanLink247[2] , \ScanLink247[1] , \ScanLink247[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_120[31] , 
        \wRegOut_7_120[30] , \wRegOut_7_120[29] , \wRegOut_7_120[28] , 
        \wRegOut_7_120[27] , \wRegOut_7_120[26] , \wRegOut_7_120[25] , 
        \wRegOut_7_120[24] , \wRegOut_7_120[23] , \wRegOut_7_120[22] , 
        \wRegOut_7_120[21] , \wRegOut_7_120[20] , \wRegOut_7_120[19] , 
        \wRegOut_7_120[18] , \wRegOut_7_120[17] , \wRegOut_7_120[16] , 
        \wRegOut_7_120[15] , \wRegOut_7_120[14] , \wRegOut_7_120[13] , 
        \wRegOut_7_120[12] , \wRegOut_7_120[11] , \wRegOut_7_120[10] , 
        \wRegOut_7_120[9] , \wRegOut_7_120[8] , \wRegOut_7_120[7] , 
        \wRegOut_7_120[6] , \wRegOut_7_120[5] , \wRegOut_7_120[4] , 
        \wRegOut_7_120[3] , \wRegOut_7_120[2] , \wRegOut_7_120[1] , 
        \wRegOut_7_120[0] }), .Enable1(\wRegEnTop_7_120[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_120[31] , \wRegInTop_7_120[30] , 
        \wRegInTop_7_120[29] , \wRegInTop_7_120[28] , \wRegInTop_7_120[27] , 
        \wRegInTop_7_120[26] , \wRegInTop_7_120[25] , \wRegInTop_7_120[24] , 
        \wRegInTop_7_120[23] , \wRegInTop_7_120[22] , \wRegInTop_7_120[21] , 
        \wRegInTop_7_120[20] , \wRegInTop_7_120[19] , \wRegInTop_7_120[18] , 
        \wRegInTop_7_120[17] , \wRegInTop_7_120[16] , \wRegInTop_7_120[15] , 
        \wRegInTop_7_120[14] , \wRegInTop_7_120[13] , \wRegInTop_7_120[12] , 
        \wRegInTop_7_120[11] , \wRegInTop_7_120[10] , \wRegInTop_7_120[9] , 
        \wRegInTop_7_120[8] , \wRegInTop_7_120[7] , \wRegInTop_7_120[6] , 
        \wRegInTop_7_120[5] , \wRegInTop_7_120[4] , \wRegInTop_7_120[3] , 
        \wRegInTop_7_120[2] , \wRegInTop_7_120[1] , \wRegInTop_7_120[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_83 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink211[31] , \ScanLink211[30] , \ScanLink211[29] , 
        \ScanLink211[28] , \ScanLink211[27] , \ScanLink211[26] , 
        \ScanLink211[25] , \ScanLink211[24] , \ScanLink211[23] , 
        \ScanLink211[22] , \ScanLink211[21] , \ScanLink211[20] , 
        \ScanLink211[19] , \ScanLink211[18] , \ScanLink211[17] , 
        \ScanLink211[16] , \ScanLink211[15] , \ScanLink211[14] , 
        \ScanLink211[13] , \ScanLink211[12] , \ScanLink211[11] , 
        \ScanLink211[10] , \ScanLink211[9] , \ScanLink211[8] , 
        \ScanLink211[7] , \ScanLink211[6] , \ScanLink211[5] , \ScanLink211[4] , 
        \ScanLink211[3] , \ScanLink211[2] , \ScanLink211[1] , \ScanLink211[0] 
        }), .ScanOut({\ScanLink210[31] , \ScanLink210[30] , \ScanLink210[29] , 
        \ScanLink210[28] , \ScanLink210[27] , \ScanLink210[26] , 
        \ScanLink210[25] , \ScanLink210[24] , \ScanLink210[23] , 
        \ScanLink210[22] , \ScanLink210[21] , \ScanLink210[20] , 
        \ScanLink210[19] , \ScanLink210[18] , \ScanLink210[17] , 
        \ScanLink210[16] , \ScanLink210[15] , \ScanLink210[14] , 
        \ScanLink210[13] , \ScanLink210[12] , \ScanLink210[11] , 
        \ScanLink210[10] , \ScanLink210[9] , \ScanLink210[8] , 
        \ScanLink210[7] , \ScanLink210[6] , \ScanLink210[5] , \ScanLink210[4] , 
        \ScanLink210[3] , \ScanLink210[2] , \ScanLink210[1] , \ScanLink210[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_83[31] , 
        \wRegOut_7_83[30] , \wRegOut_7_83[29] , \wRegOut_7_83[28] , 
        \wRegOut_7_83[27] , \wRegOut_7_83[26] , \wRegOut_7_83[25] , 
        \wRegOut_7_83[24] , \wRegOut_7_83[23] , \wRegOut_7_83[22] , 
        \wRegOut_7_83[21] , \wRegOut_7_83[20] , \wRegOut_7_83[19] , 
        \wRegOut_7_83[18] , \wRegOut_7_83[17] , \wRegOut_7_83[16] , 
        \wRegOut_7_83[15] , \wRegOut_7_83[14] , \wRegOut_7_83[13] , 
        \wRegOut_7_83[12] , \wRegOut_7_83[11] , \wRegOut_7_83[10] , 
        \wRegOut_7_83[9] , \wRegOut_7_83[8] , \wRegOut_7_83[7] , 
        \wRegOut_7_83[6] , \wRegOut_7_83[5] , \wRegOut_7_83[4] , 
        \wRegOut_7_83[3] , \wRegOut_7_83[2] , \wRegOut_7_83[1] , 
        \wRegOut_7_83[0] }), .Enable1(\wRegEnTop_7_83[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_83[31] , \wRegInTop_7_83[30] , \wRegInTop_7_83[29] , 
        \wRegInTop_7_83[28] , \wRegInTop_7_83[27] , \wRegInTop_7_83[26] , 
        \wRegInTop_7_83[25] , \wRegInTop_7_83[24] , \wRegInTop_7_83[23] , 
        \wRegInTop_7_83[22] , \wRegInTop_7_83[21] , \wRegInTop_7_83[20] , 
        \wRegInTop_7_83[19] , \wRegInTop_7_83[18] , \wRegInTop_7_83[17] , 
        \wRegInTop_7_83[16] , \wRegInTop_7_83[15] , \wRegInTop_7_83[14] , 
        \wRegInTop_7_83[13] , \wRegInTop_7_83[12] , \wRegInTop_7_83[11] , 
        \wRegInTop_7_83[10] , \wRegInTop_7_83[9] , \wRegInTop_7_83[8] , 
        \wRegInTop_7_83[7] , \wRegInTop_7_83[6] , \wRegInTop_7_83[5] , 
        \wRegInTop_7_83[4] , \wRegInTop_7_83[3] , \wRegInTop_7_83[2] , 
        \wRegInTop_7_83[1] , \wRegInTop_7_83[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_3[0] ), .P_In({\wRegOut_3_3[31] , 
        \wRegOut_3_3[30] , \wRegOut_3_3[29] , \wRegOut_3_3[28] , 
        \wRegOut_3_3[27] , \wRegOut_3_3[26] , \wRegOut_3_3[25] , 
        \wRegOut_3_3[24] , \wRegOut_3_3[23] , \wRegOut_3_3[22] , 
        \wRegOut_3_3[21] , \wRegOut_3_3[20] , \wRegOut_3_3[19] , 
        \wRegOut_3_3[18] , \wRegOut_3_3[17] , \wRegOut_3_3[16] , 
        \wRegOut_3_3[15] , \wRegOut_3_3[14] , \wRegOut_3_3[13] , 
        \wRegOut_3_3[12] , \wRegOut_3_3[11] , \wRegOut_3_3[10] , 
        \wRegOut_3_3[9] , \wRegOut_3_3[8] , \wRegOut_3_3[7] , \wRegOut_3_3[6] , 
        \wRegOut_3_3[5] , \wRegOut_3_3[4] , \wRegOut_3_3[3] , \wRegOut_3_3[2] , 
        \wRegOut_3_3[1] , \wRegOut_3_3[0] }), .P_Out({\wRegInBot_3_3[31] , 
        \wRegInBot_3_3[30] , \wRegInBot_3_3[29] , \wRegInBot_3_3[28] , 
        \wRegInBot_3_3[27] , \wRegInBot_3_3[26] , \wRegInBot_3_3[25] , 
        \wRegInBot_3_3[24] , \wRegInBot_3_3[23] , \wRegInBot_3_3[22] , 
        \wRegInBot_3_3[21] , \wRegInBot_3_3[20] , \wRegInBot_3_3[19] , 
        \wRegInBot_3_3[18] , \wRegInBot_3_3[17] , \wRegInBot_3_3[16] , 
        \wRegInBot_3_3[15] , \wRegInBot_3_3[14] , \wRegInBot_3_3[13] , 
        \wRegInBot_3_3[12] , \wRegInBot_3_3[11] , \wRegInBot_3_3[10] , 
        \wRegInBot_3_3[9] , \wRegInBot_3_3[8] , \wRegInBot_3_3[7] , 
        \wRegInBot_3_3[6] , \wRegInBot_3_3[5] , \wRegInBot_3_3[4] , 
        \wRegInBot_3_3[3] , \wRegInBot_3_3[2] , \wRegInBot_3_3[1] , 
        \wRegInBot_3_3[0] }), .L_WR(\wRegEnTop_4_6[0] ), .L_In({
        \wRegOut_4_6[31] , \wRegOut_4_6[30] , \wRegOut_4_6[29] , 
        \wRegOut_4_6[28] , \wRegOut_4_6[27] , \wRegOut_4_6[26] , 
        \wRegOut_4_6[25] , \wRegOut_4_6[24] , \wRegOut_4_6[23] , 
        \wRegOut_4_6[22] , \wRegOut_4_6[21] , \wRegOut_4_6[20] , 
        \wRegOut_4_6[19] , \wRegOut_4_6[18] , \wRegOut_4_6[17] , 
        \wRegOut_4_6[16] , \wRegOut_4_6[15] , \wRegOut_4_6[14] , 
        \wRegOut_4_6[13] , \wRegOut_4_6[12] , \wRegOut_4_6[11] , 
        \wRegOut_4_6[10] , \wRegOut_4_6[9] , \wRegOut_4_6[8] , 
        \wRegOut_4_6[7] , \wRegOut_4_6[6] , \wRegOut_4_6[5] , \wRegOut_4_6[4] , 
        \wRegOut_4_6[3] , \wRegOut_4_6[2] , \wRegOut_4_6[1] , \wRegOut_4_6[0] 
        }), .L_Out({\wRegInTop_4_6[31] , \wRegInTop_4_6[30] , 
        \wRegInTop_4_6[29] , \wRegInTop_4_6[28] , \wRegInTop_4_6[27] , 
        \wRegInTop_4_6[26] , \wRegInTop_4_6[25] , \wRegInTop_4_6[24] , 
        \wRegInTop_4_6[23] , \wRegInTop_4_6[22] , \wRegInTop_4_6[21] , 
        \wRegInTop_4_6[20] , \wRegInTop_4_6[19] , \wRegInTop_4_6[18] , 
        \wRegInTop_4_6[17] , \wRegInTop_4_6[16] , \wRegInTop_4_6[15] , 
        \wRegInTop_4_6[14] , \wRegInTop_4_6[13] , \wRegInTop_4_6[12] , 
        \wRegInTop_4_6[11] , \wRegInTop_4_6[10] , \wRegInTop_4_6[9] , 
        \wRegInTop_4_6[8] , \wRegInTop_4_6[7] , \wRegInTop_4_6[6] , 
        \wRegInTop_4_6[5] , \wRegInTop_4_6[4] , \wRegInTop_4_6[3] , 
        \wRegInTop_4_6[2] , \wRegInTop_4_6[1] , \wRegInTop_4_6[0] }), .R_WR(
        \wRegEnTop_4_7[0] ), .R_In({\wRegOut_4_7[31] , \wRegOut_4_7[30] , 
        \wRegOut_4_7[29] , \wRegOut_4_7[28] , \wRegOut_4_7[27] , 
        \wRegOut_4_7[26] , \wRegOut_4_7[25] , \wRegOut_4_7[24] , 
        \wRegOut_4_7[23] , \wRegOut_4_7[22] , \wRegOut_4_7[21] , 
        \wRegOut_4_7[20] , \wRegOut_4_7[19] , \wRegOut_4_7[18] , 
        \wRegOut_4_7[17] , \wRegOut_4_7[16] , \wRegOut_4_7[15] , 
        \wRegOut_4_7[14] , \wRegOut_4_7[13] , \wRegOut_4_7[12] , 
        \wRegOut_4_7[11] , \wRegOut_4_7[10] , \wRegOut_4_7[9] , 
        \wRegOut_4_7[8] , \wRegOut_4_7[7] , \wRegOut_4_7[6] , \wRegOut_4_7[5] , 
        \wRegOut_4_7[4] , \wRegOut_4_7[3] , \wRegOut_4_7[2] , \wRegOut_4_7[1] , 
        \wRegOut_4_7[0] }), .R_Out({\wRegInTop_4_7[31] , \wRegInTop_4_7[30] , 
        \wRegInTop_4_7[29] , \wRegInTop_4_7[28] , \wRegInTop_4_7[27] , 
        \wRegInTop_4_7[26] , \wRegInTop_4_7[25] , \wRegInTop_4_7[24] , 
        \wRegInTop_4_7[23] , \wRegInTop_4_7[22] , \wRegInTop_4_7[21] , 
        \wRegInTop_4_7[20] , \wRegInTop_4_7[19] , \wRegInTop_4_7[18] , 
        \wRegInTop_4_7[17] , \wRegInTop_4_7[16] , \wRegInTop_4_7[15] , 
        \wRegInTop_4_7[14] , \wRegInTop_4_7[13] , \wRegInTop_4_7[12] , 
        \wRegInTop_4_7[11] , \wRegInTop_4_7[10] , \wRegInTop_4_7[9] , 
        \wRegInTop_4_7[8] , \wRegInTop_4_7[7] , \wRegInTop_4_7[6] , 
        \wRegInTop_4_7[5] , \wRegInTop_4_7[4] , \wRegInTop_4_7[3] , 
        \wRegInTop_4_7[2] , \wRegInTop_4_7[1] , \wRegInTop_4_7[0] }) );
    BHeap_Node_WIDTH32 BHN_4_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_9[0] ), .P_In({\wRegOut_4_9[31] , 
        \wRegOut_4_9[30] , \wRegOut_4_9[29] , \wRegOut_4_9[28] , 
        \wRegOut_4_9[27] , \wRegOut_4_9[26] , \wRegOut_4_9[25] , 
        \wRegOut_4_9[24] , \wRegOut_4_9[23] , \wRegOut_4_9[22] , 
        \wRegOut_4_9[21] , \wRegOut_4_9[20] , \wRegOut_4_9[19] , 
        \wRegOut_4_9[18] , \wRegOut_4_9[17] , \wRegOut_4_9[16] , 
        \wRegOut_4_9[15] , \wRegOut_4_9[14] , \wRegOut_4_9[13] , 
        \wRegOut_4_9[12] , \wRegOut_4_9[11] , \wRegOut_4_9[10] , 
        \wRegOut_4_9[9] , \wRegOut_4_9[8] , \wRegOut_4_9[7] , \wRegOut_4_9[6] , 
        \wRegOut_4_9[5] , \wRegOut_4_9[4] , \wRegOut_4_9[3] , \wRegOut_4_9[2] , 
        \wRegOut_4_9[1] , \wRegOut_4_9[0] }), .P_Out({\wRegInBot_4_9[31] , 
        \wRegInBot_4_9[30] , \wRegInBot_4_9[29] , \wRegInBot_4_9[28] , 
        \wRegInBot_4_9[27] , \wRegInBot_4_9[26] , \wRegInBot_4_9[25] , 
        \wRegInBot_4_9[24] , \wRegInBot_4_9[23] , \wRegInBot_4_9[22] , 
        \wRegInBot_4_9[21] , \wRegInBot_4_9[20] , \wRegInBot_4_9[19] , 
        \wRegInBot_4_9[18] , \wRegInBot_4_9[17] , \wRegInBot_4_9[16] , 
        \wRegInBot_4_9[15] , \wRegInBot_4_9[14] , \wRegInBot_4_9[13] , 
        \wRegInBot_4_9[12] , \wRegInBot_4_9[11] , \wRegInBot_4_9[10] , 
        \wRegInBot_4_9[9] , \wRegInBot_4_9[8] , \wRegInBot_4_9[7] , 
        \wRegInBot_4_9[6] , \wRegInBot_4_9[5] , \wRegInBot_4_9[4] , 
        \wRegInBot_4_9[3] , \wRegInBot_4_9[2] , \wRegInBot_4_9[1] , 
        \wRegInBot_4_9[0] }), .L_WR(\wRegEnTop_5_18[0] ), .L_In({
        \wRegOut_5_18[31] , \wRegOut_5_18[30] , \wRegOut_5_18[29] , 
        \wRegOut_5_18[28] , \wRegOut_5_18[27] , \wRegOut_5_18[26] , 
        \wRegOut_5_18[25] , \wRegOut_5_18[24] , \wRegOut_5_18[23] , 
        \wRegOut_5_18[22] , \wRegOut_5_18[21] , \wRegOut_5_18[20] , 
        \wRegOut_5_18[19] , \wRegOut_5_18[18] , \wRegOut_5_18[17] , 
        \wRegOut_5_18[16] , \wRegOut_5_18[15] , \wRegOut_5_18[14] , 
        \wRegOut_5_18[13] , \wRegOut_5_18[12] , \wRegOut_5_18[11] , 
        \wRegOut_5_18[10] , \wRegOut_5_18[9] , \wRegOut_5_18[8] , 
        \wRegOut_5_18[7] , \wRegOut_5_18[6] , \wRegOut_5_18[5] , 
        \wRegOut_5_18[4] , \wRegOut_5_18[3] , \wRegOut_5_18[2] , 
        \wRegOut_5_18[1] , \wRegOut_5_18[0] }), .L_Out({\wRegInTop_5_18[31] , 
        \wRegInTop_5_18[30] , \wRegInTop_5_18[29] , \wRegInTop_5_18[28] , 
        \wRegInTop_5_18[27] , \wRegInTop_5_18[26] , \wRegInTop_5_18[25] , 
        \wRegInTop_5_18[24] , \wRegInTop_5_18[23] , \wRegInTop_5_18[22] , 
        \wRegInTop_5_18[21] , \wRegInTop_5_18[20] , \wRegInTop_5_18[19] , 
        \wRegInTop_5_18[18] , \wRegInTop_5_18[17] , \wRegInTop_5_18[16] , 
        \wRegInTop_5_18[15] , \wRegInTop_5_18[14] , \wRegInTop_5_18[13] , 
        \wRegInTop_5_18[12] , \wRegInTop_5_18[11] , \wRegInTop_5_18[10] , 
        \wRegInTop_5_18[9] , \wRegInTop_5_18[8] , \wRegInTop_5_18[7] , 
        \wRegInTop_5_18[6] , \wRegInTop_5_18[5] , \wRegInTop_5_18[4] , 
        \wRegInTop_5_18[3] , \wRegInTop_5_18[2] , \wRegInTop_5_18[1] , 
        \wRegInTop_5_18[0] }), .R_WR(\wRegEnTop_5_19[0] ), .R_In({
        \wRegOut_5_19[31] , \wRegOut_5_19[30] , \wRegOut_5_19[29] , 
        \wRegOut_5_19[28] , \wRegOut_5_19[27] , \wRegOut_5_19[26] , 
        \wRegOut_5_19[25] , \wRegOut_5_19[24] , \wRegOut_5_19[23] , 
        \wRegOut_5_19[22] , \wRegOut_5_19[21] , \wRegOut_5_19[20] , 
        \wRegOut_5_19[19] , \wRegOut_5_19[18] , \wRegOut_5_19[17] , 
        \wRegOut_5_19[16] , \wRegOut_5_19[15] , \wRegOut_5_19[14] , 
        \wRegOut_5_19[13] , \wRegOut_5_19[12] , \wRegOut_5_19[11] , 
        \wRegOut_5_19[10] , \wRegOut_5_19[9] , \wRegOut_5_19[8] , 
        \wRegOut_5_19[7] , \wRegOut_5_19[6] , \wRegOut_5_19[5] , 
        \wRegOut_5_19[4] , \wRegOut_5_19[3] , \wRegOut_5_19[2] , 
        \wRegOut_5_19[1] , \wRegOut_5_19[0] }), .R_Out({\wRegInTop_5_19[31] , 
        \wRegInTop_5_19[30] , \wRegInTop_5_19[29] , \wRegInTop_5_19[28] , 
        \wRegInTop_5_19[27] , \wRegInTop_5_19[26] , \wRegInTop_5_19[25] , 
        \wRegInTop_5_19[24] , \wRegInTop_5_19[23] , \wRegInTop_5_19[22] , 
        \wRegInTop_5_19[21] , \wRegInTop_5_19[20] , \wRegInTop_5_19[19] , 
        \wRegInTop_5_19[18] , \wRegInTop_5_19[17] , \wRegInTop_5_19[16] , 
        \wRegInTop_5_19[15] , \wRegInTop_5_19[14] , \wRegInTop_5_19[13] , 
        \wRegInTop_5_19[12] , \wRegInTop_5_19[11] , \wRegInTop_5_19[10] , 
        \wRegInTop_5_19[9] , \wRegInTop_5_19[8] , \wRegInTop_5_19[7] , 
        \wRegInTop_5_19[6] , \wRegInTop_5_19[5] , \wRegInTop_5_19[4] , 
        \wRegInTop_5_19[3] , \wRegInTop_5_19[2] , \wRegInTop_5_19[1] , 
        \wRegInTop_5_19[0] }) );
    BHeap_Node_WIDTH32 BHN_4_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_10[0] ), .P_In({\wRegOut_4_10[31] , 
        \wRegOut_4_10[30] , \wRegOut_4_10[29] , \wRegOut_4_10[28] , 
        \wRegOut_4_10[27] , \wRegOut_4_10[26] , \wRegOut_4_10[25] , 
        \wRegOut_4_10[24] , \wRegOut_4_10[23] , \wRegOut_4_10[22] , 
        \wRegOut_4_10[21] , \wRegOut_4_10[20] , \wRegOut_4_10[19] , 
        \wRegOut_4_10[18] , \wRegOut_4_10[17] , \wRegOut_4_10[16] , 
        \wRegOut_4_10[15] , \wRegOut_4_10[14] , \wRegOut_4_10[13] , 
        \wRegOut_4_10[12] , \wRegOut_4_10[11] , \wRegOut_4_10[10] , 
        \wRegOut_4_10[9] , \wRegOut_4_10[8] , \wRegOut_4_10[7] , 
        \wRegOut_4_10[6] , \wRegOut_4_10[5] , \wRegOut_4_10[4] , 
        \wRegOut_4_10[3] , \wRegOut_4_10[2] , \wRegOut_4_10[1] , 
        \wRegOut_4_10[0] }), .P_Out({\wRegInBot_4_10[31] , 
        \wRegInBot_4_10[30] , \wRegInBot_4_10[29] , \wRegInBot_4_10[28] , 
        \wRegInBot_4_10[27] , \wRegInBot_4_10[26] , \wRegInBot_4_10[25] , 
        \wRegInBot_4_10[24] , \wRegInBot_4_10[23] , \wRegInBot_4_10[22] , 
        \wRegInBot_4_10[21] , \wRegInBot_4_10[20] , \wRegInBot_4_10[19] , 
        \wRegInBot_4_10[18] , \wRegInBot_4_10[17] , \wRegInBot_4_10[16] , 
        \wRegInBot_4_10[15] , \wRegInBot_4_10[14] , \wRegInBot_4_10[13] , 
        \wRegInBot_4_10[12] , \wRegInBot_4_10[11] , \wRegInBot_4_10[10] , 
        \wRegInBot_4_10[9] , \wRegInBot_4_10[8] , \wRegInBot_4_10[7] , 
        \wRegInBot_4_10[6] , \wRegInBot_4_10[5] , \wRegInBot_4_10[4] , 
        \wRegInBot_4_10[3] , \wRegInBot_4_10[2] , \wRegInBot_4_10[1] , 
        \wRegInBot_4_10[0] }), .L_WR(\wRegEnTop_5_20[0] ), .L_In({
        \wRegOut_5_20[31] , \wRegOut_5_20[30] , \wRegOut_5_20[29] , 
        \wRegOut_5_20[28] , \wRegOut_5_20[27] , \wRegOut_5_20[26] , 
        \wRegOut_5_20[25] , \wRegOut_5_20[24] , \wRegOut_5_20[23] , 
        \wRegOut_5_20[22] , \wRegOut_5_20[21] , \wRegOut_5_20[20] , 
        \wRegOut_5_20[19] , \wRegOut_5_20[18] , \wRegOut_5_20[17] , 
        \wRegOut_5_20[16] , \wRegOut_5_20[15] , \wRegOut_5_20[14] , 
        \wRegOut_5_20[13] , \wRegOut_5_20[12] , \wRegOut_5_20[11] , 
        \wRegOut_5_20[10] , \wRegOut_5_20[9] , \wRegOut_5_20[8] , 
        \wRegOut_5_20[7] , \wRegOut_5_20[6] , \wRegOut_5_20[5] , 
        \wRegOut_5_20[4] , \wRegOut_5_20[3] , \wRegOut_5_20[2] , 
        \wRegOut_5_20[1] , \wRegOut_5_20[0] }), .L_Out({\wRegInTop_5_20[31] , 
        \wRegInTop_5_20[30] , \wRegInTop_5_20[29] , \wRegInTop_5_20[28] , 
        \wRegInTop_5_20[27] , \wRegInTop_5_20[26] , \wRegInTop_5_20[25] , 
        \wRegInTop_5_20[24] , \wRegInTop_5_20[23] , \wRegInTop_5_20[22] , 
        \wRegInTop_5_20[21] , \wRegInTop_5_20[20] , \wRegInTop_5_20[19] , 
        \wRegInTop_5_20[18] , \wRegInTop_5_20[17] , \wRegInTop_5_20[16] , 
        \wRegInTop_5_20[15] , \wRegInTop_5_20[14] , \wRegInTop_5_20[13] , 
        \wRegInTop_5_20[12] , \wRegInTop_5_20[11] , \wRegInTop_5_20[10] , 
        \wRegInTop_5_20[9] , \wRegInTop_5_20[8] , \wRegInTop_5_20[7] , 
        \wRegInTop_5_20[6] , \wRegInTop_5_20[5] , \wRegInTop_5_20[4] , 
        \wRegInTop_5_20[3] , \wRegInTop_5_20[2] , \wRegInTop_5_20[1] , 
        \wRegInTop_5_20[0] }), .R_WR(\wRegEnTop_5_21[0] ), .R_In({
        \wRegOut_5_21[31] , \wRegOut_5_21[30] , \wRegOut_5_21[29] , 
        \wRegOut_5_21[28] , \wRegOut_5_21[27] , \wRegOut_5_21[26] , 
        \wRegOut_5_21[25] , \wRegOut_5_21[24] , \wRegOut_5_21[23] , 
        \wRegOut_5_21[22] , \wRegOut_5_21[21] , \wRegOut_5_21[20] , 
        \wRegOut_5_21[19] , \wRegOut_5_21[18] , \wRegOut_5_21[17] , 
        \wRegOut_5_21[16] , \wRegOut_5_21[15] , \wRegOut_5_21[14] , 
        \wRegOut_5_21[13] , \wRegOut_5_21[12] , \wRegOut_5_21[11] , 
        \wRegOut_5_21[10] , \wRegOut_5_21[9] , \wRegOut_5_21[8] , 
        \wRegOut_5_21[7] , \wRegOut_5_21[6] , \wRegOut_5_21[5] , 
        \wRegOut_5_21[4] , \wRegOut_5_21[3] , \wRegOut_5_21[2] , 
        \wRegOut_5_21[1] , \wRegOut_5_21[0] }), .R_Out({\wRegInTop_5_21[31] , 
        \wRegInTop_5_21[30] , \wRegInTop_5_21[29] , \wRegInTop_5_21[28] , 
        \wRegInTop_5_21[27] , \wRegInTop_5_21[26] , \wRegInTop_5_21[25] , 
        \wRegInTop_5_21[24] , \wRegInTop_5_21[23] , \wRegInTop_5_21[22] , 
        \wRegInTop_5_21[21] , \wRegInTop_5_21[20] , \wRegInTop_5_21[19] , 
        \wRegInTop_5_21[18] , \wRegInTop_5_21[17] , \wRegInTop_5_21[16] , 
        \wRegInTop_5_21[15] , \wRegInTop_5_21[14] , \wRegInTop_5_21[13] , 
        \wRegInTop_5_21[12] , \wRegInTop_5_21[11] , \wRegInTop_5_21[10] , 
        \wRegInTop_5_21[9] , \wRegInTop_5_21[8] , \wRegInTop_5_21[7] , 
        \wRegInTop_5_21[6] , \wRegInTop_5_21[5] , \wRegInTop_5_21[4] , 
        \wRegInTop_5_21[3] , \wRegInTop_5_21[2] , \wRegInTop_5_21[1] , 
        \wRegInTop_5_21[0] }) );
    BHeap_Node_WIDTH32 BHN_6_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_54[0] ), .P_In({\wRegOut_6_54[31] , 
        \wRegOut_6_54[30] , \wRegOut_6_54[29] , \wRegOut_6_54[28] , 
        \wRegOut_6_54[27] , \wRegOut_6_54[26] , \wRegOut_6_54[25] , 
        \wRegOut_6_54[24] , \wRegOut_6_54[23] , \wRegOut_6_54[22] , 
        \wRegOut_6_54[21] , \wRegOut_6_54[20] , \wRegOut_6_54[19] , 
        \wRegOut_6_54[18] , \wRegOut_6_54[17] , \wRegOut_6_54[16] , 
        \wRegOut_6_54[15] , \wRegOut_6_54[14] , \wRegOut_6_54[13] , 
        \wRegOut_6_54[12] , \wRegOut_6_54[11] , \wRegOut_6_54[10] , 
        \wRegOut_6_54[9] , \wRegOut_6_54[8] , \wRegOut_6_54[7] , 
        \wRegOut_6_54[6] , \wRegOut_6_54[5] , \wRegOut_6_54[4] , 
        \wRegOut_6_54[3] , \wRegOut_6_54[2] , \wRegOut_6_54[1] , 
        \wRegOut_6_54[0] }), .P_Out({\wRegInBot_6_54[31] , 
        \wRegInBot_6_54[30] , \wRegInBot_6_54[29] , \wRegInBot_6_54[28] , 
        \wRegInBot_6_54[27] , \wRegInBot_6_54[26] , \wRegInBot_6_54[25] , 
        \wRegInBot_6_54[24] , \wRegInBot_6_54[23] , \wRegInBot_6_54[22] , 
        \wRegInBot_6_54[21] , \wRegInBot_6_54[20] , \wRegInBot_6_54[19] , 
        \wRegInBot_6_54[18] , \wRegInBot_6_54[17] , \wRegInBot_6_54[16] , 
        \wRegInBot_6_54[15] , \wRegInBot_6_54[14] , \wRegInBot_6_54[13] , 
        \wRegInBot_6_54[12] , \wRegInBot_6_54[11] , \wRegInBot_6_54[10] , 
        \wRegInBot_6_54[9] , \wRegInBot_6_54[8] , \wRegInBot_6_54[7] , 
        \wRegInBot_6_54[6] , \wRegInBot_6_54[5] , \wRegInBot_6_54[4] , 
        \wRegInBot_6_54[3] , \wRegInBot_6_54[2] , \wRegInBot_6_54[1] , 
        \wRegInBot_6_54[0] }), .L_WR(\wRegEnTop_7_108[0] ), .L_In({
        \wRegOut_7_108[31] , \wRegOut_7_108[30] , \wRegOut_7_108[29] , 
        \wRegOut_7_108[28] , \wRegOut_7_108[27] , \wRegOut_7_108[26] , 
        \wRegOut_7_108[25] , \wRegOut_7_108[24] , \wRegOut_7_108[23] , 
        \wRegOut_7_108[22] , \wRegOut_7_108[21] , \wRegOut_7_108[20] , 
        \wRegOut_7_108[19] , \wRegOut_7_108[18] , \wRegOut_7_108[17] , 
        \wRegOut_7_108[16] , \wRegOut_7_108[15] , \wRegOut_7_108[14] , 
        \wRegOut_7_108[13] , \wRegOut_7_108[12] , \wRegOut_7_108[11] , 
        \wRegOut_7_108[10] , \wRegOut_7_108[9] , \wRegOut_7_108[8] , 
        \wRegOut_7_108[7] , \wRegOut_7_108[6] , \wRegOut_7_108[5] , 
        \wRegOut_7_108[4] , \wRegOut_7_108[3] , \wRegOut_7_108[2] , 
        \wRegOut_7_108[1] , \wRegOut_7_108[0] }), .L_Out({
        \wRegInTop_7_108[31] , \wRegInTop_7_108[30] , \wRegInTop_7_108[29] , 
        \wRegInTop_7_108[28] , \wRegInTop_7_108[27] , \wRegInTop_7_108[26] , 
        \wRegInTop_7_108[25] , \wRegInTop_7_108[24] , \wRegInTop_7_108[23] , 
        \wRegInTop_7_108[22] , \wRegInTop_7_108[21] , \wRegInTop_7_108[20] , 
        \wRegInTop_7_108[19] , \wRegInTop_7_108[18] , \wRegInTop_7_108[17] , 
        \wRegInTop_7_108[16] , \wRegInTop_7_108[15] , \wRegInTop_7_108[14] , 
        \wRegInTop_7_108[13] , \wRegInTop_7_108[12] , \wRegInTop_7_108[11] , 
        \wRegInTop_7_108[10] , \wRegInTop_7_108[9] , \wRegInTop_7_108[8] , 
        \wRegInTop_7_108[7] , \wRegInTop_7_108[6] , \wRegInTop_7_108[5] , 
        \wRegInTop_7_108[4] , \wRegInTop_7_108[3] , \wRegInTop_7_108[2] , 
        \wRegInTop_7_108[1] , \wRegInTop_7_108[0] }), .R_WR(
        \wRegEnTop_7_109[0] ), .R_In({\wRegOut_7_109[31] , \wRegOut_7_109[30] , 
        \wRegOut_7_109[29] , \wRegOut_7_109[28] , \wRegOut_7_109[27] , 
        \wRegOut_7_109[26] , \wRegOut_7_109[25] , \wRegOut_7_109[24] , 
        \wRegOut_7_109[23] , \wRegOut_7_109[22] , \wRegOut_7_109[21] , 
        \wRegOut_7_109[20] , \wRegOut_7_109[19] , \wRegOut_7_109[18] , 
        \wRegOut_7_109[17] , \wRegOut_7_109[16] , \wRegOut_7_109[15] , 
        \wRegOut_7_109[14] , \wRegOut_7_109[13] , \wRegOut_7_109[12] , 
        \wRegOut_7_109[11] , \wRegOut_7_109[10] , \wRegOut_7_109[9] , 
        \wRegOut_7_109[8] , \wRegOut_7_109[7] , \wRegOut_7_109[6] , 
        \wRegOut_7_109[5] , \wRegOut_7_109[4] , \wRegOut_7_109[3] , 
        \wRegOut_7_109[2] , \wRegOut_7_109[1] , \wRegOut_7_109[0] }), .R_Out({
        \wRegInTop_7_109[31] , \wRegInTop_7_109[30] , \wRegInTop_7_109[29] , 
        \wRegInTop_7_109[28] , \wRegInTop_7_109[27] , \wRegInTop_7_109[26] , 
        \wRegInTop_7_109[25] , \wRegInTop_7_109[24] , \wRegInTop_7_109[23] , 
        \wRegInTop_7_109[22] , \wRegInTop_7_109[21] , \wRegInTop_7_109[20] , 
        \wRegInTop_7_109[19] , \wRegInTop_7_109[18] , \wRegInTop_7_109[17] , 
        \wRegInTop_7_109[16] , \wRegInTop_7_109[15] , \wRegInTop_7_109[14] , 
        \wRegInTop_7_109[13] , \wRegInTop_7_109[12] , \wRegInTop_7_109[11] , 
        \wRegInTop_7_109[10] , \wRegInTop_7_109[9] , \wRegInTop_7_109[8] , 
        \wRegInTop_7_109[7] , \wRegInTop_7_109[6] , \wRegInTop_7_109[5] , 
        \wRegInTop_7_109[4] , \wRegInTop_7_109[3] , \wRegInTop_7_109[2] , 
        \wRegInTop_7_109[1] , \wRegInTop_7_109[0] }) );
    BHeap_Node_WIDTH32 BHN_6_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_5[0] ), .P_In({\wRegOut_6_5[31] , 
        \wRegOut_6_5[30] , \wRegOut_6_5[29] , \wRegOut_6_5[28] , 
        \wRegOut_6_5[27] , \wRegOut_6_5[26] , \wRegOut_6_5[25] , 
        \wRegOut_6_5[24] , \wRegOut_6_5[23] , \wRegOut_6_5[22] , 
        \wRegOut_6_5[21] , \wRegOut_6_5[20] , \wRegOut_6_5[19] , 
        \wRegOut_6_5[18] , \wRegOut_6_5[17] , \wRegOut_6_5[16] , 
        \wRegOut_6_5[15] , \wRegOut_6_5[14] , \wRegOut_6_5[13] , 
        \wRegOut_6_5[12] , \wRegOut_6_5[11] , \wRegOut_6_5[10] , 
        \wRegOut_6_5[9] , \wRegOut_6_5[8] , \wRegOut_6_5[7] , \wRegOut_6_5[6] , 
        \wRegOut_6_5[5] , \wRegOut_6_5[4] , \wRegOut_6_5[3] , \wRegOut_6_5[2] , 
        \wRegOut_6_5[1] , \wRegOut_6_5[0] }), .P_Out({\wRegInBot_6_5[31] , 
        \wRegInBot_6_5[30] , \wRegInBot_6_5[29] , \wRegInBot_6_5[28] , 
        \wRegInBot_6_5[27] , \wRegInBot_6_5[26] , \wRegInBot_6_5[25] , 
        \wRegInBot_6_5[24] , \wRegInBot_6_5[23] , \wRegInBot_6_5[22] , 
        \wRegInBot_6_5[21] , \wRegInBot_6_5[20] , \wRegInBot_6_5[19] , 
        \wRegInBot_6_5[18] , \wRegInBot_6_5[17] , \wRegInBot_6_5[16] , 
        \wRegInBot_6_5[15] , \wRegInBot_6_5[14] , \wRegInBot_6_5[13] , 
        \wRegInBot_6_5[12] , \wRegInBot_6_5[11] , \wRegInBot_6_5[10] , 
        \wRegInBot_6_5[9] , \wRegInBot_6_5[8] , \wRegInBot_6_5[7] , 
        \wRegInBot_6_5[6] , \wRegInBot_6_5[5] , \wRegInBot_6_5[4] , 
        \wRegInBot_6_5[3] , \wRegInBot_6_5[2] , \wRegInBot_6_5[1] , 
        \wRegInBot_6_5[0] }), .L_WR(\wRegEnTop_7_10[0] ), .L_In({
        \wRegOut_7_10[31] , \wRegOut_7_10[30] , \wRegOut_7_10[29] , 
        \wRegOut_7_10[28] , \wRegOut_7_10[27] , \wRegOut_7_10[26] , 
        \wRegOut_7_10[25] , \wRegOut_7_10[24] , \wRegOut_7_10[23] , 
        \wRegOut_7_10[22] , \wRegOut_7_10[21] , \wRegOut_7_10[20] , 
        \wRegOut_7_10[19] , \wRegOut_7_10[18] , \wRegOut_7_10[17] , 
        \wRegOut_7_10[16] , \wRegOut_7_10[15] , \wRegOut_7_10[14] , 
        \wRegOut_7_10[13] , \wRegOut_7_10[12] , \wRegOut_7_10[11] , 
        \wRegOut_7_10[10] , \wRegOut_7_10[9] , \wRegOut_7_10[8] , 
        \wRegOut_7_10[7] , \wRegOut_7_10[6] , \wRegOut_7_10[5] , 
        \wRegOut_7_10[4] , \wRegOut_7_10[3] , \wRegOut_7_10[2] , 
        \wRegOut_7_10[1] , \wRegOut_7_10[0] }), .L_Out({\wRegInTop_7_10[31] , 
        \wRegInTop_7_10[30] , \wRegInTop_7_10[29] , \wRegInTop_7_10[28] , 
        \wRegInTop_7_10[27] , \wRegInTop_7_10[26] , \wRegInTop_7_10[25] , 
        \wRegInTop_7_10[24] , \wRegInTop_7_10[23] , \wRegInTop_7_10[22] , 
        \wRegInTop_7_10[21] , \wRegInTop_7_10[20] , \wRegInTop_7_10[19] , 
        \wRegInTop_7_10[18] , \wRegInTop_7_10[17] , \wRegInTop_7_10[16] , 
        \wRegInTop_7_10[15] , \wRegInTop_7_10[14] , \wRegInTop_7_10[13] , 
        \wRegInTop_7_10[12] , \wRegInTop_7_10[11] , \wRegInTop_7_10[10] , 
        \wRegInTop_7_10[9] , \wRegInTop_7_10[8] , \wRegInTop_7_10[7] , 
        \wRegInTop_7_10[6] , \wRegInTop_7_10[5] , \wRegInTop_7_10[4] , 
        \wRegInTop_7_10[3] , \wRegInTop_7_10[2] , \wRegInTop_7_10[1] , 
        \wRegInTop_7_10[0] }), .R_WR(\wRegEnTop_7_11[0] ), .R_In({
        \wRegOut_7_11[31] , \wRegOut_7_11[30] , \wRegOut_7_11[29] , 
        \wRegOut_7_11[28] , \wRegOut_7_11[27] , \wRegOut_7_11[26] , 
        \wRegOut_7_11[25] , \wRegOut_7_11[24] , \wRegOut_7_11[23] , 
        \wRegOut_7_11[22] , \wRegOut_7_11[21] , \wRegOut_7_11[20] , 
        \wRegOut_7_11[19] , \wRegOut_7_11[18] , \wRegOut_7_11[17] , 
        \wRegOut_7_11[16] , \wRegOut_7_11[15] , \wRegOut_7_11[14] , 
        \wRegOut_7_11[13] , \wRegOut_7_11[12] , \wRegOut_7_11[11] , 
        \wRegOut_7_11[10] , \wRegOut_7_11[9] , \wRegOut_7_11[8] , 
        \wRegOut_7_11[7] , \wRegOut_7_11[6] , \wRegOut_7_11[5] , 
        \wRegOut_7_11[4] , \wRegOut_7_11[3] , \wRegOut_7_11[2] , 
        \wRegOut_7_11[1] , \wRegOut_7_11[0] }), .R_Out({\wRegInTop_7_11[31] , 
        \wRegInTop_7_11[30] , \wRegInTop_7_11[29] , \wRegInTop_7_11[28] , 
        \wRegInTop_7_11[27] , \wRegInTop_7_11[26] , \wRegInTop_7_11[25] , 
        \wRegInTop_7_11[24] , \wRegInTop_7_11[23] , \wRegInTop_7_11[22] , 
        \wRegInTop_7_11[21] , \wRegInTop_7_11[20] , \wRegInTop_7_11[19] , 
        \wRegInTop_7_11[18] , \wRegInTop_7_11[17] , \wRegInTop_7_11[16] , 
        \wRegInTop_7_11[15] , \wRegInTop_7_11[14] , \wRegInTop_7_11[13] , 
        \wRegInTop_7_11[12] , \wRegInTop_7_11[11] , \wRegInTop_7_11[10] , 
        \wRegInTop_7_11[9] , \wRegInTop_7_11[8] , \wRegInTop_7_11[7] , 
        \wRegInTop_7_11[6] , \wRegInTop_7_11[5] , \wRegInTop_7_11[4] , 
        \wRegInTop_7_11[3] , \wRegInTop_7_11[2] , \wRegInTop_7_11[1] , 
        \wRegInTop_7_11[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink19[31] , \ScanLink19[30] , \ScanLink19[29] , 
        \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , \ScanLink19[25] , 
        \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , \ScanLink19[21] , 
        \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , \ScanLink19[17] , 
        \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , \ScanLink19[13] , 
        \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , \ScanLink19[9] , 
        \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , \ScanLink19[5] , 
        \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , \ScanLink19[1] , 
        \ScanLink19[0] }), .ScanOut({\ScanLink18[31] , \ScanLink18[30] , 
        \ScanLink18[29] , \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , 
        \ScanLink18[25] , \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , 
        \ScanLink18[21] , \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , 
        \ScanLink18[17] , \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , 
        \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , 
        \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , 
        \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , 
        \ScanLink18[1] , \ScanLink18[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_3[31] , \wRegOut_4_3[30] , \wRegOut_4_3[29] , 
        \wRegOut_4_3[28] , \wRegOut_4_3[27] , \wRegOut_4_3[26] , 
        \wRegOut_4_3[25] , \wRegOut_4_3[24] , \wRegOut_4_3[23] , 
        \wRegOut_4_3[22] , \wRegOut_4_3[21] , \wRegOut_4_3[20] , 
        \wRegOut_4_3[19] , \wRegOut_4_3[18] , \wRegOut_4_3[17] , 
        \wRegOut_4_3[16] , \wRegOut_4_3[15] , \wRegOut_4_3[14] , 
        \wRegOut_4_3[13] , \wRegOut_4_3[12] , \wRegOut_4_3[11] , 
        \wRegOut_4_3[10] , \wRegOut_4_3[9] , \wRegOut_4_3[8] , 
        \wRegOut_4_3[7] , \wRegOut_4_3[6] , \wRegOut_4_3[5] , \wRegOut_4_3[4] , 
        \wRegOut_4_3[3] , \wRegOut_4_3[2] , \wRegOut_4_3[1] , \wRegOut_4_3[0] 
        }), .Enable1(\wRegEnTop_4_3[0] ), .Enable2(\wRegEnBot_4_3[0] ), .In1({
        \wRegInTop_4_3[31] , \wRegInTop_4_3[30] , \wRegInTop_4_3[29] , 
        \wRegInTop_4_3[28] , \wRegInTop_4_3[27] , \wRegInTop_4_3[26] , 
        \wRegInTop_4_3[25] , \wRegInTop_4_3[24] , \wRegInTop_4_3[23] , 
        \wRegInTop_4_3[22] , \wRegInTop_4_3[21] , \wRegInTop_4_3[20] , 
        \wRegInTop_4_3[19] , \wRegInTop_4_3[18] , \wRegInTop_4_3[17] , 
        \wRegInTop_4_3[16] , \wRegInTop_4_3[15] , \wRegInTop_4_3[14] , 
        \wRegInTop_4_3[13] , \wRegInTop_4_3[12] , \wRegInTop_4_3[11] , 
        \wRegInTop_4_3[10] , \wRegInTop_4_3[9] , \wRegInTop_4_3[8] , 
        \wRegInTop_4_3[7] , \wRegInTop_4_3[6] , \wRegInTop_4_3[5] , 
        \wRegInTop_4_3[4] , \wRegInTop_4_3[3] , \wRegInTop_4_3[2] , 
        \wRegInTop_4_3[1] , \wRegInTop_4_3[0] }), .In2({\wRegInBot_4_3[31] , 
        \wRegInBot_4_3[30] , \wRegInBot_4_3[29] , \wRegInBot_4_3[28] , 
        \wRegInBot_4_3[27] , \wRegInBot_4_3[26] , \wRegInBot_4_3[25] , 
        \wRegInBot_4_3[24] , \wRegInBot_4_3[23] , \wRegInBot_4_3[22] , 
        \wRegInBot_4_3[21] , \wRegInBot_4_3[20] , \wRegInBot_4_3[19] , 
        \wRegInBot_4_3[18] , \wRegInBot_4_3[17] , \wRegInBot_4_3[16] , 
        \wRegInBot_4_3[15] , \wRegInBot_4_3[14] , \wRegInBot_4_3[13] , 
        \wRegInBot_4_3[12] , \wRegInBot_4_3[11] , \wRegInBot_4_3[10] , 
        \wRegInBot_4_3[9] , \wRegInBot_4_3[8] , \wRegInBot_4_3[7] , 
        \wRegInBot_4_3[6] , \wRegInBot_4_3[5] , \wRegInBot_4_3[4] , 
        \wRegInBot_4_3[3] , \wRegInBot_4_3[2] , \wRegInBot_4_3[1] , 
        \wRegInBot_4_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink35[31] , \ScanLink35[30] , \ScanLink35[29] , 
        \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , \ScanLink35[25] , 
        \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , \ScanLink35[21] , 
        \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , \ScanLink35[17] , 
        \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , \ScanLink35[13] , 
        \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , \ScanLink35[9] , 
        \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , \ScanLink35[5] , 
        \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , \ScanLink35[1] , 
        \ScanLink35[0] }), .ScanOut({\ScanLink34[31] , \ScanLink34[30] , 
        \ScanLink34[29] , \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , 
        \ScanLink34[25] , \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , 
        \ScanLink34[21] , \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , 
        \ScanLink34[17] , \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , 
        \ScanLink34[13] , \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , 
        \ScanLink34[9] , \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , 
        \ScanLink34[5] , \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , 
        \ScanLink34[1] , \ScanLink34[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_3[31] , \wRegOut_5_3[30] , \wRegOut_5_3[29] , 
        \wRegOut_5_3[28] , \wRegOut_5_3[27] , \wRegOut_5_3[26] , 
        \wRegOut_5_3[25] , \wRegOut_5_3[24] , \wRegOut_5_3[23] , 
        \wRegOut_5_3[22] , \wRegOut_5_3[21] , \wRegOut_5_3[20] , 
        \wRegOut_5_3[19] , \wRegOut_5_3[18] , \wRegOut_5_3[17] , 
        \wRegOut_5_3[16] , \wRegOut_5_3[15] , \wRegOut_5_3[14] , 
        \wRegOut_5_3[13] , \wRegOut_5_3[12] , \wRegOut_5_3[11] , 
        \wRegOut_5_3[10] , \wRegOut_5_3[9] , \wRegOut_5_3[8] , 
        \wRegOut_5_3[7] , \wRegOut_5_3[6] , \wRegOut_5_3[5] , \wRegOut_5_3[4] , 
        \wRegOut_5_3[3] , \wRegOut_5_3[2] , \wRegOut_5_3[1] , \wRegOut_5_3[0] 
        }), .Enable1(\wRegEnTop_5_3[0] ), .Enable2(\wRegEnBot_5_3[0] ), .In1({
        \wRegInTop_5_3[31] , \wRegInTop_5_3[30] , \wRegInTop_5_3[29] , 
        \wRegInTop_5_3[28] , \wRegInTop_5_3[27] , \wRegInTop_5_3[26] , 
        \wRegInTop_5_3[25] , \wRegInTop_5_3[24] , \wRegInTop_5_3[23] , 
        \wRegInTop_5_3[22] , \wRegInTop_5_3[21] , \wRegInTop_5_3[20] , 
        \wRegInTop_5_3[19] , \wRegInTop_5_3[18] , \wRegInTop_5_3[17] , 
        \wRegInTop_5_3[16] , \wRegInTop_5_3[15] , \wRegInTop_5_3[14] , 
        \wRegInTop_5_3[13] , \wRegInTop_5_3[12] , \wRegInTop_5_3[11] , 
        \wRegInTop_5_3[10] , \wRegInTop_5_3[9] , \wRegInTop_5_3[8] , 
        \wRegInTop_5_3[7] , \wRegInTop_5_3[6] , \wRegInTop_5_3[5] , 
        \wRegInTop_5_3[4] , \wRegInTop_5_3[3] , \wRegInTop_5_3[2] , 
        \wRegInTop_5_3[1] , \wRegInTop_5_3[0] }), .In2({\wRegInBot_5_3[31] , 
        \wRegInBot_5_3[30] , \wRegInBot_5_3[29] , \wRegInBot_5_3[28] , 
        \wRegInBot_5_3[27] , \wRegInBot_5_3[26] , \wRegInBot_5_3[25] , 
        \wRegInBot_5_3[24] , \wRegInBot_5_3[23] , \wRegInBot_5_3[22] , 
        \wRegInBot_5_3[21] , \wRegInBot_5_3[20] , \wRegInBot_5_3[19] , 
        \wRegInBot_5_3[18] , \wRegInBot_5_3[17] , \wRegInBot_5_3[16] , 
        \wRegInBot_5_3[15] , \wRegInBot_5_3[14] , \wRegInBot_5_3[13] , 
        \wRegInBot_5_3[12] , \wRegInBot_5_3[11] , \wRegInBot_5_3[10] , 
        \wRegInBot_5_3[9] , \wRegInBot_5_3[8] , \wRegInBot_5_3[7] , 
        \wRegInBot_5_3[6] , \wRegInBot_5_3[5] , \wRegInBot_5_3[4] , 
        \wRegInBot_5_3[3] , \wRegInBot_5_3[2] , \wRegInBot_5_3[1] , 
        \wRegInBot_5_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_22 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink54[31] , \ScanLink54[30] , \ScanLink54[29] , 
        \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , \ScanLink54[25] , 
        \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , \ScanLink54[21] , 
        \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , \ScanLink54[17] , 
        \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , \ScanLink54[13] , 
        \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , \ScanLink54[9] , 
        \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , \ScanLink54[5] , 
        \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , \ScanLink54[1] , 
        \ScanLink54[0] }), .ScanOut({\ScanLink53[31] , \ScanLink53[30] , 
        \ScanLink53[29] , \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , 
        \ScanLink53[25] , \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , 
        \ScanLink53[21] , \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , 
        \ScanLink53[17] , \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , 
        \ScanLink53[13] , \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , 
        \ScanLink53[9] , \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , 
        \ScanLink53[5] , \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , 
        \ScanLink53[1] , \ScanLink53[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_22[31] , \wRegOut_5_22[30] , 
        \wRegOut_5_22[29] , \wRegOut_5_22[28] , \wRegOut_5_22[27] , 
        \wRegOut_5_22[26] , \wRegOut_5_22[25] , \wRegOut_5_22[24] , 
        \wRegOut_5_22[23] , \wRegOut_5_22[22] , \wRegOut_5_22[21] , 
        \wRegOut_5_22[20] , \wRegOut_5_22[19] , \wRegOut_5_22[18] , 
        \wRegOut_5_22[17] , \wRegOut_5_22[16] , \wRegOut_5_22[15] , 
        \wRegOut_5_22[14] , \wRegOut_5_22[13] , \wRegOut_5_22[12] , 
        \wRegOut_5_22[11] , \wRegOut_5_22[10] , \wRegOut_5_22[9] , 
        \wRegOut_5_22[8] , \wRegOut_5_22[7] , \wRegOut_5_22[6] , 
        \wRegOut_5_22[5] , \wRegOut_5_22[4] , \wRegOut_5_22[3] , 
        \wRegOut_5_22[2] , \wRegOut_5_22[1] , \wRegOut_5_22[0] }), .Enable1(
        \wRegEnTop_5_22[0] ), .Enable2(\wRegEnBot_5_22[0] ), .In1({
        \wRegInTop_5_22[31] , \wRegInTop_5_22[30] , \wRegInTop_5_22[29] , 
        \wRegInTop_5_22[28] , \wRegInTop_5_22[27] , \wRegInTop_5_22[26] , 
        \wRegInTop_5_22[25] , \wRegInTop_5_22[24] , \wRegInTop_5_22[23] , 
        \wRegInTop_5_22[22] , \wRegInTop_5_22[21] , \wRegInTop_5_22[20] , 
        \wRegInTop_5_22[19] , \wRegInTop_5_22[18] , \wRegInTop_5_22[17] , 
        \wRegInTop_5_22[16] , \wRegInTop_5_22[15] , \wRegInTop_5_22[14] , 
        \wRegInTop_5_22[13] , \wRegInTop_5_22[12] , \wRegInTop_5_22[11] , 
        \wRegInTop_5_22[10] , \wRegInTop_5_22[9] , \wRegInTop_5_22[8] , 
        \wRegInTop_5_22[7] , \wRegInTop_5_22[6] , \wRegInTop_5_22[5] , 
        \wRegInTop_5_22[4] , \wRegInTop_5_22[3] , \wRegInTop_5_22[2] , 
        \wRegInTop_5_22[1] , \wRegInTop_5_22[0] }), .In2({\wRegInBot_5_22[31] , 
        \wRegInBot_5_22[30] , \wRegInBot_5_22[29] , \wRegInBot_5_22[28] , 
        \wRegInBot_5_22[27] , \wRegInBot_5_22[26] , \wRegInBot_5_22[25] , 
        \wRegInBot_5_22[24] , \wRegInBot_5_22[23] , \wRegInBot_5_22[22] , 
        \wRegInBot_5_22[21] , \wRegInBot_5_22[20] , \wRegInBot_5_22[19] , 
        \wRegInBot_5_22[18] , \wRegInBot_5_22[17] , \wRegInBot_5_22[16] , 
        \wRegInBot_5_22[15] , \wRegInBot_5_22[14] , \wRegInBot_5_22[13] , 
        \wRegInBot_5_22[12] , \wRegInBot_5_22[11] , \wRegInBot_5_22[10] , 
        \wRegInBot_5_22[9] , \wRegInBot_5_22[8] , \wRegInBot_5_22[7] , 
        \wRegInBot_5_22[6] , \wRegInBot_5_22[5] , \wRegInBot_5_22[4] , 
        \wRegInBot_5_22[3] , \wRegInBot_5_22[2] , \wRegInBot_5_22[1] , 
        \wRegInBot_5_22[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_66 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink194[31] , \ScanLink194[30] , \ScanLink194[29] , 
        \ScanLink194[28] , \ScanLink194[27] , \ScanLink194[26] , 
        \ScanLink194[25] , \ScanLink194[24] , \ScanLink194[23] , 
        \ScanLink194[22] , \ScanLink194[21] , \ScanLink194[20] , 
        \ScanLink194[19] , \ScanLink194[18] , \ScanLink194[17] , 
        \ScanLink194[16] , \ScanLink194[15] , \ScanLink194[14] , 
        \ScanLink194[13] , \ScanLink194[12] , \ScanLink194[11] , 
        \ScanLink194[10] , \ScanLink194[9] , \ScanLink194[8] , 
        \ScanLink194[7] , \ScanLink194[6] , \ScanLink194[5] , \ScanLink194[4] , 
        \ScanLink194[3] , \ScanLink194[2] , \ScanLink194[1] , \ScanLink194[0] 
        }), .ScanOut({\ScanLink193[31] , \ScanLink193[30] , \ScanLink193[29] , 
        \ScanLink193[28] , \ScanLink193[27] , \ScanLink193[26] , 
        \ScanLink193[25] , \ScanLink193[24] , \ScanLink193[23] , 
        \ScanLink193[22] , \ScanLink193[21] , \ScanLink193[20] , 
        \ScanLink193[19] , \ScanLink193[18] , \ScanLink193[17] , 
        \ScanLink193[16] , \ScanLink193[15] , \ScanLink193[14] , 
        \ScanLink193[13] , \ScanLink193[12] , \ScanLink193[11] , 
        \ScanLink193[10] , \ScanLink193[9] , \ScanLink193[8] , 
        \ScanLink193[7] , \ScanLink193[6] , \ScanLink193[5] , \ScanLink193[4] , 
        \ScanLink193[3] , \ScanLink193[2] , \ScanLink193[1] , \ScanLink193[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_66[31] , 
        \wRegOut_7_66[30] , \wRegOut_7_66[29] , \wRegOut_7_66[28] , 
        \wRegOut_7_66[27] , \wRegOut_7_66[26] , \wRegOut_7_66[25] , 
        \wRegOut_7_66[24] , \wRegOut_7_66[23] , \wRegOut_7_66[22] , 
        \wRegOut_7_66[21] , \wRegOut_7_66[20] , \wRegOut_7_66[19] , 
        \wRegOut_7_66[18] , \wRegOut_7_66[17] , \wRegOut_7_66[16] , 
        \wRegOut_7_66[15] , \wRegOut_7_66[14] , \wRegOut_7_66[13] , 
        \wRegOut_7_66[12] , \wRegOut_7_66[11] , \wRegOut_7_66[10] , 
        \wRegOut_7_66[9] , \wRegOut_7_66[8] , \wRegOut_7_66[7] , 
        \wRegOut_7_66[6] , \wRegOut_7_66[5] , \wRegOut_7_66[4] , 
        \wRegOut_7_66[3] , \wRegOut_7_66[2] , \wRegOut_7_66[1] , 
        \wRegOut_7_66[0] }), .Enable1(\wRegEnTop_7_66[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_66[31] , \wRegInTop_7_66[30] , \wRegInTop_7_66[29] , 
        \wRegInTop_7_66[28] , \wRegInTop_7_66[27] , \wRegInTop_7_66[26] , 
        \wRegInTop_7_66[25] , \wRegInTop_7_66[24] , \wRegInTop_7_66[23] , 
        \wRegInTop_7_66[22] , \wRegInTop_7_66[21] , \wRegInTop_7_66[20] , 
        \wRegInTop_7_66[19] , \wRegInTop_7_66[18] , \wRegInTop_7_66[17] , 
        \wRegInTop_7_66[16] , \wRegInTop_7_66[15] , \wRegInTop_7_66[14] , 
        \wRegInTop_7_66[13] , \wRegInTop_7_66[12] , \wRegInTop_7_66[11] , 
        \wRegInTop_7_66[10] , \wRegInTop_7_66[9] , \wRegInTop_7_66[8] , 
        \wRegInTop_7_66[7] , \wRegInTop_7_66[6] , \wRegInTop_7_66[5] , 
        \wRegInTop_7_66[4] , \wRegInTop_7_66[3] , \wRegInTop_7_66[2] , 
        \wRegInTop_7_66[1] , \wRegInTop_7_66[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink76[31] , \ScanLink76[30] , \ScanLink76[29] , 
        \ScanLink76[28] , \ScanLink76[27] , \ScanLink76[26] , \ScanLink76[25] , 
        \ScanLink76[24] , \ScanLink76[23] , \ScanLink76[22] , \ScanLink76[21] , 
        \ScanLink76[20] , \ScanLink76[19] , \ScanLink76[18] , \ScanLink76[17] , 
        \ScanLink76[16] , \ScanLink76[15] , \ScanLink76[14] , \ScanLink76[13] , 
        \ScanLink76[12] , \ScanLink76[11] , \ScanLink76[10] , \ScanLink76[9] , 
        \ScanLink76[8] , \ScanLink76[7] , \ScanLink76[6] , \ScanLink76[5] , 
        \ScanLink76[4] , \ScanLink76[3] , \ScanLink76[2] , \ScanLink76[1] , 
        \ScanLink76[0] }), .ScanOut({\ScanLink75[31] , \ScanLink75[30] , 
        \ScanLink75[29] , \ScanLink75[28] , \ScanLink75[27] , \ScanLink75[26] , 
        \ScanLink75[25] , \ScanLink75[24] , \ScanLink75[23] , \ScanLink75[22] , 
        \ScanLink75[21] , \ScanLink75[20] , \ScanLink75[19] , \ScanLink75[18] , 
        \ScanLink75[17] , \ScanLink75[16] , \ScanLink75[15] , \ScanLink75[14] , 
        \ScanLink75[13] , \ScanLink75[12] , \ScanLink75[11] , \ScanLink75[10] , 
        \ScanLink75[9] , \ScanLink75[8] , \ScanLink75[7] , \ScanLink75[6] , 
        \ScanLink75[5] , \ScanLink75[4] , \ScanLink75[3] , \ScanLink75[2] , 
        \ScanLink75[1] , \ScanLink75[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_12[31] , \wRegOut_6_12[30] , 
        \wRegOut_6_12[29] , \wRegOut_6_12[28] , \wRegOut_6_12[27] , 
        \wRegOut_6_12[26] , \wRegOut_6_12[25] , \wRegOut_6_12[24] , 
        \wRegOut_6_12[23] , \wRegOut_6_12[22] , \wRegOut_6_12[21] , 
        \wRegOut_6_12[20] , \wRegOut_6_12[19] , \wRegOut_6_12[18] , 
        \wRegOut_6_12[17] , \wRegOut_6_12[16] , \wRegOut_6_12[15] , 
        \wRegOut_6_12[14] , \wRegOut_6_12[13] , \wRegOut_6_12[12] , 
        \wRegOut_6_12[11] , \wRegOut_6_12[10] , \wRegOut_6_12[9] , 
        \wRegOut_6_12[8] , \wRegOut_6_12[7] , \wRegOut_6_12[6] , 
        \wRegOut_6_12[5] , \wRegOut_6_12[4] , \wRegOut_6_12[3] , 
        \wRegOut_6_12[2] , \wRegOut_6_12[1] , \wRegOut_6_12[0] }), .Enable1(
        \wRegEnTop_6_12[0] ), .Enable2(\wRegEnBot_6_12[0] ), .In1({
        \wRegInTop_6_12[31] , \wRegInTop_6_12[30] , \wRegInTop_6_12[29] , 
        \wRegInTop_6_12[28] , \wRegInTop_6_12[27] , \wRegInTop_6_12[26] , 
        \wRegInTop_6_12[25] , \wRegInTop_6_12[24] , \wRegInTop_6_12[23] , 
        \wRegInTop_6_12[22] , \wRegInTop_6_12[21] , \wRegInTop_6_12[20] , 
        \wRegInTop_6_12[19] , \wRegInTop_6_12[18] , \wRegInTop_6_12[17] , 
        \wRegInTop_6_12[16] , \wRegInTop_6_12[15] , \wRegInTop_6_12[14] , 
        \wRegInTop_6_12[13] , \wRegInTop_6_12[12] , \wRegInTop_6_12[11] , 
        \wRegInTop_6_12[10] , \wRegInTop_6_12[9] , \wRegInTop_6_12[8] , 
        \wRegInTop_6_12[7] , \wRegInTop_6_12[6] , \wRegInTop_6_12[5] , 
        \wRegInTop_6_12[4] , \wRegInTop_6_12[3] , \wRegInTop_6_12[2] , 
        \wRegInTop_6_12[1] , \wRegInTop_6_12[0] }), .In2({\wRegInBot_6_12[31] , 
        \wRegInBot_6_12[30] , \wRegInBot_6_12[29] , \wRegInBot_6_12[28] , 
        \wRegInBot_6_12[27] , \wRegInBot_6_12[26] , \wRegInBot_6_12[25] , 
        \wRegInBot_6_12[24] , \wRegInBot_6_12[23] , \wRegInBot_6_12[22] , 
        \wRegInBot_6_12[21] , \wRegInBot_6_12[20] , \wRegInBot_6_12[19] , 
        \wRegInBot_6_12[18] , \wRegInBot_6_12[17] , \wRegInBot_6_12[16] , 
        \wRegInBot_6_12[15] , \wRegInBot_6_12[14] , \wRegInBot_6_12[13] , 
        \wRegInBot_6_12[12] , \wRegInBot_6_12[11] , \wRegInBot_6_12[10] , 
        \wRegInBot_6_12[9] , \wRegInBot_6_12[8] , \wRegInBot_6_12[7] , 
        \wRegInBot_6_12[6] , \wRegInBot_6_12[5] , \wRegInBot_6_12[4] , 
        \wRegInBot_6_12[3] , \wRegInBot_6_12[2] , \wRegInBot_6_12[1] , 
        \wRegInBot_6_12[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_35 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink99[31] , \ScanLink99[30] , \ScanLink99[29] , 
        \ScanLink99[28] , \ScanLink99[27] , \ScanLink99[26] , \ScanLink99[25] , 
        \ScanLink99[24] , \ScanLink99[23] , \ScanLink99[22] , \ScanLink99[21] , 
        \ScanLink99[20] , \ScanLink99[19] , \ScanLink99[18] , \ScanLink99[17] , 
        \ScanLink99[16] , \ScanLink99[15] , \ScanLink99[14] , \ScanLink99[13] , 
        \ScanLink99[12] , \ScanLink99[11] , \ScanLink99[10] , \ScanLink99[9] , 
        \ScanLink99[8] , \ScanLink99[7] , \ScanLink99[6] , \ScanLink99[5] , 
        \ScanLink99[4] , \ScanLink99[3] , \ScanLink99[2] , \ScanLink99[1] , 
        \ScanLink99[0] }), .ScanOut({\ScanLink98[31] , \ScanLink98[30] , 
        \ScanLink98[29] , \ScanLink98[28] , \ScanLink98[27] , \ScanLink98[26] , 
        \ScanLink98[25] , \ScanLink98[24] , \ScanLink98[23] , \ScanLink98[22] , 
        \ScanLink98[21] , \ScanLink98[20] , \ScanLink98[19] , \ScanLink98[18] , 
        \ScanLink98[17] , \ScanLink98[16] , \ScanLink98[15] , \ScanLink98[14] , 
        \ScanLink98[13] , \ScanLink98[12] , \ScanLink98[11] , \ScanLink98[10] , 
        \ScanLink98[9] , \ScanLink98[8] , \ScanLink98[7] , \ScanLink98[6] , 
        \ScanLink98[5] , \ScanLink98[4] , \ScanLink98[3] , \ScanLink98[2] , 
        \ScanLink98[1] , \ScanLink98[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_35[31] , \wRegOut_6_35[30] , 
        \wRegOut_6_35[29] , \wRegOut_6_35[28] , \wRegOut_6_35[27] , 
        \wRegOut_6_35[26] , \wRegOut_6_35[25] , \wRegOut_6_35[24] , 
        \wRegOut_6_35[23] , \wRegOut_6_35[22] , \wRegOut_6_35[21] , 
        \wRegOut_6_35[20] , \wRegOut_6_35[19] , \wRegOut_6_35[18] , 
        \wRegOut_6_35[17] , \wRegOut_6_35[16] , \wRegOut_6_35[15] , 
        \wRegOut_6_35[14] , \wRegOut_6_35[13] , \wRegOut_6_35[12] , 
        \wRegOut_6_35[11] , \wRegOut_6_35[10] , \wRegOut_6_35[9] , 
        \wRegOut_6_35[8] , \wRegOut_6_35[7] , \wRegOut_6_35[6] , 
        \wRegOut_6_35[5] , \wRegOut_6_35[4] , \wRegOut_6_35[3] , 
        \wRegOut_6_35[2] , \wRegOut_6_35[1] , \wRegOut_6_35[0] }), .Enable1(
        \wRegEnTop_6_35[0] ), .Enable2(\wRegEnBot_6_35[0] ), .In1({
        \wRegInTop_6_35[31] , \wRegInTop_6_35[30] , \wRegInTop_6_35[29] , 
        \wRegInTop_6_35[28] , \wRegInTop_6_35[27] , \wRegInTop_6_35[26] , 
        \wRegInTop_6_35[25] , \wRegInTop_6_35[24] , \wRegInTop_6_35[23] , 
        \wRegInTop_6_35[22] , \wRegInTop_6_35[21] , \wRegInTop_6_35[20] , 
        \wRegInTop_6_35[19] , \wRegInTop_6_35[18] , \wRegInTop_6_35[17] , 
        \wRegInTop_6_35[16] , \wRegInTop_6_35[15] , \wRegInTop_6_35[14] , 
        \wRegInTop_6_35[13] , \wRegInTop_6_35[12] , \wRegInTop_6_35[11] , 
        \wRegInTop_6_35[10] , \wRegInTop_6_35[9] , \wRegInTop_6_35[8] , 
        \wRegInTop_6_35[7] , \wRegInTop_6_35[6] , \wRegInTop_6_35[5] , 
        \wRegInTop_6_35[4] , \wRegInTop_6_35[3] , \wRegInTop_6_35[2] , 
        \wRegInTop_6_35[1] , \wRegInTop_6_35[0] }), .In2({\wRegInBot_6_35[31] , 
        \wRegInBot_6_35[30] , \wRegInBot_6_35[29] , \wRegInBot_6_35[28] , 
        \wRegInBot_6_35[27] , \wRegInBot_6_35[26] , \wRegInBot_6_35[25] , 
        \wRegInBot_6_35[24] , \wRegInBot_6_35[23] , \wRegInBot_6_35[22] , 
        \wRegInBot_6_35[21] , \wRegInBot_6_35[20] , \wRegInBot_6_35[19] , 
        \wRegInBot_6_35[18] , \wRegInBot_6_35[17] , \wRegInBot_6_35[16] , 
        \wRegInBot_6_35[15] , \wRegInBot_6_35[14] , \wRegInBot_6_35[13] , 
        \wRegInBot_6_35[12] , \wRegInBot_6_35[11] , \wRegInBot_6_35[10] , 
        \wRegInBot_6_35[9] , \wRegInBot_6_35[8] , \wRegInBot_6_35[7] , 
        \wRegInBot_6_35[6] , \wRegInBot_6_35[5] , \wRegInBot_6_35[4] , 
        \wRegInBot_6_35[3] , \wRegInBot_6_35[2] , \wRegInBot_6_35[1] , 
        \wRegInBot_6_35[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink135[31] , \ScanLink135[30] , \ScanLink135[29] , 
        \ScanLink135[28] , \ScanLink135[27] , \ScanLink135[26] , 
        \ScanLink135[25] , \ScanLink135[24] , \ScanLink135[23] , 
        \ScanLink135[22] , \ScanLink135[21] , \ScanLink135[20] , 
        \ScanLink135[19] , \ScanLink135[18] , \ScanLink135[17] , 
        \ScanLink135[16] , \ScanLink135[15] , \ScanLink135[14] , 
        \ScanLink135[13] , \ScanLink135[12] , \ScanLink135[11] , 
        \ScanLink135[10] , \ScanLink135[9] , \ScanLink135[8] , 
        \ScanLink135[7] , \ScanLink135[6] , \ScanLink135[5] , \ScanLink135[4] , 
        \ScanLink135[3] , \ScanLink135[2] , \ScanLink135[1] , \ScanLink135[0] 
        }), .ScanOut({\ScanLink134[31] , \ScanLink134[30] , \ScanLink134[29] , 
        \ScanLink134[28] , \ScanLink134[27] , \ScanLink134[26] , 
        \ScanLink134[25] , \ScanLink134[24] , \ScanLink134[23] , 
        \ScanLink134[22] , \ScanLink134[21] , \ScanLink134[20] , 
        \ScanLink134[19] , \ScanLink134[18] , \ScanLink134[17] , 
        \ScanLink134[16] , \ScanLink134[15] , \ScanLink134[14] , 
        \ScanLink134[13] , \ScanLink134[12] , \ScanLink134[11] , 
        \ScanLink134[10] , \ScanLink134[9] , \ScanLink134[8] , 
        \ScanLink134[7] , \ScanLink134[6] , \ScanLink134[5] , \ScanLink134[4] , 
        \ScanLink134[3] , \ScanLink134[2] , \ScanLink134[1] , \ScanLink134[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_7[31] , 
        \wRegOut_7_7[30] , \wRegOut_7_7[29] , \wRegOut_7_7[28] , 
        \wRegOut_7_7[27] , \wRegOut_7_7[26] , \wRegOut_7_7[25] , 
        \wRegOut_7_7[24] , \wRegOut_7_7[23] , \wRegOut_7_7[22] , 
        \wRegOut_7_7[21] , \wRegOut_7_7[20] , \wRegOut_7_7[19] , 
        \wRegOut_7_7[18] , \wRegOut_7_7[17] , \wRegOut_7_7[16] , 
        \wRegOut_7_7[15] , \wRegOut_7_7[14] , \wRegOut_7_7[13] , 
        \wRegOut_7_7[12] , \wRegOut_7_7[11] , \wRegOut_7_7[10] , 
        \wRegOut_7_7[9] , \wRegOut_7_7[8] , \wRegOut_7_7[7] , \wRegOut_7_7[6] , 
        \wRegOut_7_7[5] , \wRegOut_7_7[4] , \wRegOut_7_7[3] , \wRegOut_7_7[2] , 
        \wRegOut_7_7[1] , \wRegOut_7_7[0] }), .Enable1(\wRegEnTop_7_7[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_7[31] , \wRegInTop_7_7[30] , 
        \wRegInTop_7_7[29] , \wRegInTop_7_7[28] , \wRegInTop_7_7[27] , 
        \wRegInTop_7_7[26] , \wRegInTop_7_7[25] , \wRegInTop_7_7[24] , 
        \wRegInTop_7_7[23] , \wRegInTop_7_7[22] , \wRegInTop_7_7[21] , 
        \wRegInTop_7_7[20] , \wRegInTop_7_7[19] , \wRegInTop_7_7[18] , 
        \wRegInTop_7_7[17] , \wRegInTop_7_7[16] , \wRegInTop_7_7[15] , 
        \wRegInTop_7_7[14] , \wRegInTop_7_7[13] , \wRegInTop_7_7[12] , 
        \wRegInTop_7_7[11] , \wRegInTop_7_7[10] , \wRegInTop_7_7[9] , 
        \wRegInTop_7_7[8] , \wRegInTop_7_7[7] , \wRegInTop_7_7[6] , 
        \wRegInTop_7_7[5] , \wRegInTop_7_7[4] , \wRegInTop_7_7[3] , 
        \wRegInTop_7_7[2] , \wRegInTop_7_7[1] , \wRegInTop_7_7[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_41 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink169[31] , \ScanLink169[30] , \ScanLink169[29] , 
        \ScanLink169[28] , \ScanLink169[27] , \ScanLink169[26] , 
        \ScanLink169[25] , \ScanLink169[24] , \ScanLink169[23] , 
        \ScanLink169[22] , \ScanLink169[21] , \ScanLink169[20] , 
        \ScanLink169[19] , \ScanLink169[18] , \ScanLink169[17] , 
        \ScanLink169[16] , \ScanLink169[15] , \ScanLink169[14] , 
        \ScanLink169[13] , \ScanLink169[12] , \ScanLink169[11] , 
        \ScanLink169[10] , \ScanLink169[9] , \ScanLink169[8] , 
        \ScanLink169[7] , \ScanLink169[6] , \ScanLink169[5] , \ScanLink169[4] , 
        \ScanLink169[3] , \ScanLink169[2] , \ScanLink169[1] , \ScanLink169[0] 
        }), .ScanOut({\ScanLink168[31] , \ScanLink168[30] , \ScanLink168[29] , 
        \ScanLink168[28] , \ScanLink168[27] , \ScanLink168[26] , 
        \ScanLink168[25] , \ScanLink168[24] , \ScanLink168[23] , 
        \ScanLink168[22] , \ScanLink168[21] , \ScanLink168[20] , 
        \ScanLink168[19] , \ScanLink168[18] , \ScanLink168[17] , 
        \ScanLink168[16] , \ScanLink168[15] , \ScanLink168[14] , 
        \ScanLink168[13] , \ScanLink168[12] , \ScanLink168[11] , 
        \ScanLink168[10] , \ScanLink168[9] , \ScanLink168[8] , 
        \ScanLink168[7] , \ScanLink168[6] , \ScanLink168[5] , \ScanLink168[4] , 
        \ScanLink168[3] , \ScanLink168[2] , \ScanLink168[1] , \ScanLink168[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_41[31] , 
        \wRegOut_7_41[30] , \wRegOut_7_41[29] , \wRegOut_7_41[28] , 
        \wRegOut_7_41[27] , \wRegOut_7_41[26] , \wRegOut_7_41[25] , 
        \wRegOut_7_41[24] , \wRegOut_7_41[23] , \wRegOut_7_41[22] , 
        \wRegOut_7_41[21] , \wRegOut_7_41[20] , \wRegOut_7_41[19] , 
        \wRegOut_7_41[18] , \wRegOut_7_41[17] , \wRegOut_7_41[16] , 
        \wRegOut_7_41[15] , \wRegOut_7_41[14] , \wRegOut_7_41[13] , 
        \wRegOut_7_41[12] , \wRegOut_7_41[11] , \wRegOut_7_41[10] , 
        \wRegOut_7_41[9] , \wRegOut_7_41[8] , \wRegOut_7_41[7] , 
        \wRegOut_7_41[6] , \wRegOut_7_41[5] , \wRegOut_7_41[4] , 
        \wRegOut_7_41[3] , \wRegOut_7_41[2] , \wRegOut_7_41[1] , 
        \wRegOut_7_41[0] }), .Enable1(\wRegEnTop_7_41[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_41[31] , \wRegInTop_7_41[30] , \wRegInTop_7_41[29] , 
        \wRegInTop_7_41[28] , \wRegInTop_7_41[27] , \wRegInTop_7_41[26] , 
        \wRegInTop_7_41[25] , \wRegInTop_7_41[24] , \wRegInTop_7_41[23] , 
        \wRegInTop_7_41[22] , \wRegInTop_7_41[21] , \wRegInTop_7_41[20] , 
        \wRegInTop_7_41[19] , \wRegInTop_7_41[18] , \wRegInTop_7_41[17] , 
        \wRegInTop_7_41[16] , \wRegInTop_7_41[15] , \wRegInTop_7_41[14] , 
        \wRegInTop_7_41[13] , \wRegInTop_7_41[12] , \wRegInTop_7_41[11] , 
        \wRegInTop_7_41[10] , \wRegInTop_7_41[9] , \wRegInTop_7_41[8] , 
        \wRegInTop_7_41[7] , \wRegInTop_7_41[6] , \wRegInTop_7_41[5] , 
        \wRegInTop_7_41[4] , \wRegInTop_7_41[3] , \wRegInTop_7_41[2] , 
        \wRegInTop_7_41[1] , \wRegInTop_7_41[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_48 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink112[31] , \ScanLink112[30] , \ScanLink112[29] , 
        \ScanLink112[28] , \ScanLink112[27] , \ScanLink112[26] , 
        \ScanLink112[25] , \ScanLink112[24] , \ScanLink112[23] , 
        \ScanLink112[22] , \ScanLink112[21] , \ScanLink112[20] , 
        \ScanLink112[19] , \ScanLink112[18] , \ScanLink112[17] , 
        \ScanLink112[16] , \ScanLink112[15] , \ScanLink112[14] , 
        \ScanLink112[13] , \ScanLink112[12] , \ScanLink112[11] , 
        \ScanLink112[10] , \ScanLink112[9] , \ScanLink112[8] , 
        \ScanLink112[7] , \ScanLink112[6] , \ScanLink112[5] , \ScanLink112[4] , 
        \ScanLink112[3] , \ScanLink112[2] , \ScanLink112[1] , \ScanLink112[0] 
        }), .ScanOut({\ScanLink111[31] , \ScanLink111[30] , \ScanLink111[29] , 
        \ScanLink111[28] , \ScanLink111[27] , \ScanLink111[26] , 
        \ScanLink111[25] , \ScanLink111[24] , \ScanLink111[23] , 
        \ScanLink111[22] , \ScanLink111[21] , \ScanLink111[20] , 
        \ScanLink111[19] , \ScanLink111[18] , \ScanLink111[17] , 
        \ScanLink111[16] , \ScanLink111[15] , \ScanLink111[14] , 
        \ScanLink111[13] , \ScanLink111[12] , \ScanLink111[11] , 
        \ScanLink111[10] , \ScanLink111[9] , \ScanLink111[8] , 
        \ScanLink111[7] , \ScanLink111[6] , \ScanLink111[5] , \ScanLink111[4] , 
        \ScanLink111[3] , \ScanLink111[2] , \ScanLink111[1] , \ScanLink111[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_48[31] , 
        \wRegOut_6_48[30] , \wRegOut_6_48[29] , \wRegOut_6_48[28] , 
        \wRegOut_6_48[27] , \wRegOut_6_48[26] , \wRegOut_6_48[25] , 
        \wRegOut_6_48[24] , \wRegOut_6_48[23] , \wRegOut_6_48[22] , 
        \wRegOut_6_48[21] , \wRegOut_6_48[20] , \wRegOut_6_48[19] , 
        \wRegOut_6_48[18] , \wRegOut_6_48[17] , \wRegOut_6_48[16] , 
        \wRegOut_6_48[15] , \wRegOut_6_48[14] , \wRegOut_6_48[13] , 
        \wRegOut_6_48[12] , \wRegOut_6_48[11] , \wRegOut_6_48[10] , 
        \wRegOut_6_48[9] , \wRegOut_6_48[8] , \wRegOut_6_48[7] , 
        \wRegOut_6_48[6] , \wRegOut_6_48[5] , \wRegOut_6_48[4] , 
        \wRegOut_6_48[3] , \wRegOut_6_48[2] , \wRegOut_6_48[1] , 
        \wRegOut_6_48[0] }), .Enable1(\wRegEnTop_6_48[0] ), .Enable2(
        \wRegEnBot_6_48[0] ), .In1({\wRegInTop_6_48[31] , \wRegInTop_6_48[30] , 
        \wRegInTop_6_48[29] , \wRegInTop_6_48[28] , \wRegInTop_6_48[27] , 
        \wRegInTop_6_48[26] , \wRegInTop_6_48[25] , \wRegInTop_6_48[24] , 
        \wRegInTop_6_48[23] , \wRegInTop_6_48[22] , \wRegInTop_6_48[21] , 
        \wRegInTop_6_48[20] , \wRegInTop_6_48[19] , \wRegInTop_6_48[18] , 
        \wRegInTop_6_48[17] , \wRegInTop_6_48[16] , \wRegInTop_6_48[15] , 
        \wRegInTop_6_48[14] , \wRegInTop_6_48[13] , \wRegInTop_6_48[12] , 
        \wRegInTop_6_48[11] , \wRegInTop_6_48[10] , \wRegInTop_6_48[9] , 
        \wRegInTop_6_48[8] , \wRegInTop_6_48[7] , \wRegInTop_6_48[6] , 
        \wRegInTop_6_48[5] , \wRegInTop_6_48[4] , \wRegInTop_6_48[3] , 
        \wRegInTop_6_48[2] , \wRegInTop_6_48[1] , \wRegInTop_6_48[0] }), .In2(
        {\wRegInBot_6_48[31] , \wRegInBot_6_48[30] , \wRegInBot_6_48[29] , 
        \wRegInBot_6_48[28] , \wRegInBot_6_48[27] , \wRegInBot_6_48[26] , 
        \wRegInBot_6_48[25] , \wRegInBot_6_48[24] , \wRegInBot_6_48[23] , 
        \wRegInBot_6_48[22] , \wRegInBot_6_48[21] , \wRegInBot_6_48[20] , 
        \wRegInBot_6_48[19] , \wRegInBot_6_48[18] , \wRegInBot_6_48[17] , 
        \wRegInBot_6_48[16] , \wRegInBot_6_48[15] , \wRegInBot_6_48[14] , 
        \wRegInBot_6_48[13] , \wRegInBot_6_48[12] , \wRegInBot_6_48[11] , 
        \wRegInBot_6_48[10] , \wRegInBot_6_48[9] , \wRegInBot_6_48[8] , 
        \wRegInBot_6_48[7] , \wRegInBot_6_48[6] , \wRegInBot_6_48[5] , 
        \wRegInBot_6_48[4] , \wRegInBot_6_48[3] , \wRegInBot_6_48[2] , 
        \wRegInBot_6_48[1] , \wRegInBot_6_48[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_53 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink117[31] , \ScanLink117[30] , \ScanLink117[29] , 
        \ScanLink117[28] , \ScanLink117[27] , \ScanLink117[26] , 
        \ScanLink117[25] , \ScanLink117[24] , \ScanLink117[23] , 
        \ScanLink117[22] , \ScanLink117[21] , \ScanLink117[20] , 
        \ScanLink117[19] , \ScanLink117[18] , \ScanLink117[17] , 
        \ScanLink117[16] , \ScanLink117[15] , \ScanLink117[14] , 
        \ScanLink117[13] , \ScanLink117[12] , \ScanLink117[11] , 
        \ScanLink117[10] , \ScanLink117[9] , \ScanLink117[8] , 
        \ScanLink117[7] , \ScanLink117[6] , \ScanLink117[5] , \ScanLink117[4] , 
        \ScanLink117[3] , \ScanLink117[2] , \ScanLink117[1] , \ScanLink117[0] 
        }), .ScanOut({\ScanLink116[31] , \ScanLink116[30] , \ScanLink116[29] , 
        \ScanLink116[28] , \ScanLink116[27] , \ScanLink116[26] , 
        \ScanLink116[25] , \ScanLink116[24] , \ScanLink116[23] , 
        \ScanLink116[22] , \ScanLink116[21] , \ScanLink116[20] , 
        \ScanLink116[19] , \ScanLink116[18] , \ScanLink116[17] , 
        \ScanLink116[16] , \ScanLink116[15] , \ScanLink116[14] , 
        \ScanLink116[13] , \ScanLink116[12] , \ScanLink116[11] , 
        \ScanLink116[10] , \ScanLink116[9] , \ScanLink116[8] , 
        \ScanLink116[7] , \ScanLink116[6] , \ScanLink116[5] , \ScanLink116[4] , 
        \ScanLink116[3] , \ScanLink116[2] , \ScanLink116[1] , \ScanLink116[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_53[31] , 
        \wRegOut_6_53[30] , \wRegOut_6_53[29] , \wRegOut_6_53[28] , 
        \wRegOut_6_53[27] , \wRegOut_6_53[26] , \wRegOut_6_53[25] , 
        \wRegOut_6_53[24] , \wRegOut_6_53[23] , \wRegOut_6_53[22] , 
        \wRegOut_6_53[21] , \wRegOut_6_53[20] , \wRegOut_6_53[19] , 
        \wRegOut_6_53[18] , \wRegOut_6_53[17] , \wRegOut_6_53[16] , 
        \wRegOut_6_53[15] , \wRegOut_6_53[14] , \wRegOut_6_53[13] , 
        \wRegOut_6_53[12] , \wRegOut_6_53[11] , \wRegOut_6_53[10] , 
        \wRegOut_6_53[9] , \wRegOut_6_53[8] , \wRegOut_6_53[7] , 
        \wRegOut_6_53[6] , \wRegOut_6_53[5] , \wRegOut_6_53[4] , 
        \wRegOut_6_53[3] , \wRegOut_6_53[2] , \wRegOut_6_53[1] , 
        \wRegOut_6_53[0] }), .Enable1(\wRegEnTop_6_53[0] ), .Enable2(
        \wRegEnBot_6_53[0] ), .In1({\wRegInTop_6_53[31] , \wRegInTop_6_53[30] , 
        \wRegInTop_6_53[29] , \wRegInTop_6_53[28] , \wRegInTop_6_53[27] , 
        \wRegInTop_6_53[26] , \wRegInTop_6_53[25] , \wRegInTop_6_53[24] , 
        \wRegInTop_6_53[23] , \wRegInTop_6_53[22] , \wRegInTop_6_53[21] , 
        \wRegInTop_6_53[20] , \wRegInTop_6_53[19] , \wRegInTop_6_53[18] , 
        \wRegInTop_6_53[17] , \wRegInTop_6_53[16] , \wRegInTop_6_53[15] , 
        \wRegInTop_6_53[14] , \wRegInTop_6_53[13] , \wRegInTop_6_53[12] , 
        \wRegInTop_6_53[11] , \wRegInTop_6_53[10] , \wRegInTop_6_53[9] , 
        \wRegInTop_6_53[8] , \wRegInTop_6_53[7] , \wRegInTop_6_53[6] , 
        \wRegInTop_6_53[5] , \wRegInTop_6_53[4] , \wRegInTop_6_53[3] , 
        \wRegInTop_6_53[2] , \wRegInTop_6_53[1] , \wRegInTop_6_53[0] }), .In2(
        {\wRegInBot_6_53[31] , \wRegInBot_6_53[30] , \wRegInBot_6_53[29] , 
        \wRegInBot_6_53[28] , \wRegInBot_6_53[27] , \wRegInBot_6_53[26] , 
        \wRegInBot_6_53[25] , \wRegInBot_6_53[24] , \wRegInBot_6_53[23] , 
        \wRegInBot_6_53[22] , \wRegInBot_6_53[21] , \wRegInBot_6_53[20] , 
        \wRegInBot_6_53[19] , \wRegInBot_6_53[18] , \wRegInBot_6_53[17] , 
        \wRegInBot_6_53[16] , \wRegInBot_6_53[15] , \wRegInBot_6_53[14] , 
        \wRegInBot_6_53[13] , \wRegInBot_6_53[12] , \wRegInBot_6_53[11] , 
        \wRegInBot_6_53[10] , \wRegInBot_6_53[9] , \wRegInBot_6_53[8] , 
        \wRegInBot_6_53[7] , \wRegInBot_6_53[6] , \wRegInBot_6_53[5] , 
        \wRegInBot_6_53[4] , \wRegInBot_6_53[3] , \wRegInBot_6_53[2] , 
        \wRegInBot_6_53[1] , \wRegInBot_6_53[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_27 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink155[31] , \ScanLink155[30] , \ScanLink155[29] , 
        \ScanLink155[28] , \ScanLink155[27] , \ScanLink155[26] , 
        \ScanLink155[25] , \ScanLink155[24] , \ScanLink155[23] , 
        \ScanLink155[22] , \ScanLink155[21] , \ScanLink155[20] , 
        \ScanLink155[19] , \ScanLink155[18] , \ScanLink155[17] , 
        \ScanLink155[16] , \ScanLink155[15] , \ScanLink155[14] , 
        \ScanLink155[13] , \ScanLink155[12] , \ScanLink155[11] , 
        \ScanLink155[10] , \ScanLink155[9] , \ScanLink155[8] , 
        \ScanLink155[7] , \ScanLink155[6] , \ScanLink155[5] , \ScanLink155[4] , 
        \ScanLink155[3] , \ScanLink155[2] , \ScanLink155[1] , \ScanLink155[0] 
        }), .ScanOut({\ScanLink154[31] , \ScanLink154[30] , \ScanLink154[29] , 
        \ScanLink154[28] , \ScanLink154[27] , \ScanLink154[26] , 
        \ScanLink154[25] , \ScanLink154[24] , \ScanLink154[23] , 
        \ScanLink154[22] , \ScanLink154[21] , \ScanLink154[20] , 
        \ScanLink154[19] , \ScanLink154[18] , \ScanLink154[17] , 
        \ScanLink154[16] , \ScanLink154[15] , \ScanLink154[14] , 
        \ScanLink154[13] , \ScanLink154[12] , \ScanLink154[11] , 
        \ScanLink154[10] , \ScanLink154[9] , \ScanLink154[8] , 
        \ScanLink154[7] , \ScanLink154[6] , \ScanLink154[5] , \ScanLink154[4] , 
        \ScanLink154[3] , \ScanLink154[2] , \ScanLink154[1] , \ScanLink154[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_27[31] , 
        \wRegOut_7_27[30] , \wRegOut_7_27[29] , \wRegOut_7_27[28] , 
        \wRegOut_7_27[27] , \wRegOut_7_27[26] , \wRegOut_7_27[25] , 
        \wRegOut_7_27[24] , \wRegOut_7_27[23] , \wRegOut_7_27[22] , 
        \wRegOut_7_27[21] , \wRegOut_7_27[20] , \wRegOut_7_27[19] , 
        \wRegOut_7_27[18] , \wRegOut_7_27[17] , \wRegOut_7_27[16] , 
        \wRegOut_7_27[15] , \wRegOut_7_27[14] , \wRegOut_7_27[13] , 
        \wRegOut_7_27[12] , \wRegOut_7_27[11] , \wRegOut_7_27[10] , 
        \wRegOut_7_27[9] , \wRegOut_7_27[8] , \wRegOut_7_27[7] , 
        \wRegOut_7_27[6] , \wRegOut_7_27[5] , \wRegOut_7_27[4] , 
        \wRegOut_7_27[3] , \wRegOut_7_27[2] , \wRegOut_7_27[1] , 
        \wRegOut_7_27[0] }), .Enable1(\wRegEnTop_7_27[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_27[31] , \wRegInTop_7_27[30] , \wRegInTop_7_27[29] , 
        \wRegInTop_7_27[28] , \wRegInTop_7_27[27] , \wRegInTop_7_27[26] , 
        \wRegInTop_7_27[25] , \wRegInTop_7_27[24] , \wRegInTop_7_27[23] , 
        \wRegInTop_7_27[22] , \wRegInTop_7_27[21] , \wRegInTop_7_27[20] , 
        \wRegInTop_7_27[19] , \wRegInTop_7_27[18] , \wRegInTop_7_27[17] , 
        \wRegInTop_7_27[16] , \wRegInTop_7_27[15] , \wRegInTop_7_27[14] , 
        \wRegInTop_7_27[13] , \wRegInTop_7_27[12] , \wRegInTop_7_27[11] , 
        \wRegInTop_7_27[10] , \wRegInTop_7_27[9] , \wRegInTop_7_27[8] , 
        \wRegInTop_7_27[7] , \wRegInTop_7_27[6] , \wRegInTop_7_27[5] , 
        \wRegInTop_7_27[4] , \wRegInTop_7_27[3] , \wRegInTop_7_27[2] , 
        \wRegInTop_7_27[1] , \wRegInTop_7_27[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_49 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink177[31] , \ScanLink177[30] , \ScanLink177[29] , 
        \ScanLink177[28] , \ScanLink177[27] , \ScanLink177[26] , 
        \ScanLink177[25] , \ScanLink177[24] , \ScanLink177[23] , 
        \ScanLink177[22] , \ScanLink177[21] , \ScanLink177[20] , 
        \ScanLink177[19] , \ScanLink177[18] , \ScanLink177[17] , 
        \ScanLink177[16] , \ScanLink177[15] , \ScanLink177[14] , 
        \ScanLink177[13] , \ScanLink177[12] , \ScanLink177[11] , 
        \ScanLink177[10] , \ScanLink177[9] , \ScanLink177[8] , 
        \ScanLink177[7] , \ScanLink177[6] , \ScanLink177[5] , \ScanLink177[4] , 
        \ScanLink177[3] , \ScanLink177[2] , \ScanLink177[1] , \ScanLink177[0] 
        }), .ScanOut({\ScanLink176[31] , \ScanLink176[30] , \ScanLink176[29] , 
        \ScanLink176[28] , \ScanLink176[27] , \ScanLink176[26] , 
        \ScanLink176[25] , \ScanLink176[24] , \ScanLink176[23] , 
        \ScanLink176[22] , \ScanLink176[21] , \ScanLink176[20] , 
        \ScanLink176[19] , \ScanLink176[18] , \ScanLink176[17] , 
        \ScanLink176[16] , \ScanLink176[15] , \ScanLink176[14] , 
        \ScanLink176[13] , \ScanLink176[12] , \ScanLink176[11] , 
        \ScanLink176[10] , \ScanLink176[9] , \ScanLink176[8] , 
        \ScanLink176[7] , \ScanLink176[6] , \ScanLink176[5] , \ScanLink176[4] , 
        \ScanLink176[3] , \ScanLink176[2] , \ScanLink176[1] , \ScanLink176[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_49[31] , 
        \wRegOut_7_49[30] , \wRegOut_7_49[29] , \wRegOut_7_49[28] , 
        \wRegOut_7_49[27] , \wRegOut_7_49[26] , \wRegOut_7_49[25] , 
        \wRegOut_7_49[24] , \wRegOut_7_49[23] , \wRegOut_7_49[22] , 
        \wRegOut_7_49[21] , \wRegOut_7_49[20] , \wRegOut_7_49[19] , 
        \wRegOut_7_49[18] , \wRegOut_7_49[17] , \wRegOut_7_49[16] , 
        \wRegOut_7_49[15] , \wRegOut_7_49[14] , \wRegOut_7_49[13] , 
        \wRegOut_7_49[12] , \wRegOut_7_49[11] , \wRegOut_7_49[10] , 
        \wRegOut_7_49[9] , \wRegOut_7_49[8] , \wRegOut_7_49[7] , 
        \wRegOut_7_49[6] , \wRegOut_7_49[5] , \wRegOut_7_49[4] , 
        \wRegOut_7_49[3] , \wRegOut_7_49[2] , \wRegOut_7_49[1] , 
        \wRegOut_7_49[0] }), .Enable1(\wRegEnTop_7_49[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_49[31] , \wRegInTop_7_49[30] , \wRegInTop_7_49[29] , 
        \wRegInTop_7_49[28] , \wRegInTop_7_49[27] , \wRegInTop_7_49[26] , 
        \wRegInTop_7_49[25] , \wRegInTop_7_49[24] , \wRegInTop_7_49[23] , 
        \wRegInTop_7_49[22] , \wRegInTop_7_49[21] , \wRegInTop_7_49[20] , 
        \wRegInTop_7_49[19] , \wRegInTop_7_49[18] , \wRegInTop_7_49[17] , 
        \wRegInTop_7_49[16] , \wRegInTop_7_49[15] , \wRegInTop_7_49[14] , 
        \wRegInTop_7_49[13] , \wRegInTop_7_49[12] , \wRegInTop_7_49[11] , 
        \wRegInTop_7_49[10] , \wRegInTop_7_49[9] , \wRegInTop_7_49[8] , 
        \wRegInTop_7_49[7] , \wRegInTop_7_49[6] , \wRegInTop_7_49[5] , 
        \wRegInTop_7_49[4] , \wRegInTop_7_49[3] , \wRegInTop_7_49[2] , 
        \wRegInTop_7_49[1] , \wRegInTop_7_49[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_114 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink242[31] , \ScanLink242[30] , \ScanLink242[29] , 
        \ScanLink242[28] , \ScanLink242[27] , \ScanLink242[26] , 
        \ScanLink242[25] , \ScanLink242[24] , \ScanLink242[23] , 
        \ScanLink242[22] , \ScanLink242[21] , \ScanLink242[20] , 
        \ScanLink242[19] , \ScanLink242[18] , \ScanLink242[17] , 
        \ScanLink242[16] , \ScanLink242[15] , \ScanLink242[14] , 
        \ScanLink242[13] , \ScanLink242[12] , \ScanLink242[11] , 
        \ScanLink242[10] , \ScanLink242[9] , \ScanLink242[8] , 
        \ScanLink242[7] , \ScanLink242[6] , \ScanLink242[5] , \ScanLink242[4] , 
        \ScanLink242[3] , \ScanLink242[2] , \ScanLink242[1] , \ScanLink242[0] 
        }), .ScanOut({\ScanLink241[31] , \ScanLink241[30] , \ScanLink241[29] , 
        \ScanLink241[28] , \ScanLink241[27] , \ScanLink241[26] , 
        \ScanLink241[25] , \ScanLink241[24] , \ScanLink241[23] , 
        \ScanLink241[22] , \ScanLink241[21] , \ScanLink241[20] , 
        \ScanLink241[19] , \ScanLink241[18] , \ScanLink241[17] , 
        \ScanLink241[16] , \ScanLink241[15] , \ScanLink241[14] , 
        \ScanLink241[13] , \ScanLink241[12] , \ScanLink241[11] , 
        \ScanLink241[10] , \ScanLink241[9] , \ScanLink241[8] , 
        \ScanLink241[7] , \ScanLink241[6] , \ScanLink241[5] , \ScanLink241[4] , 
        \ScanLink241[3] , \ScanLink241[2] , \ScanLink241[1] , \ScanLink241[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_114[31] , 
        \wRegOut_7_114[30] , \wRegOut_7_114[29] , \wRegOut_7_114[28] , 
        \wRegOut_7_114[27] , \wRegOut_7_114[26] , \wRegOut_7_114[25] , 
        \wRegOut_7_114[24] , \wRegOut_7_114[23] , \wRegOut_7_114[22] , 
        \wRegOut_7_114[21] , \wRegOut_7_114[20] , \wRegOut_7_114[19] , 
        \wRegOut_7_114[18] , \wRegOut_7_114[17] , \wRegOut_7_114[16] , 
        \wRegOut_7_114[15] , \wRegOut_7_114[14] , \wRegOut_7_114[13] , 
        \wRegOut_7_114[12] , \wRegOut_7_114[11] , \wRegOut_7_114[10] , 
        \wRegOut_7_114[9] , \wRegOut_7_114[8] , \wRegOut_7_114[7] , 
        \wRegOut_7_114[6] , \wRegOut_7_114[5] , \wRegOut_7_114[4] , 
        \wRegOut_7_114[3] , \wRegOut_7_114[2] , \wRegOut_7_114[1] , 
        \wRegOut_7_114[0] }), .Enable1(\wRegEnTop_7_114[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_114[31] , \wRegInTop_7_114[30] , 
        \wRegInTop_7_114[29] , \wRegInTop_7_114[28] , \wRegInTop_7_114[27] , 
        \wRegInTop_7_114[26] , \wRegInTop_7_114[25] , \wRegInTop_7_114[24] , 
        \wRegInTop_7_114[23] , \wRegInTop_7_114[22] , \wRegInTop_7_114[21] , 
        \wRegInTop_7_114[20] , \wRegInTop_7_114[19] , \wRegInTop_7_114[18] , 
        \wRegInTop_7_114[17] , \wRegInTop_7_114[16] , \wRegInTop_7_114[15] , 
        \wRegInTop_7_114[14] , \wRegInTop_7_114[13] , \wRegInTop_7_114[12] , 
        \wRegInTop_7_114[11] , \wRegInTop_7_114[10] , \wRegInTop_7_114[9] , 
        \wRegInTop_7_114[8] , \wRegInTop_7_114[7] , \wRegInTop_7_114[6] , 
        \wRegInTop_7_114[5] , \wRegInTop_7_114[4] , \wRegInTop_7_114[3] , 
        \wRegInTop_7_114[2] , \wRegInTop_7_114[1] , \wRegInTop_7_114[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_25[0] ), .P_In({\wRegOut_5_25[31] , 
        \wRegOut_5_25[30] , \wRegOut_5_25[29] , \wRegOut_5_25[28] , 
        \wRegOut_5_25[27] , \wRegOut_5_25[26] , \wRegOut_5_25[25] , 
        \wRegOut_5_25[24] , \wRegOut_5_25[23] , \wRegOut_5_25[22] , 
        \wRegOut_5_25[21] , \wRegOut_5_25[20] , \wRegOut_5_25[19] , 
        \wRegOut_5_25[18] , \wRegOut_5_25[17] , \wRegOut_5_25[16] , 
        \wRegOut_5_25[15] , \wRegOut_5_25[14] , \wRegOut_5_25[13] , 
        \wRegOut_5_25[12] , \wRegOut_5_25[11] , \wRegOut_5_25[10] , 
        \wRegOut_5_25[9] , \wRegOut_5_25[8] , \wRegOut_5_25[7] , 
        \wRegOut_5_25[6] , \wRegOut_5_25[5] , \wRegOut_5_25[4] , 
        \wRegOut_5_25[3] , \wRegOut_5_25[2] , \wRegOut_5_25[1] , 
        \wRegOut_5_25[0] }), .P_Out({\wRegInBot_5_25[31] , 
        \wRegInBot_5_25[30] , \wRegInBot_5_25[29] , \wRegInBot_5_25[28] , 
        \wRegInBot_5_25[27] , \wRegInBot_5_25[26] , \wRegInBot_5_25[25] , 
        \wRegInBot_5_25[24] , \wRegInBot_5_25[23] , \wRegInBot_5_25[22] , 
        \wRegInBot_5_25[21] , \wRegInBot_5_25[20] , \wRegInBot_5_25[19] , 
        \wRegInBot_5_25[18] , \wRegInBot_5_25[17] , \wRegInBot_5_25[16] , 
        \wRegInBot_5_25[15] , \wRegInBot_5_25[14] , \wRegInBot_5_25[13] , 
        \wRegInBot_5_25[12] , \wRegInBot_5_25[11] , \wRegInBot_5_25[10] , 
        \wRegInBot_5_25[9] , \wRegInBot_5_25[8] , \wRegInBot_5_25[7] , 
        \wRegInBot_5_25[6] , \wRegInBot_5_25[5] , \wRegInBot_5_25[4] , 
        \wRegInBot_5_25[3] , \wRegInBot_5_25[2] , \wRegInBot_5_25[1] , 
        \wRegInBot_5_25[0] }), .L_WR(\wRegEnTop_6_50[0] ), .L_In({
        \wRegOut_6_50[31] , \wRegOut_6_50[30] , \wRegOut_6_50[29] , 
        \wRegOut_6_50[28] , \wRegOut_6_50[27] , \wRegOut_6_50[26] , 
        \wRegOut_6_50[25] , \wRegOut_6_50[24] , \wRegOut_6_50[23] , 
        \wRegOut_6_50[22] , \wRegOut_6_50[21] , \wRegOut_6_50[20] , 
        \wRegOut_6_50[19] , \wRegOut_6_50[18] , \wRegOut_6_50[17] , 
        \wRegOut_6_50[16] , \wRegOut_6_50[15] , \wRegOut_6_50[14] , 
        \wRegOut_6_50[13] , \wRegOut_6_50[12] , \wRegOut_6_50[11] , 
        \wRegOut_6_50[10] , \wRegOut_6_50[9] , \wRegOut_6_50[8] , 
        \wRegOut_6_50[7] , \wRegOut_6_50[6] , \wRegOut_6_50[5] , 
        \wRegOut_6_50[4] , \wRegOut_6_50[3] , \wRegOut_6_50[2] , 
        \wRegOut_6_50[1] , \wRegOut_6_50[0] }), .L_Out({\wRegInTop_6_50[31] , 
        \wRegInTop_6_50[30] , \wRegInTop_6_50[29] , \wRegInTop_6_50[28] , 
        \wRegInTop_6_50[27] , \wRegInTop_6_50[26] , \wRegInTop_6_50[25] , 
        \wRegInTop_6_50[24] , \wRegInTop_6_50[23] , \wRegInTop_6_50[22] , 
        \wRegInTop_6_50[21] , \wRegInTop_6_50[20] , \wRegInTop_6_50[19] , 
        \wRegInTop_6_50[18] , \wRegInTop_6_50[17] , \wRegInTop_6_50[16] , 
        \wRegInTop_6_50[15] , \wRegInTop_6_50[14] , \wRegInTop_6_50[13] , 
        \wRegInTop_6_50[12] , \wRegInTop_6_50[11] , \wRegInTop_6_50[10] , 
        \wRegInTop_6_50[9] , \wRegInTop_6_50[8] , \wRegInTop_6_50[7] , 
        \wRegInTop_6_50[6] , \wRegInTop_6_50[5] , \wRegInTop_6_50[4] , 
        \wRegInTop_6_50[3] , \wRegInTop_6_50[2] , \wRegInTop_6_50[1] , 
        \wRegInTop_6_50[0] }), .R_WR(\wRegEnTop_6_51[0] ), .R_In({
        \wRegOut_6_51[31] , \wRegOut_6_51[30] , \wRegOut_6_51[29] , 
        \wRegOut_6_51[28] , \wRegOut_6_51[27] , \wRegOut_6_51[26] , 
        \wRegOut_6_51[25] , \wRegOut_6_51[24] , \wRegOut_6_51[23] , 
        \wRegOut_6_51[22] , \wRegOut_6_51[21] , \wRegOut_6_51[20] , 
        \wRegOut_6_51[19] , \wRegOut_6_51[18] , \wRegOut_6_51[17] , 
        \wRegOut_6_51[16] , \wRegOut_6_51[15] , \wRegOut_6_51[14] , 
        \wRegOut_6_51[13] , \wRegOut_6_51[12] , \wRegOut_6_51[11] , 
        \wRegOut_6_51[10] , \wRegOut_6_51[9] , \wRegOut_6_51[8] , 
        \wRegOut_6_51[7] , \wRegOut_6_51[6] , \wRegOut_6_51[5] , 
        \wRegOut_6_51[4] , \wRegOut_6_51[3] , \wRegOut_6_51[2] , 
        \wRegOut_6_51[1] , \wRegOut_6_51[0] }), .R_Out({\wRegInTop_6_51[31] , 
        \wRegInTop_6_51[30] , \wRegInTop_6_51[29] , \wRegInTop_6_51[28] , 
        \wRegInTop_6_51[27] , \wRegInTop_6_51[26] , \wRegInTop_6_51[25] , 
        \wRegInTop_6_51[24] , \wRegInTop_6_51[23] , \wRegInTop_6_51[22] , 
        \wRegInTop_6_51[21] , \wRegInTop_6_51[20] , \wRegInTop_6_51[19] , 
        \wRegInTop_6_51[18] , \wRegInTop_6_51[17] , \wRegInTop_6_51[16] , 
        \wRegInTop_6_51[15] , \wRegInTop_6_51[14] , \wRegInTop_6_51[13] , 
        \wRegInTop_6_51[12] , \wRegInTop_6_51[11] , \wRegInTop_6_51[10] , 
        \wRegInTop_6_51[9] , \wRegInTop_6_51[8] , \wRegInTop_6_51[7] , 
        \wRegInTop_6_51[6] , \wRegInTop_6_51[5] , \wRegInTop_6_51[4] , 
        \wRegInTop_6_51[3] , \wRegInTop_6_51[2] , \wRegInTop_6_51[1] , 
        \wRegInTop_6_51[0] }) );
    BHeap_Node_WIDTH32 BHN_6_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_15[0] ), .P_In({\wRegOut_6_15[31] , 
        \wRegOut_6_15[30] , \wRegOut_6_15[29] , \wRegOut_6_15[28] , 
        \wRegOut_6_15[27] , \wRegOut_6_15[26] , \wRegOut_6_15[25] , 
        \wRegOut_6_15[24] , \wRegOut_6_15[23] , \wRegOut_6_15[22] , 
        \wRegOut_6_15[21] , \wRegOut_6_15[20] , \wRegOut_6_15[19] , 
        \wRegOut_6_15[18] , \wRegOut_6_15[17] , \wRegOut_6_15[16] , 
        \wRegOut_6_15[15] , \wRegOut_6_15[14] , \wRegOut_6_15[13] , 
        \wRegOut_6_15[12] , \wRegOut_6_15[11] , \wRegOut_6_15[10] , 
        \wRegOut_6_15[9] , \wRegOut_6_15[8] , \wRegOut_6_15[7] , 
        \wRegOut_6_15[6] , \wRegOut_6_15[5] , \wRegOut_6_15[4] , 
        \wRegOut_6_15[3] , \wRegOut_6_15[2] , \wRegOut_6_15[1] , 
        \wRegOut_6_15[0] }), .P_Out({\wRegInBot_6_15[31] , 
        \wRegInBot_6_15[30] , \wRegInBot_6_15[29] , \wRegInBot_6_15[28] , 
        \wRegInBot_6_15[27] , \wRegInBot_6_15[26] , \wRegInBot_6_15[25] , 
        \wRegInBot_6_15[24] , \wRegInBot_6_15[23] , \wRegInBot_6_15[22] , 
        \wRegInBot_6_15[21] , \wRegInBot_6_15[20] , \wRegInBot_6_15[19] , 
        \wRegInBot_6_15[18] , \wRegInBot_6_15[17] , \wRegInBot_6_15[16] , 
        \wRegInBot_6_15[15] , \wRegInBot_6_15[14] , \wRegInBot_6_15[13] , 
        \wRegInBot_6_15[12] , \wRegInBot_6_15[11] , \wRegInBot_6_15[10] , 
        \wRegInBot_6_15[9] , \wRegInBot_6_15[8] , \wRegInBot_6_15[7] , 
        \wRegInBot_6_15[6] , \wRegInBot_6_15[5] , \wRegInBot_6_15[4] , 
        \wRegInBot_6_15[3] , \wRegInBot_6_15[2] , \wRegInBot_6_15[1] , 
        \wRegInBot_6_15[0] }), .L_WR(\wRegEnTop_7_30[0] ), .L_In({
        \wRegOut_7_30[31] , \wRegOut_7_30[30] , \wRegOut_7_30[29] , 
        \wRegOut_7_30[28] , \wRegOut_7_30[27] , \wRegOut_7_30[26] , 
        \wRegOut_7_30[25] , \wRegOut_7_30[24] , \wRegOut_7_30[23] , 
        \wRegOut_7_30[22] , \wRegOut_7_30[21] , \wRegOut_7_30[20] , 
        \wRegOut_7_30[19] , \wRegOut_7_30[18] , \wRegOut_7_30[17] , 
        \wRegOut_7_30[16] , \wRegOut_7_30[15] , \wRegOut_7_30[14] , 
        \wRegOut_7_30[13] , \wRegOut_7_30[12] , \wRegOut_7_30[11] , 
        \wRegOut_7_30[10] , \wRegOut_7_30[9] , \wRegOut_7_30[8] , 
        \wRegOut_7_30[7] , \wRegOut_7_30[6] , \wRegOut_7_30[5] , 
        \wRegOut_7_30[4] , \wRegOut_7_30[3] , \wRegOut_7_30[2] , 
        \wRegOut_7_30[1] , \wRegOut_7_30[0] }), .L_Out({\wRegInTop_7_30[31] , 
        \wRegInTop_7_30[30] , \wRegInTop_7_30[29] , \wRegInTop_7_30[28] , 
        \wRegInTop_7_30[27] , \wRegInTop_7_30[26] , \wRegInTop_7_30[25] , 
        \wRegInTop_7_30[24] , \wRegInTop_7_30[23] , \wRegInTop_7_30[22] , 
        \wRegInTop_7_30[21] , \wRegInTop_7_30[20] , \wRegInTop_7_30[19] , 
        \wRegInTop_7_30[18] , \wRegInTop_7_30[17] , \wRegInTop_7_30[16] , 
        \wRegInTop_7_30[15] , \wRegInTop_7_30[14] , \wRegInTop_7_30[13] , 
        \wRegInTop_7_30[12] , \wRegInTop_7_30[11] , \wRegInTop_7_30[10] , 
        \wRegInTop_7_30[9] , \wRegInTop_7_30[8] , \wRegInTop_7_30[7] , 
        \wRegInTop_7_30[6] , \wRegInTop_7_30[5] , \wRegInTop_7_30[4] , 
        \wRegInTop_7_30[3] , \wRegInTop_7_30[2] , \wRegInTop_7_30[1] , 
        \wRegInTop_7_30[0] }), .R_WR(\wRegEnTop_7_31[0] ), .R_In({
        \wRegOut_7_31[31] , \wRegOut_7_31[30] , \wRegOut_7_31[29] , 
        \wRegOut_7_31[28] , \wRegOut_7_31[27] , \wRegOut_7_31[26] , 
        \wRegOut_7_31[25] , \wRegOut_7_31[24] , \wRegOut_7_31[23] , 
        \wRegOut_7_31[22] , \wRegOut_7_31[21] , \wRegOut_7_31[20] , 
        \wRegOut_7_31[19] , \wRegOut_7_31[18] , \wRegOut_7_31[17] , 
        \wRegOut_7_31[16] , \wRegOut_7_31[15] , \wRegOut_7_31[14] , 
        \wRegOut_7_31[13] , \wRegOut_7_31[12] , \wRegOut_7_31[11] , 
        \wRegOut_7_31[10] , \wRegOut_7_31[9] , \wRegOut_7_31[8] , 
        \wRegOut_7_31[7] , \wRegOut_7_31[6] , \wRegOut_7_31[5] , 
        \wRegOut_7_31[4] , \wRegOut_7_31[3] , \wRegOut_7_31[2] , 
        \wRegOut_7_31[1] , \wRegOut_7_31[0] }), .R_Out({\wRegInTop_7_31[31] , 
        \wRegInTop_7_31[30] , \wRegInTop_7_31[29] , \wRegInTop_7_31[28] , 
        \wRegInTop_7_31[27] , \wRegInTop_7_31[26] , \wRegInTop_7_31[25] , 
        \wRegInTop_7_31[24] , \wRegInTop_7_31[23] , \wRegInTop_7_31[22] , 
        \wRegInTop_7_31[21] , \wRegInTop_7_31[20] , \wRegInTop_7_31[19] , 
        \wRegInTop_7_31[18] , \wRegInTop_7_31[17] , \wRegInTop_7_31[16] , 
        \wRegInTop_7_31[15] , \wRegInTop_7_31[14] , \wRegInTop_7_31[13] , 
        \wRegInTop_7_31[12] , \wRegInTop_7_31[11] , \wRegInTop_7_31[10] , 
        \wRegInTop_7_31[9] , \wRegInTop_7_31[8] , \wRegInTop_7_31[7] , 
        \wRegInTop_7_31[6] , \wRegInTop_7_31[5] , \wRegInTop_7_31[4] , 
        \wRegInTop_7_31[3] , \wRegInTop_7_31[2] , \wRegInTop_7_31[1] , 
        \wRegInTop_7_31[0] }) );
    BHeap_Node_WIDTH32 BHN_6_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_32[0] ), .P_In({\wRegOut_6_32[31] , 
        \wRegOut_6_32[30] , \wRegOut_6_32[29] , \wRegOut_6_32[28] , 
        \wRegOut_6_32[27] , \wRegOut_6_32[26] , \wRegOut_6_32[25] , 
        \wRegOut_6_32[24] , \wRegOut_6_32[23] , \wRegOut_6_32[22] , 
        \wRegOut_6_32[21] , \wRegOut_6_32[20] , \wRegOut_6_32[19] , 
        \wRegOut_6_32[18] , \wRegOut_6_32[17] , \wRegOut_6_32[16] , 
        \wRegOut_6_32[15] , \wRegOut_6_32[14] , \wRegOut_6_32[13] , 
        \wRegOut_6_32[12] , \wRegOut_6_32[11] , \wRegOut_6_32[10] , 
        \wRegOut_6_32[9] , \wRegOut_6_32[8] , \wRegOut_6_32[7] , 
        \wRegOut_6_32[6] , \wRegOut_6_32[5] , \wRegOut_6_32[4] , 
        \wRegOut_6_32[3] , \wRegOut_6_32[2] , \wRegOut_6_32[1] , 
        \wRegOut_6_32[0] }), .P_Out({\wRegInBot_6_32[31] , 
        \wRegInBot_6_32[30] , \wRegInBot_6_32[29] , \wRegInBot_6_32[28] , 
        \wRegInBot_6_32[27] , \wRegInBot_6_32[26] , \wRegInBot_6_32[25] , 
        \wRegInBot_6_32[24] , \wRegInBot_6_32[23] , \wRegInBot_6_32[22] , 
        \wRegInBot_6_32[21] , \wRegInBot_6_32[20] , \wRegInBot_6_32[19] , 
        \wRegInBot_6_32[18] , \wRegInBot_6_32[17] , \wRegInBot_6_32[16] , 
        \wRegInBot_6_32[15] , \wRegInBot_6_32[14] , \wRegInBot_6_32[13] , 
        \wRegInBot_6_32[12] , \wRegInBot_6_32[11] , \wRegInBot_6_32[10] , 
        \wRegInBot_6_32[9] , \wRegInBot_6_32[8] , \wRegInBot_6_32[7] , 
        \wRegInBot_6_32[6] , \wRegInBot_6_32[5] , \wRegInBot_6_32[4] , 
        \wRegInBot_6_32[3] , \wRegInBot_6_32[2] , \wRegInBot_6_32[1] , 
        \wRegInBot_6_32[0] }), .L_WR(\wRegEnTop_7_64[0] ), .L_In({
        \wRegOut_7_64[31] , \wRegOut_7_64[30] , \wRegOut_7_64[29] , 
        \wRegOut_7_64[28] , \wRegOut_7_64[27] , \wRegOut_7_64[26] , 
        \wRegOut_7_64[25] , \wRegOut_7_64[24] , \wRegOut_7_64[23] , 
        \wRegOut_7_64[22] , \wRegOut_7_64[21] , \wRegOut_7_64[20] , 
        \wRegOut_7_64[19] , \wRegOut_7_64[18] , \wRegOut_7_64[17] , 
        \wRegOut_7_64[16] , \wRegOut_7_64[15] , \wRegOut_7_64[14] , 
        \wRegOut_7_64[13] , \wRegOut_7_64[12] , \wRegOut_7_64[11] , 
        \wRegOut_7_64[10] , \wRegOut_7_64[9] , \wRegOut_7_64[8] , 
        \wRegOut_7_64[7] , \wRegOut_7_64[6] , \wRegOut_7_64[5] , 
        \wRegOut_7_64[4] , \wRegOut_7_64[3] , \wRegOut_7_64[2] , 
        \wRegOut_7_64[1] , \wRegOut_7_64[0] }), .L_Out({\wRegInTop_7_64[31] , 
        \wRegInTop_7_64[30] , \wRegInTop_7_64[29] , \wRegInTop_7_64[28] , 
        \wRegInTop_7_64[27] , \wRegInTop_7_64[26] , \wRegInTop_7_64[25] , 
        \wRegInTop_7_64[24] , \wRegInTop_7_64[23] , \wRegInTop_7_64[22] , 
        \wRegInTop_7_64[21] , \wRegInTop_7_64[20] , \wRegInTop_7_64[19] , 
        \wRegInTop_7_64[18] , \wRegInTop_7_64[17] , \wRegInTop_7_64[16] , 
        \wRegInTop_7_64[15] , \wRegInTop_7_64[14] , \wRegInTop_7_64[13] , 
        \wRegInTop_7_64[12] , \wRegInTop_7_64[11] , \wRegInTop_7_64[10] , 
        \wRegInTop_7_64[9] , \wRegInTop_7_64[8] , \wRegInTop_7_64[7] , 
        \wRegInTop_7_64[6] , \wRegInTop_7_64[5] , \wRegInTop_7_64[4] , 
        \wRegInTop_7_64[3] , \wRegInTop_7_64[2] , \wRegInTop_7_64[1] , 
        \wRegInTop_7_64[0] }), .R_WR(\wRegEnTop_7_65[0] ), .R_In({
        \wRegOut_7_65[31] , \wRegOut_7_65[30] , \wRegOut_7_65[29] , 
        \wRegOut_7_65[28] , \wRegOut_7_65[27] , \wRegOut_7_65[26] , 
        \wRegOut_7_65[25] , \wRegOut_7_65[24] , \wRegOut_7_65[23] , 
        \wRegOut_7_65[22] , \wRegOut_7_65[21] , \wRegOut_7_65[20] , 
        \wRegOut_7_65[19] , \wRegOut_7_65[18] , \wRegOut_7_65[17] , 
        \wRegOut_7_65[16] , \wRegOut_7_65[15] , \wRegOut_7_65[14] , 
        \wRegOut_7_65[13] , \wRegOut_7_65[12] , \wRegOut_7_65[11] , 
        \wRegOut_7_65[10] , \wRegOut_7_65[9] , \wRegOut_7_65[8] , 
        \wRegOut_7_65[7] , \wRegOut_7_65[6] , \wRegOut_7_65[5] , 
        \wRegOut_7_65[4] , \wRegOut_7_65[3] , \wRegOut_7_65[2] , 
        \wRegOut_7_65[1] , \wRegOut_7_65[0] }), .R_Out({\wRegInTop_7_65[31] , 
        \wRegInTop_7_65[30] , \wRegInTop_7_65[29] , \wRegInTop_7_65[28] , 
        \wRegInTop_7_65[27] , \wRegInTop_7_65[26] , \wRegInTop_7_65[25] , 
        \wRegInTop_7_65[24] , \wRegInTop_7_65[23] , \wRegInTop_7_65[22] , 
        \wRegInTop_7_65[21] , \wRegInTop_7_65[20] , \wRegInTop_7_65[19] , 
        \wRegInTop_7_65[18] , \wRegInTop_7_65[17] , \wRegInTop_7_65[16] , 
        \wRegInTop_7_65[15] , \wRegInTop_7_65[14] , \wRegInTop_7_65[13] , 
        \wRegInTop_7_65[12] , \wRegInTop_7_65[11] , \wRegInTop_7_65[10] , 
        \wRegInTop_7_65[9] , \wRegInTop_7_65[8] , \wRegInTop_7_65[7] , 
        \wRegInTop_7_65[6] , \wRegInTop_7_65[5] , \wRegInTop_7_65[4] , 
        \wRegInTop_7_65[3] , \wRegInTop_7_65[2] , \wRegInTop_7_65[1] , 
        \wRegInTop_7_65[0] }) );
    BHeap_Node_WIDTH32 BHN_4_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_1[0] ), .P_In({\wRegOut_4_1[31] , 
        \wRegOut_4_1[30] , \wRegOut_4_1[29] , \wRegOut_4_1[28] , 
        \wRegOut_4_1[27] , \wRegOut_4_1[26] , \wRegOut_4_1[25] , 
        \wRegOut_4_1[24] , \wRegOut_4_1[23] , \wRegOut_4_1[22] , 
        \wRegOut_4_1[21] , \wRegOut_4_1[20] , \wRegOut_4_1[19] , 
        \wRegOut_4_1[18] , \wRegOut_4_1[17] , \wRegOut_4_1[16] , 
        \wRegOut_4_1[15] , \wRegOut_4_1[14] , \wRegOut_4_1[13] , 
        \wRegOut_4_1[12] , \wRegOut_4_1[11] , \wRegOut_4_1[10] , 
        \wRegOut_4_1[9] , \wRegOut_4_1[8] , \wRegOut_4_1[7] , \wRegOut_4_1[6] , 
        \wRegOut_4_1[5] , \wRegOut_4_1[4] , \wRegOut_4_1[3] , \wRegOut_4_1[2] , 
        \wRegOut_4_1[1] , \wRegOut_4_1[0] }), .P_Out({\wRegInBot_4_1[31] , 
        \wRegInBot_4_1[30] , \wRegInBot_4_1[29] , \wRegInBot_4_1[28] , 
        \wRegInBot_4_1[27] , \wRegInBot_4_1[26] , \wRegInBot_4_1[25] , 
        \wRegInBot_4_1[24] , \wRegInBot_4_1[23] , \wRegInBot_4_1[22] , 
        \wRegInBot_4_1[21] , \wRegInBot_4_1[20] , \wRegInBot_4_1[19] , 
        \wRegInBot_4_1[18] , \wRegInBot_4_1[17] , \wRegInBot_4_1[16] , 
        \wRegInBot_4_1[15] , \wRegInBot_4_1[14] , \wRegInBot_4_1[13] , 
        \wRegInBot_4_1[12] , \wRegInBot_4_1[11] , \wRegInBot_4_1[10] , 
        \wRegInBot_4_1[9] , \wRegInBot_4_1[8] , \wRegInBot_4_1[7] , 
        \wRegInBot_4_1[6] , \wRegInBot_4_1[5] , \wRegInBot_4_1[4] , 
        \wRegInBot_4_1[3] , \wRegInBot_4_1[2] , \wRegInBot_4_1[1] , 
        \wRegInBot_4_1[0] }), .L_WR(\wRegEnTop_5_2[0] ), .L_In({
        \wRegOut_5_2[31] , \wRegOut_5_2[30] , \wRegOut_5_2[29] , 
        \wRegOut_5_2[28] , \wRegOut_5_2[27] , \wRegOut_5_2[26] , 
        \wRegOut_5_2[25] , \wRegOut_5_2[24] , \wRegOut_5_2[23] , 
        \wRegOut_5_2[22] , \wRegOut_5_2[21] , \wRegOut_5_2[20] , 
        \wRegOut_5_2[19] , \wRegOut_5_2[18] , \wRegOut_5_2[17] , 
        \wRegOut_5_2[16] , \wRegOut_5_2[15] , \wRegOut_5_2[14] , 
        \wRegOut_5_2[13] , \wRegOut_5_2[12] , \wRegOut_5_2[11] , 
        \wRegOut_5_2[10] , \wRegOut_5_2[9] , \wRegOut_5_2[8] , 
        \wRegOut_5_2[7] , \wRegOut_5_2[6] , \wRegOut_5_2[5] , \wRegOut_5_2[4] , 
        \wRegOut_5_2[3] , \wRegOut_5_2[2] , \wRegOut_5_2[1] , \wRegOut_5_2[0] 
        }), .L_Out({\wRegInTop_5_2[31] , \wRegInTop_5_2[30] , 
        \wRegInTop_5_2[29] , \wRegInTop_5_2[28] , \wRegInTop_5_2[27] , 
        \wRegInTop_5_2[26] , \wRegInTop_5_2[25] , \wRegInTop_5_2[24] , 
        \wRegInTop_5_2[23] , \wRegInTop_5_2[22] , \wRegInTop_5_2[21] , 
        \wRegInTop_5_2[20] , \wRegInTop_5_2[19] , \wRegInTop_5_2[18] , 
        \wRegInTop_5_2[17] , \wRegInTop_5_2[16] , \wRegInTop_5_2[15] , 
        \wRegInTop_5_2[14] , \wRegInTop_5_2[13] , \wRegInTop_5_2[12] , 
        \wRegInTop_5_2[11] , \wRegInTop_5_2[10] , \wRegInTop_5_2[9] , 
        \wRegInTop_5_2[8] , \wRegInTop_5_2[7] , \wRegInTop_5_2[6] , 
        \wRegInTop_5_2[5] , \wRegInTop_5_2[4] , \wRegInTop_5_2[3] , 
        \wRegInTop_5_2[2] , \wRegInTop_5_2[1] , \wRegInTop_5_2[0] }), .R_WR(
        \wRegEnTop_5_3[0] ), .R_In({\wRegOut_5_3[31] , \wRegOut_5_3[30] , 
        \wRegOut_5_3[29] , \wRegOut_5_3[28] , \wRegOut_5_3[27] , 
        \wRegOut_5_3[26] , \wRegOut_5_3[25] , \wRegOut_5_3[24] , 
        \wRegOut_5_3[23] , \wRegOut_5_3[22] , \wRegOut_5_3[21] , 
        \wRegOut_5_3[20] , \wRegOut_5_3[19] , \wRegOut_5_3[18] , 
        \wRegOut_5_3[17] , \wRegOut_5_3[16] , \wRegOut_5_3[15] , 
        \wRegOut_5_3[14] , \wRegOut_5_3[13] , \wRegOut_5_3[12] , 
        \wRegOut_5_3[11] , \wRegOut_5_3[10] , \wRegOut_5_3[9] , 
        \wRegOut_5_3[8] , \wRegOut_5_3[7] , \wRegOut_5_3[6] , \wRegOut_5_3[5] , 
        \wRegOut_5_3[4] , \wRegOut_5_3[3] , \wRegOut_5_3[2] , \wRegOut_5_3[1] , 
        \wRegOut_5_3[0] }), .R_Out({\wRegInTop_5_3[31] , \wRegInTop_5_3[30] , 
        \wRegInTop_5_3[29] , \wRegInTop_5_3[28] , \wRegInTop_5_3[27] , 
        \wRegInTop_5_3[26] , \wRegInTop_5_3[25] , \wRegInTop_5_3[24] , 
        \wRegInTop_5_3[23] , \wRegInTop_5_3[22] , \wRegInTop_5_3[21] , 
        \wRegInTop_5_3[20] , \wRegInTop_5_3[19] , \wRegInTop_5_3[18] , 
        \wRegInTop_5_3[17] , \wRegInTop_5_3[16] , \wRegInTop_5_3[15] , 
        \wRegInTop_5_3[14] , \wRegInTop_5_3[13] , \wRegInTop_5_3[12] , 
        \wRegInTop_5_3[11] , \wRegInTop_5_3[10] , \wRegInTop_5_3[9] , 
        \wRegInTop_5_3[8] , \wRegInTop_5_3[7] , \wRegInTop_5_3[6] , 
        \wRegInTop_5_3[5] , \wRegInTop_5_3[4] , \wRegInTop_5_3[3] , 
        \wRegInTop_5_3[2] , \wRegInTop_5_3[1] , \wRegInTop_5_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_90 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink218[31] , \ScanLink218[30] , \ScanLink218[29] , 
        \ScanLink218[28] , \ScanLink218[27] , \ScanLink218[26] , 
        \ScanLink218[25] , \ScanLink218[24] , \ScanLink218[23] , 
        \ScanLink218[22] , \ScanLink218[21] , \ScanLink218[20] , 
        \ScanLink218[19] , \ScanLink218[18] , \ScanLink218[17] , 
        \ScanLink218[16] , \ScanLink218[15] , \ScanLink218[14] , 
        \ScanLink218[13] , \ScanLink218[12] , \ScanLink218[11] , 
        \ScanLink218[10] , \ScanLink218[9] , \ScanLink218[8] , 
        \ScanLink218[7] , \ScanLink218[6] , \ScanLink218[5] , \ScanLink218[4] , 
        \ScanLink218[3] , \ScanLink218[2] , \ScanLink218[1] , \ScanLink218[0] 
        }), .ScanOut({\ScanLink217[31] , \ScanLink217[30] , \ScanLink217[29] , 
        \ScanLink217[28] , \ScanLink217[27] , \ScanLink217[26] , 
        \ScanLink217[25] , \ScanLink217[24] , \ScanLink217[23] , 
        \ScanLink217[22] , \ScanLink217[21] , \ScanLink217[20] , 
        \ScanLink217[19] , \ScanLink217[18] , \ScanLink217[17] , 
        \ScanLink217[16] , \ScanLink217[15] , \ScanLink217[14] , 
        \ScanLink217[13] , \ScanLink217[12] , \ScanLink217[11] , 
        \ScanLink217[10] , \ScanLink217[9] , \ScanLink217[8] , 
        \ScanLink217[7] , \ScanLink217[6] , \ScanLink217[5] , \ScanLink217[4] , 
        \ScanLink217[3] , \ScanLink217[2] , \ScanLink217[1] , \ScanLink217[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_90[31] , 
        \wRegOut_7_90[30] , \wRegOut_7_90[29] , \wRegOut_7_90[28] , 
        \wRegOut_7_90[27] , \wRegOut_7_90[26] , \wRegOut_7_90[25] , 
        \wRegOut_7_90[24] , \wRegOut_7_90[23] , \wRegOut_7_90[22] , 
        \wRegOut_7_90[21] , \wRegOut_7_90[20] , \wRegOut_7_90[19] , 
        \wRegOut_7_90[18] , \wRegOut_7_90[17] , \wRegOut_7_90[16] , 
        \wRegOut_7_90[15] , \wRegOut_7_90[14] , \wRegOut_7_90[13] , 
        \wRegOut_7_90[12] , \wRegOut_7_90[11] , \wRegOut_7_90[10] , 
        \wRegOut_7_90[9] , \wRegOut_7_90[8] , \wRegOut_7_90[7] , 
        \wRegOut_7_90[6] , \wRegOut_7_90[5] , \wRegOut_7_90[4] , 
        \wRegOut_7_90[3] , \wRegOut_7_90[2] , \wRegOut_7_90[1] , 
        \wRegOut_7_90[0] }), .Enable1(\wRegEnTop_7_90[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_90[31] , \wRegInTop_7_90[30] , \wRegInTop_7_90[29] , 
        \wRegInTop_7_90[28] , \wRegInTop_7_90[27] , \wRegInTop_7_90[26] , 
        \wRegInTop_7_90[25] , \wRegInTop_7_90[24] , \wRegInTop_7_90[23] , 
        \wRegInTop_7_90[22] , \wRegInTop_7_90[21] , \wRegInTop_7_90[20] , 
        \wRegInTop_7_90[19] , \wRegInTop_7_90[18] , \wRegInTop_7_90[17] , 
        \wRegInTop_7_90[16] , \wRegInTop_7_90[15] , \wRegInTop_7_90[14] , 
        \wRegInTop_7_90[13] , \wRegInTop_7_90[12] , \wRegInTop_7_90[11] , 
        \wRegInTop_7_90[10] , \wRegInTop_7_90[9] , \wRegInTop_7_90[8] , 
        \wRegInTop_7_90[7] , \wRegInTop_7_90[6] , \wRegInTop_7_90[5] , 
        \wRegInTop_7_90[4] , \wRegInTop_7_90[3] , \wRegInTop_7_90[2] , 
        \wRegInTop_7_90[1] , \wRegInTop_7_90[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_1[0] ), .P_In({\wRegOut_5_1[31] , 
        \wRegOut_5_1[30] , \wRegOut_5_1[29] , \wRegOut_5_1[28] , 
        \wRegOut_5_1[27] , \wRegOut_5_1[26] , \wRegOut_5_1[25] , 
        \wRegOut_5_1[24] , \wRegOut_5_1[23] , \wRegOut_5_1[22] , 
        \wRegOut_5_1[21] , \wRegOut_5_1[20] , \wRegOut_5_1[19] , 
        \wRegOut_5_1[18] , \wRegOut_5_1[17] , \wRegOut_5_1[16] , 
        \wRegOut_5_1[15] , \wRegOut_5_1[14] , \wRegOut_5_1[13] , 
        \wRegOut_5_1[12] , \wRegOut_5_1[11] , \wRegOut_5_1[10] , 
        \wRegOut_5_1[9] , \wRegOut_5_1[8] , \wRegOut_5_1[7] , \wRegOut_5_1[6] , 
        \wRegOut_5_1[5] , \wRegOut_5_1[4] , \wRegOut_5_1[3] , \wRegOut_5_1[2] , 
        \wRegOut_5_1[1] , \wRegOut_5_1[0] }), .P_Out({\wRegInBot_5_1[31] , 
        \wRegInBot_5_1[30] , \wRegInBot_5_1[29] , \wRegInBot_5_1[28] , 
        \wRegInBot_5_1[27] , \wRegInBot_5_1[26] , \wRegInBot_5_1[25] , 
        \wRegInBot_5_1[24] , \wRegInBot_5_1[23] , \wRegInBot_5_1[22] , 
        \wRegInBot_5_1[21] , \wRegInBot_5_1[20] , \wRegInBot_5_1[19] , 
        \wRegInBot_5_1[18] , \wRegInBot_5_1[17] , \wRegInBot_5_1[16] , 
        \wRegInBot_5_1[15] , \wRegInBot_5_1[14] , \wRegInBot_5_1[13] , 
        \wRegInBot_5_1[12] , \wRegInBot_5_1[11] , \wRegInBot_5_1[10] , 
        \wRegInBot_5_1[9] , \wRegInBot_5_1[8] , \wRegInBot_5_1[7] , 
        \wRegInBot_5_1[6] , \wRegInBot_5_1[5] , \wRegInBot_5_1[4] , 
        \wRegInBot_5_1[3] , \wRegInBot_5_1[2] , \wRegInBot_5_1[1] , 
        \wRegInBot_5_1[0] }), .L_WR(\wRegEnTop_6_2[0] ), .L_In({
        \wRegOut_6_2[31] , \wRegOut_6_2[30] , \wRegOut_6_2[29] , 
        \wRegOut_6_2[28] , \wRegOut_6_2[27] , \wRegOut_6_2[26] , 
        \wRegOut_6_2[25] , \wRegOut_6_2[24] , \wRegOut_6_2[23] , 
        \wRegOut_6_2[22] , \wRegOut_6_2[21] , \wRegOut_6_2[20] , 
        \wRegOut_6_2[19] , \wRegOut_6_2[18] , \wRegOut_6_2[17] , 
        \wRegOut_6_2[16] , \wRegOut_6_2[15] , \wRegOut_6_2[14] , 
        \wRegOut_6_2[13] , \wRegOut_6_2[12] , \wRegOut_6_2[11] , 
        \wRegOut_6_2[10] , \wRegOut_6_2[9] , \wRegOut_6_2[8] , 
        \wRegOut_6_2[7] , \wRegOut_6_2[6] , \wRegOut_6_2[5] , \wRegOut_6_2[4] , 
        \wRegOut_6_2[3] , \wRegOut_6_2[2] , \wRegOut_6_2[1] , \wRegOut_6_2[0] 
        }), .L_Out({\wRegInTop_6_2[31] , \wRegInTop_6_2[30] , 
        \wRegInTop_6_2[29] , \wRegInTop_6_2[28] , \wRegInTop_6_2[27] , 
        \wRegInTop_6_2[26] , \wRegInTop_6_2[25] , \wRegInTop_6_2[24] , 
        \wRegInTop_6_2[23] , \wRegInTop_6_2[22] , \wRegInTop_6_2[21] , 
        \wRegInTop_6_2[20] , \wRegInTop_6_2[19] , \wRegInTop_6_2[18] , 
        \wRegInTop_6_2[17] , \wRegInTop_6_2[16] , \wRegInTop_6_2[15] , 
        \wRegInTop_6_2[14] , \wRegInTop_6_2[13] , \wRegInTop_6_2[12] , 
        \wRegInTop_6_2[11] , \wRegInTop_6_2[10] , \wRegInTop_6_2[9] , 
        \wRegInTop_6_2[8] , \wRegInTop_6_2[7] , \wRegInTop_6_2[6] , 
        \wRegInTop_6_2[5] , \wRegInTop_6_2[4] , \wRegInTop_6_2[3] , 
        \wRegInTop_6_2[2] , \wRegInTop_6_2[1] , \wRegInTop_6_2[0] }), .R_WR(
        \wRegEnTop_6_3[0] ), .R_In({\wRegOut_6_3[31] , \wRegOut_6_3[30] , 
        \wRegOut_6_3[29] , \wRegOut_6_3[28] , \wRegOut_6_3[27] , 
        \wRegOut_6_3[26] , \wRegOut_6_3[25] , \wRegOut_6_3[24] , 
        \wRegOut_6_3[23] , \wRegOut_6_3[22] , \wRegOut_6_3[21] , 
        \wRegOut_6_3[20] , \wRegOut_6_3[19] , \wRegOut_6_3[18] , 
        \wRegOut_6_3[17] , \wRegOut_6_3[16] , \wRegOut_6_3[15] , 
        \wRegOut_6_3[14] , \wRegOut_6_3[13] , \wRegOut_6_3[12] , 
        \wRegOut_6_3[11] , \wRegOut_6_3[10] , \wRegOut_6_3[9] , 
        \wRegOut_6_3[8] , \wRegOut_6_3[7] , \wRegOut_6_3[6] , \wRegOut_6_3[5] , 
        \wRegOut_6_3[4] , \wRegOut_6_3[3] , \wRegOut_6_3[2] , \wRegOut_6_3[1] , 
        \wRegOut_6_3[0] }), .R_Out({\wRegInTop_6_3[31] , \wRegInTop_6_3[30] , 
        \wRegInTop_6_3[29] , \wRegInTop_6_3[28] , \wRegInTop_6_3[27] , 
        \wRegInTop_6_3[26] , \wRegInTop_6_3[25] , \wRegInTop_6_3[24] , 
        \wRegInTop_6_3[23] , \wRegInTop_6_3[22] , \wRegInTop_6_3[21] , 
        \wRegInTop_6_3[20] , \wRegInTop_6_3[19] , \wRegInTop_6_3[18] , 
        \wRegInTop_6_3[17] , \wRegInTop_6_3[16] , \wRegInTop_6_3[15] , 
        \wRegInTop_6_3[14] , \wRegInTop_6_3[13] , \wRegInTop_6_3[12] , 
        \wRegInTop_6_3[11] , \wRegInTop_6_3[10] , \wRegInTop_6_3[9] , 
        \wRegInTop_6_3[8] , \wRegInTop_6_3[7] , \wRegInTop_6_3[6] , 
        \wRegInTop_6_3[5] , \wRegInTop_6_3[4] , \wRegInTop_6_3[3] , 
        \wRegInTop_6_3[2] , \wRegInTop_6_3[1] , \wRegInTop_6_3[0] }) );
    BHeap_Node_WIDTH32 BHN_6_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_47[0] ), .P_In({\wRegOut_6_47[31] , 
        \wRegOut_6_47[30] , \wRegOut_6_47[29] , \wRegOut_6_47[28] , 
        \wRegOut_6_47[27] , \wRegOut_6_47[26] , \wRegOut_6_47[25] , 
        \wRegOut_6_47[24] , \wRegOut_6_47[23] , \wRegOut_6_47[22] , 
        \wRegOut_6_47[21] , \wRegOut_6_47[20] , \wRegOut_6_47[19] , 
        \wRegOut_6_47[18] , \wRegOut_6_47[17] , \wRegOut_6_47[16] , 
        \wRegOut_6_47[15] , \wRegOut_6_47[14] , \wRegOut_6_47[13] , 
        \wRegOut_6_47[12] , \wRegOut_6_47[11] , \wRegOut_6_47[10] , 
        \wRegOut_6_47[9] , \wRegOut_6_47[8] , \wRegOut_6_47[7] , 
        \wRegOut_6_47[6] , \wRegOut_6_47[5] , \wRegOut_6_47[4] , 
        \wRegOut_6_47[3] , \wRegOut_6_47[2] , \wRegOut_6_47[1] , 
        \wRegOut_6_47[0] }), .P_Out({\wRegInBot_6_47[31] , 
        \wRegInBot_6_47[30] , \wRegInBot_6_47[29] , \wRegInBot_6_47[28] , 
        \wRegInBot_6_47[27] , \wRegInBot_6_47[26] , \wRegInBot_6_47[25] , 
        \wRegInBot_6_47[24] , \wRegInBot_6_47[23] , \wRegInBot_6_47[22] , 
        \wRegInBot_6_47[21] , \wRegInBot_6_47[20] , \wRegInBot_6_47[19] , 
        \wRegInBot_6_47[18] , \wRegInBot_6_47[17] , \wRegInBot_6_47[16] , 
        \wRegInBot_6_47[15] , \wRegInBot_6_47[14] , \wRegInBot_6_47[13] , 
        \wRegInBot_6_47[12] , \wRegInBot_6_47[11] , \wRegInBot_6_47[10] , 
        \wRegInBot_6_47[9] , \wRegInBot_6_47[8] , \wRegInBot_6_47[7] , 
        \wRegInBot_6_47[6] , \wRegInBot_6_47[5] , \wRegInBot_6_47[4] , 
        \wRegInBot_6_47[3] , \wRegInBot_6_47[2] , \wRegInBot_6_47[1] , 
        \wRegInBot_6_47[0] }), .L_WR(\wRegEnTop_7_94[0] ), .L_In({
        \wRegOut_7_94[31] , \wRegOut_7_94[30] , \wRegOut_7_94[29] , 
        \wRegOut_7_94[28] , \wRegOut_7_94[27] , \wRegOut_7_94[26] , 
        \wRegOut_7_94[25] , \wRegOut_7_94[24] , \wRegOut_7_94[23] , 
        \wRegOut_7_94[22] , \wRegOut_7_94[21] , \wRegOut_7_94[20] , 
        \wRegOut_7_94[19] , \wRegOut_7_94[18] , \wRegOut_7_94[17] , 
        \wRegOut_7_94[16] , \wRegOut_7_94[15] , \wRegOut_7_94[14] , 
        \wRegOut_7_94[13] , \wRegOut_7_94[12] , \wRegOut_7_94[11] , 
        \wRegOut_7_94[10] , \wRegOut_7_94[9] , \wRegOut_7_94[8] , 
        \wRegOut_7_94[7] , \wRegOut_7_94[6] , \wRegOut_7_94[5] , 
        \wRegOut_7_94[4] , \wRegOut_7_94[3] , \wRegOut_7_94[2] , 
        \wRegOut_7_94[1] , \wRegOut_7_94[0] }), .L_Out({\wRegInTop_7_94[31] , 
        \wRegInTop_7_94[30] , \wRegInTop_7_94[29] , \wRegInTop_7_94[28] , 
        \wRegInTop_7_94[27] , \wRegInTop_7_94[26] , \wRegInTop_7_94[25] , 
        \wRegInTop_7_94[24] , \wRegInTop_7_94[23] , \wRegInTop_7_94[22] , 
        \wRegInTop_7_94[21] , \wRegInTop_7_94[20] , \wRegInTop_7_94[19] , 
        \wRegInTop_7_94[18] , \wRegInTop_7_94[17] , \wRegInTop_7_94[16] , 
        \wRegInTop_7_94[15] , \wRegInTop_7_94[14] , \wRegInTop_7_94[13] , 
        \wRegInTop_7_94[12] , \wRegInTop_7_94[11] , \wRegInTop_7_94[10] , 
        \wRegInTop_7_94[9] , \wRegInTop_7_94[8] , \wRegInTop_7_94[7] , 
        \wRegInTop_7_94[6] , \wRegInTop_7_94[5] , \wRegInTop_7_94[4] , 
        \wRegInTop_7_94[3] , \wRegInTop_7_94[2] , \wRegInTop_7_94[1] , 
        \wRegInTop_7_94[0] }), .R_WR(\wRegEnTop_7_95[0] ), .R_In({
        \wRegOut_7_95[31] , \wRegOut_7_95[30] , \wRegOut_7_95[29] , 
        \wRegOut_7_95[28] , \wRegOut_7_95[27] , \wRegOut_7_95[26] , 
        \wRegOut_7_95[25] , \wRegOut_7_95[24] , \wRegOut_7_95[23] , 
        \wRegOut_7_95[22] , \wRegOut_7_95[21] , \wRegOut_7_95[20] , 
        \wRegOut_7_95[19] , \wRegOut_7_95[18] , \wRegOut_7_95[17] , 
        \wRegOut_7_95[16] , \wRegOut_7_95[15] , \wRegOut_7_95[14] , 
        \wRegOut_7_95[13] , \wRegOut_7_95[12] , \wRegOut_7_95[11] , 
        \wRegOut_7_95[10] , \wRegOut_7_95[9] , \wRegOut_7_95[8] , 
        \wRegOut_7_95[7] , \wRegOut_7_95[6] , \wRegOut_7_95[5] , 
        \wRegOut_7_95[4] , \wRegOut_7_95[3] , \wRegOut_7_95[2] , 
        \wRegOut_7_95[1] , \wRegOut_7_95[0] }), .R_Out({\wRegInTop_7_95[31] , 
        \wRegInTop_7_95[30] , \wRegInTop_7_95[29] , \wRegInTop_7_95[28] , 
        \wRegInTop_7_95[27] , \wRegInTop_7_95[26] , \wRegInTop_7_95[25] , 
        \wRegInTop_7_95[24] , \wRegInTop_7_95[23] , \wRegInTop_7_95[22] , 
        \wRegInTop_7_95[21] , \wRegInTop_7_95[20] , \wRegInTop_7_95[19] , 
        \wRegInTop_7_95[18] , \wRegInTop_7_95[17] , \wRegInTop_7_95[16] , 
        \wRegInTop_7_95[15] , \wRegInTop_7_95[14] , \wRegInTop_7_95[13] , 
        \wRegInTop_7_95[12] , \wRegInTop_7_95[11] , \wRegInTop_7_95[10] , 
        \wRegInTop_7_95[9] , \wRegInTop_7_95[8] , \wRegInTop_7_95[7] , 
        \wRegInTop_7_95[6] , \wRegInTop_7_95[5] , \wRegInTop_7_95[4] , 
        \wRegInTop_7_95[3] , \wRegInTop_7_95[2] , \wRegInTop_7_95[1] , 
        \wRegInTop_7_95[0] }) );
    BHeap_Node_WIDTH32 BHN_6_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_60[0] ), .P_In({\wRegOut_6_60[31] , 
        \wRegOut_6_60[30] , \wRegOut_6_60[29] , \wRegOut_6_60[28] , 
        \wRegOut_6_60[27] , \wRegOut_6_60[26] , \wRegOut_6_60[25] , 
        \wRegOut_6_60[24] , \wRegOut_6_60[23] , \wRegOut_6_60[22] , 
        \wRegOut_6_60[21] , \wRegOut_6_60[20] , \wRegOut_6_60[19] , 
        \wRegOut_6_60[18] , \wRegOut_6_60[17] , \wRegOut_6_60[16] , 
        \wRegOut_6_60[15] , \wRegOut_6_60[14] , \wRegOut_6_60[13] , 
        \wRegOut_6_60[12] , \wRegOut_6_60[11] , \wRegOut_6_60[10] , 
        \wRegOut_6_60[9] , \wRegOut_6_60[8] , \wRegOut_6_60[7] , 
        \wRegOut_6_60[6] , \wRegOut_6_60[5] , \wRegOut_6_60[4] , 
        \wRegOut_6_60[3] , \wRegOut_6_60[2] , \wRegOut_6_60[1] , 
        \wRegOut_6_60[0] }), .P_Out({\wRegInBot_6_60[31] , 
        \wRegInBot_6_60[30] , \wRegInBot_6_60[29] , \wRegInBot_6_60[28] , 
        \wRegInBot_6_60[27] , \wRegInBot_6_60[26] , \wRegInBot_6_60[25] , 
        \wRegInBot_6_60[24] , \wRegInBot_6_60[23] , \wRegInBot_6_60[22] , 
        \wRegInBot_6_60[21] , \wRegInBot_6_60[20] , \wRegInBot_6_60[19] , 
        \wRegInBot_6_60[18] , \wRegInBot_6_60[17] , \wRegInBot_6_60[16] , 
        \wRegInBot_6_60[15] , \wRegInBot_6_60[14] , \wRegInBot_6_60[13] , 
        \wRegInBot_6_60[12] , \wRegInBot_6_60[11] , \wRegInBot_6_60[10] , 
        \wRegInBot_6_60[9] , \wRegInBot_6_60[8] , \wRegInBot_6_60[7] , 
        \wRegInBot_6_60[6] , \wRegInBot_6_60[5] , \wRegInBot_6_60[4] , 
        \wRegInBot_6_60[3] , \wRegInBot_6_60[2] , \wRegInBot_6_60[1] , 
        \wRegInBot_6_60[0] }), .L_WR(\wRegEnTop_7_120[0] ), .L_In({
        \wRegOut_7_120[31] , \wRegOut_7_120[30] , \wRegOut_7_120[29] , 
        \wRegOut_7_120[28] , \wRegOut_7_120[27] , \wRegOut_7_120[26] , 
        \wRegOut_7_120[25] , \wRegOut_7_120[24] , \wRegOut_7_120[23] , 
        \wRegOut_7_120[22] , \wRegOut_7_120[21] , \wRegOut_7_120[20] , 
        \wRegOut_7_120[19] , \wRegOut_7_120[18] , \wRegOut_7_120[17] , 
        \wRegOut_7_120[16] , \wRegOut_7_120[15] , \wRegOut_7_120[14] , 
        \wRegOut_7_120[13] , \wRegOut_7_120[12] , \wRegOut_7_120[11] , 
        \wRegOut_7_120[10] , \wRegOut_7_120[9] , \wRegOut_7_120[8] , 
        \wRegOut_7_120[7] , \wRegOut_7_120[6] , \wRegOut_7_120[5] , 
        \wRegOut_7_120[4] , \wRegOut_7_120[3] , \wRegOut_7_120[2] , 
        \wRegOut_7_120[1] , \wRegOut_7_120[0] }), .L_Out({
        \wRegInTop_7_120[31] , \wRegInTop_7_120[30] , \wRegInTop_7_120[29] , 
        \wRegInTop_7_120[28] , \wRegInTop_7_120[27] , \wRegInTop_7_120[26] , 
        \wRegInTop_7_120[25] , \wRegInTop_7_120[24] , \wRegInTop_7_120[23] , 
        \wRegInTop_7_120[22] , \wRegInTop_7_120[21] , \wRegInTop_7_120[20] , 
        \wRegInTop_7_120[19] , \wRegInTop_7_120[18] , \wRegInTop_7_120[17] , 
        \wRegInTop_7_120[16] , \wRegInTop_7_120[15] , \wRegInTop_7_120[14] , 
        \wRegInTop_7_120[13] , \wRegInTop_7_120[12] , \wRegInTop_7_120[11] , 
        \wRegInTop_7_120[10] , \wRegInTop_7_120[9] , \wRegInTop_7_120[8] , 
        \wRegInTop_7_120[7] , \wRegInTop_7_120[6] , \wRegInTop_7_120[5] , 
        \wRegInTop_7_120[4] , \wRegInTop_7_120[3] , \wRegInTop_7_120[2] , 
        \wRegInTop_7_120[1] , \wRegInTop_7_120[0] }), .R_WR(
        \wRegEnTop_7_121[0] ), .R_In({\wRegOut_7_121[31] , \wRegOut_7_121[30] , 
        \wRegOut_7_121[29] , \wRegOut_7_121[28] , \wRegOut_7_121[27] , 
        \wRegOut_7_121[26] , \wRegOut_7_121[25] , \wRegOut_7_121[24] , 
        \wRegOut_7_121[23] , \wRegOut_7_121[22] , \wRegOut_7_121[21] , 
        \wRegOut_7_121[20] , \wRegOut_7_121[19] , \wRegOut_7_121[18] , 
        \wRegOut_7_121[17] , \wRegOut_7_121[16] , \wRegOut_7_121[15] , 
        \wRegOut_7_121[14] , \wRegOut_7_121[13] , \wRegOut_7_121[12] , 
        \wRegOut_7_121[11] , \wRegOut_7_121[10] , \wRegOut_7_121[9] , 
        \wRegOut_7_121[8] , \wRegOut_7_121[7] , \wRegOut_7_121[6] , 
        \wRegOut_7_121[5] , \wRegOut_7_121[4] , \wRegOut_7_121[3] , 
        \wRegOut_7_121[2] , \wRegOut_7_121[1] , \wRegOut_7_121[0] }), .R_Out({
        \wRegInTop_7_121[31] , \wRegInTop_7_121[30] , \wRegInTop_7_121[29] , 
        \wRegInTop_7_121[28] , \wRegInTop_7_121[27] , \wRegInTop_7_121[26] , 
        \wRegInTop_7_121[25] , \wRegInTop_7_121[24] , \wRegInTop_7_121[23] , 
        \wRegInTop_7_121[22] , \wRegInTop_7_121[21] , \wRegInTop_7_121[20] , 
        \wRegInTop_7_121[19] , \wRegInTop_7_121[18] , \wRegInTop_7_121[17] , 
        \wRegInTop_7_121[16] , \wRegInTop_7_121[15] , \wRegInTop_7_121[14] , 
        \wRegInTop_7_121[13] , \wRegInTop_7_121[12] , \wRegInTop_7_121[11] , 
        \wRegInTop_7_121[10] , \wRegInTop_7_121[9] , \wRegInTop_7_121[8] , 
        \wRegInTop_7_121[7] , \wRegInTop_7_121[6] , \wRegInTop_7_121[5] , 
        \wRegInTop_7_121[4] , \wRegInTop_7_121[3] , \wRegInTop_7_121[2] , 
        \wRegInTop_7_121[1] , \wRegInTop_7_121[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_16 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink48[31] , \ScanLink48[30] , \ScanLink48[29] , 
        \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , \ScanLink48[25] , 
        \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , \ScanLink48[21] , 
        \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , \ScanLink48[17] , 
        \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , \ScanLink48[13] , 
        \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , \ScanLink48[9] , 
        \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , \ScanLink48[5] , 
        \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , \ScanLink48[1] , 
        \ScanLink48[0] }), .ScanOut({\ScanLink47[31] , \ScanLink47[30] , 
        \ScanLink47[29] , \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , 
        \ScanLink47[25] , \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , 
        \ScanLink47[21] , \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , 
        \ScanLink47[17] , \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , 
        \ScanLink47[13] , \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , 
        \ScanLink47[9] , \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , 
        \ScanLink47[5] , \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , 
        \ScanLink47[1] , \ScanLink47[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_16[31] , \wRegOut_5_16[30] , 
        \wRegOut_5_16[29] , \wRegOut_5_16[28] , \wRegOut_5_16[27] , 
        \wRegOut_5_16[26] , \wRegOut_5_16[25] , \wRegOut_5_16[24] , 
        \wRegOut_5_16[23] , \wRegOut_5_16[22] , \wRegOut_5_16[21] , 
        \wRegOut_5_16[20] , \wRegOut_5_16[19] , \wRegOut_5_16[18] , 
        \wRegOut_5_16[17] , \wRegOut_5_16[16] , \wRegOut_5_16[15] , 
        \wRegOut_5_16[14] , \wRegOut_5_16[13] , \wRegOut_5_16[12] , 
        \wRegOut_5_16[11] , \wRegOut_5_16[10] , \wRegOut_5_16[9] , 
        \wRegOut_5_16[8] , \wRegOut_5_16[7] , \wRegOut_5_16[6] , 
        \wRegOut_5_16[5] , \wRegOut_5_16[4] , \wRegOut_5_16[3] , 
        \wRegOut_5_16[2] , \wRegOut_5_16[1] , \wRegOut_5_16[0] }), .Enable1(
        \wRegEnTop_5_16[0] ), .Enable2(\wRegEnBot_5_16[0] ), .In1({
        \wRegInTop_5_16[31] , \wRegInTop_5_16[30] , \wRegInTop_5_16[29] , 
        \wRegInTop_5_16[28] , \wRegInTop_5_16[27] , \wRegInTop_5_16[26] , 
        \wRegInTop_5_16[25] , \wRegInTop_5_16[24] , \wRegInTop_5_16[23] , 
        \wRegInTop_5_16[22] , \wRegInTop_5_16[21] , \wRegInTop_5_16[20] , 
        \wRegInTop_5_16[19] , \wRegInTop_5_16[18] , \wRegInTop_5_16[17] , 
        \wRegInTop_5_16[16] , \wRegInTop_5_16[15] , \wRegInTop_5_16[14] , 
        \wRegInTop_5_16[13] , \wRegInTop_5_16[12] , \wRegInTop_5_16[11] , 
        \wRegInTop_5_16[10] , \wRegInTop_5_16[9] , \wRegInTop_5_16[8] , 
        \wRegInTop_5_16[7] , \wRegInTop_5_16[6] , \wRegInTop_5_16[5] , 
        \wRegInTop_5_16[4] , \wRegInTop_5_16[3] , \wRegInTop_5_16[2] , 
        \wRegInTop_5_16[1] , \wRegInTop_5_16[0] }), .In2({\wRegInBot_5_16[31] , 
        \wRegInBot_5_16[30] , \wRegInBot_5_16[29] , \wRegInBot_5_16[28] , 
        \wRegInBot_5_16[27] , \wRegInBot_5_16[26] , \wRegInBot_5_16[25] , 
        \wRegInBot_5_16[24] , \wRegInBot_5_16[23] , \wRegInBot_5_16[22] , 
        \wRegInBot_5_16[21] , \wRegInBot_5_16[20] , \wRegInBot_5_16[19] , 
        \wRegInBot_5_16[18] , \wRegInBot_5_16[17] , \wRegInBot_5_16[16] , 
        \wRegInBot_5_16[15] , \wRegInBot_5_16[14] , \wRegInBot_5_16[13] , 
        \wRegInBot_5_16[12] , \wRegInBot_5_16[11] , \wRegInBot_5_16[10] , 
        \wRegInBot_5_16[9] , \wRegInBot_5_16[8] , \wRegInBot_5_16[7] , 
        \wRegInBot_5_16[6] , \wRegInBot_5_16[5] , \wRegInBot_5_16[4] , 
        \wRegInBot_5_16[3] , \wRegInBot_5_16[2] , \wRegInBot_5_16[1] , 
        \wRegInBot_5_16[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_31 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink63[31] , \ScanLink63[30] , \ScanLink63[29] , 
        \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , \ScanLink63[25] , 
        \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , \ScanLink63[21] , 
        \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , \ScanLink63[17] , 
        \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , \ScanLink63[13] , 
        \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , \ScanLink63[9] , 
        \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , \ScanLink63[5] , 
        \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , \ScanLink63[1] , 
        \ScanLink63[0] }), .ScanOut({\ScanLink62[31] , \ScanLink62[30] , 
        \ScanLink62[29] , \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , 
        \ScanLink62[25] , \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , 
        \ScanLink62[21] , \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , 
        \ScanLink62[17] , \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , 
        \ScanLink62[13] , \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , 
        \ScanLink62[9] , \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , 
        \ScanLink62[5] , \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , 
        \ScanLink62[1] , \ScanLink62[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_31[31] , \wRegOut_5_31[30] , 
        \wRegOut_5_31[29] , \wRegOut_5_31[28] , \wRegOut_5_31[27] , 
        \wRegOut_5_31[26] , \wRegOut_5_31[25] , \wRegOut_5_31[24] , 
        \wRegOut_5_31[23] , \wRegOut_5_31[22] , \wRegOut_5_31[21] , 
        \wRegOut_5_31[20] , \wRegOut_5_31[19] , \wRegOut_5_31[18] , 
        \wRegOut_5_31[17] , \wRegOut_5_31[16] , \wRegOut_5_31[15] , 
        \wRegOut_5_31[14] , \wRegOut_5_31[13] , \wRegOut_5_31[12] , 
        \wRegOut_5_31[11] , \wRegOut_5_31[10] , \wRegOut_5_31[9] , 
        \wRegOut_5_31[8] , \wRegOut_5_31[7] , \wRegOut_5_31[6] , 
        \wRegOut_5_31[5] , \wRegOut_5_31[4] , \wRegOut_5_31[3] , 
        \wRegOut_5_31[2] , \wRegOut_5_31[1] , \wRegOut_5_31[0] }), .Enable1(
        \wRegEnTop_5_31[0] ), .Enable2(\wRegEnBot_5_31[0] ), .In1({
        \wRegInTop_5_31[31] , \wRegInTop_5_31[30] , \wRegInTop_5_31[29] , 
        \wRegInTop_5_31[28] , \wRegInTop_5_31[27] , \wRegInTop_5_31[26] , 
        \wRegInTop_5_31[25] , \wRegInTop_5_31[24] , \wRegInTop_5_31[23] , 
        \wRegInTop_5_31[22] , \wRegInTop_5_31[21] , \wRegInTop_5_31[20] , 
        \wRegInTop_5_31[19] , \wRegInTop_5_31[18] , \wRegInTop_5_31[17] , 
        \wRegInTop_5_31[16] , \wRegInTop_5_31[15] , \wRegInTop_5_31[14] , 
        \wRegInTop_5_31[13] , \wRegInTop_5_31[12] , \wRegInTop_5_31[11] , 
        \wRegInTop_5_31[10] , \wRegInTop_5_31[9] , \wRegInTop_5_31[8] , 
        \wRegInTop_5_31[7] , \wRegInTop_5_31[6] , \wRegInTop_5_31[5] , 
        \wRegInTop_5_31[4] , \wRegInTop_5_31[3] , \wRegInTop_5_31[2] , 
        \wRegInTop_5_31[1] , \wRegInTop_5_31[0] }), .In2({\wRegInBot_5_31[31] , 
        \wRegInBot_5_31[30] , \wRegInBot_5_31[29] , \wRegInBot_5_31[28] , 
        \wRegInBot_5_31[27] , \wRegInBot_5_31[26] , \wRegInBot_5_31[25] , 
        \wRegInBot_5_31[24] , \wRegInBot_5_31[23] , \wRegInBot_5_31[22] , 
        \wRegInBot_5_31[21] , \wRegInBot_5_31[20] , \wRegInBot_5_31[19] , 
        \wRegInBot_5_31[18] , \wRegInBot_5_31[17] , \wRegInBot_5_31[16] , 
        \wRegInBot_5_31[15] , \wRegInBot_5_31[14] , \wRegInBot_5_31[13] , 
        \wRegInBot_5_31[12] , \wRegInBot_5_31[11] , \wRegInBot_5_31[10] , 
        \wRegInBot_5_31[9] , \wRegInBot_5_31[8] , \wRegInBot_5_31[7] , 
        \wRegInBot_5_31[6] , \wRegInBot_5_31[5] , \wRegInBot_5_31[4] , 
        \wRegInBot_5_31[3] , \wRegInBot_5_31[2] , \wRegInBot_5_31[1] , 
        \wRegInBot_5_31[0] }) );
    BHeap_Node_WIDTH32 BHN_5_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_19[0] ), .P_In({\wRegOut_5_19[31] , 
        \wRegOut_5_19[30] , \wRegOut_5_19[29] , \wRegOut_5_19[28] , 
        \wRegOut_5_19[27] , \wRegOut_5_19[26] , \wRegOut_5_19[25] , 
        \wRegOut_5_19[24] , \wRegOut_5_19[23] , \wRegOut_5_19[22] , 
        \wRegOut_5_19[21] , \wRegOut_5_19[20] , \wRegOut_5_19[19] , 
        \wRegOut_5_19[18] , \wRegOut_5_19[17] , \wRegOut_5_19[16] , 
        \wRegOut_5_19[15] , \wRegOut_5_19[14] , \wRegOut_5_19[13] , 
        \wRegOut_5_19[12] , \wRegOut_5_19[11] , \wRegOut_5_19[10] , 
        \wRegOut_5_19[9] , \wRegOut_5_19[8] , \wRegOut_5_19[7] , 
        \wRegOut_5_19[6] , \wRegOut_5_19[5] , \wRegOut_5_19[4] , 
        \wRegOut_5_19[3] , \wRegOut_5_19[2] , \wRegOut_5_19[1] , 
        \wRegOut_5_19[0] }), .P_Out({\wRegInBot_5_19[31] , 
        \wRegInBot_5_19[30] , \wRegInBot_5_19[29] , \wRegInBot_5_19[28] , 
        \wRegInBot_5_19[27] , \wRegInBot_5_19[26] , \wRegInBot_5_19[25] , 
        \wRegInBot_5_19[24] , \wRegInBot_5_19[23] , \wRegInBot_5_19[22] , 
        \wRegInBot_5_19[21] , \wRegInBot_5_19[20] , \wRegInBot_5_19[19] , 
        \wRegInBot_5_19[18] , \wRegInBot_5_19[17] , \wRegInBot_5_19[16] , 
        \wRegInBot_5_19[15] , \wRegInBot_5_19[14] , \wRegInBot_5_19[13] , 
        \wRegInBot_5_19[12] , \wRegInBot_5_19[11] , \wRegInBot_5_19[10] , 
        \wRegInBot_5_19[9] , \wRegInBot_5_19[8] , \wRegInBot_5_19[7] , 
        \wRegInBot_5_19[6] , \wRegInBot_5_19[5] , \wRegInBot_5_19[4] , 
        \wRegInBot_5_19[3] , \wRegInBot_5_19[2] , \wRegInBot_5_19[1] , 
        \wRegInBot_5_19[0] }), .L_WR(\wRegEnTop_6_38[0] ), .L_In({
        \wRegOut_6_38[31] , \wRegOut_6_38[30] , \wRegOut_6_38[29] , 
        \wRegOut_6_38[28] , \wRegOut_6_38[27] , \wRegOut_6_38[26] , 
        \wRegOut_6_38[25] , \wRegOut_6_38[24] , \wRegOut_6_38[23] , 
        \wRegOut_6_38[22] , \wRegOut_6_38[21] , \wRegOut_6_38[20] , 
        \wRegOut_6_38[19] , \wRegOut_6_38[18] , \wRegOut_6_38[17] , 
        \wRegOut_6_38[16] , \wRegOut_6_38[15] , \wRegOut_6_38[14] , 
        \wRegOut_6_38[13] , \wRegOut_6_38[12] , \wRegOut_6_38[11] , 
        \wRegOut_6_38[10] , \wRegOut_6_38[9] , \wRegOut_6_38[8] , 
        \wRegOut_6_38[7] , \wRegOut_6_38[6] , \wRegOut_6_38[5] , 
        \wRegOut_6_38[4] , \wRegOut_6_38[3] , \wRegOut_6_38[2] , 
        \wRegOut_6_38[1] , \wRegOut_6_38[0] }), .L_Out({\wRegInTop_6_38[31] , 
        \wRegInTop_6_38[30] , \wRegInTop_6_38[29] , \wRegInTop_6_38[28] , 
        \wRegInTop_6_38[27] , \wRegInTop_6_38[26] , \wRegInTop_6_38[25] , 
        \wRegInTop_6_38[24] , \wRegInTop_6_38[23] , \wRegInTop_6_38[22] , 
        \wRegInTop_6_38[21] , \wRegInTop_6_38[20] , \wRegInTop_6_38[19] , 
        \wRegInTop_6_38[18] , \wRegInTop_6_38[17] , \wRegInTop_6_38[16] , 
        \wRegInTop_6_38[15] , \wRegInTop_6_38[14] , \wRegInTop_6_38[13] , 
        \wRegInTop_6_38[12] , \wRegInTop_6_38[11] , \wRegInTop_6_38[10] , 
        \wRegInTop_6_38[9] , \wRegInTop_6_38[8] , \wRegInTop_6_38[7] , 
        \wRegInTop_6_38[6] , \wRegInTop_6_38[5] , \wRegInTop_6_38[4] , 
        \wRegInTop_6_38[3] , \wRegInTop_6_38[2] , \wRegInTop_6_38[1] , 
        \wRegInTop_6_38[0] }), .R_WR(\wRegEnTop_6_39[0] ), .R_In({
        \wRegOut_6_39[31] , \wRegOut_6_39[30] , \wRegOut_6_39[29] , 
        \wRegOut_6_39[28] , \wRegOut_6_39[27] , \wRegOut_6_39[26] , 
        \wRegOut_6_39[25] , \wRegOut_6_39[24] , \wRegOut_6_39[23] , 
        \wRegOut_6_39[22] , \wRegOut_6_39[21] , \wRegOut_6_39[20] , 
        \wRegOut_6_39[19] , \wRegOut_6_39[18] , \wRegOut_6_39[17] , 
        \wRegOut_6_39[16] , \wRegOut_6_39[15] , \wRegOut_6_39[14] , 
        \wRegOut_6_39[13] , \wRegOut_6_39[12] , \wRegOut_6_39[11] , 
        \wRegOut_6_39[10] , \wRegOut_6_39[9] , \wRegOut_6_39[8] , 
        \wRegOut_6_39[7] , \wRegOut_6_39[6] , \wRegOut_6_39[5] , 
        \wRegOut_6_39[4] , \wRegOut_6_39[3] , \wRegOut_6_39[2] , 
        \wRegOut_6_39[1] , \wRegOut_6_39[0] }), .R_Out({\wRegInTop_6_39[31] , 
        \wRegInTop_6_39[30] , \wRegInTop_6_39[29] , \wRegInTop_6_39[28] , 
        \wRegInTop_6_39[27] , \wRegInTop_6_39[26] , \wRegInTop_6_39[25] , 
        \wRegInTop_6_39[24] , \wRegInTop_6_39[23] , \wRegInTop_6_39[22] , 
        \wRegInTop_6_39[21] , \wRegInTop_6_39[20] , \wRegInTop_6_39[19] , 
        \wRegInTop_6_39[18] , \wRegInTop_6_39[17] , \wRegInTop_6_39[16] , 
        \wRegInTop_6_39[15] , \wRegInTop_6_39[14] , \wRegInTop_6_39[13] , 
        \wRegInTop_6_39[12] , \wRegInTop_6_39[11] , \wRegInTop_6_39[10] , 
        \wRegInTop_6_39[9] , \wRegInTop_6_39[8] , \wRegInTop_6_39[7] , 
        \wRegInTop_6_39[6] , \wRegInTop_6_39[5] , \wRegInTop_6_39[4] , 
        \wRegInTop_6_39[3] , \wRegInTop_6_39[2] , \wRegInTop_6_39[1] , 
        \wRegInTop_6_39[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_26 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink90[31] , \ScanLink90[30] , \ScanLink90[29] , 
        \ScanLink90[28] , \ScanLink90[27] , \ScanLink90[26] , \ScanLink90[25] , 
        \ScanLink90[24] , \ScanLink90[23] , \ScanLink90[22] , \ScanLink90[21] , 
        \ScanLink90[20] , \ScanLink90[19] , \ScanLink90[18] , \ScanLink90[17] , 
        \ScanLink90[16] , \ScanLink90[15] , \ScanLink90[14] , \ScanLink90[13] , 
        \ScanLink90[12] , \ScanLink90[11] , \ScanLink90[10] , \ScanLink90[9] , 
        \ScanLink90[8] , \ScanLink90[7] , \ScanLink90[6] , \ScanLink90[5] , 
        \ScanLink90[4] , \ScanLink90[3] , \ScanLink90[2] , \ScanLink90[1] , 
        \ScanLink90[0] }), .ScanOut({\ScanLink89[31] , \ScanLink89[30] , 
        \ScanLink89[29] , \ScanLink89[28] , \ScanLink89[27] , \ScanLink89[26] , 
        \ScanLink89[25] , \ScanLink89[24] , \ScanLink89[23] , \ScanLink89[22] , 
        \ScanLink89[21] , \ScanLink89[20] , \ScanLink89[19] , \ScanLink89[18] , 
        \ScanLink89[17] , \ScanLink89[16] , \ScanLink89[15] , \ScanLink89[14] , 
        \ScanLink89[13] , \ScanLink89[12] , \ScanLink89[11] , \ScanLink89[10] , 
        \ScanLink89[9] , \ScanLink89[8] , \ScanLink89[7] , \ScanLink89[6] , 
        \ScanLink89[5] , \ScanLink89[4] , \ScanLink89[3] , \ScanLink89[2] , 
        \ScanLink89[1] , \ScanLink89[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_26[31] , \wRegOut_6_26[30] , 
        \wRegOut_6_26[29] , \wRegOut_6_26[28] , \wRegOut_6_26[27] , 
        \wRegOut_6_26[26] , \wRegOut_6_26[25] , \wRegOut_6_26[24] , 
        \wRegOut_6_26[23] , \wRegOut_6_26[22] , \wRegOut_6_26[21] , 
        \wRegOut_6_26[20] , \wRegOut_6_26[19] , \wRegOut_6_26[18] , 
        \wRegOut_6_26[17] , \wRegOut_6_26[16] , \wRegOut_6_26[15] , 
        \wRegOut_6_26[14] , \wRegOut_6_26[13] , \wRegOut_6_26[12] , 
        \wRegOut_6_26[11] , \wRegOut_6_26[10] , \wRegOut_6_26[9] , 
        \wRegOut_6_26[8] , \wRegOut_6_26[7] , \wRegOut_6_26[6] , 
        \wRegOut_6_26[5] , \wRegOut_6_26[4] , \wRegOut_6_26[3] , 
        \wRegOut_6_26[2] , \wRegOut_6_26[1] , \wRegOut_6_26[0] }), .Enable1(
        \wRegEnTop_6_26[0] ), .Enable2(\wRegEnBot_6_26[0] ), .In1({
        \wRegInTop_6_26[31] , \wRegInTop_6_26[30] , \wRegInTop_6_26[29] , 
        \wRegInTop_6_26[28] , \wRegInTop_6_26[27] , \wRegInTop_6_26[26] , 
        \wRegInTop_6_26[25] , \wRegInTop_6_26[24] , \wRegInTop_6_26[23] , 
        \wRegInTop_6_26[22] , \wRegInTop_6_26[21] , \wRegInTop_6_26[20] , 
        \wRegInTop_6_26[19] , \wRegInTop_6_26[18] , \wRegInTop_6_26[17] , 
        \wRegInTop_6_26[16] , \wRegInTop_6_26[15] , \wRegInTop_6_26[14] , 
        \wRegInTop_6_26[13] , \wRegInTop_6_26[12] , \wRegInTop_6_26[11] , 
        \wRegInTop_6_26[10] , \wRegInTop_6_26[9] , \wRegInTop_6_26[8] , 
        \wRegInTop_6_26[7] , \wRegInTop_6_26[6] , \wRegInTop_6_26[5] , 
        \wRegInTop_6_26[4] , \wRegInTop_6_26[3] , \wRegInTop_6_26[2] , 
        \wRegInTop_6_26[1] , \wRegInTop_6_26[0] }), .In2({\wRegInBot_6_26[31] , 
        \wRegInBot_6_26[30] , \wRegInBot_6_26[29] , \wRegInBot_6_26[28] , 
        \wRegInBot_6_26[27] , \wRegInBot_6_26[26] , \wRegInBot_6_26[25] , 
        \wRegInBot_6_26[24] , \wRegInBot_6_26[23] , \wRegInBot_6_26[22] , 
        \wRegInBot_6_26[21] , \wRegInBot_6_26[20] , \wRegInBot_6_26[19] , 
        \wRegInBot_6_26[18] , \wRegInBot_6_26[17] , \wRegInBot_6_26[16] , 
        \wRegInBot_6_26[15] , \wRegInBot_6_26[14] , \wRegInBot_6_26[13] , 
        \wRegInBot_6_26[12] , \wRegInBot_6_26[11] , \wRegInBot_6_26[10] , 
        \wRegInBot_6_26[9] , \wRegInBot_6_26[8] , \wRegInBot_6_26[7] , 
        \wRegInBot_6_26[6] , \wRegInBot_6_26[5] , \wRegInBot_6_26[4] , 
        \wRegInBot_6_26[3] , \wRegInBot_6_26[2] , \wRegInBot_6_26[1] , 
        \wRegInBot_6_26[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_75 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink203[31] , \ScanLink203[30] , \ScanLink203[29] , 
        \ScanLink203[28] , \ScanLink203[27] , \ScanLink203[26] , 
        \ScanLink203[25] , \ScanLink203[24] , \ScanLink203[23] , 
        \ScanLink203[22] , \ScanLink203[21] , \ScanLink203[20] , 
        \ScanLink203[19] , \ScanLink203[18] , \ScanLink203[17] , 
        \ScanLink203[16] , \ScanLink203[15] , \ScanLink203[14] , 
        \ScanLink203[13] , \ScanLink203[12] , \ScanLink203[11] , 
        \ScanLink203[10] , \ScanLink203[9] , \ScanLink203[8] , 
        \ScanLink203[7] , \ScanLink203[6] , \ScanLink203[5] , \ScanLink203[4] , 
        \ScanLink203[3] , \ScanLink203[2] , \ScanLink203[1] , \ScanLink203[0] 
        }), .ScanOut({\ScanLink202[31] , \ScanLink202[30] , \ScanLink202[29] , 
        \ScanLink202[28] , \ScanLink202[27] , \ScanLink202[26] , 
        \ScanLink202[25] , \ScanLink202[24] , \ScanLink202[23] , 
        \ScanLink202[22] , \ScanLink202[21] , \ScanLink202[20] , 
        \ScanLink202[19] , \ScanLink202[18] , \ScanLink202[17] , 
        \ScanLink202[16] , \ScanLink202[15] , \ScanLink202[14] , 
        \ScanLink202[13] , \ScanLink202[12] , \ScanLink202[11] , 
        \ScanLink202[10] , \ScanLink202[9] , \ScanLink202[8] , 
        \ScanLink202[7] , \ScanLink202[6] , \ScanLink202[5] , \ScanLink202[4] , 
        \ScanLink202[3] , \ScanLink202[2] , \ScanLink202[1] , \ScanLink202[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_75[31] , 
        \wRegOut_7_75[30] , \wRegOut_7_75[29] , \wRegOut_7_75[28] , 
        \wRegOut_7_75[27] , \wRegOut_7_75[26] , \wRegOut_7_75[25] , 
        \wRegOut_7_75[24] , \wRegOut_7_75[23] , \wRegOut_7_75[22] , 
        \wRegOut_7_75[21] , \wRegOut_7_75[20] , \wRegOut_7_75[19] , 
        \wRegOut_7_75[18] , \wRegOut_7_75[17] , \wRegOut_7_75[16] , 
        \wRegOut_7_75[15] , \wRegOut_7_75[14] , \wRegOut_7_75[13] , 
        \wRegOut_7_75[12] , \wRegOut_7_75[11] , \wRegOut_7_75[10] , 
        \wRegOut_7_75[9] , \wRegOut_7_75[8] , \wRegOut_7_75[7] , 
        \wRegOut_7_75[6] , \wRegOut_7_75[5] , \wRegOut_7_75[4] , 
        \wRegOut_7_75[3] , \wRegOut_7_75[2] , \wRegOut_7_75[1] , 
        \wRegOut_7_75[0] }), .Enable1(\wRegEnTop_7_75[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_75[31] , \wRegInTop_7_75[30] , \wRegInTop_7_75[29] , 
        \wRegInTop_7_75[28] , \wRegInTop_7_75[27] , \wRegInTop_7_75[26] , 
        \wRegInTop_7_75[25] , \wRegInTop_7_75[24] , \wRegInTop_7_75[23] , 
        \wRegInTop_7_75[22] , \wRegInTop_7_75[21] , \wRegInTop_7_75[20] , 
        \wRegInTop_7_75[19] , \wRegInTop_7_75[18] , \wRegInTop_7_75[17] , 
        \wRegInTop_7_75[16] , \wRegInTop_7_75[15] , \wRegInTop_7_75[14] , 
        \wRegInTop_7_75[13] , \wRegInTop_7_75[12] , \wRegInTop_7_75[11] , 
        \wRegInTop_7_75[10] , \wRegInTop_7_75[9] , \wRegInTop_7_75[8] , 
        \wRegInTop_7_75[7] , \wRegInTop_7_75[6] , \wRegInTop_7_75[5] , 
        \wRegInTop_7_75[4] , \wRegInTop_7_75[3] , \wRegInTop_7_75[2] , 
        \wRegInTop_7_75[1] , \wRegInTop_7_75[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_29[0] ), .P_In({\wRegOut_6_29[31] , 
        \wRegOut_6_29[30] , \wRegOut_6_29[29] , \wRegOut_6_29[28] , 
        \wRegOut_6_29[27] , \wRegOut_6_29[26] , \wRegOut_6_29[25] , 
        \wRegOut_6_29[24] , \wRegOut_6_29[23] , \wRegOut_6_29[22] , 
        \wRegOut_6_29[21] , \wRegOut_6_29[20] , \wRegOut_6_29[19] , 
        \wRegOut_6_29[18] , \wRegOut_6_29[17] , \wRegOut_6_29[16] , 
        \wRegOut_6_29[15] , \wRegOut_6_29[14] , \wRegOut_6_29[13] , 
        \wRegOut_6_29[12] , \wRegOut_6_29[11] , \wRegOut_6_29[10] , 
        \wRegOut_6_29[9] , \wRegOut_6_29[8] , \wRegOut_6_29[7] , 
        \wRegOut_6_29[6] , \wRegOut_6_29[5] , \wRegOut_6_29[4] , 
        \wRegOut_6_29[3] , \wRegOut_6_29[2] , \wRegOut_6_29[1] , 
        \wRegOut_6_29[0] }), .P_Out({\wRegInBot_6_29[31] , 
        \wRegInBot_6_29[30] , \wRegInBot_6_29[29] , \wRegInBot_6_29[28] , 
        \wRegInBot_6_29[27] , \wRegInBot_6_29[26] , \wRegInBot_6_29[25] , 
        \wRegInBot_6_29[24] , \wRegInBot_6_29[23] , \wRegInBot_6_29[22] , 
        \wRegInBot_6_29[21] , \wRegInBot_6_29[20] , \wRegInBot_6_29[19] , 
        \wRegInBot_6_29[18] , \wRegInBot_6_29[17] , \wRegInBot_6_29[16] , 
        \wRegInBot_6_29[15] , \wRegInBot_6_29[14] , \wRegInBot_6_29[13] , 
        \wRegInBot_6_29[12] , \wRegInBot_6_29[11] , \wRegInBot_6_29[10] , 
        \wRegInBot_6_29[9] , \wRegInBot_6_29[8] , \wRegInBot_6_29[7] , 
        \wRegInBot_6_29[6] , \wRegInBot_6_29[5] , \wRegInBot_6_29[4] , 
        \wRegInBot_6_29[3] , \wRegInBot_6_29[2] , \wRegInBot_6_29[1] , 
        \wRegInBot_6_29[0] }), .L_WR(\wRegEnTop_7_58[0] ), .L_In({
        \wRegOut_7_58[31] , \wRegOut_7_58[30] , \wRegOut_7_58[29] , 
        \wRegOut_7_58[28] , \wRegOut_7_58[27] , \wRegOut_7_58[26] , 
        \wRegOut_7_58[25] , \wRegOut_7_58[24] , \wRegOut_7_58[23] , 
        \wRegOut_7_58[22] , \wRegOut_7_58[21] , \wRegOut_7_58[20] , 
        \wRegOut_7_58[19] , \wRegOut_7_58[18] , \wRegOut_7_58[17] , 
        \wRegOut_7_58[16] , \wRegOut_7_58[15] , \wRegOut_7_58[14] , 
        \wRegOut_7_58[13] , \wRegOut_7_58[12] , \wRegOut_7_58[11] , 
        \wRegOut_7_58[10] , \wRegOut_7_58[9] , \wRegOut_7_58[8] , 
        \wRegOut_7_58[7] , \wRegOut_7_58[6] , \wRegOut_7_58[5] , 
        \wRegOut_7_58[4] , \wRegOut_7_58[3] , \wRegOut_7_58[2] , 
        \wRegOut_7_58[1] , \wRegOut_7_58[0] }), .L_Out({\wRegInTop_7_58[31] , 
        \wRegInTop_7_58[30] , \wRegInTop_7_58[29] , \wRegInTop_7_58[28] , 
        \wRegInTop_7_58[27] , \wRegInTop_7_58[26] , \wRegInTop_7_58[25] , 
        \wRegInTop_7_58[24] , \wRegInTop_7_58[23] , \wRegInTop_7_58[22] , 
        \wRegInTop_7_58[21] , \wRegInTop_7_58[20] , \wRegInTop_7_58[19] , 
        \wRegInTop_7_58[18] , \wRegInTop_7_58[17] , \wRegInTop_7_58[16] , 
        \wRegInTop_7_58[15] , \wRegInTop_7_58[14] , \wRegInTop_7_58[13] , 
        \wRegInTop_7_58[12] , \wRegInTop_7_58[11] , \wRegInTop_7_58[10] , 
        \wRegInTop_7_58[9] , \wRegInTop_7_58[8] , \wRegInTop_7_58[7] , 
        \wRegInTop_7_58[6] , \wRegInTop_7_58[5] , \wRegInTop_7_58[4] , 
        \wRegInTop_7_58[3] , \wRegInTop_7_58[2] , \wRegInTop_7_58[1] , 
        \wRegInTop_7_58[0] }), .R_WR(\wRegEnTop_7_59[0] ), .R_In({
        \wRegOut_7_59[31] , \wRegOut_7_59[30] , \wRegOut_7_59[29] , 
        \wRegOut_7_59[28] , \wRegOut_7_59[27] , \wRegOut_7_59[26] , 
        \wRegOut_7_59[25] , \wRegOut_7_59[24] , \wRegOut_7_59[23] , 
        \wRegOut_7_59[22] , \wRegOut_7_59[21] , \wRegOut_7_59[20] , 
        \wRegOut_7_59[19] , \wRegOut_7_59[18] , \wRegOut_7_59[17] , 
        \wRegOut_7_59[16] , \wRegOut_7_59[15] , \wRegOut_7_59[14] , 
        \wRegOut_7_59[13] , \wRegOut_7_59[12] , \wRegOut_7_59[11] , 
        \wRegOut_7_59[10] , \wRegOut_7_59[9] , \wRegOut_7_59[8] , 
        \wRegOut_7_59[7] , \wRegOut_7_59[6] , \wRegOut_7_59[5] , 
        \wRegOut_7_59[4] , \wRegOut_7_59[3] , \wRegOut_7_59[2] , 
        \wRegOut_7_59[1] , \wRegOut_7_59[0] }), .R_Out({\wRegInTop_7_59[31] , 
        \wRegInTop_7_59[30] , \wRegInTop_7_59[29] , \wRegInTop_7_59[28] , 
        \wRegInTop_7_59[27] , \wRegInTop_7_59[26] , \wRegInTop_7_59[25] , 
        \wRegInTop_7_59[24] , \wRegInTop_7_59[23] , \wRegInTop_7_59[22] , 
        \wRegInTop_7_59[21] , \wRegInTop_7_59[20] , \wRegInTop_7_59[19] , 
        \wRegInTop_7_59[18] , \wRegInTop_7_59[17] , \wRegInTop_7_59[16] , 
        \wRegInTop_7_59[15] , \wRegInTop_7_59[14] , \wRegInTop_7_59[13] , 
        \wRegInTop_7_59[12] , \wRegInTop_7_59[11] , \wRegInTop_7_59[10] , 
        \wRegInTop_7_59[9] , \wRegInTop_7_59[8] , \wRegInTop_7_59[7] , 
        \wRegInTop_7_59[6] , \wRegInTop_7_59[5] , \wRegInTop_7_59[4] , 
        \wRegInTop_7_59[3] , \wRegInTop_7_59[2] , \wRegInTop_7_59[1] , 
        \wRegInTop_7_59[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_52 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink180[31] , \ScanLink180[30] , \ScanLink180[29] , 
        \ScanLink180[28] , \ScanLink180[27] , \ScanLink180[26] , 
        \ScanLink180[25] , \ScanLink180[24] , \ScanLink180[23] , 
        \ScanLink180[22] , \ScanLink180[21] , \ScanLink180[20] , 
        \ScanLink180[19] , \ScanLink180[18] , \ScanLink180[17] , 
        \ScanLink180[16] , \ScanLink180[15] , \ScanLink180[14] , 
        \ScanLink180[13] , \ScanLink180[12] , \ScanLink180[11] , 
        \ScanLink180[10] , \ScanLink180[9] , \ScanLink180[8] , 
        \ScanLink180[7] , \ScanLink180[6] , \ScanLink180[5] , \ScanLink180[4] , 
        \ScanLink180[3] , \ScanLink180[2] , \ScanLink180[1] , \ScanLink180[0] 
        }), .ScanOut({\ScanLink179[31] , \ScanLink179[30] , \ScanLink179[29] , 
        \ScanLink179[28] , \ScanLink179[27] , \ScanLink179[26] , 
        \ScanLink179[25] , \ScanLink179[24] , \ScanLink179[23] , 
        \ScanLink179[22] , \ScanLink179[21] , \ScanLink179[20] , 
        \ScanLink179[19] , \ScanLink179[18] , \ScanLink179[17] , 
        \ScanLink179[16] , \ScanLink179[15] , \ScanLink179[14] , 
        \ScanLink179[13] , \ScanLink179[12] , \ScanLink179[11] , 
        \ScanLink179[10] , \ScanLink179[9] , \ScanLink179[8] , 
        \ScanLink179[7] , \ScanLink179[6] , \ScanLink179[5] , \ScanLink179[4] , 
        \ScanLink179[3] , \ScanLink179[2] , \ScanLink179[1] , \ScanLink179[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_52[31] , 
        \wRegOut_7_52[30] , \wRegOut_7_52[29] , \wRegOut_7_52[28] , 
        \wRegOut_7_52[27] , \wRegOut_7_52[26] , \wRegOut_7_52[25] , 
        \wRegOut_7_52[24] , \wRegOut_7_52[23] , \wRegOut_7_52[22] , 
        \wRegOut_7_52[21] , \wRegOut_7_52[20] , \wRegOut_7_52[19] , 
        \wRegOut_7_52[18] , \wRegOut_7_52[17] , \wRegOut_7_52[16] , 
        \wRegOut_7_52[15] , \wRegOut_7_52[14] , \wRegOut_7_52[13] , 
        \wRegOut_7_52[12] , \wRegOut_7_52[11] , \wRegOut_7_52[10] , 
        \wRegOut_7_52[9] , \wRegOut_7_52[8] , \wRegOut_7_52[7] , 
        \wRegOut_7_52[6] , \wRegOut_7_52[5] , \wRegOut_7_52[4] , 
        \wRegOut_7_52[3] , \wRegOut_7_52[2] , \wRegOut_7_52[1] , 
        \wRegOut_7_52[0] }), .Enable1(\wRegEnTop_7_52[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_52[31] , \wRegInTop_7_52[30] , \wRegInTop_7_52[29] , 
        \wRegInTop_7_52[28] , \wRegInTop_7_52[27] , \wRegInTop_7_52[26] , 
        \wRegInTop_7_52[25] , \wRegInTop_7_52[24] , \wRegInTop_7_52[23] , 
        \wRegInTop_7_52[22] , \wRegInTop_7_52[21] , \wRegInTop_7_52[20] , 
        \wRegInTop_7_52[19] , \wRegInTop_7_52[18] , \wRegInTop_7_52[17] , 
        \wRegInTop_7_52[16] , \wRegInTop_7_52[15] , \wRegInTop_7_52[14] , 
        \wRegInTop_7_52[13] , \wRegInTop_7_52[12] , \wRegInTop_7_52[11] , 
        \wRegInTop_7_52[10] , \wRegInTop_7_52[9] , \wRegInTop_7_52[8] , 
        \wRegInTop_7_52[7] , \wRegInTop_7_52[6] , \wRegInTop_7_52[5] , 
        \wRegInTop_7_52[4] , \wRegInTop_7_52[3] , \wRegInTop_7_52[2] , 
        \wRegInTop_7_52[1] , \wRegInTop_7_52[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink8[31] , \ScanLink8[30] , \ScanLink8[29] , 
        \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , \ScanLink8[25] , 
        \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , \ScanLink8[21] , 
        \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , \ScanLink8[17] , 
        \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , \ScanLink8[13] , 
        \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , \ScanLink8[9] , 
        \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , \ScanLink8[5] , 
        \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , \ScanLink8[1] , 
        \ScanLink8[0] }), .ScanOut({\ScanLink7[31] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , 
        \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , 
        \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , 
        \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , 
        \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , 
        \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_0[31] , \wRegOut_3_0[30] , \wRegOut_3_0[29] , 
        \wRegOut_3_0[28] , \wRegOut_3_0[27] , \wRegOut_3_0[26] , 
        \wRegOut_3_0[25] , \wRegOut_3_0[24] , \wRegOut_3_0[23] , 
        \wRegOut_3_0[22] , \wRegOut_3_0[21] , \wRegOut_3_0[20] , 
        \wRegOut_3_0[19] , \wRegOut_3_0[18] , \wRegOut_3_0[17] , 
        \wRegOut_3_0[16] , \wRegOut_3_0[15] , \wRegOut_3_0[14] , 
        \wRegOut_3_0[13] , \wRegOut_3_0[12] , \wRegOut_3_0[11] , 
        \wRegOut_3_0[10] , \wRegOut_3_0[9] , \wRegOut_3_0[8] , 
        \wRegOut_3_0[7] , \wRegOut_3_0[6] , \wRegOut_3_0[5] , \wRegOut_3_0[4] , 
        \wRegOut_3_0[3] , \wRegOut_3_0[2] , \wRegOut_3_0[1] , \wRegOut_3_0[0] 
        }), .Enable1(\wRegEnTop_3_0[0] ), .Enable2(\wRegEnBot_3_0[0] ), .In1({
        \wRegInTop_3_0[31] , \wRegInTop_3_0[30] , \wRegInTop_3_0[29] , 
        \wRegInTop_3_0[28] , \wRegInTop_3_0[27] , \wRegInTop_3_0[26] , 
        \wRegInTop_3_0[25] , \wRegInTop_3_0[24] , \wRegInTop_3_0[23] , 
        \wRegInTop_3_0[22] , \wRegInTop_3_0[21] , \wRegInTop_3_0[20] , 
        \wRegInTop_3_0[19] , \wRegInTop_3_0[18] , \wRegInTop_3_0[17] , 
        \wRegInTop_3_0[16] , \wRegInTop_3_0[15] , \wRegInTop_3_0[14] , 
        \wRegInTop_3_0[13] , \wRegInTop_3_0[12] , \wRegInTop_3_0[11] , 
        \wRegInTop_3_0[10] , \wRegInTop_3_0[9] , \wRegInTop_3_0[8] , 
        \wRegInTop_3_0[7] , \wRegInTop_3_0[6] , \wRegInTop_3_0[5] , 
        \wRegInTop_3_0[4] , \wRegInTop_3_0[3] , \wRegInTop_3_0[2] , 
        \wRegInTop_3_0[1] , \wRegInTop_3_0[0] }), .In2({\wRegInBot_3_0[31] , 
        \wRegInBot_3_0[30] , \wRegInBot_3_0[29] , \wRegInBot_3_0[28] , 
        \wRegInBot_3_0[27] , \wRegInBot_3_0[26] , \wRegInBot_3_0[25] , 
        \wRegInBot_3_0[24] , \wRegInBot_3_0[23] , \wRegInBot_3_0[22] , 
        \wRegInBot_3_0[21] , \wRegInBot_3_0[20] , \wRegInBot_3_0[19] , 
        \wRegInBot_3_0[18] , \wRegInBot_3_0[17] , \wRegInBot_3_0[16] , 
        \wRegInBot_3_0[15] , \wRegInBot_3_0[14] , \wRegInBot_3_0[13] , 
        \wRegInBot_3_0[12] , \wRegInBot_3_0[11] , \wRegInBot_3_0[10] , 
        \wRegInBot_3_0[9] , \wRegInBot_3_0[8] , \wRegInBot_3_0[7] , 
        \wRegInBot_3_0[6] , \wRegInBot_3_0[5] , \wRegInBot_3_0[4] , 
        \wRegInBot_3_0[3] , \wRegInBot_3_0[2] , \wRegInBot_3_0[1] , 
        \wRegInBot_3_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_23 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink55[31] , \ScanLink55[30] , \ScanLink55[29] , 
        \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , \ScanLink55[25] , 
        \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , \ScanLink55[21] , 
        \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , \ScanLink55[17] , 
        \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , \ScanLink55[13] , 
        \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , \ScanLink55[9] , 
        \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , \ScanLink55[5] , 
        \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , \ScanLink55[1] , 
        \ScanLink55[0] }), .ScanOut({\ScanLink54[31] , \ScanLink54[30] , 
        \ScanLink54[29] , \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , 
        \ScanLink54[25] , \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , 
        \ScanLink54[21] , \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , 
        \ScanLink54[17] , \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , 
        \ScanLink54[13] , \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , 
        \ScanLink54[9] , \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , 
        \ScanLink54[5] , \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , 
        \ScanLink54[1] , \ScanLink54[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_23[31] , \wRegOut_5_23[30] , 
        \wRegOut_5_23[29] , \wRegOut_5_23[28] , \wRegOut_5_23[27] , 
        \wRegOut_5_23[26] , \wRegOut_5_23[25] , \wRegOut_5_23[24] , 
        \wRegOut_5_23[23] , \wRegOut_5_23[22] , \wRegOut_5_23[21] , 
        \wRegOut_5_23[20] , \wRegOut_5_23[19] , \wRegOut_5_23[18] , 
        \wRegOut_5_23[17] , \wRegOut_5_23[16] , \wRegOut_5_23[15] , 
        \wRegOut_5_23[14] , \wRegOut_5_23[13] , \wRegOut_5_23[12] , 
        \wRegOut_5_23[11] , \wRegOut_5_23[10] , \wRegOut_5_23[9] , 
        \wRegOut_5_23[8] , \wRegOut_5_23[7] , \wRegOut_5_23[6] , 
        \wRegOut_5_23[5] , \wRegOut_5_23[4] , \wRegOut_5_23[3] , 
        \wRegOut_5_23[2] , \wRegOut_5_23[1] , \wRegOut_5_23[0] }), .Enable1(
        \wRegEnTop_5_23[0] ), .Enable2(\wRegEnBot_5_23[0] ), .In1({
        \wRegInTop_5_23[31] , \wRegInTop_5_23[30] , \wRegInTop_5_23[29] , 
        \wRegInTop_5_23[28] , \wRegInTop_5_23[27] , \wRegInTop_5_23[26] , 
        \wRegInTop_5_23[25] , \wRegInTop_5_23[24] , \wRegInTop_5_23[23] , 
        \wRegInTop_5_23[22] , \wRegInTop_5_23[21] , \wRegInTop_5_23[20] , 
        \wRegInTop_5_23[19] , \wRegInTop_5_23[18] , \wRegInTop_5_23[17] , 
        \wRegInTop_5_23[16] , \wRegInTop_5_23[15] , \wRegInTop_5_23[14] , 
        \wRegInTop_5_23[13] , \wRegInTop_5_23[12] , \wRegInTop_5_23[11] , 
        \wRegInTop_5_23[10] , \wRegInTop_5_23[9] , \wRegInTop_5_23[8] , 
        \wRegInTop_5_23[7] , \wRegInTop_5_23[6] , \wRegInTop_5_23[5] , 
        \wRegInTop_5_23[4] , \wRegInTop_5_23[3] , \wRegInTop_5_23[2] , 
        \wRegInTop_5_23[1] , \wRegInTop_5_23[0] }), .In2({\wRegInBot_5_23[31] , 
        \wRegInBot_5_23[30] , \wRegInBot_5_23[29] , \wRegInBot_5_23[28] , 
        \wRegInBot_5_23[27] , \wRegInBot_5_23[26] , \wRegInBot_5_23[25] , 
        \wRegInBot_5_23[24] , \wRegInBot_5_23[23] , \wRegInBot_5_23[22] , 
        \wRegInBot_5_23[21] , \wRegInBot_5_23[20] , \wRegInBot_5_23[19] , 
        \wRegInBot_5_23[18] , \wRegInBot_5_23[17] , \wRegInBot_5_23[16] , 
        \wRegInBot_5_23[15] , \wRegInBot_5_23[14] , \wRegInBot_5_23[13] , 
        \wRegInBot_5_23[12] , \wRegInBot_5_23[11] , \wRegInBot_5_23[10] , 
        \wRegInBot_5_23[9] , \wRegInBot_5_23[8] , \wRegInBot_5_23[7] , 
        \wRegInBot_5_23[6] , \wRegInBot_5_23[5] , \wRegInBot_5_23[4] , 
        \wRegInBot_5_23[3] , \wRegInBot_5_23[2] , \wRegInBot_5_23[1] , 
        \wRegInBot_5_23[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink77[31] , \ScanLink77[30] , \ScanLink77[29] , 
        \ScanLink77[28] , \ScanLink77[27] , \ScanLink77[26] , \ScanLink77[25] , 
        \ScanLink77[24] , \ScanLink77[23] , \ScanLink77[22] , \ScanLink77[21] , 
        \ScanLink77[20] , \ScanLink77[19] , \ScanLink77[18] , \ScanLink77[17] , 
        \ScanLink77[16] , \ScanLink77[15] , \ScanLink77[14] , \ScanLink77[13] , 
        \ScanLink77[12] , \ScanLink77[11] , \ScanLink77[10] , \ScanLink77[9] , 
        \ScanLink77[8] , \ScanLink77[7] , \ScanLink77[6] , \ScanLink77[5] , 
        \ScanLink77[4] , \ScanLink77[3] , \ScanLink77[2] , \ScanLink77[1] , 
        \ScanLink77[0] }), .ScanOut({\ScanLink76[31] , \ScanLink76[30] , 
        \ScanLink76[29] , \ScanLink76[28] , \ScanLink76[27] , \ScanLink76[26] , 
        \ScanLink76[25] , \ScanLink76[24] , \ScanLink76[23] , \ScanLink76[22] , 
        \ScanLink76[21] , \ScanLink76[20] , \ScanLink76[19] , \ScanLink76[18] , 
        \ScanLink76[17] , \ScanLink76[16] , \ScanLink76[15] , \ScanLink76[14] , 
        \ScanLink76[13] , \ScanLink76[12] , \ScanLink76[11] , \ScanLink76[10] , 
        \ScanLink76[9] , \ScanLink76[8] , \ScanLink76[7] , \ScanLink76[6] , 
        \ScanLink76[5] , \ScanLink76[4] , \ScanLink76[3] , \ScanLink76[2] , 
        \ScanLink76[1] , \ScanLink76[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_13[31] , \wRegOut_6_13[30] , 
        \wRegOut_6_13[29] , \wRegOut_6_13[28] , \wRegOut_6_13[27] , 
        \wRegOut_6_13[26] , \wRegOut_6_13[25] , \wRegOut_6_13[24] , 
        \wRegOut_6_13[23] , \wRegOut_6_13[22] , \wRegOut_6_13[21] , 
        \wRegOut_6_13[20] , \wRegOut_6_13[19] , \wRegOut_6_13[18] , 
        \wRegOut_6_13[17] , \wRegOut_6_13[16] , \wRegOut_6_13[15] , 
        \wRegOut_6_13[14] , \wRegOut_6_13[13] , \wRegOut_6_13[12] , 
        \wRegOut_6_13[11] , \wRegOut_6_13[10] , \wRegOut_6_13[9] , 
        \wRegOut_6_13[8] , \wRegOut_6_13[7] , \wRegOut_6_13[6] , 
        \wRegOut_6_13[5] , \wRegOut_6_13[4] , \wRegOut_6_13[3] , 
        \wRegOut_6_13[2] , \wRegOut_6_13[1] , \wRegOut_6_13[0] }), .Enable1(
        \wRegEnTop_6_13[0] ), .Enable2(\wRegEnBot_6_13[0] ), .In1({
        \wRegInTop_6_13[31] , \wRegInTop_6_13[30] , \wRegInTop_6_13[29] , 
        \wRegInTop_6_13[28] , \wRegInTop_6_13[27] , \wRegInTop_6_13[26] , 
        \wRegInTop_6_13[25] , \wRegInTop_6_13[24] , \wRegInTop_6_13[23] , 
        \wRegInTop_6_13[22] , \wRegInTop_6_13[21] , \wRegInTop_6_13[20] , 
        \wRegInTop_6_13[19] , \wRegInTop_6_13[18] , \wRegInTop_6_13[17] , 
        \wRegInTop_6_13[16] , \wRegInTop_6_13[15] , \wRegInTop_6_13[14] , 
        \wRegInTop_6_13[13] , \wRegInTop_6_13[12] , \wRegInTop_6_13[11] , 
        \wRegInTop_6_13[10] , \wRegInTop_6_13[9] , \wRegInTop_6_13[8] , 
        \wRegInTop_6_13[7] , \wRegInTop_6_13[6] , \wRegInTop_6_13[5] , 
        \wRegInTop_6_13[4] , \wRegInTop_6_13[3] , \wRegInTop_6_13[2] , 
        \wRegInTop_6_13[1] , \wRegInTop_6_13[0] }), .In2({\wRegInBot_6_13[31] , 
        \wRegInBot_6_13[30] , \wRegInBot_6_13[29] , \wRegInBot_6_13[28] , 
        \wRegInBot_6_13[27] , \wRegInBot_6_13[26] , \wRegInBot_6_13[25] , 
        \wRegInBot_6_13[24] , \wRegInBot_6_13[23] , \wRegInBot_6_13[22] , 
        \wRegInBot_6_13[21] , \wRegInBot_6_13[20] , \wRegInBot_6_13[19] , 
        \wRegInBot_6_13[18] , \wRegInBot_6_13[17] , \wRegInBot_6_13[16] , 
        \wRegInBot_6_13[15] , \wRegInBot_6_13[14] , \wRegInBot_6_13[13] , 
        \wRegInBot_6_13[12] , \wRegInBot_6_13[11] , \wRegInBot_6_13[10] , 
        \wRegInBot_6_13[9] , \wRegInBot_6_13[8] , \wRegInBot_6_13[7] , 
        \wRegInBot_6_13[6] , \wRegInBot_6_13[5] , \wRegInBot_6_13[4] , 
        \wRegInBot_6_13[3] , \wRegInBot_6_13[2] , \wRegInBot_6_13[1] , 
        \wRegInBot_6_13[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_67 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink195[31] , \ScanLink195[30] , \ScanLink195[29] , 
        \ScanLink195[28] , \ScanLink195[27] , \ScanLink195[26] , 
        \ScanLink195[25] , \ScanLink195[24] , \ScanLink195[23] , 
        \ScanLink195[22] , \ScanLink195[21] , \ScanLink195[20] , 
        \ScanLink195[19] , \ScanLink195[18] , \ScanLink195[17] , 
        \ScanLink195[16] , \ScanLink195[15] , \ScanLink195[14] , 
        \ScanLink195[13] , \ScanLink195[12] , \ScanLink195[11] , 
        \ScanLink195[10] , \ScanLink195[9] , \ScanLink195[8] , 
        \ScanLink195[7] , \ScanLink195[6] , \ScanLink195[5] , \ScanLink195[4] , 
        \ScanLink195[3] , \ScanLink195[2] , \ScanLink195[1] , \ScanLink195[0] 
        }), .ScanOut({\ScanLink194[31] , \ScanLink194[30] , \ScanLink194[29] , 
        \ScanLink194[28] , \ScanLink194[27] , \ScanLink194[26] , 
        \ScanLink194[25] , \ScanLink194[24] , \ScanLink194[23] , 
        \ScanLink194[22] , \ScanLink194[21] , \ScanLink194[20] , 
        \ScanLink194[19] , \ScanLink194[18] , \ScanLink194[17] , 
        \ScanLink194[16] , \ScanLink194[15] , \ScanLink194[14] , 
        \ScanLink194[13] , \ScanLink194[12] , \ScanLink194[11] , 
        \ScanLink194[10] , \ScanLink194[9] , \ScanLink194[8] , 
        \ScanLink194[7] , \ScanLink194[6] , \ScanLink194[5] , \ScanLink194[4] , 
        \ScanLink194[3] , \ScanLink194[2] , \ScanLink194[1] , \ScanLink194[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_67[31] , 
        \wRegOut_7_67[30] , \wRegOut_7_67[29] , \wRegOut_7_67[28] , 
        \wRegOut_7_67[27] , \wRegOut_7_67[26] , \wRegOut_7_67[25] , 
        \wRegOut_7_67[24] , \wRegOut_7_67[23] , \wRegOut_7_67[22] , 
        \wRegOut_7_67[21] , \wRegOut_7_67[20] , \wRegOut_7_67[19] , 
        \wRegOut_7_67[18] , \wRegOut_7_67[17] , \wRegOut_7_67[16] , 
        \wRegOut_7_67[15] , \wRegOut_7_67[14] , \wRegOut_7_67[13] , 
        \wRegOut_7_67[12] , \wRegOut_7_67[11] , \wRegOut_7_67[10] , 
        \wRegOut_7_67[9] , \wRegOut_7_67[8] , \wRegOut_7_67[7] , 
        \wRegOut_7_67[6] , \wRegOut_7_67[5] , \wRegOut_7_67[4] , 
        \wRegOut_7_67[3] , \wRegOut_7_67[2] , \wRegOut_7_67[1] , 
        \wRegOut_7_67[0] }), .Enable1(\wRegEnTop_7_67[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_67[31] , \wRegInTop_7_67[30] , \wRegInTop_7_67[29] , 
        \wRegInTop_7_67[28] , \wRegInTop_7_67[27] , \wRegInTop_7_67[26] , 
        \wRegInTop_7_67[25] , \wRegInTop_7_67[24] , \wRegInTop_7_67[23] , 
        \wRegInTop_7_67[22] , \wRegInTop_7_67[21] , \wRegInTop_7_67[20] , 
        \wRegInTop_7_67[19] , \wRegInTop_7_67[18] , \wRegInTop_7_67[17] , 
        \wRegInTop_7_67[16] , \wRegInTop_7_67[15] , \wRegInTop_7_67[14] , 
        \wRegInTop_7_67[13] , \wRegInTop_7_67[12] , \wRegInTop_7_67[11] , 
        \wRegInTop_7_67[10] , \wRegInTop_7_67[9] , \wRegInTop_7_67[8] , 
        \wRegInTop_7_67[7] , \wRegInTop_7_67[6] , \wRegInTop_7_67[5] , 
        \wRegInTop_7_67[4] , \wRegInTop_7_67[3] , \wRegInTop_7_67[2] , 
        \wRegInTop_7_67[1] , \wRegInTop_7_67[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink70[31] , \ScanLink70[30] , \ScanLink70[29] , 
        \ScanLink70[28] , \ScanLink70[27] , \ScanLink70[26] , \ScanLink70[25] , 
        \ScanLink70[24] , \ScanLink70[23] , \ScanLink70[22] , \ScanLink70[21] , 
        \ScanLink70[20] , \ScanLink70[19] , \ScanLink70[18] , \ScanLink70[17] , 
        \ScanLink70[16] , \ScanLink70[15] , \ScanLink70[14] , \ScanLink70[13] , 
        \ScanLink70[12] , \ScanLink70[11] , \ScanLink70[10] , \ScanLink70[9] , 
        \ScanLink70[8] , \ScanLink70[7] , \ScanLink70[6] , \ScanLink70[5] , 
        \ScanLink70[4] , \ScanLink70[3] , \ScanLink70[2] , \ScanLink70[1] , 
        \ScanLink70[0] }), .ScanOut({\ScanLink69[31] , \ScanLink69[30] , 
        \ScanLink69[29] , \ScanLink69[28] , \ScanLink69[27] , \ScanLink69[26] , 
        \ScanLink69[25] , \ScanLink69[24] , \ScanLink69[23] , \ScanLink69[22] , 
        \ScanLink69[21] , \ScanLink69[20] , \ScanLink69[19] , \ScanLink69[18] , 
        \ScanLink69[17] , \ScanLink69[16] , \ScanLink69[15] , \ScanLink69[14] , 
        \ScanLink69[13] , \ScanLink69[12] , \ScanLink69[11] , \ScanLink69[10] , 
        \ScanLink69[9] , \ScanLink69[8] , \ScanLink69[7] , \ScanLink69[6] , 
        \ScanLink69[5] , \ScanLink69[4] , \ScanLink69[3] , \ScanLink69[2] , 
        \ScanLink69[1] , \ScanLink69[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_6[31] , \wRegOut_6_6[30] , \wRegOut_6_6[29] , 
        \wRegOut_6_6[28] , \wRegOut_6_6[27] , \wRegOut_6_6[26] , 
        \wRegOut_6_6[25] , \wRegOut_6_6[24] , \wRegOut_6_6[23] , 
        \wRegOut_6_6[22] , \wRegOut_6_6[21] , \wRegOut_6_6[20] , 
        \wRegOut_6_6[19] , \wRegOut_6_6[18] , \wRegOut_6_6[17] , 
        \wRegOut_6_6[16] , \wRegOut_6_6[15] , \wRegOut_6_6[14] , 
        \wRegOut_6_6[13] , \wRegOut_6_6[12] , \wRegOut_6_6[11] , 
        \wRegOut_6_6[10] , \wRegOut_6_6[9] , \wRegOut_6_6[8] , 
        \wRegOut_6_6[7] , \wRegOut_6_6[6] , \wRegOut_6_6[5] , \wRegOut_6_6[4] , 
        \wRegOut_6_6[3] , \wRegOut_6_6[2] , \wRegOut_6_6[1] , \wRegOut_6_6[0] 
        }), .Enable1(\wRegEnTop_6_6[0] ), .Enable2(\wRegEnBot_6_6[0] ), .In1({
        \wRegInTop_6_6[31] , \wRegInTop_6_6[30] , \wRegInTop_6_6[29] , 
        \wRegInTop_6_6[28] , \wRegInTop_6_6[27] , \wRegInTop_6_6[26] , 
        \wRegInTop_6_6[25] , \wRegInTop_6_6[24] , \wRegInTop_6_6[23] , 
        \wRegInTop_6_6[22] , \wRegInTop_6_6[21] , \wRegInTop_6_6[20] , 
        \wRegInTop_6_6[19] , \wRegInTop_6_6[18] , \wRegInTop_6_6[17] , 
        \wRegInTop_6_6[16] , \wRegInTop_6_6[15] , \wRegInTop_6_6[14] , 
        \wRegInTop_6_6[13] , \wRegInTop_6_6[12] , \wRegInTop_6_6[11] , 
        \wRegInTop_6_6[10] , \wRegInTop_6_6[9] , \wRegInTop_6_6[8] , 
        \wRegInTop_6_6[7] , \wRegInTop_6_6[6] , \wRegInTop_6_6[5] , 
        \wRegInTop_6_6[4] , \wRegInTop_6_6[3] , \wRegInTop_6_6[2] , 
        \wRegInTop_6_6[1] , \wRegInTop_6_6[0] }), .In2({\wRegInBot_6_6[31] , 
        \wRegInBot_6_6[30] , \wRegInBot_6_6[29] , \wRegInBot_6_6[28] , 
        \wRegInBot_6_6[27] , \wRegInBot_6_6[26] , \wRegInBot_6_6[25] , 
        \wRegInBot_6_6[24] , \wRegInBot_6_6[23] , \wRegInBot_6_6[22] , 
        \wRegInBot_6_6[21] , \wRegInBot_6_6[20] , \wRegInBot_6_6[19] , 
        \wRegInBot_6_6[18] , \wRegInBot_6_6[17] , \wRegInBot_6_6[16] , 
        \wRegInBot_6_6[15] , \wRegInBot_6_6[14] , \wRegInBot_6_6[13] , 
        \wRegInBot_6_6[12] , \wRegInBot_6_6[11] , \wRegInBot_6_6[10] , 
        \wRegInBot_6_6[9] , \wRegInBot_6_6[8] , \wRegInBot_6_6[7] , 
        \wRegInBot_6_6[6] , \wRegInBot_6_6[5] , \wRegInBot_6_6[4] , 
        \wRegInBot_6_6[3] , \wRegInBot_6_6[2] , \wRegInBot_6_6[1] , 
        \wRegInBot_6_6[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_34 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink98[31] , \ScanLink98[30] , \ScanLink98[29] , 
        \ScanLink98[28] , \ScanLink98[27] , \ScanLink98[26] , \ScanLink98[25] , 
        \ScanLink98[24] , \ScanLink98[23] , \ScanLink98[22] , \ScanLink98[21] , 
        \ScanLink98[20] , \ScanLink98[19] , \ScanLink98[18] , \ScanLink98[17] , 
        \ScanLink98[16] , \ScanLink98[15] , \ScanLink98[14] , \ScanLink98[13] , 
        \ScanLink98[12] , \ScanLink98[11] , \ScanLink98[10] , \ScanLink98[9] , 
        \ScanLink98[8] , \ScanLink98[7] , \ScanLink98[6] , \ScanLink98[5] , 
        \ScanLink98[4] , \ScanLink98[3] , \ScanLink98[2] , \ScanLink98[1] , 
        \ScanLink98[0] }), .ScanOut({\ScanLink97[31] , \ScanLink97[30] , 
        \ScanLink97[29] , \ScanLink97[28] , \ScanLink97[27] , \ScanLink97[26] , 
        \ScanLink97[25] , \ScanLink97[24] , \ScanLink97[23] , \ScanLink97[22] , 
        \ScanLink97[21] , \ScanLink97[20] , \ScanLink97[19] , \ScanLink97[18] , 
        \ScanLink97[17] , \ScanLink97[16] , \ScanLink97[15] , \ScanLink97[14] , 
        \ScanLink97[13] , \ScanLink97[12] , \ScanLink97[11] , \ScanLink97[10] , 
        \ScanLink97[9] , \ScanLink97[8] , \ScanLink97[7] , \ScanLink97[6] , 
        \ScanLink97[5] , \ScanLink97[4] , \ScanLink97[3] , \ScanLink97[2] , 
        \ScanLink97[1] , \ScanLink97[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_34[31] , \wRegOut_6_34[30] , 
        \wRegOut_6_34[29] , \wRegOut_6_34[28] , \wRegOut_6_34[27] , 
        \wRegOut_6_34[26] , \wRegOut_6_34[25] , \wRegOut_6_34[24] , 
        \wRegOut_6_34[23] , \wRegOut_6_34[22] , \wRegOut_6_34[21] , 
        \wRegOut_6_34[20] , \wRegOut_6_34[19] , \wRegOut_6_34[18] , 
        \wRegOut_6_34[17] , \wRegOut_6_34[16] , \wRegOut_6_34[15] , 
        \wRegOut_6_34[14] , \wRegOut_6_34[13] , \wRegOut_6_34[12] , 
        \wRegOut_6_34[11] , \wRegOut_6_34[10] , \wRegOut_6_34[9] , 
        \wRegOut_6_34[8] , \wRegOut_6_34[7] , \wRegOut_6_34[6] , 
        \wRegOut_6_34[5] , \wRegOut_6_34[4] , \wRegOut_6_34[3] , 
        \wRegOut_6_34[2] , \wRegOut_6_34[1] , \wRegOut_6_34[0] }), .Enable1(
        \wRegEnTop_6_34[0] ), .Enable2(\wRegEnBot_6_34[0] ), .In1({
        \wRegInTop_6_34[31] , \wRegInTop_6_34[30] , \wRegInTop_6_34[29] , 
        \wRegInTop_6_34[28] , \wRegInTop_6_34[27] , \wRegInTop_6_34[26] , 
        \wRegInTop_6_34[25] , \wRegInTop_6_34[24] , \wRegInTop_6_34[23] , 
        \wRegInTop_6_34[22] , \wRegInTop_6_34[21] , \wRegInTop_6_34[20] , 
        \wRegInTop_6_34[19] , \wRegInTop_6_34[18] , \wRegInTop_6_34[17] , 
        \wRegInTop_6_34[16] , \wRegInTop_6_34[15] , \wRegInTop_6_34[14] , 
        \wRegInTop_6_34[13] , \wRegInTop_6_34[12] , \wRegInTop_6_34[11] , 
        \wRegInTop_6_34[10] , \wRegInTop_6_34[9] , \wRegInTop_6_34[8] , 
        \wRegInTop_6_34[7] , \wRegInTop_6_34[6] , \wRegInTop_6_34[5] , 
        \wRegInTop_6_34[4] , \wRegInTop_6_34[3] , \wRegInTop_6_34[2] , 
        \wRegInTop_6_34[1] , \wRegInTop_6_34[0] }), .In2({\wRegInBot_6_34[31] , 
        \wRegInBot_6_34[30] , \wRegInBot_6_34[29] , \wRegInBot_6_34[28] , 
        \wRegInBot_6_34[27] , \wRegInBot_6_34[26] , \wRegInBot_6_34[25] , 
        \wRegInBot_6_34[24] , \wRegInBot_6_34[23] , \wRegInBot_6_34[22] , 
        \wRegInBot_6_34[21] , \wRegInBot_6_34[20] , \wRegInBot_6_34[19] , 
        \wRegInBot_6_34[18] , \wRegInBot_6_34[17] , \wRegInBot_6_34[16] , 
        \wRegInBot_6_34[15] , \wRegInBot_6_34[14] , \wRegInBot_6_34[13] , 
        \wRegInBot_6_34[12] , \wRegInBot_6_34[11] , \wRegInBot_6_34[10] , 
        \wRegInBot_6_34[9] , \wRegInBot_6_34[8] , \wRegInBot_6_34[7] , 
        \wRegInBot_6_34[6] , \wRegInBot_6_34[5] , \wRegInBot_6_34[4] , 
        \wRegInBot_6_34[3] , \wRegInBot_6_34[2] , \wRegInBot_6_34[1] , 
        \wRegInBot_6_34[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_41 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink105[31] , \ScanLink105[30] , \ScanLink105[29] , 
        \ScanLink105[28] , \ScanLink105[27] , \ScanLink105[26] , 
        \ScanLink105[25] , \ScanLink105[24] , \ScanLink105[23] , 
        \ScanLink105[22] , \ScanLink105[21] , \ScanLink105[20] , 
        \ScanLink105[19] , \ScanLink105[18] , \ScanLink105[17] , 
        \ScanLink105[16] , \ScanLink105[15] , \ScanLink105[14] , 
        \ScanLink105[13] , \ScanLink105[12] , \ScanLink105[11] , 
        \ScanLink105[10] , \ScanLink105[9] , \ScanLink105[8] , 
        \ScanLink105[7] , \ScanLink105[6] , \ScanLink105[5] , \ScanLink105[4] , 
        \ScanLink105[3] , \ScanLink105[2] , \ScanLink105[1] , \ScanLink105[0] 
        }), .ScanOut({\ScanLink104[31] , \ScanLink104[30] , \ScanLink104[29] , 
        \ScanLink104[28] , \ScanLink104[27] , \ScanLink104[26] , 
        \ScanLink104[25] , \ScanLink104[24] , \ScanLink104[23] , 
        \ScanLink104[22] , \ScanLink104[21] , \ScanLink104[20] , 
        \ScanLink104[19] , \ScanLink104[18] , \ScanLink104[17] , 
        \ScanLink104[16] , \ScanLink104[15] , \ScanLink104[14] , 
        \ScanLink104[13] , \ScanLink104[12] , \ScanLink104[11] , 
        \ScanLink104[10] , \ScanLink104[9] , \ScanLink104[8] , 
        \ScanLink104[7] , \ScanLink104[6] , \ScanLink104[5] , \ScanLink104[4] , 
        \ScanLink104[3] , \ScanLink104[2] , \ScanLink104[1] , \ScanLink104[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_41[31] , 
        \wRegOut_6_41[30] , \wRegOut_6_41[29] , \wRegOut_6_41[28] , 
        \wRegOut_6_41[27] , \wRegOut_6_41[26] , \wRegOut_6_41[25] , 
        \wRegOut_6_41[24] , \wRegOut_6_41[23] , \wRegOut_6_41[22] , 
        \wRegOut_6_41[21] , \wRegOut_6_41[20] , \wRegOut_6_41[19] , 
        \wRegOut_6_41[18] , \wRegOut_6_41[17] , \wRegOut_6_41[16] , 
        \wRegOut_6_41[15] , \wRegOut_6_41[14] , \wRegOut_6_41[13] , 
        \wRegOut_6_41[12] , \wRegOut_6_41[11] , \wRegOut_6_41[10] , 
        \wRegOut_6_41[9] , \wRegOut_6_41[8] , \wRegOut_6_41[7] , 
        \wRegOut_6_41[6] , \wRegOut_6_41[5] , \wRegOut_6_41[4] , 
        \wRegOut_6_41[3] , \wRegOut_6_41[2] , \wRegOut_6_41[1] , 
        \wRegOut_6_41[0] }), .Enable1(\wRegEnTop_6_41[0] ), .Enable2(
        \wRegEnBot_6_41[0] ), .In1({\wRegInTop_6_41[31] , \wRegInTop_6_41[30] , 
        \wRegInTop_6_41[29] , \wRegInTop_6_41[28] , \wRegInTop_6_41[27] , 
        \wRegInTop_6_41[26] , \wRegInTop_6_41[25] , \wRegInTop_6_41[24] , 
        \wRegInTop_6_41[23] , \wRegInTop_6_41[22] , \wRegInTop_6_41[21] , 
        \wRegInTop_6_41[20] , \wRegInTop_6_41[19] , \wRegInTop_6_41[18] , 
        \wRegInTop_6_41[17] , \wRegInTop_6_41[16] , \wRegInTop_6_41[15] , 
        \wRegInTop_6_41[14] , \wRegInTop_6_41[13] , \wRegInTop_6_41[12] , 
        \wRegInTop_6_41[11] , \wRegInTop_6_41[10] , \wRegInTop_6_41[9] , 
        \wRegInTop_6_41[8] , \wRegInTop_6_41[7] , \wRegInTop_6_41[6] , 
        \wRegInTop_6_41[5] , \wRegInTop_6_41[4] , \wRegInTop_6_41[3] , 
        \wRegInTop_6_41[2] , \wRegInTop_6_41[1] , \wRegInTop_6_41[0] }), .In2(
        {\wRegInBot_6_41[31] , \wRegInBot_6_41[30] , \wRegInBot_6_41[29] , 
        \wRegInBot_6_41[28] , \wRegInBot_6_41[27] , \wRegInBot_6_41[26] , 
        \wRegInBot_6_41[25] , \wRegInBot_6_41[24] , \wRegInBot_6_41[23] , 
        \wRegInBot_6_41[22] , \wRegInBot_6_41[21] , \wRegInBot_6_41[20] , 
        \wRegInBot_6_41[19] , \wRegInBot_6_41[18] , \wRegInBot_6_41[17] , 
        \wRegInBot_6_41[16] , \wRegInBot_6_41[15] , \wRegInBot_6_41[14] , 
        \wRegInBot_6_41[13] , \wRegInBot_6_41[12] , \wRegInBot_6_41[11] , 
        \wRegInBot_6_41[10] , \wRegInBot_6_41[9] , \wRegInBot_6_41[8] , 
        \wRegInBot_6_41[7] , \wRegInBot_6_41[6] , \wRegInBot_6_41[5] , 
        \wRegInBot_6_41[4] , \wRegInBot_6_41[3] , \wRegInBot_6_41[2] , 
        \wRegInBot_6_41[1] , \wRegInBot_6_41[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink134[31] , \ScanLink134[30] , \ScanLink134[29] , 
        \ScanLink134[28] , \ScanLink134[27] , \ScanLink134[26] , 
        \ScanLink134[25] , \ScanLink134[24] , \ScanLink134[23] , 
        \ScanLink134[22] , \ScanLink134[21] , \ScanLink134[20] , 
        \ScanLink134[19] , \ScanLink134[18] , \ScanLink134[17] , 
        \ScanLink134[16] , \ScanLink134[15] , \ScanLink134[14] , 
        \ScanLink134[13] , \ScanLink134[12] , \ScanLink134[11] , 
        \ScanLink134[10] , \ScanLink134[9] , \ScanLink134[8] , 
        \ScanLink134[7] , \ScanLink134[6] , \ScanLink134[5] , \ScanLink134[4] , 
        \ScanLink134[3] , \ScanLink134[2] , \ScanLink134[1] , \ScanLink134[0] 
        }), .ScanOut({\ScanLink133[31] , \ScanLink133[30] , \ScanLink133[29] , 
        \ScanLink133[28] , \ScanLink133[27] , \ScanLink133[26] , 
        \ScanLink133[25] , \ScanLink133[24] , \ScanLink133[23] , 
        \ScanLink133[22] , \ScanLink133[21] , \ScanLink133[20] , 
        \ScanLink133[19] , \ScanLink133[18] , \ScanLink133[17] , 
        \ScanLink133[16] , \ScanLink133[15] , \ScanLink133[14] , 
        \ScanLink133[13] , \ScanLink133[12] , \ScanLink133[11] , 
        \ScanLink133[10] , \ScanLink133[9] , \ScanLink133[8] , 
        \ScanLink133[7] , \ScanLink133[6] , \ScanLink133[5] , \ScanLink133[4] , 
        \ScanLink133[3] , \ScanLink133[2] , \ScanLink133[1] , \ScanLink133[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_6[31] , 
        \wRegOut_7_6[30] , \wRegOut_7_6[29] , \wRegOut_7_6[28] , 
        \wRegOut_7_6[27] , \wRegOut_7_6[26] , \wRegOut_7_6[25] , 
        \wRegOut_7_6[24] , \wRegOut_7_6[23] , \wRegOut_7_6[22] , 
        \wRegOut_7_6[21] , \wRegOut_7_6[20] , \wRegOut_7_6[19] , 
        \wRegOut_7_6[18] , \wRegOut_7_6[17] , \wRegOut_7_6[16] , 
        \wRegOut_7_6[15] , \wRegOut_7_6[14] , \wRegOut_7_6[13] , 
        \wRegOut_7_6[12] , \wRegOut_7_6[11] , \wRegOut_7_6[10] , 
        \wRegOut_7_6[9] , \wRegOut_7_6[8] , \wRegOut_7_6[7] , \wRegOut_7_6[6] , 
        \wRegOut_7_6[5] , \wRegOut_7_6[4] , \wRegOut_7_6[3] , \wRegOut_7_6[2] , 
        \wRegOut_7_6[1] , \wRegOut_7_6[0] }), .Enable1(\wRegEnTop_7_6[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_6[31] , \wRegInTop_7_6[30] , 
        \wRegInTop_7_6[29] , \wRegInTop_7_6[28] , \wRegInTop_7_6[27] , 
        \wRegInTop_7_6[26] , \wRegInTop_7_6[25] , \wRegInTop_7_6[24] , 
        \wRegInTop_7_6[23] , \wRegInTop_7_6[22] , \wRegInTop_7_6[21] , 
        \wRegInTop_7_6[20] , \wRegInTop_7_6[19] , \wRegInTop_7_6[18] , 
        \wRegInTop_7_6[17] , \wRegInTop_7_6[16] , \wRegInTop_7_6[15] , 
        \wRegInTop_7_6[14] , \wRegInTop_7_6[13] , \wRegInTop_7_6[12] , 
        \wRegInTop_7_6[11] , \wRegInTop_7_6[10] , \wRegInTop_7_6[9] , 
        \wRegInTop_7_6[8] , \wRegInTop_7_6[7] , \wRegInTop_7_6[6] , 
        \wRegInTop_7_6[5] , \wRegInTop_7_6[4] , \wRegInTop_7_6[3] , 
        \wRegInTop_7_6[2] , \wRegInTop_7_6[1] , \wRegInTop_7_6[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_40 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink168[31] , \ScanLink168[30] , \ScanLink168[29] , 
        \ScanLink168[28] , \ScanLink168[27] , \ScanLink168[26] , 
        \ScanLink168[25] , \ScanLink168[24] , \ScanLink168[23] , 
        \ScanLink168[22] , \ScanLink168[21] , \ScanLink168[20] , 
        \ScanLink168[19] , \ScanLink168[18] , \ScanLink168[17] , 
        \ScanLink168[16] , \ScanLink168[15] , \ScanLink168[14] , 
        \ScanLink168[13] , \ScanLink168[12] , \ScanLink168[11] , 
        \ScanLink168[10] , \ScanLink168[9] , \ScanLink168[8] , 
        \ScanLink168[7] , \ScanLink168[6] , \ScanLink168[5] , \ScanLink168[4] , 
        \ScanLink168[3] , \ScanLink168[2] , \ScanLink168[1] , \ScanLink168[0] 
        }), .ScanOut({\ScanLink167[31] , \ScanLink167[30] , \ScanLink167[29] , 
        \ScanLink167[28] , \ScanLink167[27] , \ScanLink167[26] , 
        \ScanLink167[25] , \ScanLink167[24] , \ScanLink167[23] , 
        \ScanLink167[22] , \ScanLink167[21] , \ScanLink167[20] , 
        \ScanLink167[19] , \ScanLink167[18] , \ScanLink167[17] , 
        \ScanLink167[16] , \ScanLink167[15] , \ScanLink167[14] , 
        \ScanLink167[13] , \ScanLink167[12] , \ScanLink167[11] , 
        \ScanLink167[10] , \ScanLink167[9] , \ScanLink167[8] , 
        \ScanLink167[7] , \ScanLink167[6] , \ScanLink167[5] , \ScanLink167[4] , 
        \ScanLink167[3] , \ScanLink167[2] , \ScanLink167[1] , \ScanLink167[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_40[31] , 
        \wRegOut_7_40[30] , \wRegOut_7_40[29] , \wRegOut_7_40[28] , 
        \wRegOut_7_40[27] , \wRegOut_7_40[26] , \wRegOut_7_40[25] , 
        \wRegOut_7_40[24] , \wRegOut_7_40[23] , \wRegOut_7_40[22] , 
        \wRegOut_7_40[21] , \wRegOut_7_40[20] , \wRegOut_7_40[19] , 
        \wRegOut_7_40[18] , \wRegOut_7_40[17] , \wRegOut_7_40[16] , 
        \wRegOut_7_40[15] , \wRegOut_7_40[14] , \wRegOut_7_40[13] , 
        \wRegOut_7_40[12] , \wRegOut_7_40[11] , \wRegOut_7_40[10] , 
        \wRegOut_7_40[9] , \wRegOut_7_40[8] , \wRegOut_7_40[7] , 
        \wRegOut_7_40[6] , \wRegOut_7_40[5] , \wRegOut_7_40[4] , 
        \wRegOut_7_40[3] , \wRegOut_7_40[2] , \wRegOut_7_40[1] , 
        \wRegOut_7_40[0] }), .Enable1(\wRegEnTop_7_40[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_40[31] , \wRegInTop_7_40[30] , \wRegInTop_7_40[29] , 
        \wRegInTop_7_40[28] , \wRegInTop_7_40[27] , \wRegInTop_7_40[26] , 
        \wRegInTop_7_40[25] , \wRegInTop_7_40[24] , \wRegInTop_7_40[23] , 
        \wRegInTop_7_40[22] , \wRegInTop_7_40[21] , \wRegInTop_7_40[20] , 
        \wRegInTop_7_40[19] , \wRegInTop_7_40[18] , \wRegInTop_7_40[17] , 
        \wRegInTop_7_40[16] , \wRegInTop_7_40[15] , \wRegInTop_7_40[14] , 
        \wRegInTop_7_40[13] , \wRegInTop_7_40[12] , \wRegInTop_7_40[11] , 
        \wRegInTop_7_40[10] , \wRegInTop_7_40[9] , \wRegInTop_7_40[8] , 
        \wRegInTop_7_40[7] , \wRegInTop_7_40[6] , \wRegInTop_7_40[5] , 
        \wRegInTop_7_40[4] , \wRegInTop_7_40[3] , \wRegInTop_7_40[2] , 
        \wRegInTop_7_40[1] , \wRegInTop_7_40[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink140[31] , \ScanLink140[30] , \ScanLink140[29] , 
        \ScanLink140[28] , \ScanLink140[27] , \ScanLink140[26] , 
        \ScanLink140[25] , \ScanLink140[24] , \ScanLink140[23] , 
        \ScanLink140[22] , \ScanLink140[21] , \ScanLink140[20] , 
        \ScanLink140[19] , \ScanLink140[18] , \ScanLink140[17] , 
        \ScanLink140[16] , \ScanLink140[15] , \ScanLink140[14] , 
        \ScanLink140[13] , \ScanLink140[12] , \ScanLink140[11] , 
        \ScanLink140[10] , \ScanLink140[9] , \ScanLink140[8] , 
        \ScanLink140[7] , \ScanLink140[6] , \ScanLink140[5] , \ScanLink140[4] , 
        \ScanLink140[3] , \ScanLink140[2] , \ScanLink140[1] , \ScanLink140[0] 
        }), .ScanOut({\ScanLink139[31] , \ScanLink139[30] , \ScanLink139[29] , 
        \ScanLink139[28] , \ScanLink139[27] , \ScanLink139[26] , 
        \ScanLink139[25] , \ScanLink139[24] , \ScanLink139[23] , 
        \ScanLink139[22] , \ScanLink139[21] , \ScanLink139[20] , 
        \ScanLink139[19] , \ScanLink139[18] , \ScanLink139[17] , 
        \ScanLink139[16] , \ScanLink139[15] , \ScanLink139[14] , 
        \ScanLink139[13] , \ScanLink139[12] , \ScanLink139[11] , 
        \ScanLink139[10] , \ScanLink139[9] , \ScanLink139[8] , 
        \ScanLink139[7] , \ScanLink139[6] , \ScanLink139[5] , \ScanLink139[4] , 
        \ScanLink139[3] , \ScanLink139[2] , \ScanLink139[1] , \ScanLink139[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_12[31] , 
        \wRegOut_7_12[30] , \wRegOut_7_12[29] , \wRegOut_7_12[28] , 
        \wRegOut_7_12[27] , \wRegOut_7_12[26] , \wRegOut_7_12[25] , 
        \wRegOut_7_12[24] , \wRegOut_7_12[23] , \wRegOut_7_12[22] , 
        \wRegOut_7_12[21] , \wRegOut_7_12[20] , \wRegOut_7_12[19] , 
        \wRegOut_7_12[18] , \wRegOut_7_12[17] , \wRegOut_7_12[16] , 
        \wRegOut_7_12[15] , \wRegOut_7_12[14] , \wRegOut_7_12[13] , 
        \wRegOut_7_12[12] , \wRegOut_7_12[11] , \wRegOut_7_12[10] , 
        \wRegOut_7_12[9] , \wRegOut_7_12[8] , \wRegOut_7_12[7] , 
        \wRegOut_7_12[6] , \wRegOut_7_12[5] , \wRegOut_7_12[4] , 
        \wRegOut_7_12[3] , \wRegOut_7_12[2] , \wRegOut_7_12[1] , 
        \wRegOut_7_12[0] }), .Enable1(\wRegEnTop_7_12[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_12[31] , \wRegInTop_7_12[30] , \wRegInTop_7_12[29] , 
        \wRegInTop_7_12[28] , \wRegInTop_7_12[27] , \wRegInTop_7_12[26] , 
        \wRegInTop_7_12[25] , \wRegInTop_7_12[24] , \wRegInTop_7_12[23] , 
        \wRegInTop_7_12[22] , \wRegInTop_7_12[21] , \wRegInTop_7_12[20] , 
        \wRegInTop_7_12[19] , \wRegInTop_7_12[18] , \wRegInTop_7_12[17] , 
        \wRegInTop_7_12[16] , \wRegInTop_7_12[15] , \wRegInTop_7_12[14] , 
        \wRegInTop_7_12[13] , \wRegInTop_7_12[12] , \wRegInTop_7_12[11] , 
        \wRegInTop_7_12[10] , \wRegInTop_7_12[9] , \wRegInTop_7_12[8] , 
        \wRegInTop_7_12[7] , \wRegInTop_7_12[6] , \wRegInTop_7_12[5] , 
        \wRegInTop_7_12[4] , \wRegInTop_7_12[3] , \wRegInTop_7_12[2] , 
        \wRegInTop_7_12[1] , \wRegInTop_7_12[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_82 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink210[31] , \ScanLink210[30] , \ScanLink210[29] , 
        \ScanLink210[28] , \ScanLink210[27] , \ScanLink210[26] , 
        \ScanLink210[25] , \ScanLink210[24] , \ScanLink210[23] , 
        \ScanLink210[22] , \ScanLink210[21] , \ScanLink210[20] , 
        \ScanLink210[19] , \ScanLink210[18] , \ScanLink210[17] , 
        \ScanLink210[16] , \ScanLink210[15] , \ScanLink210[14] , 
        \ScanLink210[13] , \ScanLink210[12] , \ScanLink210[11] , 
        \ScanLink210[10] , \ScanLink210[9] , \ScanLink210[8] , 
        \ScanLink210[7] , \ScanLink210[6] , \ScanLink210[5] , \ScanLink210[4] , 
        \ScanLink210[3] , \ScanLink210[2] , \ScanLink210[1] , \ScanLink210[0] 
        }), .ScanOut({\ScanLink209[31] , \ScanLink209[30] , \ScanLink209[29] , 
        \ScanLink209[28] , \ScanLink209[27] , \ScanLink209[26] , 
        \ScanLink209[25] , \ScanLink209[24] , \ScanLink209[23] , 
        \ScanLink209[22] , \ScanLink209[21] , \ScanLink209[20] , 
        \ScanLink209[19] , \ScanLink209[18] , \ScanLink209[17] , 
        \ScanLink209[16] , \ScanLink209[15] , \ScanLink209[14] , 
        \ScanLink209[13] , \ScanLink209[12] , \ScanLink209[11] , 
        \ScanLink209[10] , \ScanLink209[9] , \ScanLink209[8] , 
        \ScanLink209[7] , \ScanLink209[6] , \ScanLink209[5] , \ScanLink209[4] , 
        \ScanLink209[3] , \ScanLink209[2] , \ScanLink209[1] , \ScanLink209[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_82[31] , 
        \wRegOut_7_82[30] , \wRegOut_7_82[29] , \wRegOut_7_82[28] , 
        \wRegOut_7_82[27] , \wRegOut_7_82[26] , \wRegOut_7_82[25] , 
        \wRegOut_7_82[24] , \wRegOut_7_82[23] , \wRegOut_7_82[22] , 
        \wRegOut_7_82[21] , \wRegOut_7_82[20] , \wRegOut_7_82[19] , 
        \wRegOut_7_82[18] , \wRegOut_7_82[17] , \wRegOut_7_82[16] , 
        \wRegOut_7_82[15] , \wRegOut_7_82[14] , \wRegOut_7_82[13] , 
        \wRegOut_7_82[12] , \wRegOut_7_82[11] , \wRegOut_7_82[10] , 
        \wRegOut_7_82[9] , \wRegOut_7_82[8] , \wRegOut_7_82[7] , 
        \wRegOut_7_82[6] , \wRegOut_7_82[5] , \wRegOut_7_82[4] , 
        \wRegOut_7_82[3] , \wRegOut_7_82[2] , \wRegOut_7_82[1] , 
        \wRegOut_7_82[0] }), .Enable1(\wRegEnTop_7_82[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_82[31] , \wRegInTop_7_82[30] , \wRegInTop_7_82[29] , 
        \wRegInTop_7_82[28] , \wRegInTop_7_82[27] , \wRegInTop_7_82[26] , 
        \wRegInTop_7_82[25] , \wRegInTop_7_82[24] , \wRegInTop_7_82[23] , 
        \wRegInTop_7_82[22] , \wRegInTop_7_82[21] , \wRegInTop_7_82[20] , 
        \wRegInTop_7_82[19] , \wRegInTop_7_82[18] , \wRegInTop_7_82[17] , 
        \wRegInTop_7_82[16] , \wRegInTop_7_82[15] , \wRegInTop_7_82[14] , 
        \wRegInTop_7_82[13] , \wRegInTop_7_82[12] , \wRegInTop_7_82[11] , 
        \wRegInTop_7_82[10] , \wRegInTop_7_82[9] , \wRegInTop_7_82[8] , 
        \wRegInTop_7_82[7] , \wRegInTop_7_82[6] , \wRegInTop_7_82[5] , 
        \wRegInTop_7_82[4] , \wRegInTop_7_82[3] , \wRegInTop_7_82[2] , 
        \wRegInTop_7_82[1] , \wRegInTop_7_82[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_2[0] ), .P_In({\wRegOut_3_2[31] , 
        \wRegOut_3_2[30] , \wRegOut_3_2[29] , \wRegOut_3_2[28] , 
        \wRegOut_3_2[27] , \wRegOut_3_2[26] , \wRegOut_3_2[25] , 
        \wRegOut_3_2[24] , \wRegOut_3_2[23] , \wRegOut_3_2[22] , 
        \wRegOut_3_2[21] , \wRegOut_3_2[20] , \wRegOut_3_2[19] , 
        \wRegOut_3_2[18] , \wRegOut_3_2[17] , \wRegOut_3_2[16] , 
        \wRegOut_3_2[15] , \wRegOut_3_2[14] , \wRegOut_3_2[13] , 
        \wRegOut_3_2[12] , \wRegOut_3_2[11] , \wRegOut_3_2[10] , 
        \wRegOut_3_2[9] , \wRegOut_3_2[8] , \wRegOut_3_2[7] , \wRegOut_3_2[6] , 
        \wRegOut_3_2[5] , \wRegOut_3_2[4] , \wRegOut_3_2[3] , \wRegOut_3_2[2] , 
        \wRegOut_3_2[1] , \wRegOut_3_2[0] }), .P_Out({\wRegInBot_3_2[31] , 
        \wRegInBot_3_2[30] , \wRegInBot_3_2[29] , \wRegInBot_3_2[28] , 
        \wRegInBot_3_2[27] , \wRegInBot_3_2[26] , \wRegInBot_3_2[25] , 
        \wRegInBot_3_2[24] , \wRegInBot_3_2[23] , \wRegInBot_3_2[22] , 
        \wRegInBot_3_2[21] , \wRegInBot_3_2[20] , \wRegInBot_3_2[19] , 
        \wRegInBot_3_2[18] , \wRegInBot_3_2[17] , \wRegInBot_3_2[16] , 
        \wRegInBot_3_2[15] , \wRegInBot_3_2[14] , \wRegInBot_3_2[13] , 
        \wRegInBot_3_2[12] , \wRegInBot_3_2[11] , \wRegInBot_3_2[10] , 
        \wRegInBot_3_2[9] , \wRegInBot_3_2[8] , \wRegInBot_3_2[7] , 
        \wRegInBot_3_2[6] , \wRegInBot_3_2[5] , \wRegInBot_3_2[4] , 
        \wRegInBot_3_2[3] , \wRegInBot_3_2[2] , \wRegInBot_3_2[1] , 
        \wRegInBot_3_2[0] }), .L_WR(\wRegEnTop_4_4[0] ), .L_In({
        \wRegOut_4_4[31] , \wRegOut_4_4[30] , \wRegOut_4_4[29] , 
        \wRegOut_4_4[28] , \wRegOut_4_4[27] , \wRegOut_4_4[26] , 
        \wRegOut_4_4[25] , \wRegOut_4_4[24] , \wRegOut_4_4[23] , 
        \wRegOut_4_4[22] , \wRegOut_4_4[21] , \wRegOut_4_4[20] , 
        \wRegOut_4_4[19] , \wRegOut_4_4[18] , \wRegOut_4_4[17] , 
        \wRegOut_4_4[16] , \wRegOut_4_4[15] , \wRegOut_4_4[14] , 
        \wRegOut_4_4[13] , \wRegOut_4_4[12] , \wRegOut_4_4[11] , 
        \wRegOut_4_4[10] , \wRegOut_4_4[9] , \wRegOut_4_4[8] , 
        \wRegOut_4_4[7] , \wRegOut_4_4[6] , \wRegOut_4_4[5] , \wRegOut_4_4[4] , 
        \wRegOut_4_4[3] , \wRegOut_4_4[2] , \wRegOut_4_4[1] , \wRegOut_4_4[0] 
        }), .L_Out({\wRegInTop_4_4[31] , \wRegInTop_4_4[30] , 
        \wRegInTop_4_4[29] , \wRegInTop_4_4[28] , \wRegInTop_4_4[27] , 
        \wRegInTop_4_4[26] , \wRegInTop_4_4[25] , \wRegInTop_4_4[24] , 
        \wRegInTop_4_4[23] , \wRegInTop_4_4[22] , \wRegInTop_4_4[21] , 
        \wRegInTop_4_4[20] , \wRegInTop_4_4[19] , \wRegInTop_4_4[18] , 
        \wRegInTop_4_4[17] , \wRegInTop_4_4[16] , \wRegInTop_4_4[15] , 
        \wRegInTop_4_4[14] , \wRegInTop_4_4[13] , \wRegInTop_4_4[12] , 
        \wRegInTop_4_4[11] , \wRegInTop_4_4[10] , \wRegInTop_4_4[9] , 
        \wRegInTop_4_4[8] , \wRegInTop_4_4[7] , \wRegInTop_4_4[6] , 
        \wRegInTop_4_4[5] , \wRegInTop_4_4[4] , \wRegInTop_4_4[3] , 
        \wRegInTop_4_4[2] , \wRegInTop_4_4[1] , \wRegInTop_4_4[0] }), .R_WR(
        \wRegEnTop_4_5[0] ), .R_In({\wRegOut_4_5[31] , \wRegOut_4_5[30] , 
        \wRegOut_4_5[29] , \wRegOut_4_5[28] , \wRegOut_4_5[27] , 
        \wRegOut_4_5[26] , \wRegOut_4_5[25] , \wRegOut_4_5[24] , 
        \wRegOut_4_5[23] , \wRegOut_4_5[22] , \wRegOut_4_5[21] , 
        \wRegOut_4_5[20] , \wRegOut_4_5[19] , \wRegOut_4_5[18] , 
        \wRegOut_4_5[17] , \wRegOut_4_5[16] , \wRegOut_4_5[15] , 
        \wRegOut_4_5[14] , \wRegOut_4_5[13] , \wRegOut_4_5[12] , 
        \wRegOut_4_5[11] , \wRegOut_4_5[10] , \wRegOut_4_5[9] , 
        \wRegOut_4_5[8] , \wRegOut_4_5[7] , \wRegOut_4_5[6] , \wRegOut_4_5[5] , 
        \wRegOut_4_5[4] , \wRegOut_4_5[3] , \wRegOut_4_5[2] , \wRegOut_4_5[1] , 
        \wRegOut_4_5[0] }), .R_Out({\wRegInTop_4_5[31] , \wRegInTop_4_5[30] , 
        \wRegInTop_4_5[29] , \wRegInTop_4_5[28] , \wRegInTop_4_5[27] , 
        \wRegInTop_4_5[26] , \wRegInTop_4_5[25] , \wRegInTop_4_5[24] , 
        \wRegInTop_4_5[23] , \wRegInTop_4_5[22] , \wRegInTop_4_5[21] , 
        \wRegInTop_4_5[20] , \wRegInTop_4_5[19] , \wRegInTop_4_5[18] , 
        \wRegInTop_4_5[17] , \wRegInTop_4_5[16] , \wRegInTop_4_5[15] , 
        \wRegInTop_4_5[14] , \wRegInTop_4_5[13] , \wRegInTop_4_5[12] , 
        \wRegInTop_4_5[11] , \wRegInTop_4_5[10] , \wRegInTop_4_5[9] , 
        \wRegInTop_4_5[8] , \wRegInTop_4_5[7] , \wRegInTop_4_5[6] , 
        \wRegInTop_4_5[5] , \wRegInTop_4_5[4] , \wRegInTop_4_5[3] , 
        \wRegInTop_4_5[2] , \wRegInTop_4_5[1] , \wRegInTop_4_5[0] }) );
    BHeap_Node_WIDTH32 BHN_4_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_8[0] ), .P_In({\wRegOut_4_8[31] , 
        \wRegOut_4_8[30] , \wRegOut_4_8[29] , \wRegOut_4_8[28] , 
        \wRegOut_4_8[27] , \wRegOut_4_8[26] , \wRegOut_4_8[25] , 
        \wRegOut_4_8[24] , \wRegOut_4_8[23] , \wRegOut_4_8[22] , 
        \wRegOut_4_8[21] , \wRegOut_4_8[20] , \wRegOut_4_8[19] , 
        \wRegOut_4_8[18] , \wRegOut_4_8[17] , \wRegOut_4_8[16] , 
        \wRegOut_4_8[15] , \wRegOut_4_8[14] , \wRegOut_4_8[13] , 
        \wRegOut_4_8[12] , \wRegOut_4_8[11] , \wRegOut_4_8[10] , 
        \wRegOut_4_8[9] , \wRegOut_4_8[8] , \wRegOut_4_8[7] , \wRegOut_4_8[6] , 
        \wRegOut_4_8[5] , \wRegOut_4_8[4] , \wRegOut_4_8[3] , \wRegOut_4_8[2] , 
        \wRegOut_4_8[1] , \wRegOut_4_8[0] }), .P_Out({\wRegInBot_4_8[31] , 
        \wRegInBot_4_8[30] , \wRegInBot_4_8[29] , \wRegInBot_4_8[28] , 
        \wRegInBot_4_8[27] , \wRegInBot_4_8[26] , \wRegInBot_4_8[25] , 
        \wRegInBot_4_8[24] , \wRegInBot_4_8[23] , \wRegInBot_4_8[22] , 
        \wRegInBot_4_8[21] , \wRegInBot_4_8[20] , \wRegInBot_4_8[19] , 
        \wRegInBot_4_8[18] , \wRegInBot_4_8[17] , \wRegInBot_4_8[16] , 
        \wRegInBot_4_8[15] , \wRegInBot_4_8[14] , \wRegInBot_4_8[13] , 
        \wRegInBot_4_8[12] , \wRegInBot_4_8[11] , \wRegInBot_4_8[10] , 
        \wRegInBot_4_8[9] , \wRegInBot_4_8[8] , \wRegInBot_4_8[7] , 
        \wRegInBot_4_8[6] , \wRegInBot_4_8[5] , \wRegInBot_4_8[4] , 
        \wRegInBot_4_8[3] , \wRegInBot_4_8[2] , \wRegInBot_4_8[1] , 
        \wRegInBot_4_8[0] }), .L_WR(\wRegEnTop_5_16[0] ), .L_In({
        \wRegOut_5_16[31] , \wRegOut_5_16[30] , \wRegOut_5_16[29] , 
        \wRegOut_5_16[28] , \wRegOut_5_16[27] , \wRegOut_5_16[26] , 
        \wRegOut_5_16[25] , \wRegOut_5_16[24] , \wRegOut_5_16[23] , 
        \wRegOut_5_16[22] , \wRegOut_5_16[21] , \wRegOut_5_16[20] , 
        \wRegOut_5_16[19] , \wRegOut_5_16[18] , \wRegOut_5_16[17] , 
        \wRegOut_5_16[16] , \wRegOut_5_16[15] , \wRegOut_5_16[14] , 
        \wRegOut_5_16[13] , \wRegOut_5_16[12] , \wRegOut_5_16[11] , 
        \wRegOut_5_16[10] , \wRegOut_5_16[9] , \wRegOut_5_16[8] , 
        \wRegOut_5_16[7] , \wRegOut_5_16[6] , \wRegOut_5_16[5] , 
        \wRegOut_5_16[4] , \wRegOut_5_16[3] , \wRegOut_5_16[2] , 
        \wRegOut_5_16[1] , \wRegOut_5_16[0] }), .L_Out({\wRegInTop_5_16[31] , 
        \wRegInTop_5_16[30] , \wRegInTop_5_16[29] , \wRegInTop_5_16[28] , 
        \wRegInTop_5_16[27] , \wRegInTop_5_16[26] , \wRegInTop_5_16[25] , 
        \wRegInTop_5_16[24] , \wRegInTop_5_16[23] , \wRegInTop_5_16[22] , 
        \wRegInTop_5_16[21] , \wRegInTop_5_16[20] , \wRegInTop_5_16[19] , 
        \wRegInTop_5_16[18] , \wRegInTop_5_16[17] , \wRegInTop_5_16[16] , 
        \wRegInTop_5_16[15] , \wRegInTop_5_16[14] , \wRegInTop_5_16[13] , 
        \wRegInTop_5_16[12] , \wRegInTop_5_16[11] , \wRegInTop_5_16[10] , 
        \wRegInTop_5_16[9] , \wRegInTop_5_16[8] , \wRegInTop_5_16[7] , 
        \wRegInTop_5_16[6] , \wRegInTop_5_16[5] , \wRegInTop_5_16[4] , 
        \wRegInTop_5_16[3] , \wRegInTop_5_16[2] , \wRegInTop_5_16[1] , 
        \wRegInTop_5_16[0] }), .R_WR(\wRegEnTop_5_17[0] ), .R_In({
        \wRegOut_5_17[31] , \wRegOut_5_17[30] , \wRegOut_5_17[29] , 
        \wRegOut_5_17[28] , \wRegOut_5_17[27] , \wRegOut_5_17[26] , 
        \wRegOut_5_17[25] , \wRegOut_5_17[24] , \wRegOut_5_17[23] , 
        \wRegOut_5_17[22] , \wRegOut_5_17[21] , \wRegOut_5_17[20] , 
        \wRegOut_5_17[19] , \wRegOut_5_17[18] , \wRegOut_5_17[17] , 
        \wRegOut_5_17[16] , \wRegOut_5_17[15] , \wRegOut_5_17[14] , 
        \wRegOut_5_17[13] , \wRegOut_5_17[12] , \wRegOut_5_17[11] , 
        \wRegOut_5_17[10] , \wRegOut_5_17[9] , \wRegOut_5_17[8] , 
        \wRegOut_5_17[7] , \wRegOut_5_17[6] , \wRegOut_5_17[5] , 
        \wRegOut_5_17[4] , \wRegOut_5_17[3] , \wRegOut_5_17[2] , 
        \wRegOut_5_17[1] , \wRegOut_5_17[0] }), .R_Out({\wRegInTop_5_17[31] , 
        \wRegInTop_5_17[30] , \wRegInTop_5_17[29] , \wRegInTop_5_17[28] , 
        \wRegInTop_5_17[27] , \wRegInTop_5_17[26] , \wRegInTop_5_17[25] , 
        \wRegInTop_5_17[24] , \wRegInTop_5_17[23] , \wRegInTop_5_17[22] , 
        \wRegInTop_5_17[21] , \wRegInTop_5_17[20] , \wRegInTop_5_17[19] , 
        \wRegInTop_5_17[18] , \wRegInTop_5_17[17] , \wRegInTop_5_17[16] , 
        \wRegInTop_5_17[15] , \wRegInTop_5_17[14] , \wRegInTop_5_17[13] , 
        \wRegInTop_5_17[12] , \wRegInTop_5_17[11] , \wRegInTop_5_17[10] , 
        \wRegInTop_5_17[9] , \wRegInTop_5_17[8] , \wRegInTop_5_17[7] , 
        \wRegInTop_5_17[6] , \wRegInTop_5_17[5] , \wRegInTop_5_17[4] , 
        \wRegInTop_5_17[3] , \wRegInTop_5_17[2] , \wRegInTop_5_17[1] , 
        \wRegInTop_5_17[0] }) );
    BHeap_Node_WIDTH32 BHN_4_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_11[0] ), .P_In({\wRegOut_4_11[31] , 
        \wRegOut_4_11[30] , \wRegOut_4_11[29] , \wRegOut_4_11[28] , 
        \wRegOut_4_11[27] , \wRegOut_4_11[26] , \wRegOut_4_11[25] , 
        \wRegOut_4_11[24] , \wRegOut_4_11[23] , \wRegOut_4_11[22] , 
        \wRegOut_4_11[21] , \wRegOut_4_11[20] , \wRegOut_4_11[19] , 
        \wRegOut_4_11[18] , \wRegOut_4_11[17] , \wRegOut_4_11[16] , 
        \wRegOut_4_11[15] , \wRegOut_4_11[14] , \wRegOut_4_11[13] , 
        \wRegOut_4_11[12] , \wRegOut_4_11[11] , \wRegOut_4_11[10] , 
        \wRegOut_4_11[9] , \wRegOut_4_11[8] , \wRegOut_4_11[7] , 
        \wRegOut_4_11[6] , \wRegOut_4_11[5] , \wRegOut_4_11[4] , 
        \wRegOut_4_11[3] , \wRegOut_4_11[2] , \wRegOut_4_11[1] , 
        \wRegOut_4_11[0] }), .P_Out({\wRegInBot_4_11[31] , 
        \wRegInBot_4_11[30] , \wRegInBot_4_11[29] , \wRegInBot_4_11[28] , 
        \wRegInBot_4_11[27] , \wRegInBot_4_11[26] , \wRegInBot_4_11[25] , 
        \wRegInBot_4_11[24] , \wRegInBot_4_11[23] , \wRegInBot_4_11[22] , 
        \wRegInBot_4_11[21] , \wRegInBot_4_11[20] , \wRegInBot_4_11[19] , 
        \wRegInBot_4_11[18] , \wRegInBot_4_11[17] , \wRegInBot_4_11[16] , 
        \wRegInBot_4_11[15] , \wRegInBot_4_11[14] , \wRegInBot_4_11[13] , 
        \wRegInBot_4_11[12] , \wRegInBot_4_11[11] , \wRegInBot_4_11[10] , 
        \wRegInBot_4_11[9] , \wRegInBot_4_11[8] , \wRegInBot_4_11[7] , 
        \wRegInBot_4_11[6] , \wRegInBot_4_11[5] , \wRegInBot_4_11[4] , 
        \wRegInBot_4_11[3] , \wRegInBot_4_11[2] , \wRegInBot_4_11[1] , 
        \wRegInBot_4_11[0] }), .L_WR(\wRegEnTop_5_22[0] ), .L_In({
        \wRegOut_5_22[31] , \wRegOut_5_22[30] , \wRegOut_5_22[29] , 
        \wRegOut_5_22[28] , \wRegOut_5_22[27] , \wRegOut_5_22[26] , 
        \wRegOut_5_22[25] , \wRegOut_5_22[24] , \wRegOut_5_22[23] , 
        \wRegOut_5_22[22] , \wRegOut_5_22[21] , \wRegOut_5_22[20] , 
        \wRegOut_5_22[19] , \wRegOut_5_22[18] , \wRegOut_5_22[17] , 
        \wRegOut_5_22[16] , \wRegOut_5_22[15] , \wRegOut_5_22[14] , 
        \wRegOut_5_22[13] , \wRegOut_5_22[12] , \wRegOut_5_22[11] , 
        \wRegOut_5_22[10] , \wRegOut_5_22[9] , \wRegOut_5_22[8] , 
        \wRegOut_5_22[7] , \wRegOut_5_22[6] , \wRegOut_5_22[5] , 
        \wRegOut_5_22[4] , \wRegOut_5_22[3] , \wRegOut_5_22[2] , 
        \wRegOut_5_22[1] , \wRegOut_5_22[0] }), .L_Out({\wRegInTop_5_22[31] , 
        \wRegInTop_5_22[30] , \wRegInTop_5_22[29] , \wRegInTop_5_22[28] , 
        \wRegInTop_5_22[27] , \wRegInTop_5_22[26] , \wRegInTop_5_22[25] , 
        \wRegInTop_5_22[24] , \wRegInTop_5_22[23] , \wRegInTop_5_22[22] , 
        \wRegInTop_5_22[21] , \wRegInTop_5_22[20] , \wRegInTop_5_22[19] , 
        \wRegInTop_5_22[18] , \wRegInTop_5_22[17] , \wRegInTop_5_22[16] , 
        \wRegInTop_5_22[15] , \wRegInTop_5_22[14] , \wRegInTop_5_22[13] , 
        \wRegInTop_5_22[12] , \wRegInTop_5_22[11] , \wRegInTop_5_22[10] , 
        \wRegInTop_5_22[9] , \wRegInTop_5_22[8] , \wRegInTop_5_22[7] , 
        \wRegInTop_5_22[6] , \wRegInTop_5_22[5] , \wRegInTop_5_22[4] , 
        \wRegInTop_5_22[3] , \wRegInTop_5_22[2] , \wRegInTop_5_22[1] , 
        \wRegInTop_5_22[0] }), .R_WR(\wRegEnTop_5_23[0] ), .R_In({
        \wRegOut_5_23[31] , \wRegOut_5_23[30] , \wRegOut_5_23[29] , 
        \wRegOut_5_23[28] , \wRegOut_5_23[27] , \wRegOut_5_23[26] , 
        \wRegOut_5_23[25] , \wRegOut_5_23[24] , \wRegOut_5_23[23] , 
        \wRegOut_5_23[22] , \wRegOut_5_23[21] , \wRegOut_5_23[20] , 
        \wRegOut_5_23[19] , \wRegOut_5_23[18] , \wRegOut_5_23[17] , 
        \wRegOut_5_23[16] , \wRegOut_5_23[15] , \wRegOut_5_23[14] , 
        \wRegOut_5_23[13] , \wRegOut_5_23[12] , \wRegOut_5_23[11] , 
        \wRegOut_5_23[10] , \wRegOut_5_23[9] , \wRegOut_5_23[8] , 
        \wRegOut_5_23[7] , \wRegOut_5_23[6] , \wRegOut_5_23[5] , 
        \wRegOut_5_23[4] , \wRegOut_5_23[3] , \wRegOut_5_23[2] , 
        \wRegOut_5_23[1] , \wRegOut_5_23[0] }), .R_Out({\wRegInTop_5_23[31] , 
        \wRegInTop_5_23[30] , \wRegInTop_5_23[29] , \wRegInTop_5_23[28] , 
        \wRegInTop_5_23[27] , \wRegInTop_5_23[26] , \wRegInTop_5_23[25] , 
        \wRegInTop_5_23[24] , \wRegInTop_5_23[23] , \wRegInTop_5_23[22] , 
        \wRegInTop_5_23[21] , \wRegInTop_5_23[20] , \wRegInTop_5_23[19] , 
        \wRegInTop_5_23[18] , \wRegInTop_5_23[17] , \wRegInTop_5_23[16] , 
        \wRegInTop_5_23[15] , \wRegInTop_5_23[14] , \wRegInTop_5_23[13] , 
        \wRegInTop_5_23[12] , \wRegInTop_5_23[11] , \wRegInTop_5_23[10] , 
        \wRegInTop_5_23[9] , \wRegInTop_5_23[8] , \wRegInTop_5_23[7] , 
        \wRegInTop_5_23[6] , \wRegInTop_5_23[5] , \wRegInTop_5_23[4] , 
        \wRegInTop_5_23[3] , \wRegInTop_5_23[2] , \wRegInTop_5_23[1] , 
        \wRegInTop_5_23[0] }) );
    BHeap_Node_WIDTH32 BHN_6_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_55[0] ), .P_In({\wRegOut_6_55[31] , 
        \wRegOut_6_55[30] , \wRegOut_6_55[29] , \wRegOut_6_55[28] , 
        \wRegOut_6_55[27] , \wRegOut_6_55[26] , \wRegOut_6_55[25] , 
        \wRegOut_6_55[24] , \wRegOut_6_55[23] , \wRegOut_6_55[22] , 
        \wRegOut_6_55[21] , \wRegOut_6_55[20] , \wRegOut_6_55[19] , 
        \wRegOut_6_55[18] , \wRegOut_6_55[17] , \wRegOut_6_55[16] , 
        \wRegOut_6_55[15] , \wRegOut_6_55[14] , \wRegOut_6_55[13] , 
        \wRegOut_6_55[12] , \wRegOut_6_55[11] , \wRegOut_6_55[10] , 
        \wRegOut_6_55[9] , \wRegOut_6_55[8] , \wRegOut_6_55[7] , 
        \wRegOut_6_55[6] , \wRegOut_6_55[5] , \wRegOut_6_55[4] , 
        \wRegOut_6_55[3] , \wRegOut_6_55[2] , \wRegOut_6_55[1] , 
        \wRegOut_6_55[0] }), .P_Out({\wRegInBot_6_55[31] , 
        \wRegInBot_6_55[30] , \wRegInBot_6_55[29] , \wRegInBot_6_55[28] , 
        \wRegInBot_6_55[27] , \wRegInBot_6_55[26] , \wRegInBot_6_55[25] , 
        \wRegInBot_6_55[24] , \wRegInBot_6_55[23] , \wRegInBot_6_55[22] , 
        \wRegInBot_6_55[21] , \wRegInBot_6_55[20] , \wRegInBot_6_55[19] , 
        \wRegInBot_6_55[18] , \wRegInBot_6_55[17] , \wRegInBot_6_55[16] , 
        \wRegInBot_6_55[15] , \wRegInBot_6_55[14] , \wRegInBot_6_55[13] , 
        \wRegInBot_6_55[12] , \wRegInBot_6_55[11] , \wRegInBot_6_55[10] , 
        \wRegInBot_6_55[9] , \wRegInBot_6_55[8] , \wRegInBot_6_55[7] , 
        \wRegInBot_6_55[6] , \wRegInBot_6_55[5] , \wRegInBot_6_55[4] , 
        \wRegInBot_6_55[3] , \wRegInBot_6_55[2] , \wRegInBot_6_55[1] , 
        \wRegInBot_6_55[0] }), .L_WR(\wRegEnTop_7_110[0] ), .L_In({
        \wRegOut_7_110[31] , \wRegOut_7_110[30] , \wRegOut_7_110[29] , 
        \wRegOut_7_110[28] , \wRegOut_7_110[27] , \wRegOut_7_110[26] , 
        \wRegOut_7_110[25] , \wRegOut_7_110[24] , \wRegOut_7_110[23] , 
        \wRegOut_7_110[22] , \wRegOut_7_110[21] , \wRegOut_7_110[20] , 
        \wRegOut_7_110[19] , \wRegOut_7_110[18] , \wRegOut_7_110[17] , 
        \wRegOut_7_110[16] , \wRegOut_7_110[15] , \wRegOut_7_110[14] , 
        \wRegOut_7_110[13] , \wRegOut_7_110[12] , \wRegOut_7_110[11] , 
        \wRegOut_7_110[10] , \wRegOut_7_110[9] , \wRegOut_7_110[8] , 
        \wRegOut_7_110[7] , \wRegOut_7_110[6] , \wRegOut_7_110[5] , 
        \wRegOut_7_110[4] , \wRegOut_7_110[3] , \wRegOut_7_110[2] , 
        \wRegOut_7_110[1] , \wRegOut_7_110[0] }), .L_Out({
        \wRegInTop_7_110[31] , \wRegInTop_7_110[30] , \wRegInTop_7_110[29] , 
        \wRegInTop_7_110[28] , \wRegInTop_7_110[27] , \wRegInTop_7_110[26] , 
        \wRegInTop_7_110[25] , \wRegInTop_7_110[24] , \wRegInTop_7_110[23] , 
        \wRegInTop_7_110[22] , \wRegInTop_7_110[21] , \wRegInTop_7_110[20] , 
        \wRegInTop_7_110[19] , \wRegInTop_7_110[18] , \wRegInTop_7_110[17] , 
        \wRegInTop_7_110[16] , \wRegInTop_7_110[15] , \wRegInTop_7_110[14] , 
        \wRegInTop_7_110[13] , \wRegInTop_7_110[12] , \wRegInTop_7_110[11] , 
        \wRegInTop_7_110[10] , \wRegInTop_7_110[9] , \wRegInTop_7_110[8] , 
        \wRegInTop_7_110[7] , \wRegInTop_7_110[6] , \wRegInTop_7_110[5] , 
        \wRegInTop_7_110[4] , \wRegInTop_7_110[3] , \wRegInTop_7_110[2] , 
        \wRegInTop_7_110[1] , \wRegInTop_7_110[0] }), .R_WR(
        \wRegEnTop_7_111[0] ), .R_In({\wRegOut_7_111[31] , \wRegOut_7_111[30] , 
        \wRegOut_7_111[29] , \wRegOut_7_111[28] , \wRegOut_7_111[27] , 
        \wRegOut_7_111[26] , \wRegOut_7_111[25] , \wRegOut_7_111[24] , 
        \wRegOut_7_111[23] , \wRegOut_7_111[22] , \wRegOut_7_111[21] , 
        \wRegOut_7_111[20] , \wRegOut_7_111[19] , \wRegOut_7_111[18] , 
        \wRegOut_7_111[17] , \wRegOut_7_111[16] , \wRegOut_7_111[15] , 
        \wRegOut_7_111[14] , \wRegOut_7_111[13] , \wRegOut_7_111[12] , 
        \wRegOut_7_111[11] , \wRegOut_7_111[10] , \wRegOut_7_111[9] , 
        \wRegOut_7_111[8] , \wRegOut_7_111[7] , \wRegOut_7_111[6] , 
        \wRegOut_7_111[5] , \wRegOut_7_111[4] , \wRegOut_7_111[3] , 
        \wRegOut_7_111[2] , \wRegOut_7_111[1] , \wRegOut_7_111[0] }), .R_Out({
        \wRegInTop_7_111[31] , \wRegInTop_7_111[30] , \wRegInTop_7_111[29] , 
        \wRegInTop_7_111[28] , \wRegInTop_7_111[27] , \wRegInTop_7_111[26] , 
        \wRegInTop_7_111[25] , \wRegInTop_7_111[24] , \wRegInTop_7_111[23] , 
        \wRegInTop_7_111[22] , \wRegInTop_7_111[21] , \wRegInTop_7_111[20] , 
        \wRegInTop_7_111[19] , \wRegInTop_7_111[18] , \wRegInTop_7_111[17] , 
        \wRegInTop_7_111[16] , \wRegInTop_7_111[15] , \wRegInTop_7_111[14] , 
        \wRegInTop_7_111[13] , \wRegInTop_7_111[12] , \wRegInTop_7_111[11] , 
        \wRegInTop_7_111[10] , \wRegInTop_7_111[9] , \wRegInTop_7_111[8] , 
        \wRegInTop_7_111[7] , \wRegInTop_7_111[6] , \wRegInTop_7_111[5] , 
        \wRegInTop_7_111[4] , \wRegInTop_7_111[3] , \wRegInTop_7_111[2] , 
        \wRegInTop_7_111[1] , \wRegInTop_7_111[0] }) );
    BHeap_Node_WIDTH32 BHN_6_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_4[0] ), .P_In({\wRegOut_6_4[31] , 
        \wRegOut_6_4[30] , \wRegOut_6_4[29] , \wRegOut_6_4[28] , 
        \wRegOut_6_4[27] , \wRegOut_6_4[26] , \wRegOut_6_4[25] , 
        \wRegOut_6_4[24] , \wRegOut_6_4[23] , \wRegOut_6_4[22] , 
        \wRegOut_6_4[21] , \wRegOut_6_4[20] , \wRegOut_6_4[19] , 
        \wRegOut_6_4[18] , \wRegOut_6_4[17] , \wRegOut_6_4[16] , 
        \wRegOut_6_4[15] , \wRegOut_6_4[14] , \wRegOut_6_4[13] , 
        \wRegOut_6_4[12] , \wRegOut_6_4[11] , \wRegOut_6_4[10] , 
        \wRegOut_6_4[9] , \wRegOut_6_4[8] , \wRegOut_6_4[7] , \wRegOut_6_4[6] , 
        \wRegOut_6_4[5] , \wRegOut_6_4[4] , \wRegOut_6_4[3] , \wRegOut_6_4[2] , 
        \wRegOut_6_4[1] , \wRegOut_6_4[0] }), .P_Out({\wRegInBot_6_4[31] , 
        \wRegInBot_6_4[30] , \wRegInBot_6_4[29] , \wRegInBot_6_4[28] , 
        \wRegInBot_6_4[27] , \wRegInBot_6_4[26] , \wRegInBot_6_4[25] , 
        \wRegInBot_6_4[24] , \wRegInBot_6_4[23] , \wRegInBot_6_4[22] , 
        \wRegInBot_6_4[21] , \wRegInBot_6_4[20] , \wRegInBot_6_4[19] , 
        \wRegInBot_6_4[18] , \wRegInBot_6_4[17] , \wRegInBot_6_4[16] , 
        \wRegInBot_6_4[15] , \wRegInBot_6_4[14] , \wRegInBot_6_4[13] , 
        \wRegInBot_6_4[12] , \wRegInBot_6_4[11] , \wRegInBot_6_4[10] , 
        \wRegInBot_6_4[9] , \wRegInBot_6_4[8] , \wRegInBot_6_4[7] , 
        \wRegInBot_6_4[6] , \wRegInBot_6_4[5] , \wRegInBot_6_4[4] , 
        \wRegInBot_6_4[3] , \wRegInBot_6_4[2] , \wRegInBot_6_4[1] , 
        \wRegInBot_6_4[0] }), .L_WR(\wRegEnTop_7_8[0] ), .L_In({
        \wRegOut_7_8[31] , \wRegOut_7_8[30] , \wRegOut_7_8[29] , 
        \wRegOut_7_8[28] , \wRegOut_7_8[27] , \wRegOut_7_8[26] , 
        \wRegOut_7_8[25] , \wRegOut_7_8[24] , \wRegOut_7_8[23] , 
        \wRegOut_7_8[22] , \wRegOut_7_8[21] , \wRegOut_7_8[20] , 
        \wRegOut_7_8[19] , \wRegOut_7_8[18] , \wRegOut_7_8[17] , 
        \wRegOut_7_8[16] , \wRegOut_7_8[15] , \wRegOut_7_8[14] , 
        \wRegOut_7_8[13] , \wRegOut_7_8[12] , \wRegOut_7_8[11] , 
        \wRegOut_7_8[10] , \wRegOut_7_8[9] , \wRegOut_7_8[8] , 
        \wRegOut_7_8[7] , \wRegOut_7_8[6] , \wRegOut_7_8[5] , \wRegOut_7_8[4] , 
        \wRegOut_7_8[3] , \wRegOut_7_8[2] , \wRegOut_7_8[1] , \wRegOut_7_8[0] 
        }), .L_Out({\wRegInTop_7_8[31] , \wRegInTop_7_8[30] , 
        \wRegInTop_7_8[29] , \wRegInTop_7_8[28] , \wRegInTop_7_8[27] , 
        \wRegInTop_7_8[26] , \wRegInTop_7_8[25] , \wRegInTop_7_8[24] , 
        \wRegInTop_7_8[23] , \wRegInTop_7_8[22] , \wRegInTop_7_8[21] , 
        \wRegInTop_7_8[20] , \wRegInTop_7_8[19] , \wRegInTop_7_8[18] , 
        \wRegInTop_7_8[17] , \wRegInTop_7_8[16] , \wRegInTop_7_8[15] , 
        \wRegInTop_7_8[14] , \wRegInTop_7_8[13] , \wRegInTop_7_8[12] , 
        \wRegInTop_7_8[11] , \wRegInTop_7_8[10] , \wRegInTop_7_8[9] , 
        \wRegInTop_7_8[8] , \wRegInTop_7_8[7] , \wRegInTop_7_8[6] , 
        \wRegInTop_7_8[5] , \wRegInTop_7_8[4] , \wRegInTop_7_8[3] , 
        \wRegInTop_7_8[2] , \wRegInTop_7_8[1] , \wRegInTop_7_8[0] }), .R_WR(
        \wRegEnTop_7_9[0] ), .R_In({\wRegOut_7_9[31] , \wRegOut_7_9[30] , 
        \wRegOut_7_9[29] , \wRegOut_7_9[28] , \wRegOut_7_9[27] , 
        \wRegOut_7_9[26] , \wRegOut_7_9[25] , \wRegOut_7_9[24] , 
        \wRegOut_7_9[23] , \wRegOut_7_9[22] , \wRegOut_7_9[21] , 
        \wRegOut_7_9[20] , \wRegOut_7_9[19] , \wRegOut_7_9[18] , 
        \wRegOut_7_9[17] , \wRegOut_7_9[16] , \wRegOut_7_9[15] , 
        \wRegOut_7_9[14] , \wRegOut_7_9[13] , \wRegOut_7_9[12] , 
        \wRegOut_7_9[11] , \wRegOut_7_9[10] , \wRegOut_7_9[9] , 
        \wRegOut_7_9[8] , \wRegOut_7_9[7] , \wRegOut_7_9[6] , \wRegOut_7_9[5] , 
        \wRegOut_7_9[4] , \wRegOut_7_9[3] , \wRegOut_7_9[2] , \wRegOut_7_9[1] , 
        \wRegOut_7_9[0] }), .R_Out({\wRegInTop_7_9[31] , \wRegInTop_7_9[30] , 
        \wRegInTop_7_9[29] , \wRegInTop_7_9[28] , \wRegInTop_7_9[27] , 
        \wRegInTop_7_9[26] , \wRegInTop_7_9[25] , \wRegInTop_7_9[24] , 
        \wRegInTop_7_9[23] , \wRegInTop_7_9[22] , \wRegInTop_7_9[21] , 
        \wRegInTop_7_9[20] , \wRegInTop_7_9[19] , \wRegInTop_7_9[18] , 
        \wRegInTop_7_9[17] , \wRegInTop_7_9[16] , \wRegInTop_7_9[15] , 
        \wRegInTop_7_9[14] , \wRegInTop_7_9[13] , \wRegInTop_7_9[12] , 
        \wRegInTop_7_9[11] , \wRegInTop_7_9[10] , \wRegInTop_7_9[9] , 
        \wRegInTop_7_9[8] , \wRegInTop_7_9[7] , \wRegInTop_7_9[6] , 
        \wRegInTop_7_9[5] , \wRegInTop_7_9[4] , \wRegInTop_7_9[3] , 
        \wRegInTop_7_9[2] , \wRegInTop_7_9[1] , \wRegInTop_7_9[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_99 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink227[31] , \ScanLink227[30] , \ScanLink227[29] , 
        \ScanLink227[28] , \ScanLink227[27] , \ScanLink227[26] , 
        \ScanLink227[25] , \ScanLink227[24] , \ScanLink227[23] , 
        \ScanLink227[22] , \ScanLink227[21] , \ScanLink227[20] , 
        \ScanLink227[19] , \ScanLink227[18] , \ScanLink227[17] , 
        \ScanLink227[16] , \ScanLink227[15] , \ScanLink227[14] , 
        \ScanLink227[13] , \ScanLink227[12] , \ScanLink227[11] , 
        \ScanLink227[10] , \ScanLink227[9] , \ScanLink227[8] , 
        \ScanLink227[7] , \ScanLink227[6] , \ScanLink227[5] , \ScanLink227[4] , 
        \ScanLink227[3] , \ScanLink227[2] , \ScanLink227[1] , \ScanLink227[0] 
        }), .ScanOut({\ScanLink226[31] , \ScanLink226[30] , \ScanLink226[29] , 
        \ScanLink226[28] , \ScanLink226[27] , \ScanLink226[26] , 
        \ScanLink226[25] , \ScanLink226[24] , \ScanLink226[23] , 
        \ScanLink226[22] , \ScanLink226[21] , \ScanLink226[20] , 
        \ScanLink226[19] , \ScanLink226[18] , \ScanLink226[17] , 
        \ScanLink226[16] , \ScanLink226[15] , \ScanLink226[14] , 
        \ScanLink226[13] , \ScanLink226[12] , \ScanLink226[11] , 
        \ScanLink226[10] , \ScanLink226[9] , \ScanLink226[8] , 
        \ScanLink226[7] , \ScanLink226[6] , \ScanLink226[5] , \ScanLink226[4] , 
        \ScanLink226[3] , \ScanLink226[2] , \ScanLink226[1] , \ScanLink226[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_99[31] , 
        \wRegOut_7_99[30] , \wRegOut_7_99[29] , \wRegOut_7_99[28] , 
        \wRegOut_7_99[27] , \wRegOut_7_99[26] , \wRegOut_7_99[25] , 
        \wRegOut_7_99[24] , \wRegOut_7_99[23] , \wRegOut_7_99[22] , 
        \wRegOut_7_99[21] , \wRegOut_7_99[20] , \wRegOut_7_99[19] , 
        \wRegOut_7_99[18] , \wRegOut_7_99[17] , \wRegOut_7_99[16] , 
        \wRegOut_7_99[15] , \wRegOut_7_99[14] , \wRegOut_7_99[13] , 
        \wRegOut_7_99[12] , \wRegOut_7_99[11] , \wRegOut_7_99[10] , 
        \wRegOut_7_99[9] , \wRegOut_7_99[8] , \wRegOut_7_99[7] , 
        \wRegOut_7_99[6] , \wRegOut_7_99[5] , \wRegOut_7_99[4] , 
        \wRegOut_7_99[3] , \wRegOut_7_99[2] , \wRegOut_7_99[1] , 
        \wRegOut_7_99[0] }), .Enable1(\wRegEnTop_7_99[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_99[31] , \wRegInTop_7_99[30] , \wRegInTop_7_99[29] , 
        \wRegInTop_7_99[28] , \wRegInTop_7_99[27] , \wRegInTop_7_99[26] , 
        \wRegInTop_7_99[25] , \wRegInTop_7_99[24] , \wRegInTop_7_99[23] , 
        \wRegInTop_7_99[22] , \wRegInTop_7_99[21] , \wRegInTop_7_99[20] , 
        \wRegInTop_7_99[19] , \wRegInTop_7_99[18] , \wRegInTop_7_99[17] , 
        \wRegInTop_7_99[16] , \wRegInTop_7_99[15] , \wRegInTop_7_99[14] , 
        \wRegInTop_7_99[13] , \wRegInTop_7_99[12] , \wRegInTop_7_99[11] , 
        \wRegInTop_7_99[10] , \wRegInTop_7_99[9] , \wRegInTop_7_99[8] , 
        \wRegInTop_7_99[7] , \wRegInTop_7_99[6] , \wRegInTop_7_99[5] , 
        \wRegInTop_7_99[4] , \wRegInTop_7_99[3] , \wRegInTop_7_99[2] , 
        \wRegInTop_7_99[1] , \wRegInTop_7_99[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_8[0] ), .P_In({\wRegOut_5_8[31] , 
        \wRegOut_5_8[30] , \wRegOut_5_8[29] , \wRegOut_5_8[28] , 
        \wRegOut_5_8[27] , \wRegOut_5_8[26] , \wRegOut_5_8[25] , 
        \wRegOut_5_8[24] , \wRegOut_5_8[23] , \wRegOut_5_8[22] , 
        \wRegOut_5_8[21] , \wRegOut_5_8[20] , \wRegOut_5_8[19] , 
        \wRegOut_5_8[18] , \wRegOut_5_8[17] , \wRegOut_5_8[16] , 
        \wRegOut_5_8[15] , \wRegOut_5_8[14] , \wRegOut_5_8[13] , 
        \wRegOut_5_8[12] , \wRegOut_5_8[11] , \wRegOut_5_8[10] , 
        \wRegOut_5_8[9] , \wRegOut_5_8[8] , \wRegOut_5_8[7] , \wRegOut_5_8[6] , 
        \wRegOut_5_8[5] , \wRegOut_5_8[4] , \wRegOut_5_8[3] , \wRegOut_5_8[2] , 
        \wRegOut_5_8[1] , \wRegOut_5_8[0] }), .P_Out({\wRegInBot_5_8[31] , 
        \wRegInBot_5_8[30] , \wRegInBot_5_8[29] , \wRegInBot_5_8[28] , 
        \wRegInBot_5_8[27] , \wRegInBot_5_8[26] , \wRegInBot_5_8[25] , 
        \wRegInBot_5_8[24] , \wRegInBot_5_8[23] , \wRegInBot_5_8[22] , 
        \wRegInBot_5_8[21] , \wRegInBot_5_8[20] , \wRegInBot_5_8[19] , 
        \wRegInBot_5_8[18] , \wRegInBot_5_8[17] , \wRegInBot_5_8[16] , 
        \wRegInBot_5_8[15] , \wRegInBot_5_8[14] , \wRegInBot_5_8[13] , 
        \wRegInBot_5_8[12] , \wRegInBot_5_8[11] , \wRegInBot_5_8[10] , 
        \wRegInBot_5_8[9] , \wRegInBot_5_8[8] , \wRegInBot_5_8[7] , 
        \wRegInBot_5_8[6] , \wRegInBot_5_8[5] , \wRegInBot_5_8[4] , 
        \wRegInBot_5_8[3] , \wRegInBot_5_8[2] , \wRegInBot_5_8[1] , 
        \wRegInBot_5_8[0] }), .L_WR(\wRegEnTop_6_16[0] ), .L_In({
        \wRegOut_6_16[31] , \wRegOut_6_16[30] , \wRegOut_6_16[29] , 
        \wRegOut_6_16[28] , \wRegOut_6_16[27] , \wRegOut_6_16[26] , 
        \wRegOut_6_16[25] , \wRegOut_6_16[24] , \wRegOut_6_16[23] , 
        \wRegOut_6_16[22] , \wRegOut_6_16[21] , \wRegOut_6_16[20] , 
        \wRegOut_6_16[19] , \wRegOut_6_16[18] , \wRegOut_6_16[17] , 
        \wRegOut_6_16[16] , \wRegOut_6_16[15] , \wRegOut_6_16[14] , 
        \wRegOut_6_16[13] , \wRegOut_6_16[12] , \wRegOut_6_16[11] , 
        \wRegOut_6_16[10] , \wRegOut_6_16[9] , \wRegOut_6_16[8] , 
        \wRegOut_6_16[7] , \wRegOut_6_16[6] , \wRegOut_6_16[5] , 
        \wRegOut_6_16[4] , \wRegOut_6_16[3] , \wRegOut_6_16[2] , 
        \wRegOut_6_16[1] , \wRegOut_6_16[0] }), .L_Out({\wRegInTop_6_16[31] , 
        \wRegInTop_6_16[30] , \wRegInTop_6_16[29] , \wRegInTop_6_16[28] , 
        \wRegInTop_6_16[27] , \wRegInTop_6_16[26] , \wRegInTop_6_16[25] , 
        \wRegInTop_6_16[24] , \wRegInTop_6_16[23] , \wRegInTop_6_16[22] , 
        \wRegInTop_6_16[21] , \wRegInTop_6_16[20] , \wRegInTop_6_16[19] , 
        \wRegInTop_6_16[18] , \wRegInTop_6_16[17] , \wRegInTop_6_16[16] , 
        \wRegInTop_6_16[15] , \wRegInTop_6_16[14] , \wRegInTop_6_16[13] , 
        \wRegInTop_6_16[12] , \wRegInTop_6_16[11] , \wRegInTop_6_16[10] , 
        \wRegInTop_6_16[9] , \wRegInTop_6_16[8] , \wRegInTop_6_16[7] , 
        \wRegInTop_6_16[6] , \wRegInTop_6_16[5] , \wRegInTop_6_16[4] , 
        \wRegInTop_6_16[3] , \wRegInTop_6_16[2] , \wRegInTop_6_16[1] , 
        \wRegInTop_6_16[0] }), .R_WR(\wRegEnTop_6_17[0] ), .R_In({
        \wRegOut_6_17[31] , \wRegOut_6_17[30] , \wRegOut_6_17[29] , 
        \wRegOut_6_17[28] , \wRegOut_6_17[27] , \wRegOut_6_17[26] , 
        \wRegOut_6_17[25] , \wRegOut_6_17[24] , \wRegOut_6_17[23] , 
        \wRegOut_6_17[22] , \wRegOut_6_17[21] , \wRegOut_6_17[20] , 
        \wRegOut_6_17[19] , \wRegOut_6_17[18] , \wRegOut_6_17[17] , 
        \wRegOut_6_17[16] , \wRegOut_6_17[15] , \wRegOut_6_17[14] , 
        \wRegOut_6_17[13] , \wRegOut_6_17[12] , \wRegOut_6_17[11] , 
        \wRegOut_6_17[10] , \wRegOut_6_17[9] , \wRegOut_6_17[8] , 
        \wRegOut_6_17[7] , \wRegOut_6_17[6] , \wRegOut_6_17[5] , 
        \wRegOut_6_17[4] , \wRegOut_6_17[3] , \wRegOut_6_17[2] , 
        \wRegOut_6_17[1] , \wRegOut_6_17[0] }), .R_Out({\wRegInTop_6_17[31] , 
        \wRegInTop_6_17[30] , \wRegInTop_6_17[29] , \wRegInTop_6_17[28] , 
        \wRegInTop_6_17[27] , \wRegInTop_6_17[26] , \wRegInTop_6_17[25] , 
        \wRegInTop_6_17[24] , \wRegInTop_6_17[23] , \wRegInTop_6_17[22] , 
        \wRegInTop_6_17[21] , \wRegInTop_6_17[20] , \wRegInTop_6_17[19] , 
        \wRegInTop_6_17[18] , \wRegInTop_6_17[17] , \wRegInTop_6_17[16] , 
        \wRegInTop_6_17[15] , \wRegInTop_6_17[14] , \wRegInTop_6_17[13] , 
        \wRegInTop_6_17[12] , \wRegInTop_6_17[11] , \wRegInTop_6_17[10] , 
        \wRegInTop_6_17[9] , \wRegInTop_6_17[8] , \wRegInTop_6_17[7] , 
        \wRegInTop_6_17[6] , \wRegInTop_6_17[5] , \wRegInTop_6_17[4] , 
        \wRegInTop_6_17[3] , \wRegInTop_6_17[2] , \wRegInTop_6_17[1] , 
        \wRegInTop_6_17[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_35 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink163[31] , \ScanLink163[30] , \ScanLink163[29] , 
        \ScanLink163[28] , \ScanLink163[27] , \ScanLink163[26] , 
        \ScanLink163[25] , \ScanLink163[24] , \ScanLink163[23] , 
        \ScanLink163[22] , \ScanLink163[21] , \ScanLink163[20] , 
        \ScanLink163[19] , \ScanLink163[18] , \ScanLink163[17] , 
        \ScanLink163[16] , \ScanLink163[15] , \ScanLink163[14] , 
        \ScanLink163[13] , \ScanLink163[12] , \ScanLink163[11] , 
        \ScanLink163[10] , \ScanLink163[9] , \ScanLink163[8] , 
        \ScanLink163[7] , \ScanLink163[6] , \ScanLink163[5] , \ScanLink163[4] , 
        \ScanLink163[3] , \ScanLink163[2] , \ScanLink163[1] , \ScanLink163[0] 
        }), .ScanOut({\ScanLink162[31] , \ScanLink162[30] , \ScanLink162[29] , 
        \ScanLink162[28] , \ScanLink162[27] , \ScanLink162[26] , 
        \ScanLink162[25] , \ScanLink162[24] , \ScanLink162[23] , 
        \ScanLink162[22] , \ScanLink162[21] , \ScanLink162[20] , 
        \ScanLink162[19] , \ScanLink162[18] , \ScanLink162[17] , 
        \ScanLink162[16] , \ScanLink162[15] , \ScanLink162[14] , 
        \ScanLink162[13] , \ScanLink162[12] , \ScanLink162[11] , 
        \ScanLink162[10] , \ScanLink162[9] , \ScanLink162[8] , 
        \ScanLink162[7] , \ScanLink162[6] , \ScanLink162[5] , \ScanLink162[4] , 
        \ScanLink162[3] , \ScanLink162[2] , \ScanLink162[1] , \ScanLink162[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_35[31] , 
        \wRegOut_7_35[30] , \wRegOut_7_35[29] , \wRegOut_7_35[28] , 
        \wRegOut_7_35[27] , \wRegOut_7_35[26] , \wRegOut_7_35[25] , 
        \wRegOut_7_35[24] , \wRegOut_7_35[23] , \wRegOut_7_35[22] , 
        \wRegOut_7_35[21] , \wRegOut_7_35[20] , \wRegOut_7_35[19] , 
        \wRegOut_7_35[18] , \wRegOut_7_35[17] , \wRegOut_7_35[16] , 
        \wRegOut_7_35[15] , \wRegOut_7_35[14] , \wRegOut_7_35[13] , 
        \wRegOut_7_35[12] , \wRegOut_7_35[11] , \wRegOut_7_35[10] , 
        \wRegOut_7_35[9] , \wRegOut_7_35[8] , \wRegOut_7_35[7] , 
        \wRegOut_7_35[6] , \wRegOut_7_35[5] , \wRegOut_7_35[4] , 
        \wRegOut_7_35[3] , \wRegOut_7_35[2] , \wRegOut_7_35[1] , 
        \wRegOut_7_35[0] }), .Enable1(\wRegEnTop_7_35[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_35[31] , \wRegInTop_7_35[30] , \wRegInTop_7_35[29] , 
        \wRegInTop_7_35[28] , \wRegInTop_7_35[27] , \wRegInTop_7_35[26] , 
        \wRegInTop_7_35[25] , \wRegInTop_7_35[24] , \wRegInTop_7_35[23] , 
        \wRegInTop_7_35[22] , \wRegInTop_7_35[21] , \wRegInTop_7_35[20] , 
        \wRegInTop_7_35[19] , \wRegInTop_7_35[18] , \wRegInTop_7_35[17] , 
        \wRegInTop_7_35[16] , \wRegInTop_7_35[15] , \wRegInTop_7_35[14] , 
        \wRegInTop_7_35[13] , \wRegInTop_7_35[12] , \wRegInTop_7_35[11] , 
        \wRegInTop_7_35[10] , \wRegInTop_7_35[9] , \wRegInTop_7_35[8] , 
        \wRegInTop_7_35[7] , \wRegInTop_7_35[6] , \wRegInTop_7_35[5] , 
        \wRegInTop_7_35[4] , \wRegInTop_7_35[3] , \wRegInTop_7_35[2] , 
        \wRegInTop_7_35[1] , \wRegInTop_7_35[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_106 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink234[31] , \ScanLink234[30] , \ScanLink234[29] , 
        \ScanLink234[28] , \ScanLink234[27] , \ScanLink234[26] , 
        \ScanLink234[25] , \ScanLink234[24] , \ScanLink234[23] , 
        \ScanLink234[22] , \ScanLink234[21] , \ScanLink234[20] , 
        \ScanLink234[19] , \ScanLink234[18] , \ScanLink234[17] , 
        \ScanLink234[16] , \ScanLink234[15] , \ScanLink234[14] , 
        \ScanLink234[13] , \ScanLink234[12] , \ScanLink234[11] , 
        \ScanLink234[10] , \ScanLink234[9] , \ScanLink234[8] , 
        \ScanLink234[7] , \ScanLink234[6] , \ScanLink234[5] , \ScanLink234[4] , 
        \ScanLink234[3] , \ScanLink234[2] , \ScanLink234[1] , \ScanLink234[0] 
        }), .ScanOut({\ScanLink233[31] , \ScanLink233[30] , \ScanLink233[29] , 
        \ScanLink233[28] , \ScanLink233[27] , \ScanLink233[26] , 
        \ScanLink233[25] , \ScanLink233[24] , \ScanLink233[23] , 
        \ScanLink233[22] , \ScanLink233[21] , \ScanLink233[20] , 
        \ScanLink233[19] , \ScanLink233[18] , \ScanLink233[17] , 
        \ScanLink233[16] , \ScanLink233[15] , \ScanLink233[14] , 
        \ScanLink233[13] , \ScanLink233[12] , \ScanLink233[11] , 
        \ScanLink233[10] , \ScanLink233[9] , \ScanLink233[8] , 
        \ScanLink233[7] , \ScanLink233[6] , \ScanLink233[5] , \ScanLink233[4] , 
        \ScanLink233[3] , \ScanLink233[2] , \ScanLink233[1] , \ScanLink233[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_106[31] , 
        \wRegOut_7_106[30] , \wRegOut_7_106[29] , \wRegOut_7_106[28] , 
        \wRegOut_7_106[27] , \wRegOut_7_106[26] , \wRegOut_7_106[25] , 
        \wRegOut_7_106[24] , \wRegOut_7_106[23] , \wRegOut_7_106[22] , 
        \wRegOut_7_106[21] , \wRegOut_7_106[20] , \wRegOut_7_106[19] , 
        \wRegOut_7_106[18] , \wRegOut_7_106[17] , \wRegOut_7_106[16] , 
        \wRegOut_7_106[15] , \wRegOut_7_106[14] , \wRegOut_7_106[13] , 
        \wRegOut_7_106[12] , \wRegOut_7_106[11] , \wRegOut_7_106[10] , 
        \wRegOut_7_106[9] , \wRegOut_7_106[8] , \wRegOut_7_106[7] , 
        \wRegOut_7_106[6] , \wRegOut_7_106[5] , \wRegOut_7_106[4] , 
        \wRegOut_7_106[3] , \wRegOut_7_106[2] , \wRegOut_7_106[1] , 
        \wRegOut_7_106[0] }), .Enable1(\wRegEnTop_7_106[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_106[31] , \wRegInTop_7_106[30] , 
        \wRegInTop_7_106[29] , \wRegInTop_7_106[28] , \wRegInTop_7_106[27] , 
        \wRegInTop_7_106[26] , \wRegInTop_7_106[25] , \wRegInTop_7_106[24] , 
        \wRegInTop_7_106[23] , \wRegInTop_7_106[22] , \wRegInTop_7_106[21] , 
        \wRegInTop_7_106[20] , \wRegInTop_7_106[19] , \wRegInTop_7_106[18] , 
        \wRegInTop_7_106[17] , \wRegInTop_7_106[16] , \wRegInTop_7_106[15] , 
        \wRegInTop_7_106[14] , \wRegInTop_7_106[13] , \wRegInTop_7_106[12] , 
        \wRegInTop_7_106[11] , \wRegInTop_7_106[10] , \wRegInTop_7_106[9] , 
        \wRegInTop_7_106[8] , \wRegInTop_7_106[7] , \wRegInTop_7_106[6] , 
        \wRegInTop_7_106[5] , \wRegInTop_7_106[4] , \wRegInTop_7_106[3] , 
        \wRegInTop_7_106[2] , \wRegInTop_7_106[1] , \wRegInTop_7_106[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_2[0] ), .P_WR(\wRegEnBot_2_2[0] ), .P_In({\wRegOut_2_2[31] , 
        \wRegOut_2_2[30] , \wRegOut_2_2[29] , \wRegOut_2_2[28] , 
        \wRegOut_2_2[27] , \wRegOut_2_2[26] , \wRegOut_2_2[25] , 
        \wRegOut_2_2[24] , \wRegOut_2_2[23] , \wRegOut_2_2[22] , 
        \wRegOut_2_2[21] , \wRegOut_2_2[20] , \wRegOut_2_2[19] , 
        \wRegOut_2_2[18] , \wRegOut_2_2[17] , \wRegOut_2_2[16] , 
        \wRegOut_2_2[15] , \wRegOut_2_2[14] , \wRegOut_2_2[13] , 
        \wRegOut_2_2[12] , \wRegOut_2_2[11] , \wRegOut_2_2[10] , 
        \wRegOut_2_2[9] , \wRegOut_2_2[8] , \wRegOut_2_2[7] , \wRegOut_2_2[6] , 
        \wRegOut_2_2[5] , \wRegOut_2_2[4] , \wRegOut_2_2[3] , \wRegOut_2_2[2] , 
        \wRegOut_2_2[1] , \wRegOut_2_2[0] }), .P_Out({\wRegInBot_2_2[31] , 
        \wRegInBot_2_2[30] , \wRegInBot_2_2[29] , \wRegInBot_2_2[28] , 
        \wRegInBot_2_2[27] , \wRegInBot_2_2[26] , \wRegInBot_2_2[25] , 
        \wRegInBot_2_2[24] , \wRegInBot_2_2[23] , \wRegInBot_2_2[22] , 
        \wRegInBot_2_2[21] , \wRegInBot_2_2[20] , \wRegInBot_2_2[19] , 
        \wRegInBot_2_2[18] , \wRegInBot_2_2[17] , \wRegInBot_2_2[16] , 
        \wRegInBot_2_2[15] , \wRegInBot_2_2[14] , \wRegInBot_2_2[13] , 
        \wRegInBot_2_2[12] , \wRegInBot_2_2[11] , \wRegInBot_2_2[10] , 
        \wRegInBot_2_2[9] , \wRegInBot_2_2[8] , \wRegInBot_2_2[7] , 
        \wRegInBot_2_2[6] , \wRegInBot_2_2[5] , \wRegInBot_2_2[4] , 
        \wRegInBot_2_2[3] , \wRegInBot_2_2[2] , \wRegInBot_2_2[1] , 
        \wRegInBot_2_2[0] }), .L_WR(\wRegEnTop_3_4[0] ), .L_In({
        \wRegOut_3_4[31] , \wRegOut_3_4[30] , \wRegOut_3_4[29] , 
        \wRegOut_3_4[28] , \wRegOut_3_4[27] , \wRegOut_3_4[26] , 
        \wRegOut_3_4[25] , \wRegOut_3_4[24] , \wRegOut_3_4[23] , 
        \wRegOut_3_4[22] , \wRegOut_3_4[21] , \wRegOut_3_4[20] , 
        \wRegOut_3_4[19] , \wRegOut_3_4[18] , \wRegOut_3_4[17] , 
        \wRegOut_3_4[16] , \wRegOut_3_4[15] , \wRegOut_3_4[14] , 
        \wRegOut_3_4[13] , \wRegOut_3_4[12] , \wRegOut_3_4[11] , 
        \wRegOut_3_4[10] , \wRegOut_3_4[9] , \wRegOut_3_4[8] , 
        \wRegOut_3_4[7] , \wRegOut_3_4[6] , \wRegOut_3_4[5] , \wRegOut_3_4[4] , 
        \wRegOut_3_4[3] , \wRegOut_3_4[2] , \wRegOut_3_4[1] , \wRegOut_3_4[0] 
        }), .L_Out({\wRegInTop_3_4[31] , \wRegInTop_3_4[30] , 
        \wRegInTop_3_4[29] , \wRegInTop_3_4[28] , \wRegInTop_3_4[27] , 
        \wRegInTop_3_4[26] , \wRegInTop_3_4[25] , \wRegInTop_3_4[24] , 
        \wRegInTop_3_4[23] , \wRegInTop_3_4[22] , \wRegInTop_3_4[21] , 
        \wRegInTop_3_4[20] , \wRegInTop_3_4[19] , \wRegInTop_3_4[18] , 
        \wRegInTop_3_4[17] , \wRegInTop_3_4[16] , \wRegInTop_3_4[15] , 
        \wRegInTop_3_4[14] , \wRegInTop_3_4[13] , \wRegInTop_3_4[12] , 
        \wRegInTop_3_4[11] , \wRegInTop_3_4[10] , \wRegInTop_3_4[9] , 
        \wRegInTop_3_4[8] , \wRegInTop_3_4[7] , \wRegInTop_3_4[6] , 
        \wRegInTop_3_4[5] , \wRegInTop_3_4[4] , \wRegInTop_3_4[3] , 
        \wRegInTop_3_4[2] , \wRegInTop_3_4[1] , \wRegInTop_3_4[0] }), .R_WR(
        \wRegEnTop_3_5[0] ), .R_In({\wRegOut_3_5[31] , \wRegOut_3_5[30] , 
        \wRegOut_3_5[29] , \wRegOut_3_5[28] , \wRegOut_3_5[27] , 
        \wRegOut_3_5[26] , \wRegOut_3_5[25] , \wRegOut_3_5[24] , 
        \wRegOut_3_5[23] , \wRegOut_3_5[22] , \wRegOut_3_5[21] , 
        \wRegOut_3_5[20] , \wRegOut_3_5[19] , \wRegOut_3_5[18] , 
        \wRegOut_3_5[17] , \wRegOut_3_5[16] , \wRegOut_3_5[15] , 
        \wRegOut_3_5[14] , \wRegOut_3_5[13] , \wRegOut_3_5[12] , 
        \wRegOut_3_5[11] , \wRegOut_3_5[10] , \wRegOut_3_5[9] , 
        \wRegOut_3_5[8] , \wRegOut_3_5[7] , \wRegOut_3_5[6] , \wRegOut_3_5[5] , 
        \wRegOut_3_5[4] , \wRegOut_3_5[3] , \wRegOut_3_5[2] , \wRegOut_3_5[1] , 
        \wRegOut_3_5[0] }), .R_Out({\wRegInTop_3_5[31] , \wRegInTop_3_5[30] , 
        \wRegInTop_3_5[29] , \wRegInTop_3_5[28] , \wRegInTop_3_5[27] , 
        \wRegInTop_3_5[26] , \wRegInTop_3_5[25] , \wRegInTop_3_5[24] , 
        \wRegInTop_3_5[23] , \wRegInTop_3_5[22] , \wRegInTop_3_5[21] , 
        \wRegInTop_3_5[20] , \wRegInTop_3_5[19] , \wRegInTop_3_5[18] , 
        \wRegInTop_3_5[17] , \wRegInTop_3_5[16] , \wRegInTop_3_5[15] , 
        \wRegInTop_3_5[14] , \wRegInTop_3_5[13] , \wRegInTop_3_5[12] , 
        \wRegInTop_3_5[11] , \wRegInTop_3_5[10] , \wRegInTop_3_5[9] , 
        \wRegInTop_3_5[8] , \wRegInTop_3_5[7] , \wRegInTop_3_5[6] , 
        \wRegInTop_3_5[5] , \wRegInTop_3_5[4] , \wRegInTop_3_5[3] , 
        \wRegInTop_3_5[2] , \wRegInTop_3_5[1] , \wRegInTop_3_5[0] }) );
    BHeap_CtrlReg_WIDTH32 BHCR_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_7[0] ), 
        .Out(\wCtrlOut_6[0] ), .Enable(\wEnable_6[0] ) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_121 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink249[31] , \ScanLink249[30] , \ScanLink249[29] , 
        \ScanLink249[28] , \ScanLink249[27] , \ScanLink249[26] , 
        \ScanLink249[25] , \ScanLink249[24] , \ScanLink249[23] , 
        \ScanLink249[22] , \ScanLink249[21] , \ScanLink249[20] , 
        \ScanLink249[19] , \ScanLink249[18] , \ScanLink249[17] , 
        \ScanLink249[16] , \ScanLink249[15] , \ScanLink249[14] , 
        \ScanLink249[13] , \ScanLink249[12] , \ScanLink249[11] , 
        \ScanLink249[10] , \ScanLink249[9] , \ScanLink249[8] , 
        \ScanLink249[7] , \ScanLink249[6] , \ScanLink249[5] , \ScanLink249[4] , 
        \ScanLink249[3] , \ScanLink249[2] , \ScanLink249[1] , \ScanLink249[0] 
        }), .ScanOut({\ScanLink248[31] , \ScanLink248[30] , \ScanLink248[29] , 
        \ScanLink248[28] , \ScanLink248[27] , \ScanLink248[26] , 
        \ScanLink248[25] , \ScanLink248[24] , \ScanLink248[23] , 
        \ScanLink248[22] , \ScanLink248[21] , \ScanLink248[20] , 
        \ScanLink248[19] , \ScanLink248[18] , \ScanLink248[17] , 
        \ScanLink248[16] , \ScanLink248[15] , \ScanLink248[14] , 
        \ScanLink248[13] , \ScanLink248[12] , \ScanLink248[11] , 
        \ScanLink248[10] , \ScanLink248[9] , \ScanLink248[8] , 
        \ScanLink248[7] , \ScanLink248[6] , \ScanLink248[5] , \ScanLink248[4] , 
        \ScanLink248[3] , \ScanLink248[2] , \ScanLink248[1] , \ScanLink248[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_121[31] , 
        \wRegOut_7_121[30] , \wRegOut_7_121[29] , \wRegOut_7_121[28] , 
        \wRegOut_7_121[27] , \wRegOut_7_121[26] , \wRegOut_7_121[25] , 
        \wRegOut_7_121[24] , \wRegOut_7_121[23] , \wRegOut_7_121[22] , 
        \wRegOut_7_121[21] , \wRegOut_7_121[20] , \wRegOut_7_121[19] , 
        \wRegOut_7_121[18] , \wRegOut_7_121[17] , \wRegOut_7_121[16] , 
        \wRegOut_7_121[15] , \wRegOut_7_121[14] , \wRegOut_7_121[13] , 
        \wRegOut_7_121[12] , \wRegOut_7_121[11] , \wRegOut_7_121[10] , 
        \wRegOut_7_121[9] , \wRegOut_7_121[8] , \wRegOut_7_121[7] , 
        \wRegOut_7_121[6] , \wRegOut_7_121[5] , \wRegOut_7_121[4] , 
        \wRegOut_7_121[3] , \wRegOut_7_121[2] , \wRegOut_7_121[1] , 
        \wRegOut_7_121[0] }), .Enable1(\wRegEnTop_7_121[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_121[31] , \wRegInTop_7_121[30] , 
        \wRegInTop_7_121[29] , \wRegInTop_7_121[28] , \wRegInTop_7_121[27] , 
        \wRegInTop_7_121[26] , \wRegInTop_7_121[25] , \wRegInTop_7_121[24] , 
        \wRegInTop_7_121[23] , \wRegInTop_7_121[22] , \wRegInTop_7_121[21] , 
        \wRegInTop_7_121[20] , \wRegInTop_7_121[19] , \wRegInTop_7_121[18] , 
        \wRegInTop_7_121[17] , \wRegInTop_7_121[16] , \wRegInTop_7_121[15] , 
        \wRegInTop_7_121[14] , \wRegInTop_7_121[13] , \wRegInTop_7_121[12] , 
        \wRegInTop_7_121[11] , \wRegInTop_7_121[10] , \wRegInTop_7_121[9] , 
        \wRegInTop_7_121[8] , \wRegInTop_7_121[7] , \wRegInTop_7_121[6] , 
        \wRegInTop_7_121[5] , \wRegInTop_7_121[4] , \wRegInTop_7_121[3] , 
        \wRegInTop_7_121[2] , \wRegInTop_7_121[1] , \wRegInTop_7_121[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_5_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_10[0] ), .P_In({\wRegOut_5_10[31] , 
        \wRegOut_5_10[30] , \wRegOut_5_10[29] , \wRegOut_5_10[28] , 
        \wRegOut_5_10[27] , \wRegOut_5_10[26] , \wRegOut_5_10[25] , 
        \wRegOut_5_10[24] , \wRegOut_5_10[23] , \wRegOut_5_10[22] , 
        \wRegOut_5_10[21] , \wRegOut_5_10[20] , \wRegOut_5_10[19] , 
        \wRegOut_5_10[18] , \wRegOut_5_10[17] , \wRegOut_5_10[16] , 
        \wRegOut_5_10[15] , \wRegOut_5_10[14] , \wRegOut_5_10[13] , 
        \wRegOut_5_10[12] , \wRegOut_5_10[11] , \wRegOut_5_10[10] , 
        \wRegOut_5_10[9] , \wRegOut_5_10[8] , \wRegOut_5_10[7] , 
        \wRegOut_5_10[6] , \wRegOut_5_10[5] , \wRegOut_5_10[4] , 
        \wRegOut_5_10[3] , \wRegOut_5_10[2] , \wRegOut_5_10[1] , 
        \wRegOut_5_10[0] }), .P_Out({\wRegInBot_5_10[31] , 
        \wRegInBot_5_10[30] , \wRegInBot_5_10[29] , \wRegInBot_5_10[28] , 
        \wRegInBot_5_10[27] , \wRegInBot_5_10[26] , \wRegInBot_5_10[25] , 
        \wRegInBot_5_10[24] , \wRegInBot_5_10[23] , \wRegInBot_5_10[22] , 
        \wRegInBot_5_10[21] , \wRegInBot_5_10[20] , \wRegInBot_5_10[19] , 
        \wRegInBot_5_10[18] , \wRegInBot_5_10[17] , \wRegInBot_5_10[16] , 
        \wRegInBot_5_10[15] , \wRegInBot_5_10[14] , \wRegInBot_5_10[13] , 
        \wRegInBot_5_10[12] , \wRegInBot_5_10[11] , \wRegInBot_5_10[10] , 
        \wRegInBot_5_10[9] , \wRegInBot_5_10[8] , \wRegInBot_5_10[7] , 
        \wRegInBot_5_10[6] , \wRegInBot_5_10[5] , \wRegInBot_5_10[4] , 
        \wRegInBot_5_10[3] , \wRegInBot_5_10[2] , \wRegInBot_5_10[1] , 
        \wRegInBot_5_10[0] }), .L_WR(\wRegEnTop_6_20[0] ), .L_In({
        \wRegOut_6_20[31] , \wRegOut_6_20[30] , \wRegOut_6_20[29] , 
        \wRegOut_6_20[28] , \wRegOut_6_20[27] , \wRegOut_6_20[26] , 
        \wRegOut_6_20[25] , \wRegOut_6_20[24] , \wRegOut_6_20[23] , 
        \wRegOut_6_20[22] , \wRegOut_6_20[21] , \wRegOut_6_20[20] , 
        \wRegOut_6_20[19] , \wRegOut_6_20[18] , \wRegOut_6_20[17] , 
        \wRegOut_6_20[16] , \wRegOut_6_20[15] , \wRegOut_6_20[14] , 
        \wRegOut_6_20[13] , \wRegOut_6_20[12] , \wRegOut_6_20[11] , 
        \wRegOut_6_20[10] , \wRegOut_6_20[9] , \wRegOut_6_20[8] , 
        \wRegOut_6_20[7] , \wRegOut_6_20[6] , \wRegOut_6_20[5] , 
        \wRegOut_6_20[4] , \wRegOut_6_20[3] , \wRegOut_6_20[2] , 
        \wRegOut_6_20[1] , \wRegOut_6_20[0] }), .L_Out({\wRegInTop_6_20[31] , 
        \wRegInTop_6_20[30] , \wRegInTop_6_20[29] , \wRegInTop_6_20[28] , 
        \wRegInTop_6_20[27] , \wRegInTop_6_20[26] , \wRegInTop_6_20[25] , 
        \wRegInTop_6_20[24] , \wRegInTop_6_20[23] , \wRegInTop_6_20[22] , 
        \wRegInTop_6_20[21] , \wRegInTop_6_20[20] , \wRegInTop_6_20[19] , 
        \wRegInTop_6_20[18] , \wRegInTop_6_20[17] , \wRegInTop_6_20[16] , 
        \wRegInTop_6_20[15] , \wRegInTop_6_20[14] , \wRegInTop_6_20[13] , 
        \wRegInTop_6_20[12] , \wRegInTop_6_20[11] , \wRegInTop_6_20[10] , 
        \wRegInTop_6_20[9] , \wRegInTop_6_20[8] , \wRegInTop_6_20[7] , 
        \wRegInTop_6_20[6] , \wRegInTop_6_20[5] , \wRegInTop_6_20[4] , 
        \wRegInTop_6_20[3] , \wRegInTop_6_20[2] , \wRegInTop_6_20[1] , 
        \wRegInTop_6_20[0] }), .R_WR(\wRegEnTop_6_21[0] ), .R_In({
        \wRegOut_6_21[31] , \wRegOut_6_21[30] , \wRegOut_6_21[29] , 
        \wRegOut_6_21[28] , \wRegOut_6_21[27] , \wRegOut_6_21[26] , 
        \wRegOut_6_21[25] , \wRegOut_6_21[24] , \wRegOut_6_21[23] , 
        \wRegOut_6_21[22] , \wRegOut_6_21[21] , \wRegOut_6_21[20] , 
        \wRegOut_6_21[19] , \wRegOut_6_21[18] , \wRegOut_6_21[17] , 
        \wRegOut_6_21[16] , \wRegOut_6_21[15] , \wRegOut_6_21[14] , 
        \wRegOut_6_21[13] , \wRegOut_6_21[12] , \wRegOut_6_21[11] , 
        \wRegOut_6_21[10] , \wRegOut_6_21[9] , \wRegOut_6_21[8] , 
        \wRegOut_6_21[7] , \wRegOut_6_21[6] , \wRegOut_6_21[5] , 
        \wRegOut_6_21[4] , \wRegOut_6_21[3] , \wRegOut_6_21[2] , 
        \wRegOut_6_21[1] , \wRegOut_6_21[0] }), .R_Out({\wRegInTop_6_21[31] , 
        \wRegInTop_6_21[30] , \wRegInTop_6_21[29] , \wRegInTop_6_21[28] , 
        \wRegInTop_6_21[27] , \wRegInTop_6_21[26] , \wRegInTop_6_21[25] , 
        \wRegInTop_6_21[24] , \wRegInTop_6_21[23] , \wRegInTop_6_21[22] , 
        \wRegInTop_6_21[21] , \wRegInTop_6_21[20] , \wRegInTop_6_21[19] , 
        \wRegInTop_6_21[18] , \wRegInTop_6_21[17] , \wRegInTop_6_21[16] , 
        \wRegInTop_6_21[15] , \wRegInTop_6_21[14] , \wRegInTop_6_21[13] , 
        \wRegInTop_6_21[12] , \wRegInTop_6_21[11] , \wRegInTop_6_21[10] , 
        \wRegInTop_6_21[9] , \wRegInTop_6_21[8] , \wRegInTop_6_21[7] , 
        \wRegInTop_6_21[6] , \wRegInTop_6_21[5] , \wRegInTop_6_21[4] , 
        \wRegInTop_6_21[3] , \wRegInTop_6_21[2] , \wRegInTop_6_21[1] , 
        \wRegInTop_6_21[0] }) );
    BHeap_Node_WIDTH32 BHN_6_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_20[0] ), .P_In({\wRegOut_6_20[31] , 
        \wRegOut_6_20[30] , \wRegOut_6_20[29] , \wRegOut_6_20[28] , 
        \wRegOut_6_20[27] , \wRegOut_6_20[26] , \wRegOut_6_20[25] , 
        \wRegOut_6_20[24] , \wRegOut_6_20[23] , \wRegOut_6_20[22] , 
        \wRegOut_6_20[21] , \wRegOut_6_20[20] , \wRegOut_6_20[19] , 
        \wRegOut_6_20[18] , \wRegOut_6_20[17] , \wRegOut_6_20[16] , 
        \wRegOut_6_20[15] , \wRegOut_6_20[14] , \wRegOut_6_20[13] , 
        \wRegOut_6_20[12] , \wRegOut_6_20[11] , \wRegOut_6_20[10] , 
        \wRegOut_6_20[9] , \wRegOut_6_20[8] , \wRegOut_6_20[7] , 
        \wRegOut_6_20[6] , \wRegOut_6_20[5] , \wRegOut_6_20[4] , 
        \wRegOut_6_20[3] , \wRegOut_6_20[2] , \wRegOut_6_20[1] , 
        \wRegOut_6_20[0] }), .P_Out({\wRegInBot_6_20[31] , 
        \wRegInBot_6_20[30] , \wRegInBot_6_20[29] , \wRegInBot_6_20[28] , 
        \wRegInBot_6_20[27] , \wRegInBot_6_20[26] , \wRegInBot_6_20[25] , 
        \wRegInBot_6_20[24] , \wRegInBot_6_20[23] , \wRegInBot_6_20[22] , 
        \wRegInBot_6_20[21] , \wRegInBot_6_20[20] , \wRegInBot_6_20[19] , 
        \wRegInBot_6_20[18] , \wRegInBot_6_20[17] , \wRegInBot_6_20[16] , 
        \wRegInBot_6_20[15] , \wRegInBot_6_20[14] , \wRegInBot_6_20[13] , 
        \wRegInBot_6_20[12] , \wRegInBot_6_20[11] , \wRegInBot_6_20[10] , 
        \wRegInBot_6_20[9] , \wRegInBot_6_20[8] , \wRegInBot_6_20[7] , 
        \wRegInBot_6_20[6] , \wRegInBot_6_20[5] , \wRegInBot_6_20[4] , 
        \wRegInBot_6_20[3] , \wRegInBot_6_20[2] , \wRegInBot_6_20[1] , 
        \wRegInBot_6_20[0] }), .L_WR(\wRegEnTop_7_40[0] ), .L_In({
        \wRegOut_7_40[31] , \wRegOut_7_40[30] , \wRegOut_7_40[29] , 
        \wRegOut_7_40[28] , \wRegOut_7_40[27] , \wRegOut_7_40[26] , 
        \wRegOut_7_40[25] , \wRegOut_7_40[24] , \wRegOut_7_40[23] , 
        \wRegOut_7_40[22] , \wRegOut_7_40[21] , \wRegOut_7_40[20] , 
        \wRegOut_7_40[19] , \wRegOut_7_40[18] , \wRegOut_7_40[17] , 
        \wRegOut_7_40[16] , \wRegOut_7_40[15] , \wRegOut_7_40[14] , 
        \wRegOut_7_40[13] , \wRegOut_7_40[12] , \wRegOut_7_40[11] , 
        \wRegOut_7_40[10] , \wRegOut_7_40[9] , \wRegOut_7_40[8] , 
        \wRegOut_7_40[7] , \wRegOut_7_40[6] , \wRegOut_7_40[5] , 
        \wRegOut_7_40[4] , \wRegOut_7_40[3] , \wRegOut_7_40[2] , 
        \wRegOut_7_40[1] , \wRegOut_7_40[0] }), .L_Out({\wRegInTop_7_40[31] , 
        \wRegInTop_7_40[30] , \wRegInTop_7_40[29] , \wRegInTop_7_40[28] , 
        \wRegInTop_7_40[27] , \wRegInTop_7_40[26] , \wRegInTop_7_40[25] , 
        \wRegInTop_7_40[24] , \wRegInTop_7_40[23] , \wRegInTop_7_40[22] , 
        \wRegInTop_7_40[21] , \wRegInTop_7_40[20] , \wRegInTop_7_40[19] , 
        \wRegInTop_7_40[18] , \wRegInTop_7_40[17] , \wRegInTop_7_40[16] , 
        \wRegInTop_7_40[15] , \wRegInTop_7_40[14] , \wRegInTop_7_40[13] , 
        \wRegInTop_7_40[12] , \wRegInTop_7_40[11] , \wRegInTop_7_40[10] , 
        \wRegInTop_7_40[9] , \wRegInTop_7_40[8] , \wRegInTop_7_40[7] , 
        \wRegInTop_7_40[6] , \wRegInTop_7_40[5] , \wRegInTop_7_40[4] , 
        \wRegInTop_7_40[3] , \wRegInTop_7_40[2] , \wRegInTop_7_40[1] , 
        \wRegInTop_7_40[0] }), .R_WR(\wRegEnTop_7_41[0] ), .R_In({
        \wRegOut_7_41[31] , \wRegOut_7_41[30] , \wRegOut_7_41[29] , 
        \wRegOut_7_41[28] , \wRegOut_7_41[27] , \wRegOut_7_41[26] , 
        \wRegOut_7_41[25] , \wRegOut_7_41[24] , \wRegOut_7_41[23] , 
        \wRegOut_7_41[22] , \wRegOut_7_41[21] , \wRegOut_7_41[20] , 
        \wRegOut_7_41[19] , \wRegOut_7_41[18] , \wRegOut_7_41[17] , 
        \wRegOut_7_41[16] , \wRegOut_7_41[15] , \wRegOut_7_41[14] , 
        \wRegOut_7_41[13] , \wRegOut_7_41[12] , \wRegOut_7_41[11] , 
        \wRegOut_7_41[10] , \wRegOut_7_41[9] , \wRegOut_7_41[8] , 
        \wRegOut_7_41[7] , \wRegOut_7_41[6] , \wRegOut_7_41[5] , 
        \wRegOut_7_41[4] , \wRegOut_7_41[3] , \wRegOut_7_41[2] , 
        \wRegOut_7_41[1] , \wRegOut_7_41[0] }), .R_Out({\wRegInTop_7_41[31] , 
        \wRegInTop_7_41[30] , \wRegInTop_7_41[29] , \wRegInTop_7_41[28] , 
        \wRegInTop_7_41[27] , \wRegInTop_7_41[26] , \wRegInTop_7_41[25] , 
        \wRegInTop_7_41[24] , \wRegInTop_7_41[23] , \wRegInTop_7_41[22] , 
        \wRegInTop_7_41[21] , \wRegInTop_7_41[20] , \wRegInTop_7_41[19] , 
        \wRegInTop_7_41[18] , \wRegInTop_7_41[17] , \wRegInTop_7_41[16] , 
        \wRegInTop_7_41[15] , \wRegInTop_7_41[14] , \wRegInTop_7_41[13] , 
        \wRegInTop_7_41[12] , \wRegInTop_7_41[11] , \wRegInTop_7_41[10] , 
        \wRegInTop_7_41[9] , \wRegInTop_7_41[8] , \wRegInTop_7_41[7] , 
        \wRegInTop_7_41[6] , \wRegInTop_7_41[5] , \wRegInTop_7_41[4] , 
        \wRegInTop_7_41[3] , \wRegInTop_7_41[2] , \wRegInTop_7_41[1] , 
        \wRegInTop_7_41[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink15[31] , \ScanLink15[30] , \ScanLink15[29] , 
        \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , \ScanLink15[25] , 
        \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , \ScanLink15[21] , 
        \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , \ScanLink15[17] , 
        \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , \ScanLink15[13] , 
        \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , \ScanLink15[9] , 
        \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , \ScanLink15[5] , 
        \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , \ScanLink15[1] , 
        \ScanLink15[0] }), .ScanOut({\ScanLink14[31] , \ScanLink14[30] , 
        \ScanLink14[29] , \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , 
        \ScanLink14[25] , \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , 
        \ScanLink14[21] , \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , 
        \ScanLink14[17] , \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , 
        \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , 
        \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , 
        \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , 
        \ScanLink14[1] , \ScanLink14[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_7[31] , \wRegOut_3_7[30] , \wRegOut_3_7[29] , 
        \wRegOut_3_7[28] , \wRegOut_3_7[27] , \wRegOut_3_7[26] , 
        \wRegOut_3_7[25] , \wRegOut_3_7[24] , \wRegOut_3_7[23] , 
        \wRegOut_3_7[22] , \wRegOut_3_7[21] , \wRegOut_3_7[20] , 
        \wRegOut_3_7[19] , \wRegOut_3_7[18] , \wRegOut_3_7[17] , 
        \wRegOut_3_7[16] , \wRegOut_3_7[15] , \wRegOut_3_7[14] , 
        \wRegOut_3_7[13] , \wRegOut_3_7[12] , \wRegOut_3_7[11] , 
        \wRegOut_3_7[10] , \wRegOut_3_7[9] , \wRegOut_3_7[8] , 
        \wRegOut_3_7[7] , \wRegOut_3_7[6] , \wRegOut_3_7[5] , \wRegOut_3_7[4] , 
        \wRegOut_3_7[3] , \wRegOut_3_7[2] , \wRegOut_3_7[1] , \wRegOut_3_7[0] 
        }), .Enable1(\wRegEnTop_3_7[0] ), .Enable2(\wRegEnBot_3_7[0] ), .In1({
        \wRegInTop_3_7[31] , \wRegInTop_3_7[30] , \wRegInTop_3_7[29] , 
        \wRegInTop_3_7[28] , \wRegInTop_3_7[27] , \wRegInTop_3_7[26] , 
        \wRegInTop_3_7[25] , \wRegInTop_3_7[24] , \wRegInTop_3_7[23] , 
        \wRegInTop_3_7[22] , \wRegInTop_3_7[21] , \wRegInTop_3_7[20] , 
        \wRegInTop_3_7[19] , \wRegInTop_3_7[18] , \wRegInTop_3_7[17] , 
        \wRegInTop_3_7[16] , \wRegInTop_3_7[15] , \wRegInTop_3_7[14] , 
        \wRegInTop_3_7[13] , \wRegInTop_3_7[12] , \wRegInTop_3_7[11] , 
        \wRegInTop_3_7[10] , \wRegInTop_3_7[9] , \wRegInTop_3_7[8] , 
        \wRegInTop_3_7[7] , \wRegInTop_3_7[6] , \wRegInTop_3_7[5] , 
        \wRegInTop_3_7[4] , \wRegInTop_3_7[3] , \wRegInTop_3_7[2] , 
        \wRegInTop_3_7[1] , \wRegInTop_3_7[0] }), .In2({\wRegInBot_3_7[31] , 
        \wRegInBot_3_7[30] , \wRegInBot_3_7[29] , \wRegInBot_3_7[28] , 
        \wRegInBot_3_7[27] , \wRegInBot_3_7[26] , \wRegInBot_3_7[25] , 
        \wRegInBot_3_7[24] , \wRegInBot_3_7[23] , \wRegInBot_3_7[22] , 
        \wRegInBot_3_7[21] , \wRegInBot_3_7[20] , \wRegInBot_3_7[19] , 
        \wRegInBot_3_7[18] , \wRegInBot_3_7[17] , \wRegInBot_3_7[16] , 
        \wRegInBot_3_7[15] , \wRegInBot_3_7[14] , \wRegInBot_3_7[13] , 
        \wRegInBot_3_7[12] , \wRegInBot_3_7[11] , \wRegInBot_3_7[10] , 
        \wRegInBot_3_7[9] , \wRegInBot_3_7[8] , \wRegInBot_3_7[7] , 
        \wRegInBot_3_7[6] , \wRegInBot_3_7[5] , \wRegInBot_3_7[4] , 
        \wRegInBot_3_7[3] , \wRegInBot_3_7[2] , \wRegInBot_3_7[1] , 
        \wRegInBot_3_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_18 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink50[31] , \ScanLink50[30] , \ScanLink50[29] , 
        \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , \ScanLink50[25] , 
        \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , \ScanLink50[21] , 
        \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , \ScanLink50[17] , 
        \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , \ScanLink50[13] , 
        \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , \ScanLink50[9] , 
        \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , \ScanLink50[5] , 
        \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , \ScanLink50[1] , 
        \ScanLink50[0] }), .ScanOut({\ScanLink49[31] , \ScanLink49[30] , 
        \ScanLink49[29] , \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , 
        \ScanLink49[25] , \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , 
        \ScanLink49[21] , \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , 
        \ScanLink49[17] , \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , 
        \ScanLink49[13] , \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , 
        \ScanLink49[9] , \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , 
        \ScanLink49[5] , \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , 
        \ScanLink49[1] , \ScanLink49[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_18[31] , \wRegOut_5_18[30] , 
        \wRegOut_5_18[29] , \wRegOut_5_18[28] , \wRegOut_5_18[27] , 
        \wRegOut_5_18[26] , \wRegOut_5_18[25] , \wRegOut_5_18[24] , 
        \wRegOut_5_18[23] , \wRegOut_5_18[22] , \wRegOut_5_18[21] , 
        \wRegOut_5_18[20] , \wRegOut_5_18[19] , \wRegOut_5_18[18] , 
        \wRegOut_5_18[17] , \wRegOut_5_18[16] , \wRegOut_5_18[15] , 
        \wRegOut_5_18[14] , \wRegOut_5_18[13] , \wRegOut_5_18[12] , 
        \wRegOut_5_18[11] , \wRegOut_5_18[10] , \wRegOut_5_18[9] , 
        \wRegOut_5_18[8] , \wRegOut_5_18[7] , \wRegOut_5_18[6] , 
        \wRegOut_5_18[5] , \wRegOut_5_18[4] , \wRegOut_5_18[3] , 
        \wRegOut_5_18[2] , \wRegOut_5_18[1] , \wRegOut_5_18[0] }), .Enable1(
        \wRegEnTop_5_18[0] ), .Enable2(\wRegEnBot_5_18[0] ), .In1({
        \wRegInTop_5_18[31] , \wRegInTop_5_18[30] , \wRegInTop_5_18[29] , 
        \wRegInTop_5_18[28] , \wRegInTop_5_18[27] , \wRegInTop_5_18[26] , 
        \wRegInTop_5_18[25] , \wRegInTop_5_18[24] , \wRegInTop_5_18[23] , 
        \wRegInTop_5_18[22] , \wRegInTop_5_18[21] , \wRegInTop_5_18[20] , 
        \wRegInTop_5_18[19] , \wRegInTop_5_18[18] , \wRegInTop_5_18[17] , 
        \wRegInTop_5_18[16] , \wRegInTop_5_18[15] , \wRegInTop_5_18[14] , 
        \wRegInTop_5_18[13] , \wRegInTop_5_18[12] , \wRegInTop_5_18[11] , 
        \wRegInTop_5_18[10] , \wRegInTop_5_18[9] , \wRegInTop_5_18[8] , 
        \wRegInTop_5_18[7] , \wRegInTop_5_18[6] , \wRegInTop_5_18[5] , 
        \wRegInTop_5_18[4] , \wRegInTop_5_18[3] , \wRegInTop_5_18[2] , 
        \wRegInTop_5_18[1] , \wRegInTop_5_18[0] }), .In2({\wRegInBot_5_18[31] , 
        \wRegInBot_5_18[30] , \wRegInBot_5_18[29] , \wRegInBot_5_18[28] , 
        \wRegInBot_5_18[27] , \wRegInBot_5_18[26] , \wRegInBot_5_18[25] , 
        \wRegInBot_5_18[24] , \wRegInBot_5_18[23] , \wRegInBot_5_18[22] , 
        \wRegInBot_5_18[21] , \wRegInBot_5_18[20] , \wRegInBot_5_18[19] , 
        \wRegInBot_5_18[18] , \wRegInBot_5_18[17] , \wRegInBot_5_18[16] , 
        \wRegInBot_5_18[15] , \wRegInBot_5_18[14] , \wRegInBot_5_18[13] , 
        \wRegInBot_5_18[12] , \wRegInBot_5_18[11] , \wRegInBot_5_18[10] , 
        \wRegInBot_5_18[9] , \wRegInBot_5_18[8] , \wRegInBot_5_18[7] , 
        \wRegInBot_5_18[6] , \wRegInBot_5_18[5] , \wRegInBot_5_18[4] , 
        \wRegInBot_5_18[3] , \wRegInBot_5_18[2] , \wRegInBot_5_18[1] , 
        \wRegInBot_5_18[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_28 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink92[31] , \ScanLink92[30] , \ScanLink92[29] , 
        \ScanLink92[28] , \ScanLink92[27] , \ScanLink92[26] , \ScanLink92[25] , 
        \ScanLink92[24] , \ScanLink92[23] , \ScanLink92[22] , \ScanLink92[21] , 
        \ScanLink92[20] , \ScanLink92[19] , \ScanLink92[18] , \ScanLink92[17] , 
        \ScanLink92[16] , \ScanLink92[15] , \ScanLink92[14] , \ScanLink92[13] , 
        \ScanLink92[12] , \ScanLink92[11] , \ScanLink92[10] , \ScanLink92[9] , 
        \ScanLink92[8] , \ScanLink92[7] , \ScanLink92[6] , \ScanLink92[5] , 
        \ScanLink92[4] , \ScanLink92[3] , \ScanLink92[2] , \ScanLink92[1] , 
        \ScanLink92[0] }), .ScanOut({\ScanLink91[31] , \ScanLink91[30] , 
        \ScanLink91[29] , \ScanLink91[28] , \ScanLink91[27] , \ScanLink91[26] , 
        \ScanLink91[25] , \ScanLink91[24] , \ScanLink91[23] , \ScanLink91[22] , 
        \ScanLink91[21] , \ScanLink91[20] , \ScanLink91[19] , \ScanLink91[18] , 
        \ScanLink91[17] , \ScanLink91[16] , \ScanLink91[15] , \ScanLink91[14] , 
        \ScanLink91[13] , \ScanLink91[12] , \ScanLink91[11] , \ScanLink91[10] , 
        \ScanLink91[9] , \ScanLink91[8] , \ScanLink91[7] , \ScanLink91[6] , 
        \ScanLink91[5] , \ScanLink91[4] , \ScanLink91[3] , \ScanLink91[2] , 
        \ScanLink91[1] , \ScanLink91[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_28[31] , \wRegOut_6_28[30] , 
        \wRegOut_6_28[29] , \wRegOut_6_28[28] , \wRegOut_6_28[27] , 
        \wRegOut_6_28[26] , \wRegOut_6_28[25] , \wRegOut_6_28[24] , 
        \wRegOut_6_28[23] , \wRegOut_6_28[22] , \wRegOut_6_28[21] , 
        \wRegOut_6_28[20] , \wRegOut_6_28[19] , \wRegOut_6_28[18] , 
        \wRegOut_6_28[17] , \wRegOut_6_28[16] , \wRegOut_6_28[15] , 
        \wRegOut_6_28[14] , \wRegOut_6_28[13] , \wRegOut_6_28[12] , 
        \wRegOut_6_28[11] , \wRegOut_6_28[10] , \wRegOut_6_28[9] , 
        \wRegOut_6_28[8] , \wRegOut_6_28[7] , \wRegOut_6_28[6] , 
        \wRegOut_6_28[5] , \wRegOut_6_28[4] , \wRegOut_6_28[3] , 
        \wRegOut_6_28[2] , \wRegOut_6_28[1] , \wRegOut_6_28[0] }), .Enable1(
        \wRegEnTop_6_28[0] ), .Enable2(\wRegEnBot_6_28[0] ), .In1({
        \wRegInTop_6_28[31] , \wRegInTop_6_28[30] , \wRegInTop_6_28[29] , 
        \wRegInTop_6_28[28] , \wRegInTop_6_28[27] , \wRegInTop_6_28[26] , 
        \wRegInTop_6_28[25] , \wRegInTop_6_28[24] , \wRegInTop_6_28[23] , 
        \wRegInTop_6_28[22] , \wRegInTop_6_28[21] , \wRegInTop_6_28[20] , 
        \wRegInTop_6_28[19] , \wRegInTop_6_28[18] , \wRegInTop_6_28[17] , 
        \wRegInTop_6_28[16] , \wRegInTop_6_28[15] , \wRegInTop_6_28[14] , 
        \wRegInTop_6_28[13] , \wRegInTop_6_28[12] , \wRegInTop_6_28[11] , 
        \wRegInTop_6_28[10] , \wRegInTop_6_28[9] , \wRegInTop_6_28[8] , 
        \wRegInTop_6_28[7] , \wRegInTop_6_28[6] , \wRegInTop_6_28[5] , 
        \wRegInTop_6_28[4] , \wRegInTop_6_28[3] , \wRegInTop_6_28[2] , 
        \wRegInTop_6_28[1] , \wRegInTop_6_28[0] }), .In2({\wRegInBot_6_28[31] , 
        \wRegInBot_6_28[30] , \wRegInBot_6_28[29] , \wRegInBot_6_28[28] , 
        \wRegInBot_6_28[27] , \wRegInBot_6_28[26] , \wRegInBot_6_28[25] , 
        \wRegInBot_6_28[24] , \wRegInBot_6_28[23] , \wRegInBot_6_28[22] , 
        \wRegInBot_6_28[21] , \wRegInBot_6_28[20] , \wRegInBot_6_28[19] , 
        \wRegInBot_6_28[18] , \wRegInBot_6_28[17] , \wRegInBot_6_28[16] , 
        \wRegInBot_6_28[15] , \wRegInBot_6_28[14] , \wRegInBot_6_28[13] , 
        \wRegInBot_6_28[12] , \wRegInBot_6_28[11] , \wRegInBot_6_28[10] , 
        \wRegInBot_6_28[9] , \wRegInBot_6_28[8] , \wRegInBot_6_28[7] , 
        \wRegInBot_6_28[6] , \wRegInBot_6_28[5] , \wRegInBot_6_28[4] , 
        \wRegInBot_6_28[3] , \wRegInBot_6_28[2] , \wRegInBot_6_28[1] , 
        \wRegInBot_6_28[0] }) );
    BHeap_Node_WIDTH32 BHN_5_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_17[0] ), .P_In({\wRegOut_5_17[31] , 
        \wRegOut_5_17[30] , \wRegOut_5_17[29] , \wRegOut_5_17[28] , 
        \wRegOut_5_17[27] , \wRegOut_5_17[26] , \wRegOut_5_17[25] , 
        \wRegOut_5_17[24] , \wRegOut_5_17[23] , \wRegOut_5_17[22] , 
        \wRegOut_5_17[21] , \wRegOut_5_17[20] , \wRegOut_5_17[19] , 
        \wRegOut_5_17[18] , \wRegOut_5_17[17] , \wRegOut_5_17[16] , 
        \wRegOut_5_17[15] , \wRegOut_5_17[14] , \wRegOut_5_17[13] , 
        \wRegOut_5_17[12] , \wRegOut_5_17[11] , \wRegOut_5_17[10] , 
        \wRegOut_5_17[9] , \wRegOut_5_17[8] , \wRegOut_5_17[7] , 
        \wRegOut_5_17[6] , \wRegOut_5_17[5] , \wRegOut_5_17[4] , 
        \wRegOut_5_17[3] , \wRegOut_5_17[2] , \wRegOut_5_17[1] , 
        \wRegOut_5_17[0] }), .P_Out({\wRegInBot_5_17[31] , 
        \wRegInBot_5_17[30] , \wRegInBot_5_17[29] , \wRegInBot_5_17[28] , 
        \wRegInBot_5_17[27] , \wRegInBot_5_17[26] , \wRegInBot_5_17[25] , 
        \wRegInBot_5_17[24] , \wRegInBot_5_17[23] , \wRegInBot_5_17[22] , 
        \wRegInBot_5_17[21] , \wRegInBot_5_17[20] , \wRegInBot_5_17[19] , 
        \wRegInBot_5_17[18] , \wRegInBot_5_17[17] , \wRegInBot_5_17[16] , 
        \wRegInBot_5_17[15] , \wRegInBot_5_17[14] , \wRegInBot_5_17[13] , 
        \wRegInBot_5_17[12] , \wRegInBot_5_17[11] , \wRegInBot_5_17[10] , 
        \wRegInBot_5_17[9] , \wRegInBot_5_17[8] , \wRegInBot_5_17[7] , 
        \wRegInBot_5_17[6] , \wRegInBot_5_17[5] , \wRegInBot_5_17[4] , 
        \wRegInBot_5_17[3] , \wRegInBot_5_17[2] , \wRegInBot_5_17[1] , 
        \wRegInBot_5_17[0] }), .L_WR(\wRegEnTop_6_34[0] ), .L_In({
        \wRegOut_6_34[31] , \wRegOut_6_34[30] , \wRegOut_6_34[29] , 
        \wRegOut_6_34[28] , \wRegOut_6_34[27] , \wRegOut_6_34[26] , 
        \wRegOut_6_34[25] , \wRegOut_6_34[24] , \wRegOut_6_34[23] , 
        \wRegOut_6_34[22] , \wRegOut_6_34[21] , \wRegOut_6_34[20] , 
        \wRegOut_6_34[19] , \wRegOut_6_34[18] , \wRegOut_6_34[17] , 
        \wRegOut_6_34[16] , \wRegOut_6_34[15] , \wRegOut_6_34[14] , 
        \wRegOut_6_34[13] , \wRegOut_6_34[12] , \wRegOut_6_34[11] , 
        \wRegOut_6_34[10] , \wRegOut_6_34[9] , \wRegOut_6_34[8] , 
        \wRegOut_6_34[7] , \wRegOut_6_34[6] , \wRegOut_6_34[5] , 
        \wRegOut_6_34[4] , \wRegOut_6_34[3] , \wRegOut_6_34[2] , 
        \wRegOut_6_34[1] , \wRegOut_6_34[0] }), .L_Out({\wRegInTop_6_34[31] , 
        \wRegInTop_6_34[30] , \wRegInTop_6_34[29] , \wRegInTop_6_34[28] , 
        \wRegInTop_6_34[27] , \wRegInTop_6_34[26] , \wRegInTop_6_34[25] , 
        \wRegInTop_6_34[24] , \wRegInTop_6_34[23] , \wRegInTop_6_34[22] , 
        \wRegInTop_6_34[21] , \wRegInTop_6_34[20] , \wRegInTop_6_34[19] , 
        \wRegInTop_6_34[18] , \wRegInTop_6_34[17] , \wRegInTop_6_34[16] , 
        \wRegInTop_6_34[15] , \wRegInTop_6_34[14] , \wRegInTop_6_34[13] , 
        \wRegInTop_6_34[12] , \wRegInTop_6_34[11] , \wRegInTop_6_34[10] , 
        \wRegInTop_6_34[9] , \wRegInTop_6_34[8] , \wRegInTop_6_34[7] , 
        \wRegInTop_6_34[6] , \wRegInTop_6_34[5] , \wRegInTop_6_34[4] , 
        \wRegInTop_6_34[3] , \wRegInTop_6_34[2] , \wRegInTop_6_34[1] , 
        \wRegInTop_6_34[0] }), .R_WR(\wRegEnTop_6_35[0] ), .R_In({
        \wRegOut_6_35[31] , \wRegOut_6_35[30] , \wRegOut_6_35[29] , 
        \wRegOut_6_35[28] , \wRegOut_6_35[27] , \wRegOut_6_35[26] , 
        \wRegOut_6_35[25] , \wRegOut_6_35[24] , \wRegOut_6_35[23] , 
        \wRegOut_6_35[22] , \wRegOut_6_35[21] , \wRegOut_6_35[20] , 
        \wRegOut_6_35[19] , \wRegOut_6_35[18] , \wRegOut_6_35[17] , 
        \wRegOut_6_35[16] , \wRegOut_6_35[15] , \wRegOut_6_35[14] , 
        \wRegOut_6_35[13] , \wRegOut_6_35[12] , \wRegOut_6_35[11] , 
        \wRegOut_6_35[10] , \wRegOut_6_35[9] , \wRegOut_6_35[8] , 
        \wRegOut_6_35[7] , \wRegOut_6_35[6] , \wRegOut_6_35[5] , 
        \wRegOut_6_35[4] , \wRegOut_6_35[3] , \wRegOut_6_35[2] , 
        \wRegOut_6_35[1] , \wRegOut_6_35[0] }), .R_Out({\wRegInTop_6_35[31] , 
        \wRegInTop_6_35[30] , \wRegInTop_6_35[29] , \wRegInTop_6_35[28] , 
        \wRegInTop_6_35[27] , \wRegInTop_6_35[26] , \wRegInTop_6_35[25] , 
        \wRegInTop_6_35[24] , \wRegInTop_6_35[23] , \wRegInTop_6_35[22] , 
        \wRegInTop_6_35[21] , \wRegInTop_6_35[20] , \wRegInTop_6_35[19] , 
        \wRegInTop_6_35[18] , \wRegInTop_6_35[17] , \wRegInTop_6_35[16] , 
        \wRegInTop_6_35[15] , \wRegInTop_6_35[14] , \wRegInTop_6_35[13] , 
        \wRegInTop_6_35[12] , \wRegInTop_6_35[11] , \wRegInTop_6_35[10] , 
        \wRegInTop_6_35[9] , \wRegInTop_6_35[8] , \wRegInTop_6_35[7] , 
        \wRegInTop_6_35[6] , \wRegInTop_6_35[5] , \wRegInTop_6_35[4] , 
        \wRegInTop_6_35[3] , \wRegInTop_6_35[2] , \wRegInTop_6_35[1] , 
        \wRegInTop_6_35[0] }) );
    BHeap_Node_WIDTH32 BHN_6_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_27[0] ), .P_In({\wRegOut_6_27[31] , 
        \wRegOut_6_27[30] , \wRegOut_6_27[29] , \wRegOut_6_27[28] , 
        \wRegOut_6_27[27] , \wRegOut_6_27[26] , \wRegOut_6_27[25] , 
        \wRegOut_6_27[24] , \wRegOut_6_27[23] , \wRegOut_6_27[22] , 
        \wRegOut_6_27[21] , \wRegOut_6_27[20] , \wRegOut_6_27[19] , 
        \wRegOut_6_27[18] , \wRegOut_6_27[17] , \wRegOut_6_27[16] , 
        \wRegOut_6_27[15] , \wRegOut_6_27[14] , \wRegOut_6_27[13] , 
        \wRegOut_6_27[12] , \wRegOut_6_27[11] , \wRegOut_6_27[10] , 
        \wRegOut_6_27[9] , \wRegOut_6_27[8] , \wRegOut_6_27[7] , 
        \wRegOut_6_27[6] , \wRegOut_6_27[5] , \wRegOut_6_27[4] , 
        \wRegOut_6_27[3] , \wRegOut_6_27[2] , \wRegOut_6_27[1] , 
        \wRegOut_6_27[0] }), .P_Out({\wRegInBot_6_27[31] , 
        \wRegInBot_6_27[30] , \wRegInBot_6_27[29] , \wRegInBot_6_27[28] , 
        \wRegInBot_6_27[27] , \wRegInBot_6_27[26] , \wRegInBot_6_27[25] , 
        \wRegInBot_6_27[24] , \wRegInBot_6_27[23] , \wRegInBot_6_27[22] , 
        \wRegInBot_6_27[21] , \wRegInBot_6_27[20] , \wRegInBot_6_27[19] , 
        \wRegInBot_6_27[18] , \wRegInBot_6_27[17] , \wRegInBot_6_27[16] , 
        \wRegInBot_6_27[15] , \wRegInBot_6_27[14] , \wRegInBot_6_27[13] , 
        \wRegInBot_6_27[12] , \wRegInBot_6_27[11] , \wRegInBot_6_27[10] , 
        \wRegInBot_6_27[9] , \wRegInBot_6_27[8] , \wRegInBot_6_27[7] , 
        \wRegInBot_6_27[6] , \wRegInBot_6_27[5] , \wRegInBot_6_27[4] , 
        \wRegInBot_6_27[3] , \wRegInBot_6_27[2] , \wRegInBot_6_27[1] , 
        \wRegInBot_6_27[0] }), .L_WR(\wRegEnTop_7_54[0] ), .L_In({
        \wRegOut_7_54[31] , \wRegOut_7_54[30] , \wRegOut_7_54[29] , 
        \wRegOut_7_54[28] , \wRegOut_7_54[27] , \wRegOut_7_54[26] , 
        \wRegOut_7_54[25] , \wRegOut_7_54[24] , \wRegOut_7_54[23] , 
        \wRegOut_7_54[22] , \wRegOut_7_54[21] , \wRegOut_7_54[20] , 
        \wRegOut_7_54[19] , \wRegOut_7_54[18] , \wRegOut_7_54[17] , 
        \wRegOut_7_54[16] , \wRegOut_7_54[15] , \wRegOut_7_54[14] , 
        \wRegOut_7_54[13] , \wRegOut_7_54[12] , \wRegOut_7_54[11] , 
        \wRegOut_7_54[10] , \wRegOut_7_54[9] , \wRegOut_7_54[8] , 
        \wRegOut_7_54[7] , \wRegOut_7_54[6] , \wRegOut_7_54[5] , 
        \wRegOut_7_54[4] , \wRegOut_7_54[3] , \wRegOut_7_54[2] , 
        \wRegOut_7_54[1] , \wRegOut_7_54[0] }), .L_Out({\wRegInTop_7_54[31] , 
        \wRegInTop_7_54[30] , \wRegInTop_7_54[29] , \wRegInTop_7_54[28] , 
        \wRegInTop_7_54[27] , \wRegInTop_7_54[26] , \wRegInTop_7_54[25] , 
        \wRegInTop_7_54[24] , \wRegInTop_7_54[23] , \wRegInTop_7_54[22] , 
        \wRegInTop_7_54[21] , \wRegInTop_7_54[20] , \wRegInTop_7_54[19] , 
        \wRegInTop_7_54[18] , \wRegInTop_7_54[17] , \wRegInTop_7_54[16] , 
        \wRegInTop_7_54[15] , \wRegInTop_7_54[14] , \wRegInTop_7_54[13] , 
        \wRegInTop_7_54[12] , \wRegInTop_7_54[11] , \wRegInTop_7_54[10] , 
        \wRegInTop_7_54[9] , \wRegInTop_7_54[8] , \wRegInTop_7_54[7] , 
        \wRegInTop_7_54[6] , \wRegInTop_7_54[5] , \wRegInTop_7_54[4] , 
        \wRegInTop_7_54[3] , \wRegInTop_7_54[2] , \wRegInTop_7_54[1] , 
        \wRegInTop_7_54[0] }), .R_WR(\wRegEnTop_7_55[0] ), .R_In({
        \wRegOut_7_55[31] , \wRegOut_7_55[30] , \wRegOut_7_55[29] , 
        \wRegOut_7_55[28] , \wRegOut_7_55[27] , \wRegOut_7_55[26] , 
        \wRegOut_7_55[25] , \wRegOut_7_55[24] , \wRegOut_7_55[23] , 
        \wRegOut_7_55[22] , \wRegOut_7_55[21] , \wRegOut_7_55[20] , 
        \wRegOut_7_55[19] , \wRegOut_7_55[18] , \wRegOut_7_55[17] , 
        \wRegOut_7_55[16] , \wRegOut_7_55[15] , \wRegOut_7_55[14] , 
        \wRegOut_7_55[13] , \wRegOut_7_55[12] , \wRegOut_7_55[11] , 
        \wRegOut_7_55[10] , \wRegOut_7_55[9] , \wRegOut_7_55[8] , 
        \wRegOut_7_55[7] , \wRegOut_7_55[6] , \wRegOut_7_55[5] , 
        \wRegOut_7_55[4] , \wRegOut_7_55[3] , \wRegOut_7_55[2] , 
        \wRegOut_7_55[1] , \wRegOut_7_55[0] }), .R_Out({\wRegInTop_7_55[31] , 
        \wRegInTop_7_55[30] , \wRegInTop_7_55[29] , \wRegInTop_7_55[28] , 
        \wRegInTop_7_55[27] , \wRegInTop_7_55[26] , \wRegInTop_7_55[25] , 
        \wRegInTop_7_55[24] , \wRegInTop_7_55[23] , \wRegInTop_7_55[22] , 
        \wRegInTop_7_55[21] , \wRegInTop_7_55[20] , \wRegInTop_7_55[19] , 
        \wRegInTop_7_55[18] , \wRegInTop_7_55[17] , \wRegInTop_7_55[16] , 
        \wRegInTop_7_55[15] , \wRegInTop_7_55[14] , \wRegInTop_7_55[13] , 
        \wRegInTop_7_55[12] , \wRegInTop_7_55[11] , \wRegInTop_7_55[10] , 
        \wRegInTop_7_55[9] , \wRegInTop_7_55[8] , \wRegInTop_7_55[7] , 
        \wRegInTop_7_55[6] , \wRegInTop_7_55[5] , \wRegInTop_7_55[4] , 
        \wRegInTop_7_55[3] , \wRegInTop_7_55[2] , \wRegInTop_7_55[1] , 
        \wRegInTop_7_55[0] }) );
    BHeap_Node_WIDTH32 BHN_5_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_30[0] ), .P_In({\wRegOut_5_30[31] , 
        \wRegOut_5_30[30] , \wRegOut_5_30[29] , \wRegOut_5_30[28] , 
        \wRegOut_5_30[27] , \wRegOut_5_30[26] , \wRegOut_5_30[25] , 
        \wRegOut_5_30[24] , \wRegOut_5_30[23] , \wRegOut_5_30[22] , 
        \wRegOut_5_30[21] , \wRegOut_5_30[20] , \wRegOut_5_30[19] , 
        \wRegOut_5_30[18] , \wRegOut_5_30[17] , \wRegOut_5_30[16] , 
        \wRegOut_5_30[15] , \wRegOut_5_30[14] , \wRegOut_5_30[13] , 
        \wRegOut_5_30[12] , \wRegOut_5_30[11] , \wRegOut_5_30[10] , 
        \wRegOut_5_30[9] , \wRegOut_5_30[8] , \wRegOut_5_30[7] , 
        \wRegOut_5_30[6] , \wRegOut_5_30[5] , \wRegOut_5_30[4] , 
        \wRegOut_5_30[3] , \wRegOut_5_30[2] , \wRegOut_5_30[1] , 
        \wRegOut_5_30[0] }), .P_Out({\wRegInBot_5_30[31] , 
        \wRegInBot_5_30[30] , \wRegInBot_5_30[29] , \wRegInBot_5_30[28] , 
        \wRegInBot_5_30[27] , \wRegInBot_5_30[26] , \wRegInBot_5_30[25] , 
        \wRegInBot_5_30[24] , \wRegInBot_5_30[23] , \wRegInBot_5_30[22] , 
        \wRegInBot_5_30[21] , \wRegInBot_5_30[20] , \wRegInBot_5_30[19] , 
        \wRegInBot_5_30[18] , \wRegInBot_5_30[17] , \wRegInBot_5_30[16] , 
        \wRegInBot_5_30[15] , \wRegInBot_5_30[14] , \wRegInBot_5_30[13] , 
        \wRegInBot_5_30[12] , \wRegInBot_5_30[11] , \wRegInBot_5_30[10] , 
        \wRegInBot_5_30[9] , \wRegInBot_5_30[8] , \wRegInBot_5_30[7] , 
        \wRegInBot_5_30[6] , \wRegInBot_5_30[5] , \wRegInBot_5_30[4] , 
        \wRegInBot_5_30[3] , \wRegInBot_5_30[2] , \wRegInBot_5_30[1] , 
        \wRegInBot_5_30[0] }), .L_WR(\wRegEnTop_6_60[0] ), .L_In({
        \wRegOut_6_60[31] , \wRegOut_6_60[30] , \wRegOut_6_60[29] , 
        \wRegOut_6_60[28] , \wRegOut_6_60[27] , \wRegOut_6_60[26] , 
        \wRegOut_6_60[25] , \wRegOut_6_60[24] , \wRegOut_6_60[23] , 
        \wRegOut_6_60[22] , \wRegOut_6_60[21] , \wRegOut_6_60[20] , 
        \wRegOut_6_60[19] , \wRegOut_6_60[18] , \wRegOut_6_60[17] , 
        \wRegOut_6_60[16] , \wRegOut_6_60[15] , \wRegOut_6_60[14] , 
        \wRegOut_6_60[13] , \wRegOut_6_60[12] , \wRegOut_6_60[11] , 
        \wRegOut_6_60[10] , \wRegOut_6_60[9] , \wRegOut_6_60[8] , 
        \wRegOut_6_60[7] , \wRegOut_6_60[6] , \wRegOut_6_60[5] , 
        \wRegOut_6_60[4] , \wRegOut_6_60[3] , \wRegOut_6_60[2] , 
        \wRegOut_6_60[1] , \wRegOut_6_60[0] }), .L_Out({\wRegInTop_6_60[31] , 
        \wRegInTop_6_60[30] , \wRegInTop_6_60[29] , \wRegInTop_6_60[28] , 
        \wRegInTop_6_60[27] , \wRegInTop_6_60[26] , \wRegInTop_6_60[25] , 
        \wRegInTop_6_60[24] , \wRegInTop_6_60[23] , \wRegInTop_6_60[22] , 
        \wRegInTop_6_60[21] , \wRegInTop_6_60[20] , \wRegInTop_6_60[19] , 
        \wRegInTop_6_60[18] , \wRegInTop_6_60[17] , \wRegInTop_6_60[16] , 
        \wRegInTop_6_60[15] , \wRegInTop_6_60[14] , \wRegInTop_6_60[13] , 
        \wRegInTop_6_60[12] , \wRegInTop_6_60[11] , \wRegInTop_6_60[10] , 
        \wRegInTop_6_60[9] , \wRegInTop_6_60[8] , \wRegInTop_6_60[7] , 
        \wRegInTop_6_60[6] , \wRegInTop_6_60[5] , \wRegInTop_6_60[4] , 
        \wRegInTop_6_60[3] , \wRegInTop_6_60[2] , \wRegInTop_6_60[1] , 
        \wRegInTop_6_60[0] }), .R_WR(\wRegEnTop_6_61[0] ), .R_In({
        \wRegOut_6_61[31] , \wRegOut_6_61[30] , \wRegOut_6_61[29] , 
        \wRegOut_6_61[28] , \wRegOut_6_61[27] , \wRegOut_6_61[26] , 
        \wRegOut_6_61[25] , \wRegOut_6_61[24] , \wRegOut_6_61[23] , 
        \wRegOut_6_61[22] , \wRegOut_6_61[21] , \wRegOut_6_61[20] , 
        \wRegOut_6_61[19] , \wRegOut_6_61[18] , \wRegOut_6_61[17] , 
        \wRegOut_6_61[16] , \wRegOut_6_61[15] , \wRegOut_6_61[14] , 
        \wRegOut_6_61[13] , \wRegOut_6_61[12] , \wRegOut_6_61[11] , 
        \wRegOut_6_61[10] , \wRegOut_6_61[9] , \wRegOut_6_61[8] , 
        \wRegOut_6_61[7] , \wRegOut_6_61[6] , \wRegOut_6_61[5] , 
        \wRegOut_6_61[4] , \wRegOut_6_61[3] , \wRegOut_6_61[2] , 
        \wRegOut_6_61[1] , \wRegOut_6_61[0] }), .R_Out({\wRegInTop_6_61[31] , 
        \wRegInTop_6_61[30] , \wRegInTop_6_61[29] , \wRegInTop_6_61[28] , 
        \wRegInTop_6_61[27] , \wRegInTop_6_61[26] , \wRegInTop_6_61[25] , 
        \wRegInTop_6_61[24] , \wRegInTop_6_61[23] , \wRegInTop_6_61[22] , 
        \wRegInTop_6_61[21] , \wRegInTop_6_61[20] , \wRegInTop_6_61[19] , 
        \wRegInTop_6_61[18] , \wRegInTop_6_61[17] , \wRegInTop_6_61[16] , 
        \wRegInTop_6_61[15] , \wRegInTop_6_61[14] , \wRegInTop_6_61[13] , 
        \wRegInTop_6_61[12] , \wRegInTop_6_61[11] , \wRegInTop_6_61[10] , 
        \wRegInTop_6_61[9] , \wRegInTop_6_61[8] , \wRegInTop_6_61[7] , 
        \wRegInTop_6_61[6] , \wRegInTop_6_61[5] , \wRegInTop_6_61[4] , 
        \wRegInTop_6_61[3] , \wRegInTop_6_61[2] , \wRegInTop_6_61[1] , 
        \wRegInTop_6_61[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink20[31] , \ScanLink20[30] , \ScanLink20[29] , 
        \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , \ScanLink20[25] , 
        \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , \ScanLink20[21] , 
        \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , \ScanLink20[17] , 
        \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , \ScanLink20[13] , 
        \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , \ScanLink20[9] , 
        \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , \ScanLink20[5] , 
        \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , \ScanLink20[1] , 
        \ScanLink20[0] }), .ScanOut({\ScanLink19[31] , \ScanLink19[30] , 
        \ScanLink19[29] , \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , 
        \ScanLink19[25] , \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , 
        \ScanLink19[21] , \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , 
        \ScanLink19[17] , \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , 
        \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , 
        \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , 
        \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , 
        \ScanLink19[1] , \ScanLink19[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_4[31] , \wRegOut_4_4[30] , \wRegOut_4_4[29] , 
        \wRegOut_4_4[28] , \wRegOut_4_4[27] , \wRegOut_4_4[26] , 
        \wRegOut_4_4[25] , \wRegOut_4_4[24] , \wRegOut_4_4[23] , 
        \wRegOut_4_4[22] , \wRegOut_4_4[21] , \wRegOut_4_4[20] , 
        \wRegOut_4_4[19] , \wRegOut_4_4[18] , \wRegOut_4_4[17] , 
        \wRegOut_4_4[16] , \wRegOut_4_4[15] , \wRegOut_4_4[14] , 
        \wRegOut_4_4[13] , \wRegOut_4_4[12] , \wRegOut_4_4[11] , 
        \wRegOut_4_4[10] , \wRegOut_4_4[9] , \wRegOut_4_4[8] , 
        \wRegOut_4_4[7] , \wRegOut_4_4[6] , \wRegOut_4_4[5] , \wRegOut_4_4[4] , 
        \wRegOut_4_4[3] , \wRegOut_4_4[2] , \wRegOut_4_4[1] , \wRegOut_4_4[0] 
        }), .Enable1(\wRegEnTop_4_4[0] ), .Enable2(\wRegEnBot_4_4[0] ), .In1({
        \wRegInTop_4_4[31] , \wRegInTop_4_4[30] , \wRegInTop_4_4[29] , 
        \wRegInTop_4_4[28] , \wRegInTop_4_4[27] , \wRegInTop_4_4[26] , 
        \wRegInTop_4_4[25] , \wRegInTop_4_4[24] , \wRegInTop_4_4[23] , 
        \wRegInTop_4_4[22] , \wRegInTop_4_4[21] , \wRegInTop_4_4[20] , 
        \wRegInTop_4_4[19] , \wRegInTop_4_4[18] , \wRegInTop_4_4[17] , 
        \wRegInTop_4_4[16] , \wRegInTop_4_4[15] , \wRegInTop_4_4[14] , 
        \wRegInTop_4_4[13] , \wRegInTop_4_4[12] , \wRegInTop_4_4[11] , 
        \wRegInTop_4_4[10] , \wRegInTop_4_4[9] , \wRegInTop_4_4[8] , 
        \wRegInTop_4_4[7] , \wRegInTop_4_4[6] , \wRegInTop_4_4[5] , 
        \wRegInTop_4_4[4] , \wRegInTop_4_4[3] , \wRegInTop_4_4[2] , 
        \wRegInTop_4_4[1] , \wRegInTop_4_4[0] }), .In2({\wRegInBot_4_4[31] , 
        \wRegInBot_4_4[30] , \wRegInBot_4_4[29] , \wRegInBot_4_4[28] , 
        \wRegInBot_4_4[27] , \wRegInBot_4_4[26] , \wRegInBot_4_4[25] , 
        \wRegInBot_4_4[24] , \wRegInBot_4_4[23] , \wRegInBot_4_4[22] , 
        \wRegInBot_4_4[21] , \wRegInBot_4_4[20] , \wRegInBot_4_4[19] , 
        \wRegInBot_4_4[18] , \wRegInBot_4_4[17] , \wRegInBot_4_4[16] , 
        \wRegInBot_4_4[15] , \wRegInBot_4_4[14] , \wRegInBot_4_4[13] , 
        \wRegInBot_4_4[12] , \wRegInBot_4_4[11] , \wRegInBot_4_4[10] , 
        \wRegInBot_4_4[9] , \wRegInBot_4_4[8] , \wRegInBot_4_4[7] , 
        \wRegInBot_4_4[6] , \wRegInBot_4_4[5] , \wRegInBot_4_4[4] , 
        \wRegInBot_4_4[3] , \wRegInBot_4_4[2] , \wRegInBot_4_4[1] , 
        \wRegInBot_4_4[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink43[31] , \ScanLink43[30] , \ScanLink43[29] , 
        \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , \ScanLink43[25] , 
        \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , \ScanLink43[21] , 
        \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , \ScanLink43[17] , 
        \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , \ScanLink43[13] , 
        \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , \ScanLink43[9] , 
        \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , \ScanLink43[5] , 
        \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , \ScanLink43[1] , 
        \ScanLink43[0] }), .ScanOut({\ScanLink42[31] , \ScanLink42[30] , 
        \ScanLink42[29] , \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , 
        \ScanLink42[25] , \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , 
        \ScanLink42[21] , \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , 
        \ScanLink42[17] , \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , 
        \ScanLink42[13] , \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , 
        \ScanLink42[9] , \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , 
        \ScanLink42[5] , \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , 
        \ScanLink42[1] , \ScanLink42[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_11[31] , \wRegOut_5_11[30] , 
        \wRegOut_5_11[29] , \wRegOut_5_11[28] , \wRegOut_5_11[27] , 
        \wRegOut_5_11[26] , \wRegOut_5_11[25] , \wRegOut_5_11[24] , 
        \wRegOut_5_11[23] , \wRegOut_5_11[22] , \wRegOut_5_11[21] , 
        \wRegOut_5_11[20] , \wRegOut_5_11[19] , \wRegOut_5_11[18] , 
        \wRegOut_5_11[17] , \wRegOut_5_11[16] , \wRegOut_5_11[15] , 
        \wRegOut_5_11[14] , \wRegOut_5_11[13] , \wRegOut_5_11[12] , 
        \wRegOut_5_11[11] , \wRegOut_5_11[10] , \wRegOut_5_11[9] , 
        \wRegOut_5_11[8] , \wRegOut_5_11[7] , \wRegOut_5_11[6] , 
        \wRegOut_5_11[5] , \wRegOut_5_11[4] , \wRegOut_5_11[3] , 
        \wRegOut_5_11[2] , \wRegOut_5_11[1] , \wRegOut_5_11[0] }), .Enable1(
        \wRegEnTop_5_11[0] ), .Enable2(\wRegEnBot_5_11[0] ), .In1({
        \wRegInTop_5_11[31] , \wRegInTop_5_11[30] , \wRegInTop_5_11[29] , 
        \wRegInTop_5_11[28] , \wRegInTop_5_11[27] , \wRegInTop_5_11[26] , 
        \wRegInTop_5_11[25] , \wRegInTop_5_11[24] , \wRegInTop_5_11[23] , 
        \wRegInTop_5_11[22] , \wRegInTop_5_11[21] , \wRegInTop_5_11[20] , 
        \wRegInTop_5_11[19] , \wRegInTop_5_11[18] , \wRegInTop_5_11[17] , 
        \wRegInTop_5_11[16] , \wRegInTop_5_11[15] , \wRegInTop_5_11[14] , 
        \wRegInTop_5_11[13] , \wRegInTop_5_11[12] , \wRegInTop_5_11[11] , 
        \wRegInTop_5_11[10] , \wRegInTop_5_11[9] , \wRegInTop_5_11[8] , 
        \wRegInTop_5_11[7] , \wRegInTop_5_11[6] , \wRegInTop_5_11[5] , 
        \wRegInTop_5_11[4] , \wRegInTop_5_11[3] , \wRegInTop_5_11[2] , 
        \wRegInTop_5_11[1] , \wRegInTop_5_11[0] }), .In2({\wRegInBot_5_11[31] , 
        \wRegInBot_5_11[30] , \wRegInBot_5_11[29] , \wRegInBot_5_11[28] , 
        \wRegInBot_5_11[27] , \wRegInBot_5_11[26] , \wRegInBot_5_11[25] , 
        \wRegInBot_5_11[24] , \wRegInBot_5_11[23] , \wRegInBot_5_11[22] , 
        \wRegInBot_5_11[21] , \wRegInBot_5_11[20] , \wRegInBot_5_11[19] , 
        \wRegInBot_5_11[18] , \wRegInBot_5_11[17] , \wRegInBot_5_11[16] , 
        \wRegInBot_5_11[15] , \wRegInBot_5_11[14] , \wRegInBot_5_11[13] , 
        \wRegInBot_5_11[12] , \wRegInBot_5_11[11] , \wRegInBot_5_11[10] , 
        \wRegInBot_5_11[9] , \wRegInBot_5_11[8] , \wRegInBot_5_11[7] , 
        \wRegInBot_5_11[6] , \wRegInBot_5_11[5] , \wRegInBot_5_11[4] , 
        \wRegInBot_5_11[3] , \wRegInBot_5_11[2] , \wRegInBot_5_11[1] , 
        \wRegInBot_5_11[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_24 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink56[31] , \ScanLink56[30] , \ScanLink56[29] , 
        \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , \ScanLink56[25] , 
        \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , \ScanLink56[21] , 
        \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , \ScanLink56[17] , 
        \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , \ScanLink56[13] , 
        \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , \ScanLink56[9] , 
        \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , \ScanLink56[5] , 
        \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , \ScanLink56[1] , 
        \ScanLink56[0] }), .ScanOut({\ScanLink55[31] , \ScanLink55[30] , 
        \ScanLink55[29] , \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , 
        \ScanLink55[25] , \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , 
        \ScanLink55[21] , \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , 
        \ScanLink55[17] , \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , 
        \ScanLink55[13] , \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , 
        \ScanLink55[9] , \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , 
        \ScanLink55[5] , \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , 
        \ScanLink55[1] , \ScanLink55[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_24[31] , \wRegOut_5_24[30] , 
        \wRegOut_5_24[29] , \wRegOut_5_24[28] , \wRegOut_5_24[27] , 
        \wRegOut_5_24[26] , \wRegOut_5_24[25] , \wRegOut_5_24[24] , 
        \wRegOut_5_24[23] , \wRegOut_5_24[22] , \wRegOut_5_24[21] , 
        \wRegOut_5_24[20] , \wRegOut_5_24[19] , \wRegOut_5_24[18] , 
        \wRegOut_5_24[17] , \wRegOut_5_24[16] , \wRegOut_5_24[15] , 
        \wRegOut_5_24[14] , \wRegOut_5_24[13] , \wRegOut_5_24[12] , 
        \wRegOut_5_24[11] , \wRegOut_5_24[10] , \wRegOut_5_24[9] , 
        \wRegOut_5_24[8] , \wRegOut_5_24[7] , \wRegOut_5_24[6] , 
        \wRegOut_5_24[5] , \wRegOut_5_24[4] , \wRegOut_5_24[3] , 
        \wRegOut_5_24[2] , \wRegOut_5_24[1] , \wRegOut_5_24[0] }), .Enable1(
        \wRegEnTop_5_24[0] ), .Enable2(\wRegEnBot_5_24[0] ), .In1({
        \wRegInTop_5_24[31] , \wRegInTop_5_24[30] , \wRegInTop_5_24[29] , 
        \wRegInTop_5_24[28] , \wRegInTop_5_24[27] , \wRegInTop_5_24[26] , 
        \wRegInTop_5_24[25] , \wRegInTop_5_24[24] , \wRegInTop_5_24[23] , 
        \wRegInTop_5_24[22] , \wRegInTop_5_24[21] , \wRegInTop_5_24[20] , 
        \wRegInTop_5_24[19] , \wRegInTop_5_24[18] , \wRegInTop_5_24[17] , 
        \wRegInTop_5_24[16] , \wRegInTop_5_24[15] , \wRegInTop_5_24[14] , 
        \wRegInTop_5_24[13] , \wRegInTop_5_24[12] , \wRegInTop_5_24[11] , 
        \wRegInTop_5_24[10] , \wRegInTop_5_24[9] , \wRegInTop_5_24[8] , 
        \wRegInTop_5_24[7] , \wRegInTop_5_24[6] , \wRegInTop_5_24[5] , 
        \wRegInTop_5_24[4] , \wRegInTop_5_24[3] , \wRegInTop_5_24[2] , 
        \wRegInTop_5_24[1] , \wRegInTop_5_24[0] }), .In2({\wRegInBot_5_24[31] , 
        \wRegInBot_5_24[30] , \wRegInBot_5_24[29] , \wRegInBot_5_24[28] , 
        \wRegInBot_5_24[27] , \wRegInBot_5_24[26] , \wRegInBot_5_24[25] , 
        \wRegInBot_5_24[24] , \wRegInBot_5_24[23] , \wRegInBot_5_24[22] , 
        \wRegInBot_5_24[21] , \wRegInBot_5_24[20] , \wRegInBot_5_24[19] , 
        \wRegInBot_5_24[18] , \wRegInBot_5_24[17] , \wRegInBot_5_24[16] , 
        \wRegInBot_5_24[15] , \wRegInBot_5_24[14] , \wRegInBot_5_24[13] , 
        \wRegInBot_5_24[12] , \wRegInBot_5_24[11] , \wRegInBot_5_24[10] , 
        \wRegInBot_5_24[9] , \wRegInBot_5_24[8] , \wRegInBot_5_24[7] , 
        \wRegInBot_5_24[6] , \wRegInBot_5_24[5] , \wRegInBot_5_24[4] , 
        \wRegInBot_5_24[3] , \wRegInBot_5_24[2] , \wRegInBot_5_24[1] , 
        \wRegInBot_5_24[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink65[31] , \ScanLink65[30] , \ScanLink65[29] , 
        \ScanLink65[28] , \ScanLink65[27] , \ScanLink65[26] , \ScanLink65[25] , 
        \ScanLink65[24] , \ScanLink65[23] , \ScanLink65[22] , \ScanLink65[21] , 
        \ScanLink65[20] , \ScanLink65[19] , \ScanLink65[18] , \ScanLink65[17] , 
        \ScanLink65[16] , \ScanLink65[15] , \ScanLink65[14] , \ScanLink65[13] , 
        \ScanLink65[12] , \ScanLink65[11] , \ScanLink65[10] , \ScanLink65[9] , 
        \ScanLink65[8] , \ScanLink65[7] , \ScanLink65[6] , \ScanLink65[5] , 
        \ScanLink65[4] , \ScanLink65[3] , \ScanLink65[2] , \ScanLink65[1] , 
        \ScanLink65[0] }), .ScanOut({\ScanLink64[31] , \ScanLink64[30] , 
        \ScanLink64[29] , \ScanLink64[28] , \ScanLink64[27] , \ScanLink64[26] , 
        \ScanLink64[25] , \ScanLink64[24] , \ScanLink64[23] , \ScanLink64[22] , 
        \ScanLink64[21] , \ScanLink64[20] , \ScanLink64[19] , \ScanLink64[18] , 
        \ScanLink64[17] , \ScanLink64[16] , \ScanLink64[15] , \ScanLink64[14] , 
        \ScanLink64[13] , \ScanLink64[12] , \ScanLink64[11] , \ScanLink64[10] , 
        \ScanLink64[9] , \ScanLink64[8] , \ScanLink64[7] , \ScanLink64[6] , 
        \ScanLink64[5] , \ScanLink64[4] , \ScanLink64[3] , \ScanLink64[2] , 
        \ScanLink64[1] , \ScanLink64[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_1[31] , \wRegOut_6_1[30] , \wRegOut_6_1[29] , 
        \wRegOut_6_1[28] , \wRegOut_6_1[27] , \wRegOut_6_1[26] , 
        \wRegOut_6_1[25] , \wRegOut_6_1[24] , \wRegOut_6_1[23] , 
        \wRegOut_6_1[22] , \wRegOut_6_1[21] , \wRegOut_6_1[20] , 
        \wRegOut_6_1[19] , \wRegOut_6_1[18] , \wRegOut_6_1[17] , 
        \wRegOut_6_1[16] , \wRegOut_6_1[15] , \wRegOut_6_1[14] , 
        \wRegOut_6_1[13] , \wRegOut_6_1[12] , \wRegOut_6_1[11] , 
        \wRegOut_6_1[10] , \wRegOut_6_1[9] , \wRegOut_6_1[8] , 
        \wRegOut_6_1[7] , \wRegOut_6_1[6] , \wRegOut_6_1[5] , \wRegOut_6_1[4] , 
        \wRegOut_6_1[3] , \wRegOut_6_1[2] , \wRegOut_6_1[1] , \wRegOut_6_1[0] 
        }), .Enable1(\wRegEnTop_6_1[0] ), .Enable2(\wRegEnBot_6_1[0] ), .In1({
        \wRegInTop_6_1[31] , \wRegInTop_6_1[30] , \wRegInTop_6_1[29] , 
        \wRegInTop_6_1[28] , \wRegInTop_6_1[27] , \wRegInTop_6_1[26] , 
        \wRegInTop_6_1[25] , \wRegInTop_6_1[24] , \wRegInTop_6_1[23] , 
        \wRegInTop_6_1[22] , \wRegInTop_6_1[21] , \wRegInTop_6_1[20] , 
        \wRegInTop_6_1[19] , \wRegInTop_6_1[18] , \wRegInTop_6_1[17] , 
        \wRegInTop_6_1[16] , \wRegInTop_6_1[15] , \wRegInTop_6_1[14] , 
        \wRegInTop_6_1[13] , \wRegInTop_6_1[12] , \wRegInTop_6_1[11] , 
        \wRegInTop_6_1[10] , \wRegInTop_6_1[9] , \wRegInTop_6_1[8] , 
        \wRegInTop_6_1[7] , \wRegInTop_6_1[6] , \wRegInTop_6_1[5] , 
        \wRegInTop_6_1[4] , \wRegInTop_6_1[3] , \wRegInTop_6_1[2] , 
        \wRegInTop_6_1[1] , \wRegInTop_6_1[0] }), .In2({\wRegInBot_6_1[31] , 
        \wRegInBot_6_1[30] , \wRegInBot_6_1[29] , \wRegInBot_6_1[28] , 
        \wRegInBot_6_1[27] , \wRegInBot_6_1[26] , \wRegInBot_6_1[25] , 
        \wRegInBot_6_1[24] , \wRegInBot_6_1[23] , \wRegInBot_6_1[22] , 
        \wRegInBot_6_1[21] , \wRegInBot_6_1[20] , \wRegInBot_6_1[19] , 
        \wRegInBot_6_1[18] , \wRegInBot_6_1[17] , \wRegInBot_6_1[16] , 
        \wRegInBot_6_1[15] , \wRegInBot_6_1[14] , \wRegInBot_6_1[13] , 
        \wRegInBot_6_1[12] , \wRegInBot_6_1[11] , \wRegInBot_6_1[10] , 
        \wRegInBot_6_1[9] , \wRegInBot_6_1[8] , \wRegInBot_6_1[7] , 
        \wRegInBot_6_1[6] , \wRegInBot_6_1[5] , \wRegInBot_6_1[4] , 
        \wRegInBot_6_1[3] , \wRegInBot_6_1[2] , \wRegInBot_6_1[1] , 
        \wRegInBot_6_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_33 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink97[31] , \ScanLink97[30] , \ScanLink97[29] , 
        \ScanLink97[28] , \ScanLink97[27] , \ScanLink97[26] , \ScanLink97[25] , 
        \ScanLink97[24] , \ScanLink97[23] , \ScanLink97[22] , \ScanLink97[21] , 
        \ScanLink97[20] , \ScanLink97[19] , \ScanLink97[18] , \ScanLink97[17] , 
        \ScanLink97[16] , \ScanLink97[15] , \ScanLink97[14] , \ScanLink97[13] , 
        \ScanLink97[12] , \ScanLink97[11] , \ScanLink97[10] , \ScanLink97[9] , 
        \ScanLink97[8] , \ScanLink97[7] , \ScanLink97[6] , \ScanLink97[5] , 
        \ScanLink97[4] , \ScanLink97[3] , \ScanLink97[2] , \ScanLink97[1] , 
        \ScanLink97[0] }), .ScanOut({\ScanLink96[31] , \ScanLink96[30] , 
        \ScanLink96[29] , \ScanLink96[28] , \ScanLink96[27] , \ScanLink96[26] , 
        \ScanLink96[25] , \ScanLink96[24] , \ScanLink96[23] , \ScanLink96[22] , 
        \ScanLink96[21] , \ScanLink96[20] , \ScanLink96[19] , \ScanLink96[18] , 
        \ScanLink96[17] , \ScanLink96[16] , \ScanLink96[15] , \ScanLink96[14] , 
        \ScanLink96[13] , \ScanLink96[12] , \ScanLink96[11] , \ScanLink96[10] , 
        \ScanLink96[9] , \ScanLink96[8] , \ScanLink96[7] , \ScanLink96[6] , 
        \ScanLink96[5] , \ScanLink96[4] , \ScanLink96[3] , \ScanLink96[2] , 
        \ScanLink96[1] , \ScanLink96[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_33[31] , \wRegOut_6_33[30] , 
        \wRegOut_6_33[29] , \wRegOut_6_33[28] , \wRegOut_6_33[27] , 
        \wRegOut_6_33[26] , \wRegOut_6_33[25] , \wRegOut_6_33[24] , 
        \wRegOut_6_33[23] , \wRegOut_6_33[22] , \wRegOut_6_33[21] , 
        \wRegOut_6_33[20] , \wRegOut_6_33[19] , \wRegOut_6_33[18] , 
        \wRegOut_6_33[17] , \wRegOut_6_33[16] , \wRegOut_6_33[15] , 
        \wRegOut_6_33[14] , \wRegOut_6_33[13] , \wRegOut_6_33[12] , 
        \wRegOut_6_33[11] , \wRegOut_6_33[10] , \wRegOut_6_33[9] , 
        \wRegOut_6_33[8] , \wRegOut_6_33[7] , \wRegOut_6_33[6] , 
        \wRegOut_6_33[5] , \wRegOut_6_33[4] , \wRegOut_6_33[3] , 
        \wRegOut_6_33[2] , \wRegOut_6_33[1] , \wRegOut_6_33[0] }), .Enable1(
        \wRegEnTop_6_33[0] ), .Enable2(\wRegEnBot_6_33[0] ), .In1({
        \wRegInTop_6_33[31] , \wRegInTop_6_33[30] , \wRegInTop_6_33[29] , 
        \wRegInTop_6_33[28] , \wRegInTop_6_33[27] , \wRegInTop_6_33[26] , 
        \wRegInTop_6_33[25] , \wRegInTop_6_33[24] , \wRegInTop_6_33[23] , 
        \wRegInTop_6_33[22] , \wRegInTop_6_33[21] , \wRegInTop_6_33[20] , 
        \wRegInTop_6_33[19] , \wRegInTop_6_33[18] , \wRegInTop_6_33[17] , 
        \wRegInTop_6_33[16] , \wRegInTop_6_33[15] , \wRegInTop_6_33[14] , 
        \wRegInTop_6_33[13] , \wRegInTop_6_33[12] , \wRegInTop_6_33[11] , 
        \wRegInTop_6_33[10] , \wRegInTop_6_33[9] , \wRegInTop_6_33[8] , 
        \wRegInTop_6_33[7] , \wRegInTop_6_33[6] , \wRegInTop_6_33[5] , 
        \wRegInTop_6_33[4] , \wRegInTop_6_33[3] , \wRegInTop_6_33[2] , 
        \wRegInTop_6_33[1] , \wRegInTop_6_33[0] }), .In2({\wRegInBot_6_33[31] , 
        \wRegInBot_6_33[30] , \wRegInBot_6_33[29] , \wRegInBot_6_33[28] , 
        \wRegInBot_6_33[27] , \wRegInBot_6_33[26] , \wRegInBot_6_33[25] , 
        \wRegInBot_6_33[24] , \wRegInBot_6_33[23] , \wRegInBot_6_33[22] , 
        \wRegInBot_6_33[21] , \wRegInBot_6_33[20] , \wRegInBot_6_33[19] , 
        \wRegInBot_6_33[18] , \wRegInBot_6_33[17] , \wRegInBot_6_33[16] , 
        \wRegInBot_6_33[15] , \wRegInBot_6_33[14] , \wRegInBot_6_33[13] , 
        \wRegInBot_6_33[12] , \wRegInBot_6_33[11] , \wRegInBot_6_33[10] , 
        \wRegInBot_6_33[9] , \wRegInBot_6_33[8] , \wRegInBot_6_33[7] , 
        \wRegInBot_6_33[6] , \wRegInBot_6_33[5] , \wRegInBot_6_33[4] , 
        \wRegInBot_6_33[3] , \wRegInBot_6_33[2] , \wRegInBot_6_33[1] , 
        \wRegInBot_6_33[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_46 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink110[31] , \ScanLink110[30] , \ScanLink110[29] , 
        \ScanLink110[28] , \ScanLink110[27] , \ScanLink110[26] , 
        \ScanLink110[25] , \ScanLink110[24] , \ScanLink110[23] , 
        \ScanLink110[22] , \ScanLink110[21] , \ScanLink110[20] , 
        \ScanLink110[19] , \ScanLink110[18] , \ScanLink110[17] , 
        \ScanLink110[16] , \ScanLink110[15] , \ScanLink110[14] , 
        \ScanLink110[13] , \ScanLink110[12] , \ScanLink110[11] , 
        \ScanLink110[10] , \ScanLink110[9] , \ScanLink110[8] , 
        \ScanLink110[7] , \ScanLink110[6] , \ScanLink110[5] , \ScanLink110[4] , 
        \ScanLink110[3] , \ScanLink110[2] , \ScanLink110[1] , \ScanLink110[0] 
        }), .ScanOut({\ScanLink109[31] , \ScanLink109[30] , \ScanLink109[29] , 
        \ScanLink109[28] , \ScanLink109[27] , \ScanLink109[26] , 
        \ScanLink109[25] , \ScanLink109[24] , \ScanLink109[23] , 
        \ScanLink109[22] , \ScanLink109[21] , \ScanLink109[20] , 
        \ScanLink109[19] , \ScanLink109[18] , \ScanLink109[17] , 
        \ScanLink109[16] , \ScanLink109[15] , \ScanLink109[14] , 
        \ScanLink109[13] , \ScanLink109[12] , \ScanLink109[11] , 
        \ScanLink109[10] , \ScanLink109[9] , \ScanLink109[8] , 
        \ScanLink109[7] , \ScanLink109[6] , \ScanLink109[5] , \ScanLink109[4] , 
        \ScanLink109[3] , \ScanLink109[2] , \ScanLink109[1] , \ScanLink109[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_46[31] , 
        \wRegOut_6_46[30] , \wRegOut_6_46[29] , \wRegOut_6_46[28] , 
        \wRegOut_6_46[27] , \wRegOut_6_46[26] , \wRegOut_6_46[25] , 
        \wRegOut_6_46[24] , \wRegOut_6_46[23] , \wRegOut_6_46[22] , 
        \wRegOut_6_46[21] , \wRegOut_6_46[20] , \wRegOut_6_46[19] , 
        \wRegOut_6_46[18] , \wRegOut_6_46[17] , \wRegOut_6_46[16] , 
        \wRegOut_6_46[15] , \wRegOut_6_46[14] , \wRegOut_6_46[13] , 
        \wRegOut_6_46[12] , \wRegOut_6_46[11] , \wRegOut_6_46[10] , 
        \wRegOut_6_46[9] , \wRegOut_6_46[8] , \wRegOut_6_46[7] , 
        \wRegOut_6_46[6] , \wRegOut_6_46[5] , \wRegOut_6_46[4] , 
        \wRegOut_6_46[3] , \wRegOut_6_46[2] , \wRegOut_6_46[1] , 
        \wRegOut_6_46[0] }), .Enable1(\wRegEnTop_6_46[0] ), .Enable2(
        \wRegEnBot_6_46[0] ), .In1({\wRegInTop_6_46[31] , \wRegInTop_6_46[30] , 
        \wRegInTop_6_46[29] , \wRegInTop_6_46[28] , \wRegInTop_6_46[27] , 
        \wRegInTop_6_46[26] , \wRegInTop_6_46[25] , \wRegInTop_6_46[24] , 
        \wRegInTop_6_46[23] , \wRegInTop_6_46[22] , \wRegInTop_6_46[21] , 
        \wRegInTop_6_46[20] , \wRegInTop_6_46[19] , \wRegInTop_6_46[18] , 
        \wRegInTop_6_46[17] , \wRegInTop_6_46[16] , \wRegInTop_6_46[15] , 
        \wRegInTop_6_46[14] , \wRegInTop_6_46[13] , \wRegInTop_6_46[12] , 
        \wRegInTop_6_46[11] , \wRegInTop_6_46[10] , \wRegInTop_6_46[9] , 
        \wRegInTop_6_46[8] , \wRegInTop_6_46[7] , \wRegInTop_6_46[6] , 
        \wRegInTop_6_46[5] , \wRegInTop_6_46[4] , \wRegInTop_6_46[3] , 
        \wRegInTop_6_46[2] , \wRegInTop_6_46[1] , \wRegInTop_6_46[0] }), .In2(
        {\wRegInBot_6_46[31] , \wRegInBot_6_46[30] , \wRegInBot_6_46[29] , 
        \wRegInBot_6_46[28] , \wRegInBot_6_46[27] , \wRegInBot_6_46[26] , 
        \wRegInBot_6_46[25] , \wRegInBot_6_46[24] , \wRegInBot_6_46[23] , 
        \wRegInBot_6_46[22] , \wRegInBot_6_46[21] , \wRegInBot_6_46[20] , 
        \wRegInBot_6_46[19] , \wRegInBot_6_46[18] , \wRegInBot_6_46[17] , 
        \wRegInBot_6_46[16] , \wRegInBot_6_46[15] , \wRegInBot_6_46[14] , 
        \wRegInBot_6_46[13] , \wRegInBot_6_46[12] , \wRegInBot_6_46[11] , 
        \wRegInBot_6_46[10] , \wRegInBot_6_46[9] , \wRegInBot_6_46[8] , 
        \wRegInBot_6_46[7] , \wRegInBot_6_46[6] , \wRegInBot_6_46[5] , 
        \wRegInBot_6_46[4] , \wRegInBot_6_46[3] , \wRegInBot_6_46[2] , 
        \wRegInBot_6_46[1] , \wRegInBot_6_46[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_61 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink125[31] , \ScanLink125[30] , \ScanLink125[29] , 
        \ScanLink125[28] , \ScanLink125[27] , \ScanLink125[26] , 
        \ScanLink125[25] , \ScanLink125[24] , \ScanLink125[23] , 
        \ScanLink125[22] , \ScanLink125[21] , \ScanLink125[20] , 
        \ScanLink125[19] , \ScanLink125[18] , \ScanLink125[17] , 
        \ScanLink125[16] , \ScanLink125[15] , \ScanLink125[14] , 
        \ScanLink125[13] , \ScanLink125[12] , \ScanLink125[11] , 
        \ScanLink125[10] , \ScanLink125[9] , \ScanLink125[8] , 
        \ScanLink125[7] , \ScanLink125[6] , \ScanLink125[5] , \ScanLink125[4] , 
        \ScanLink125[3] , \ScanLink125[2] , \ScanLink125[1] , \ScanLink125[0] 
        }), .ScanOut({\ScanLink124[31] , \ScanLink124[30] , \ScanLink124[29] , 
        \ScanLink124[28] , \ScanLink124[27] , \ScanLink124[26] , 
        \ScanLink124[25] , \ScanLink124[24] , \ScanLink124[23] , 
        \ScanLink124[22] , \ScanLink124[21] , \ScanLink124[20] , 
        \ScanLink124[19] , \ScanLink124[18] , \ScanLink124[17] , 
        \ScanLink124[16] , \ScanLink124[15] , \ScanLink124[14] , 
        \ScanLink124[13] , \ScanLink124[12] , \ScanLink124[11] , 
        \ScanLink124[10] , \ScanLink124[9] , \ScanLink124[8] , 
        \ScanLink124[7] , \ScanLink124[6] , \ScanLink124[5] , \ScanLink124[4] , 
        \ScanLink124[3] , \ScanLink124[2] , \ScanLink124[1] , \ScanLink124[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_61[31] , 
        \wRegOut_6_61[30] , \wRegOut_6_61[29] , \wRegOut_6_61[28] , 
        \wRegOut_6_61[27] , \wRegOut_6_61[26] , \wRegOut_6_61[25] , 
        \wRegOut_6_61[24] , \wRegOut_6_61[23] , \wRegOut_6_61[22] , 
        \wRegOut_6_61[21] , \wRegOut_6_61[20] , \wRegOut_6_61[19] , 
        \wRegOut_6_61[18] , \wRegOut_6_61[17] , \wRegOut_6_61[16] , 
        \wRegOut_6_61[15] , \wRegOut_6_61[14] , \wRegOut_6_61[13] , 
        \wRegOut_6_61[12] , \wRegOut_6_61[11] , \wRegOut_6_61[10] , 
        \wRegOut_6_61[9] , \wRegOut_6_61[8] , \wRegOut_6_61[7] , 
        \wRegOut_6_61[6] , \wRegOut_6_61[5] , \wRegOut_6_61[4] , 
        \wRegOut_6_61[3] , \wRegOut_6_61[2] , \wRegOut_6_61[1] , 
        \wRegOut_6_61[0] }), .Enable1(\wRegEnTop_6_61[0] ), .Enable2(
        \wRegEnBot_6_61[0] ), .In1({\wRegInTop_6_61[31] , \wRegInTop_6_61[30] , 
        \wRegInTop_6_61[29] , \wRegInTop_6_61[28] , \wRegInTop_6_61[27] , 
        \wRegInTop_6_61[26] , \wRegInTop_6_61[25] , \wRegInTop_6_61[24] , 
        \wRegInTop_6_61[23] , \wRegInTop_6_61[22] , \wRegInTop_6_61[21] , 
        \wRegInTop_6_61[20] , \wRegInTop_6_61[19] , \wRegInTop_6_61[18] , 
        \wRegInTop_6_61[17] , \wRegInTop_6_61[16] , \wRegInTop_6_61[15] , 
        \wRegInTop_6_61[14] , \wRegInTop_6_61[13] , \wRegInTop_6_61[12] , 
        \wRegInTop_6_61[11] , \wRegInTop_6_61[10] , \wRegInTop_6_61[9] , 
        \wRegInTop_6_61[8] , \wRegInTop_6_61[7] , \wRegInTop_6_61[6] , 
        \wRegInTop_6_61[5] , \wRegInTop_6_61[4] , \wRegInTop_6_61[3] , 
        \wRegInTop_6_61[2] , \wRegInTop_6_61[1] , \wRegInTop_6_61[0] }), .In2(
        {\wRegInBot_6_61[31] , \wRegInBot_6_61[30] , \wRegInBot_6_61[29] , 
        \wRegInBot_6_61[28] , \wRegInBot_6_61[27] , \wRegInBot_6_61[26] , 
        \wRegInBot_6_61[25] , \wRegInBot_6_61[24] , \wRegInBot_6_61[23] , 
        \wRegInBot_6_61[22] , \wRegInBot_6_61[21] , \wRegInBot_6_61[20] , 
        \wRegInBot_6_61[19] , \wRegInBot_6_61[18] , \wRegInBot_6_61[17] , 
        \wRegInBot_6_61[16] , \wRegInBot_6_61[15] , \wRegInBot_6_61[14] , 
        \wRegInBot_6_61[13] , \wRegInBot_6_61[12] , \wRegInBot_6_61[11] , 
        \wRegInBot_6_61[10] , \wRegInBot_6_61[9] , \wRegInBot_6_61[8] , 
        \wRegInBot_6_61[7] , \wRegInBot_6_61[6] , \wRegInBot_6_61[5] , 
        \wRegInBot_6_61[4] , \wRegInBot_6_61[3] , \wRegInBot_6_61[2] , 
        \wRegInBot_6_61[1] , \wRegInBot_6_61[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_32 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink160[31] , \ScanLink160[30] , \ScanLink160[29] , 
        \ScanLink160[28] , \ScanLink160[27] , \ScanLink160[26] , 
        \ScanLink160[25] , \ScanLink160[24] , \ScanLink160[23] , 
        \ScanLink160[22] , \ScanLink160[21] , \ScanLink160[20] , 
        \ScanLink160[19] , \ScanLink160[18] , \ScanLink160[17] , 
        \ScanLink160[16] , \ScanLink160[15] , \ScanLink160[14] , 
        \ScanLink160[13] , \ScanLink160[12] , \ScanLink160[11] , 
        \ScanLink160[10] , \ScanLink160[9] , \ScanLink160[8] , 
        \ScanLink160[7] , \ScanLink160[6] , \ScanLink160[5] , \ScanLink160[4] , 
        \ScanLink160[3] , \ScanLink160[2] , \ScanLink160[1] , \ScanLink160[0] 
        }), .ScanOut({\ScanLink159[31] , \ScanLink159[30] , \ScanLink159[29] , 
        \ScanLink159[28] , \ScanLink159[27] , \ScanLink159[26] , 
        \ScanLink159[25] , \ScanLink159[24] , \ScanLink159[23] , 
        \ScanLink159[22] , \ScanLink159[21] , \ScanLink159[20] , 
        \ScanLink159[19] , \ScanLink159[18] , \ScanLink159[17] , 
        \ScanLink159[16] , \ScanLink159[15] , \ScanLink159[14] , 
        \ScanLink159[13] , \ScanLink159[12] , \ScanLink159[11] , 
        \ScanLink159[10] , \ScanLink159[9] , \ScanLink159[8] , 
        \ScanLink159[7] , \ScanLink159[6] , \ScanLink159[5] , \ScanLink159[4] , 
        \ScanLink159[3] , \ScanLink159[2] , \ScanLink159[1] , \ScanLink159[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_32[31] , 
        \wRegOut_7_32[30] , \wRegOut_7_32[29] , \wRegOut_7_32[28] , 
        \wRegOut_7_32[27] , \wRegOut_7_32[26] , \wRegOut_7_32[25] , 
        \wRegOut_7_32[24] , \wRegOut_7_32[23] , \wRegOut_7_32[22] , 
        \wRegOut_7_32[21] , \wRegOut_7_32[20] , \wRegOut_7_32[19] , 
        \wRegOut_7_32[18] , \wRegOut_7_32[17] , \wRegOut_7_32[16] , 
        \wRegOut_7_32[15] , \wRegOut_7_32[14] , \wRegOut_7_32[13] , 
        \wRegOut_7_32[12] , \wRegOut_7_32[11] , \wRegOut_7_32[10] , 
        \wRegOut_7_32[9] , \wRegOut_7_32[8] , \wRegOut_7_32[7] , 
        \wRegOut_7_32[6] , \wRegOut_7_32[5] , \wRegOut_7_32[4] , 
        \wRegOut_7_32[3] , \wRegOut_7_32[2] , \wRegOut_7_32[1] , 
        \wRegOut_7_32[0] }), .Enable1(\wRegEnTop_7_32[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_32[31] , \wRegInTop_7_32[30] , \wRegInTop_7_32[29] , 
        \wRegInTop_7_32[28] , \wRegInTop_7_32[27] , \wRegInTop_7_32[26] , 
        \wRegInTop_7_32[25] , \wRegInTop_7_32[24] , \wRegInTop_7_32[23] , 
        \wRegInTop_7_32[22] , \wRegInTop_7_32[21] , \wRegInTop_7_32[20] , 
        \wRegInTop_7_32[19] , \wRegInTop_7_32[18] , \wRegInTop_7_32[17] , 
        \wRegInTop_7_32[16] , \wRegInTop_7_32[15] , \wRegInTop_7_32[14] , 
        \wRegInTop_7_32[13] , \wRegInTop_7_32[12] , \wRegInTop_7_32[11] , 
        \wRegInTop_7_32[10] , \wRegInTop_7_32[9] , \wRegInTop_7_32[8] , 
        \wRegInTop_7_32[7] , \wRegInTop_7_32[6] , \wRegInTop_7_32[5] , 
        \wRegInTop_7_32[4] , \wRegInTop_7_32[3] , \wRegInTop_7_32[2] , 
        \wRegInTop_7_32[1] , \wRegInTop_7_32[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_126 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink254[31] , \ScanLink254[30] , \ScanLink254[29] , 
        \ScanLink254[28] , \ScanLink254[27] , \ScanLink254[26] , 
        \ScanLink254[25] , \ScanLink254[24] , \ScanLink254[23] , 
        \ScanLink254[22] , \ScanLink254[21] , \ScanLink254[20] , 
        \ScanLink254[19] , \ScanLink254[18] , \ScanLink254[17] , 
        \ScanLink254[16] , \ScanLink254[15] , \ScanLink254[14] , 
        \ScanLink254[13] , \ScanLink254[12] , \ScanLink254[11] , 
        \ScanLink254[10] , \ScanLink254[9] , \ScanLink254[8] , 
        \ScanLink254[7] , \ScanLink254[6] , \ScanLink254[5] , \ScanLink254[4] , 
        \ScanLink254[3] , \ScanLink254[2] , \ScanLink254[1] , \ScanLink254[0] 
        }), .ScanOut({\ScanLink253[31] , \ScanLink253[30] , \ScanLink253[29] , 
        \ScanLink253[28] , \ScanLink253[27] , \ScanLink253[26] , 
        \ScanLink253[25] , \ScanLink253[24] , \ScanLink253[23] , 
        \ScanLink253[22] , \ScanLink253[21] , \ScanLink253[20] , 
        \ScanLink253[19] , \ScanLink253[18] , \ScanLink253[17] , 
        \ScanLink253[16] , \ScanLink253[15] , \ScanLink253[14] , 
        \ScanLink253[13] , \ScanLink253[12] , \ScanLink253[11] , 
        \ScanLink253[10] , \ScanLink253[9] , \ScanLink253[8] , 
        \ScanLink253[7] , \ScanLink253[6] , \ScanLink253[5] , \ScanLink253[4] , 
        \ScanLink253[3] , \ScanLink253[2] , \ScanLink253[1] , \ScanLink253[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_126[31] , 
        \wRegOut_7_126[30] , \wRegOut_7_126[29] , \wRegOut_7_126[28] , 
        \wRegOut_7_126[27] , \wRegOut_7_126[26] , \wRegOut_7_126[25] , 
        \wRegOut_7_126[24] , \wRegOut_7_126[23] , \wRegOut_7_126[22] , 
        \wRegOut_7_126[21] , \wRegOut_7_126[20] , \wRegOut_7_126[19] , 
        \wRegOut_7_126[18] , \wRegOut_7_126[17] , \wRegOut_7_126[16] , 
        \wRegOut_7_126[15] , \wRegOut_7_126[14] , \wRegOut_7_126[13] , 
        \wRegOut_7_126[12] , \wRegOut_7_126[11] , \wRegOut_7_126[10] , 
        \wRegOut_7_126[9] , \wRegOut_7_126[8] , \wRegOut_7_126[7] , 
        \wRegOut_7_126[6] , \wRegOut_7_126[5] , \wRegOut_7_126[4] , 
        \wRegOut_7_126[3] , \wRegOut_7_126[2] , \wRegOut_7_126[1] , 
        \wRegOut_7_126[0] }), .Enable1(\wRegEnTop_7_126[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_126[31] , \wRegInTop_7_126[30] , 
        \wRegInTop_7_126[29] , \wRegInTop_7_126[28] , \wRegInTop_7_126[27] , 
        \wRegInTop_7_126[26] , \wRegInTop_7_126[25] , \wRegInTop_7_126[24] , 
        \wRegInTop_7_126[23] , \wRegInTop_7_126[22] , \wRegInTop_7_126[21] , 
        \wRegInTop_7_126[20] , \wRegInTop_7_126[19] , \wRegInTop_7_126[18] , 
        \wRegInTop_7_126[17] , \wRegInTop_7_126[16] , \wRegInTop_7_126[15] , 
        \wRegInTop_7_126[14] , \wRegInTop_7_126[13] , \wRegInTop_7_126[12] , 
        \wRegInTop_7_126[11] , \wRegInTop_7_126[10] , \wRegInTop_7_126[9] , 
        \wRegInTop_7_126[8] , \wRegInTop_7_126[7] , \wRegInTop_7_126[6] , 
        \wRegInTop_7_126[5] , \wRegInTop_7_126[4] , \wRegInTop_7_126[3] , 
        \wRegInTop_7_126[2] , \wRegInTop_7_126[1] , \wRegInTop_7_126[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_101 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink229[31] , \ScanLink229[30] , \ScanLink229[29] , 
        \ScanLink229[28] , \ScanLink229[27] , \ScanLink229[26] , 
        \ScanLink229[25] , \ScanLink229[24] , \ScanLink229[23] , 
        \ScanLink229[22] , \ScanLink229[21] , \ScanLink229[20] , 
        \ScanLink229[19] , \ScanLink229[18] , \ScanLink229[17] , 
        \ScanLink229[16] , \ScanLink229[15] , \ScanLink229[14] , 
        \ScanLink229[13] , \ScanLink229[12] , \ScanLink229[11] , 
        \ScanLink229[10] , \ScanLink229[9] , \ScanLink229[8] , 
        \ScanLink229[7] , \ScanLink229[6] , \ScanLink229[5] , \ScanLink229[4] , 
        \ScanLink229[3] , \ScanLink229[2] , \ScanLink229[1] , \ScanLink229[0] 
        }), .ScanOut({\ScanLink228[31] , \ScanLink228[30] , \ScanLink228[29] , 
        \ScanLink228[28] , \ScanLink228[27] , \ScanLink228[26] , 
        \ScanLink228[25] , \ScanLink228[24] , \ScanLink228[23] , 
        \ScanLink228[22] , \ScanLink228[21] , \ScanLink228[20] , 
        \ScanLink228[19] , \ScanLink228[18] , \ScanLink228[17] , 
        \ScanLink228[16] , \ScanLink228[15] , \ScanLink228[14] , 
        \ScanLink228[13] , \ScanLink228[12] , \ScanLink228[11] , 
        \ScanLink228[10] , \ScanLink228[9] , \ScanLink228[8] , 
        \ScanLink228[7] , \ScanLink228[6] , \ScanLink228[5] , \ScanLink228[4] , 
        \ScanLink228[3] , \ScanLink228[2] , \ScanLink228[1] , \ScanLink228[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_101[31] , 
        \wRegOut_7_101[30] , \wRegOut_7_101[29] , \wRegOut_7_101[28] , 
        \wRegOut_7_101[27] , \wRegOut_7_101[26] , \wRegOut_7_101[25] , 
        \wRegOut_7_101[24] , \wRegOut_7_101[23] , \wRegOut_7_101[22] , 
        \wRegOut_7_101[21] , \wRegOut_7_101[20] , \wRegOut_7_101[19] , 
        \wRegOut_7_101[18] , \wRegOut_7_101[17] , \wRegOut_7_101[16] , 
        \wRegOut_7_101[15] , \wRegOut_7_101[14] , \wRegOut_7_101[13] , 
        \wRegOut_7_101[12] , \wRegOut_7_101[11] , \wRegOut_7_101[10] , 
        \wRegOut_7_101[9] , \wRegOut_7_101[8] , \wRegOut_7_101[7] , 
        \wRegOut_7_101[6] , \wRegOut_7_101[5] , \wRegOut_7_101[4] , 
        \wRegOut_7_101[3] , \wRegOut_7_101[2] , \wRegOut_7_101[1] , 
        \wRegOut_7_101[0] }), .Enable1(\wRegEnTop_7_101[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_101[31] , \wRegInTop_7_101[30] , 
        \wRegInTop_7_101[29] , \wRegInTop_7_101[28] , \wRegInTop_7_101[27] , 
        \wRegInTop_7_101[26] , \wRegInTop_7_101[25] , \wRegInTop_7_101[24] , 
        \wRegInTop_7_101[23] , \wRegInTop_7_101[22] , \wRegInTop_7_101[21] , 
        \wRegInTop_7_101[20] , \wRegInTop_7_101[19] , \wRegInTop_7_101[18] , 
        \wRegInTop_7_101[17] , \wRegInTop_7_101[16] , \wRegInTop_7_101[15] , 
        \wRegInTop_7_101[14] , \wRegInTop_7_101[13] , \wRegInTop_7_101[12] , 
        \wRegInTop_7_101[11] , \wRegInTop_7_101[10] , \wRegInTop_7_101[9] , 
        \wRegInTop_7_101[8] , \wRegInTop_7_101[7] , \wRegInTop_7_101[6] , 
        \wRegInTop_7_101[5] , \wRegInTop_7_101[4] , \wRegInTop_7_101[3] , 
        \wRegInTop_7_101[2] , \wRegInTop_7_101[1] , \wRegInTop_7_101[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_CtrlReg_WIDTH32 BHCR_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_2[0] ), 
        .Out(\wCtrlOut_1[0] ), .Enable(\wEnable_1[0] ) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink129[31] , \ScanLink129[30] , \ScanLink129[29] , 
        \ScanLink129[28] , \ScanLink129[27] , \ScanLink129[26] , 
        \ScanLink129[25] , \ScanLink129[24] , \ScanLink129[23] , 
        \ScanLink129[22] , \ScanLink129[21] , \ScanLink129[20] , 
        \ScanLink129[19] , \ScanLink129[18] , \ScanLink129[17] , 
        \ScanLink129[16] , \ScanLink129[15] , \ScanLink129[14] , 
        \ScanLink129[13] , \ScanLink129[12] , \ScanLink129[11] , 
        \ScanLink129[10] , \ScanLink129[9] , \ScanLink129[8] , 
        \ScanLink129[7] , \ScanLink129[6] , \ScanLink129[5] , \ScanLink129[4] , 
        \ScanLink129[3] , \ScanLink129[2] , \ScanLink129[1] , \ScanLink129[0] 
        }), .ScanOut({\ScanLink128[31] , \ScanLink128[30] , \ScanLink128[29] , 
        \ScanLink128[28] , \ScanLink128[27] , \ScanLink128[26] , 
        \ScanLink128[25] , \ScanLink128[24] , \ScanLink128[23] , 
        \ScanLink128[22] , \ScanLink128[21] , \ScanLink128[20] , 
        \ScanLink128[19] , \ScanLink128[18] , \ScanLink128[17] , 
        \ScanLink128[16] , \ScanLink128[15] , \ScanLink128[14] , 
        \ScanLink128[13] , \ScanLink128[12] , \ScanLink128[11] , 
        \ScanLink128[10] , \ScanLink128[9] , \ScanLink128[8] , 
        \ScanLink128[7] , \ScanLink128[6] , \ScanLink128[5] , \ScanLink128[4] , 
        \ScanLink128[3] , \ScanLink128[2] , \ScanLink128[1] , \ScanLink128[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_1[31] , 
        \wRegOut_7_1[30] , \wRegOut_7_1[29] , \wRegOut_7_1[28] , 
        \wRegOut_7_1[27] , \wRegOut_7_1[26] , \wRegOut_7_1[25] , 
        \wRegOut_7_1[24] , \wRegOut_7_1[23] , \wRegOut_7_1[22] , 
        \wRegOut_7_1[21] , \wRegOut_7_1[20] , \wRegOut_7_1[19] , 
        \wRegOut_7_1[18] , \wRegOut_7_1[17] , \wRegOut_7_1[16] , 
        \wRegOut_7_1[15] , \wRegOut_7_1[14] , \wRegOut_7_1[13] , 
        \wRegOut_7_1[12] , \wRegOut_7_1[11] , \wRegOut_7_1[10] , 
        \wRegOut_7_1[9] , \wRegOut_7_1[8] , \wRegOut_7_1[7] , \wRegOut_7_1[6] , 
        \wRegOut_7_1[5] , \wRegOut_7_1[4] , \wRegOut_7_1[3] , \wRegOut_7_1[2] , 
        \wRegOut_7_1[1] , \wRegOut_7_1[0] }), .Enable1(\wRegEnTop_7_1[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_1[31] , \wRegInTop_7_1[30] , 
        \wRegInTop_7_1[29] , \wRegInTop_7_1[28] , \wRegInTop_7_1[27] , 
        \wRegInTop_7_1[26] , \wRegInTop_7_1[25] , \wRegInTop_7_1[24] , 
        \wRegInTop_7_1[23] , \wRegInTop_7_1[22] , \wRegInTop_7_1[21] , 
        \wRegInTop_7_1[20] , \wRegInTop_7_1[19] , \wRegInTop_7_1[18] , 
        \wRegInTop_7_1[17] , \wRegInTop_7_1[16] , \wRegInTop_7_1[15] , 
        \wRegInTop_7_1[14] , \wRegInTop_7_1[13] , \wRegInTop_7_1[12] , 
        \wRegInTop_7_1[11] , \wRegInTop_7_1[10] , \wRegInTop_7_1[9] , 
        \wRegInTop_7_1[8] , \wRegInTop_7_1[7] , \wRegInTop_7_1[6] , 
        \wRegInTop_7_1[5] , \wRegInTop_7_1[4] , \wRegInTop_7_1[3] , 
        \wRegInTop_7_1[2] , \wRegInTop_7_1[1] , \wRegInTop_7_1[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink143[31] , \ScanLink143[30] , \ScanLink143[29] , 
        \ScanLink143[28] , \ScanLink143[27] , \ScanLink143[26] , 
        \ScanLink143[25] , \ScanLink143[24] , \ScanLink143[23] , 
        \ScanLink143[22] , \ScanLink143[21] , \ScanLink143[20] , 
        \ScanLink143[19] , \ScanLink143[18] , \ScanLink143[17] , 
        \ScanLink143[16] , \ScanLink143[15] , \ScanLink143[14] , 
        \ScanLink143[13] , \ScanLink143[12] , \ScanLink143[11] , 
        \ScanLink143[10] , \ScanLink143[9] , \ScanLink143[8] , 
        \ScanLink143[7] , \ScanLink143[6] , \ScanLink143[5] , \ScanLink143[4] , 
        \ScanLink143[3] , \ScanLink143[2] , \ScanLink143[1] , \ScanLink143[0] 
        }), .ScanOut({\ScanLink142[31] , \ScanLink142[30] , \ScanLink142[29] , 
        \ScanLink142[28] , \ScanLink142[27] , \ScanLink142[26] , 
        \ScanLink142[25] , \ScanLink142[24] , \ScanLink142[23] , 
        \ScanLink142[22] , \ScanLink142[21] , \ScanLink142[20] , 
        \ScanLink142[19] , \ScanLink142[18] , \ScanLink142[17] , 
        \ScanLink142[16] , \ScanLink142[15] , \ScanLink142[14] , 
        \ScanLink142[13] , \ScanLink142[12] , \ScanLink142[11] , 
        \ScanLink142[10] , \ScanLink142[9] , \ScanLink142[8] , 
        \ScanLink142[7] , \ScanLink142[6] , \ScanLink142[5] , \ScanLink142[4] , 
        \ScanLink142[3] , \ScanLink142[2] , \ScanLink142[1] , \ScanLink142[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_15[31] , 
        \wRegOut_7_15[30] , \wRegOut_7_15[29] , \wRegOut_7_15[28] , 
        \wRegOut_7_15[27] , \wRegOut_7_15[26] , \wRegOut_7_15[25] , 
        \wRegOut_7_15[24] , \wRegOut_7_15[23] , \wRegOut_7_15[22] , 
        \wRegOut_7_15[21] , \wRegOut_7_15[20] , \wRegOut_7_15[19] , 
        \wRegOut_7_15[18] , \wRegOut_7_15[17] , \wRegOut_7_15[16] , 
        \wRegOut_7_15[15] , \wRegOut_7_15[14] , \wRegOut_7_15[13] , 
        \wRegOut_7_15[12] , \wRegOut_7_15[11] , \wRegOut_7_15[10] , 
        \wRegOut_7_15[9] , \wRegOut_7_15[8] , \wRegOut_7_15[7] , 
        \wRegOut_7_15[6] , \wRegOut_7_15[5] , \wRegOut_7_15[4] , 
        \wRegOut_7_15[3] , \wRegOut_7_15[2] , \wRegOut_7_15[1] , 
        \wRegOut_7_15[0] }), .Enable1(\wRegEnTop_7_15[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_15[31] , \wRegInTop_7_15[30] , \wRegInTop_7_15[29] , 
        \wRegInTop_7_15[28] , \wRegInTop_7_15[27] , \wRegInTop_7_15[26] , 
        \wRegInTop_7_15[25] , \wRegInTop_7_15[24] , \wRegInTop_7_15[23] , 
        \wRegInTop_7_15[22] , \wRegInTop_7_15[21] , \wRegInTop_7_15[20] , 
        \wRegInTop_7_15[19] , \wRegInTop_7_15[18] , \wRegInTop_7_15[17] , 
        \wRegInTop_7_15[16] , \wRegInTop_7_15[15] , \wRegInTop_7_15[14] , 
        \wRegInTop_7_15[13] , \wRegInTop_7_15[12] , \wRegInTop_7_15[11] , 
        \wRegInTop_7_15[10] , \wRegInTop_7_15[9] , \wRegInTop_7_15[8] , 
        \wRegInTop_7_15[7] , \wRegInTop_7_15[6] , \wRegInTop_7_15[5] , 
        \wRegInTop_7_15[4] , \wRegInTop_7_15[3] , \wRegInTop_7_15[2] , 
        \wRegInTop_7_15[1] , \wRegInTop_7_15[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_49[0] ), .P_In({\wRegOut_6_49[31] , 
        \wRegOut_6_49[30] , \wRegOut_6_49[29] , \wRegOut_6_49[28] , 
        \wRegOut_6_49[27] , \wRegOut_6_49[26] , \wRegOut_6_49[25] , 
        \wRegOut_6_49[24] , \wRegOut_6_49[23] , \wRegOut_6_49[22] , 
        \wRegOut_6_49[21] , \wRegOut_6_49[20] , \wRegOut_6_49[19] , 
        \wRegOut_6_49[18] , \wRegOut_6_49[17] , \wRegOut_6_49[16] , 
        \wRegOut_6_49[15] , \wRegOut_6_49[14] , \wRegOut_6_49[13] , 
        \wRegOut_6_49[12] , \wRegOut_6_49[11] , \wRegOut_6_49[10] , 
        \wRegOut_6_49[9] , \wRegOut_6_49[8] , \wRegOut_6_49[7] , 
        \wRegOut_6_49[6] , \wRegOut_6_49[5] , \wRegOut_6_49[4] , 
        \wRegOut_6_49[3] , \wRegOut_6_49[2] , \wRegOut_6_49[1] , 
        \wRegOut_6_49[0] }), .P_Out({\wRegInBot_6_49[31] , 
        \wRegInBot_6_49[30] , \wRegInBot_6_49[29] , \wRegInBot_6_49[28] , 
        \wRegInBot_6_49[27] , \wRegInBot_6_49[26] , \wRegInBot_6_49[25] , 
        \wRegInBot_6_49[24] , \wRegInBot_6_49[23] , \wRegInBot_6_49[22] , 
        \wRegInBot_6_49[21] , \wRegInBot_6_49[20] , \wRegInBot_6_49[19] , 
        \wRegInBot_6_49[18] , \wRegInBot_6_49[17] , \wRegInBot_6_49[16] , 
        \wRegInBot_6_49[15] , \wRegInBot_6_49[14] , \wRegInBot_6_49[13] , 
        \wRegInBot_6_49[12] , \wRegInBot_6_49[11] , \wRegInBot_6_49[10] , 
        \wRegInBot_6_49[9] , \wRegInBot_6_49[8] , \wRegInBot_6_49[7] , 
        \wRegInBot_6_49[6] , \wRegInBot_6_49[5] , \wRegInBot_6_49[4] , 
        \wRegInBot_6_49[3] , \wRegInBot_6_49[2] , \wRegInBot_6_49[1] , 
        \wRegInBot_6_49[0] }), .L_WR(\wRegEnTop_7_98[0] ), .L_In({
        \wRegOut_7_98[31] , \wRegOut_7_98[30] , \wRegOut_7_98[29] , 
        \wRegOut_7_98[28] , \wRegOut_7_98[27] , \wRegOut_7_98[26] , 
        \wRegOut_7_98[25] , \wRegOut_7_98[24] , \wRegOut_7_98[23] , 
        \wRegOut_7_98[22] , \wRegOut_7_98[21] , \wRegOut_7_98[20] , 
        \wRegOut_7_98[19] , \wRegOut_7_98[18] , \wRegOut_7_98[17] , 
        \wRegOut_7_98[16] , \wRegOut_7_98[15] , \wRegOut_7_98[14] , 
        \wRegOut_7_98[13] , \wRegOut_7_98[12] , \wRegOut_7_98[11] , 
        \wRegOut_7_98[10] , \wRegOut_7_98[9] , \wRegOut_7_98[8] , 
        \wRegOut_7_98[7] , \wRegOut_7_98[6] , \wRegOut_7_98[5] , 
        \wRegOut_7_98[4] , \wRegOut_7_98[3] , \wRegOut_7_98[2] , 
        \wRegOut_7_98[1] , \wRegOut_7_98[0] }), .L_Out({\wRegInTop_7_98[31] , 
        \wRegInTop_7_98[30] , \wRegInTop_7_98[29] , \wRegInTop_7_98[28] , 
        \wRegInTop_7_98[27] , \wRegInTop_7_98[26] , \wRegInTop_7_98[25] , 
        \wRegInTop_7_98[24] , \wRegInTop_7_98[23] , \wRegInTop_7_98[22] , 
        \wRegInTop_7_98[21] , \wRegInTop_7_98[20] , \wRegInTop_7_98[19] , 
        \wRegInTop_7_98[18] , \wRegInTop_7_98[17] , \wRegInTop_7_98[16] , 
        \wRegInTop_7_98[15] , \wRegInTop_7_98[14] , \wRegInTop_7_98[13] , 
        \wRegInTop_7_98[12] , \wRegInTop_7_98[11] , \wRegInTop_7_98[10] , 
        \wRegInTop_7_98[9] , \wRegInTop_7_98[8] , \wRegInTop_7_98[7] , 
        \wRegInTop_7_98[6] , \wRegInTop_7_98[5] , \wRegInTop_7_98[4] , 
        \wRegInTop_7_98[3] , \wRegInTop_7_98[2] , \wRegInTop_7_98[1] , 
        \wRegInTop_7_98[0] }), .R_WR(\wRegEnTop_7_99[0] ), .R_In({
        \wRegOut_7_99[31] , \wRegOut_7_99[30] , \wRegOut_7_99[29] , 
        \wRegOut_7_99[28] , \wRegOut_7_99[27] , \wRegOut_7_99[26] , 
        \wRegOut_7_99[25] , \wRegOut_7_99[24] , \wRegOut_7_99[23] , 
        \wRegOut_7_99[22] , \wRegOut_7_99[21] , \wRegOut_7_99[20] , 
        \wRegOut_7_99[19] , \wRegOut_7_99[18] , \wRegOut_7_99[17] , 
        \wRegOut_7_99[16] , \wRegOut_7_99[15] , \wRegOut_7_99[14] , 
        \wRegOut_7_99[13] , \wRegOut_7_99[12] , \wRegOut_7_99[11] , 
        \wRegOut_7_99[10] , \wRegOut_7_99[9] , \wRegOut_7_99[8] , 
        \wRegOut_7_99[7] , \wRegOut_7_99[6] , \wRegOut_7_99[5] , 
        \wRegOut_7_99[4] , \wRegOut_7_99[3] , \wRegOut_7_99[2] , 
        \wRegOut_7_99[1] , \wRegOut_7_99[0] }), .R_Out({\wRegInTop_7_99[31] , 
        \wRegInTop_7_99[30] , \wRegInTop_7_99[29] , \wRegInTop_7_99[28] , 
        \wRegInTop_7_99[27] , \wRegInTop_7_99[26] , \wRegInTop_7_99[25] , 
        \wRegInTop_7_99[24] , \wRegInTop_7_99[23] , \wRegInTop_7_99[22] , 
        \wRegInTop_7_99[21] , \wRegInTop_7_99[20] , \wRegInTop_7_99[19] , 
        \wRegInTop_7_99[18] , \wRegInTop_7_99[17] , \wRegInTop_7_99[16] , 
        \wRegInTop_7_99[15] , \wRegInTop_7_99[14] , \wRegInTop_7_99[13] , 
        \wRegInTop_7_99[12] , \wRegInTop_7_99[11] , \wRegInTop_7_99[10] , 
        \wRegInTop_7_99[9] , \wRegInTop_7_99[8] , \wRegInTop_7_99[7] , 
        \wRegInTop_7_99[6] , \wRegInTop_7_99[5] , \wRegInTop_7_99[4] , 
        \wRegInTop_7_99[3] , \wRegInTop_7_99[2] , \wRegInTop_7_99[1] , 
        \wRegInTop_7_99[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_29 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink157[31] , \ScanLink157[30] , \ScanLink157[29] , 
        \ScanLink157[28] , \ScanLink157[27] , \ScanLink157[26] , 
        \ScanLink157[25] , \ScanLink157[24] , \ScanLink157[23] , 
        \ScanLink157[22] , \ScanLink157[21] , \ScanLink157[20] , 
        \ScanLink157[19] , \ScanLink157[18] , \ScanLink157[17] , 
        \ScanLink157[16] , \ScanLink157[15] , \ScanLink157[14] , 
        \ScanLink157[13] , \ScanLink157[12] , \ScanLink157[11] , 
        \ScanLink157[10] , \ScanLink157[9] , \ScanLink157[8] , 
        \ScanLink157[7] , \ScanLink157[6] , \ScanLink157[5] , \ScanLink157[4] , 
        \ScanLink157[3] , \ScanLink157[2] , \ScanLink157[1] , \ScanLink157[0] 
        }), .ScanOut({\ScanLink156[31] , \ScanLink156[30] , \ScanLink156[29] , 
        \ScanLink156[28] , \ScanLink156[27] , \ScanLink156[26] , 
        \ScanLink156[25] , \ScanLink156[24] , \ScanLink156[23] , 
        \ScanLink156[22] , \ScanLink156[21] , \ScanLink156[20] , 
        \ScanLink156[19] , \ScanLink156[18] , \ScanLink156[17] , 
        \ScanLink156[16] , \ScanLink156[15] , \ScanLink156[14] , 
        \ScanLink156[13] , \ScanLink156[12] , \ScanLink156[11] , 
        \ScanLink156[10] , \ScanLink156[9] , \ScanLink156[8] , 
        \ScanLink156[7] , \ScanLink156[6] , \ScanLink156[5] , \ScanLink156[4] , 
        \ScanLink156[3] , \ScanLink156[2] , \ScanLink156[1] , \ScanLink156[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_29[31] , 
        \wRegOut_7_29[30] , \wRegOut_7_29[29] , \wRegOut_7_29[28] , 
        \wRegOut_7_29[27] , \wRegOut_7_29[26] , \wRegOut_7_29[25] , 
        \wRegOut_7_29[24] , \wRegOut_7_29[23] , \wRegOut_7_29[22] , 
        \wRegOut_7_29[21] , \wRegOut_7_29[20] , \wRegOut_7_29[19] , 
        \wRegOut_7_29[18] , \wRegOut_7_29[17] , \wRegOut_7_29[16] , 
        \wRegOut_7_29[15] , \wRegOut_7_29[14] , \wRegOut_7_29[13] , 
        \wRegOut_7_29[12] , \wRegOut_7_29[11] , \wRegOut_7_29[10] , 
        \wRegOut_7_29[9] , \wRegOut_7_29[8] , \wRegOut_7_29[7] , 
        \wRegOut_7_29[6] , \wRegOut_7_29[5] , \wRegOut_7_29[4] , 
        \wRegOut_7_29[3] , \wRegOut_7_29[2] , \wRegOut_7_29[1] , 
        \wRegOut_7_29[0] }), .Enable1(\wRegEnTop_7_29[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_29[31] , \wRegInTop_7_29[30] , \wRegInTop_7_29[29] , 
        \wRegInTop_7_29[28] , \wRegInTop_7_29[27] , \wRegInTop_7_29[26] , 
        \wRegInTop_7_29[25] , \wRegInTop_7_29[24] , \wRegInTop_7_29[23] , 
        \wRegInTop_7_29[22] , \wRegInTop_7_29[21] , \wRegInTop_7_29[20] , 
        \wRegInTop_7_29[19] , \wRegInTop_7_29[18] , \wRegInTop_7_29[17] , 
        \wRegInTop_7_29[16] , \wRegInTop_7_29[15] , \wRegInTop_7_29[14] , 
        \wRegInTop_7_29[13] , \wRegInTop_7_29[12] , \wRegInTop_7_29[11] , 
        \wRegInTop_7_29[10] , \wRegInTop_7_29[9] , \wRegInTop_7_29[8] , 
        \wRegInTop_7_29[7] , \wRegInTop_7_29[6] , \wRegInTop_7_29[5] , 
        \wRegInTop_7_29[4] , \wRegInTop_7_29[3] , \wRegInTop_7_29[2] , 
        \wRegInTop_7_29[1] , \wRegInTop_7_29[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_52[0] ), .P_In({\wRegOut_6_52[31] , 
        \wRegOut_6_52[30] , \wRegOut_6_52[29] , \wRegOut_6_52[28] , 
        \wRegOut_6_52[27] , \wRegOut_6_52[26] , \wRegOut_6_52[25] , 
        \wRegOut_6_52[24] , \wRegOut_6_52[23] , \wRegOut_6_52[22] , 
        \wRegOut_6_52[21] , \wRegOut_6_52[20] , \wRegOut_6_52[19] , 
        \wRegOut_6_52[18] , \wRegOut_6_52[17] , \wRegOut_6_52[16] , 
        \wRegOut_6_52[15] , \wRegOut_6_52[14] , \wRegOut_6_52[13] , 
        \wRegOut_6_52[12] , \wRegOut_6_52[11] , \wRegOut_6_52[10] , 
        \wRegOut_6_52[9] , \wRegOut_6_52[8] , \wRegOut_6_52[7] , 
        \wRegOut_6_52[6] , \wRegOut_6_52[5] , \wRegOut_6_52[4] , 
        \wRegOut_6_52[3] , \wRegOut_6_52[2] , \wRegOut_6_52[1] , 
        \wRegOut_6_52[0] }), .P_Out({\wRegInBot_6_52[31] , 
        \wRegInBot_6_52[30] , \wRegInBot_6_52[29] , \wRegInBot_6_52[28] , 
        \wRegInBot_6_52[27] , \wRegInBot_6_52[26] , \wRegInBot_6_52[25] , 
        \wRegInBot_6_52[24] , \wRegInBot_6_52[23] , \wRegInBot_6_52[22] , 
        \wRegInBot_6_52[21] , \wRegInBot_6_52[20] , \wRegInBot_6_52[19] , 
        \wRegInBot_6_52[18] , \wRegInBot_6_52[17] , \wRegInBot_6_52[16] , 
        \wRegInBot_6_52[15] , \wRegInBot_6_52[14] , \wRegInBot_6_52[13] , 
        \wRegInBot_6_52[12] , \wRegInBot_6_52[11] , \wRegInBot_6_52[10] , 
        \wRegInBot_6_52[9] , \wRegInBot_6_52[8] , \wRegInBot_6_52[7] , 
        \wRegInBot_6_52[6] , \wRegInBot_6_52[5] , \wRegInBot_6_52[4] , 
        \wRegInBot_6_52[3] , \wRegInBot_6_52[2] , \wRegInBot_6_52[1] , 
        \wRegInBot_6_52[0] }), .L_WR(\wRegEnTop_7_104[0] ), .L_In({
        \wRegOut_7_104[31] , \wRegOut_7_104[30] , \wRegOut_7_104[29] , 
        \wRegOut_7_104[28] , \wRegOut_7_104[27] , \wRegOut_7_104[26] , 
        \wRegOut_7_104[25] , \wRegOut_7_104[24] , \wRegOut_7_104[23] , 
        \wRegOut_7_104[22] , \wRegOut_7_104[21] , \wRegOut_7_104[20] , 
        \wRegOut_7_104[19] , \wRegOut_7_104[18] , \wRegOut_7_104[17] , 
        \wRegOut_7_104[16] , \wRegOut_7_104[15] , \wRegOut_7_104[14] , 
        \wRegOut_7_104[13] , \wRegOut_7_104[12] , \wRegOut_7_104[11] , 
        \wRegOut_7_104[10] , \wRegOut_7_104[9] , \wRegOut_7_104[8] , 
        \wRegOut_7_104[7] , \wRegOut_7_104[6] , \wRegOut_7_104[5] , 
        \wRegOut_7_104[4] , \wRegOut_7_104[3] , \wRegOut_7_104[2] , 
        \wRegOut_7_104[1] , \wRegOut_7_104[0] }), .L_Out({
        \wRegInTop_7_104[31] , \wRegInTop_7_104[30] , \wRegInTop_7_104[29] , 
        \wRegInTop_7_104[28] , \wRegInTop_7_104[27] , \wRegInTop_7_104[26] , 
        \wRegInTop_7_104[25] , \wRegInTop_7_104[24] , \wRegInTop_7_104[23] , 
        \wRegInTop_7_104[22] , \wRegInTop_7_104[21] , \wRegInTop_7_104[20] , 
        \wRegInTop_7_104[19] , \wRegInTop_7_104[18] , \wRegInTop_7_104[17] , 
        \wRegInTop_7_104[16] , \wRegInTop_7_104[15] , \wRegInTop_7_104[14] , 
        \wRegInTop_7_104[13] , \wRegInTop_7_104[12] , \wRegInTop_7_104[11] , 
        \wRegInTop_7_104[10] , \wRegInTop_7_104[9] , \wRegInTop_7_104[8] , 
        \wRegInTop_7_104[7] , \wRegInTop_7_104[6] , \wRegInTop_7_104[5] , 
        \wRegInTop_7_104[4] , \wRegInTop_7_104[3] , \wRegInTop_7_104[2] , 
        \wRegInTop_7_104[1] , \wRegInTop_7_104[0] }), .R_WR(
        \wRegEnTop_7_105[0] ), .R_In({\wRegOut_7_105[31] , \wRegOut_7_105[30] , 
        \wRegOut_7_105[29] , \wRegOut_7_105[28] , \wRegOut_7_105[27] , 
        \wRegOut_7_105[26] , \wRegOut_7_105[25] , \wRegOut_7_105[24] , 
        \wRegOut_7_105[23] , \wRegOut_7_105[22] , \wRegOut_7_105[21] , 
        \wRegOut_7_105[20] , \wRegOut_7_105[19] , \wRegOut_7_105[18] , 
        \wRegOut_7_105[17] , \wRegOut_7_105[16] , \wRegOut_7_105[15] , 
        \wRegOut_7_105[14] , \wRegOut_7_105[13] , \wRegOut_7_105[12] , 
        \wRegOut_7_105[11] , \wRegOut_7_105[10] , \wRegOut_7_105[9] , 
        \wRegOut_7_105[8] , \wRegOut_7_105[7] , \wRegOut_7_105[6] , 
        \wRegOut_7_105[5] , \wRegOut_7_105[4] , \wRegOut_7_105[3] , 
        \wRegOut_7_105[2] , \wRegOut_7_105[1] , \wRegOut_7_105[0] }), .R_Out({
        \wRegInTop_7_105[31] , \wRegInTop_7_105[30] , \wRegInTop_7_105[29] , 
        \wRegInTop_7_105[28] , \wRegInTop_7_105[27] , \wRegInTop_7_105[26] , 
        \wRegInTop_7_105[25] , \wRegInTop_7_105[24] , \wRegInTop_7_105[23] , 
        \wRegInTop_7_105[22] , \wRegInTop_7_105[21] , \wRegInTop_7_105[20] , 
        \wRegInTop_7_105[19] , \wRegInTop_7_105[18] , \wRegInTop_7_105[17] , 
        \wRegInTop_7_105[16] , \wRegInTop_7_105[15] , \wRegInTop_7_105[14] , 
        \wRegInTop_7_105[13] , \wRegInTop_7_105[12] , \wRegInTop_7_105[11] , 
        \wRegInTop_7_105[10] , \wRegInTop_7_105[9] , \wRegInTop_7_105[8] , 
        \wRegInTop_7_105[7] , \wRegInTop_7_105[6] , \wRegInTop_7_105[5] , 
        \wRegInTop_7_105[4] , \wRegInTop_7_105[3] , \wRegInTop_7_105[2] , 
        \wRegInTop_7_105[1] , \wRegInTop_7_105[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_85 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink213[31] , \ScanLink213[30] , \ScanLink213[29] , 
        \ScanLink213[28] , \ScanLink213[27] , \ScanLink213[26] , 
        \ScanLink213[25] , \ScanLink213[24] , \ScanLink213[23] , 
        \ScanLink213[22] , \ScanLink213[21] , \ScanLink213[20] , 
        \ScanLink213[19] , \ScanLink213[18] , \ScanLink213[17] , 
        \ScanLink213[16] , \ScanLink213[15] , \ScanLink213[14] , 
        \ScanLink213[13] , \ScanLink213[12] , \ScanLink213[11] , 
        \ScanLink213[10] , \ScanLink213[9] , \ScanLink213[8] , 
        \ScanLink213[7] , \ScanLink213[6] , \ScanLink213[5] , \ScanLink213[4] , 
        \ScanLink213[3] , \ScanLink213[2] , \ScanLink213[1] , \ScanLink213[0] 
        }), .ScanOut({\ScanLink212[31] , \ScanLink212[30] , \ScanLink212[29] , 
        \ScanLink212[28] , \ScanLink212[27] , \ScanLink212[26] , 
        \ScanLink212[25] , \ScanLink212[24] , \ScanLink212[23] , 
        \ScanLink212[22] , \ScanLink212[21] , \ScanLink212[20] , 
        \ScanLink212[19] , \ScanLink212[18] , \ScanLink212[17] , 
        \ScanLink212[16] , \ScanLink212[15] , \ScanLink212[14] , 
        \ScanLink212[13] , \ScanLink212[12] , \ScanLink212[11] , 
        \ScanLink212[10] , \ScanLink212[9] , \ScanLink212[8] , 
        \ScanLink212[7] , \ScanLink212[6] , \ScanLink212[5] , \ScanLink212[4] , 
        \ScanLink212[3] , \ScanLink212[2] , \ScanLink212[1] , \ScanLink212[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_85[31] , 
        \wRegOut_7_85[30] , \wRegOut_7_85[29] , \wRegOut_7_85[28] , 
        \wRegOut_7_85[27] , \wRegOut_7_85[26] , \wRegOut_7_85[25] , 
        \wRegOut_7_85[24] , \wRegOut_7_85[23] , \wRegOut_7_85[22] , 
        \wRegOut_7_85[21] , \wRegOut_7_85[20] , \wRegOut_7_85[19] , 
        \wRegOut_7_85[18] , \wRegOut_7_85[17] , \wRegOut_7_85[16] , 
        \wRegOut_7_85[15] , \wRegOut_7_85[14] , \wRegOut_7_85[13] , 
        \wRegOut_7_85[12] , \wRegOut_7_85[11] , \wRegOut_7_85[10] , 
        \wRegOut_7_85[9] , \wRegOut_7_85[8] , \wRegOut_7_85[7] , 
        \wRegOut_7_85[6] , \wRegOut_7_85[5] , \wRegOut_7_85[4] , 
        \wRegOut_7_85[3] , \wRegOut_7_85[2] , \wRegOut_7_85[1] , 
        \wRegOut_7_85[0] }), .Enable1(\wRegEnTop_7_85[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_85[31] , \wRegInTop_7_85[30] , \wRegInTop_7_85[29] , 
        \wRegInTop_7_85[28] , \wRegInTop_7_85[27] , \wRegInTop_7_85[26] , 
        \wRegInTop_7_85[25] , \wRegInTop_7_85[24] , \wRegInTop_7_85[23] , 
        \wRegInTop_7_85[22] , \wRegInTop_7_85[21] , \wRegInTop_7_85[20] , 
        \wRegInTop_7_85[19] , \wRegInTop_7_85[18] , \wRegInTop_7_85[17] , 
        \wRegInTop_7_85[16] , \wRegInTop_7_85[15] , \wRegInTop_7_85[14] , 
        \wRegInTop_7_85[13] , \wRegInTop_7_85[12] , \wRegInTop_7_85[11] , 
        \wRegInTop_7_85[10] , \wRegInTop_7_85[9] , \wRegInTop_7_85[8] , 
        \wRegInTop_7_85[7] , \wRegInTop_7_85[6] , \wRegInTop_7_85[5] , 
        \wRegInTop_7_85[4] , \wRegInTop_7_85[3] , \wRegInTop_7_85[2] , 
        \wRegInTop_7_85[1] , \wRegInTop_7_85[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_5[0] ), .P_In({\wRegOut_3_5[31] , 
        \wRegOut_3_5[30] , \wRegOut_3_5[29] , \wRegOut_3_5[28] , 
        \wRegOut_3_5[27] , \wRegOut_3_5[26] , \wRegOut_3_5[25] , 
        \wRegOut_3_5[24] , \wRegOut_3_5[23] , \wRegOut_3_5[22] , 
        \wRegOut_3_5[21] , \wRegOut_3_5[20] , \wRegOut_3_5[19] , 
        \wRegOut_3_5[18] , \wRegOut_3_5[17] , \wRegOut_3_5[16] , 
        \wRegOut_3_5[15] , \wRegOut_3_5[14] , \wRegOut_3_5[13] , 
        \wRegOut_3_5[12] , \wRegOut_3_5[11] , \wRegOut_3_5[10] , 
        \wRegOut_3_5[9] , \wRegOut_3_5[8] , \wRegOut_3_5[7] , \wRegOut_3_5[6] , 
        \wRegOut_3_5[5] , \wRegOut_3_5[4] , \wRegOut_3_5[3] , \wRegOut_3_5[2] , 
        \wRegOut_3_5[1] , \wRegOut_3_5[0] }), .P_Out({\wRegInBot_3_5[31] , 
        \wRegInBot_3_5[30] , \wRegInBot_3_5[29] , \wRegInBot_3_5[28] , 
        \wRegInBot_3_5[27] , \wRegInBot_3_5[26] , \wRegInBot_3_5[25] , 
        \wRegInBot_3_5[24] , \wRegInBot_3_5[23] , \wRegInBot_3_5[22] , 
        \wRegInBot_3_5[21] , \wRegInBot_3_5[20] , \wRegInBot_3_5[19] , 
        \wRegInBot_3_5[18] , \wRegInBot_3_5[17] , \wRegInBot_3_5[16] , 
        \wRegInBot_3_5[15] , \wRegInBot_3_5[14] , \wRegInBot_3_5[13] , 
        \wRegInBot_3_5[12] , \wRegInBot_3_5[11] , \wRegInBot_3_5[10] , 
        \wRegInBot_3_5[9] , \wRegInBot_3_5[8] , \wRegInBot_3_5[7] , 
        \wRegInBot_3_5[6] , \wRegInBot_3_5[5] , \wRegInBot_3_5[4] , 
        \wRegInBot_3_5[3] , \wRegInBot_3_5[2] , \wRegInBot_3_5[1] , 
        \wRegInBot_3_5[0] }), .L_WR(\wRegEnTop_4_10[0] ), .L_In({
        \wRegOut_4_10[31] , \wRegOut_4_10[30] , \wRegOut_4_10[29] , 
        \wRegOut_4_10[28] , \wRegOut_4_10[27] , \wRegOut_4_10[26] , 
        \wRegOut_4_10[25] , \wRegOut_4_10[24] , \wRegOut_4_10[23] , 
        \wRegOut_4_10[22] , \wRegOut_4_10[21] , \wRegOut_4_10[20] , 
        \wRegOut_4_10[19] , \wRegOut_4_10[18] , \wRegOut_4_10[17] , 
        \wRegOut_4_10[16] , \wRegOut_4_10[15] , \wRegOut_4_10[14] , 
        \wRegOut_4_10[13] , \wRegOut_4_10[12] , \wRegOut_4_10[11] , 
        \wRegOut_4_10[10] , \wRegOut_4_10[9] , \wRegOut_4_10[8] , 
        \wRegOut_4_10[7] , \wRegOut_4_10[6] , \wRegOut_4_10[5] , 
        \wRegOut_4_10[4] , \wRegOut_4_10[3] , \wRegOut_4_10[2] , 
        \wRegOut_4_10[1] , \wRegOut_4_10[0] }), .L_Out({\wRegInTop_4_10[31] , 
        \wRegInTop_4_10[30] , \wRegInTop_4_10[29] , \wRegInTop_4_10[28] , 
        \wRegInTop_4_10[27] , \wRegInTop_4_10[26] , \wRegInTop_4_10[25] , 
        \wRegInTop_4_10[24] , \wRegInTop_4_10[23] , \wRegInTop_4_10[22] , 
        \wRegInTop_4_10[21] , \wRegInTop_4_10[20] , \wRegInTop_4_10[19] , 
        \wRegInTop_4_10[18] , \wRegInTop_4_10[17] , \wRegInTop_4_10[16] , 
        \wRegInTop_4_10[15] , \wRegInTop_4_10[14] , \wRegInTop_4_10[13] , 
        \wRegInTop_4_10[12] , \wRegInTop_4_10[11] , \wRegInTop_4_10[10] , 
        \wRegInTop_4_10[9] , \wRegInTop_4_10[8] , \wRegInTop_4_10[7] , 
        \wRegInTop_4_10[6] , \wRegInTop_4_10[5] , \wRegInTop_4_10[4] , 
        \wRegInTop_4_10[3] , \wRegInTop_4_10[2] , \wRegInTop_4_10[1] , 
        \wRegInTop_4_10[0] }), .R_WR(\wRegEnTop_4_11[0] ), .R_In({
        \wRegOut_4_11[31] , \wRegOut_4_11[30] , \wRegOut_4_11[29] , 
        \wRegOut_4_11[28] , \wRegOut_4_11[27] , \wRegOut_4_11[26] , 
        \wRegOut_4_11[25] , \wRegOut_4_11[24] , \wRegOut_4_11[23] , 
        \wRegOut_4_11[22] , \wRegOut_4_11[21] , \wRegOut_4_11[20] , 
        \wRegOut_4_11[19] , \wRegOut_4_11[18] , \wRegOut_4_11[17] , 
        \wRegOut_4_11[16] , \wRegOut_4_11[15] , \wRegOut_4_11[14] , 
        \wRegOut_4_11[13] , \wRegOut_4_11[12] , \wRegOut_4_11[11] , 
        \wRegOut_4_11[10] , \wRegOut_4_11[9] , \wRegOut_4_11[8] , 
        \wRegOut_4_11[7] , \wRegOut_4_11[6] , \wRegOut_4_11[5] , 
        \wRegOut_4_11[4] , \wRegOut_4_11[3] , \wRegOut_4_11[2] , 
        \wRegOut_4_11[1] , \wRegOut_4_11[0] }), .R_Out({\wRegInTop_4_11[31] , 
        \wRegInTop_4_11[30] , \wRegInTop_4_11[29] , \wRegInTop_4_11[28] , 
        \wRegInTop_4_11[27] , \wRegInTop_4_11[26] , \wRegInTop_4_11[25] , 
        \wRegInTop_4_11[24] , \wRegInTop_4_11[23] , \wRegInTop_4_11[22] , 
        \wRegInTop_4_11[21] , \wRegInTop_4_11[20] , \wRegInTop_4_11[19] , 
        \wRegInTop_4_11[18] , \wRegInTop_4_11[17] , \wRegInTop_4_11[16] , 
        \wRegInTop_4_11[15] , \wRegInTop_4_11[14] , \wRegInTop_4_11[13] , 
        \wRegInTop_4_11[12] , \wRegInTop_4_11[11] , \wRegInTop_4_11[10] , 
        \wRegInTop_4_11[9] , \wRegInTop_4_11[8] , \wRegInTop_4_11[7] , 
        \wRegInTop_4_11[6] , \wRegInTop_4_11[5] , \wRegInTop_4_11[4] , 
        \wRegInTop_4_11[3] , \wRegInTop_4_11[2] , \wRegInTop_4_11[1] , 
        \wRegInTop_4_11[0] }) );
    BHeap_Node_WIDTH32 BHN_6_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_3[0] ), .P_In({\wRegOut_6_3[31] , 
        \wRegOut_6_3[30] , \wRegOut_6_3[29] , \wRegOut_6_3[28] , 
        \wRegOut_6_3[27] , \wRegOut_6_3[26] , \wRegOut_6_3[25] , 
        \wRegOut_6_3[24] , \wRegOut_6_3[23] , \wRegOut_6_3[22] , 
        \wRegOut_6_3[21] , \wRegOut_6_3[20] , \wRegOut_6_3[19] , 
        \wRegOut_6_3[18] , \wRegOut_6_3[17] , \wRegOut_6_3[16] , 
        \wRegOut_6_3[15] , \wRegOut_6_3[14] , \wRegOut_6_3[13] , 
        \wRegOut_6_3[12] , \wRegOut_6_3[11] , \wRegOut_6_3[10] , 
        \wRegOut_6_3[9] , \wRegOut_6_3[8] , \wRegOut_6_3[7] , \wRegOut_6_3[6] , 
        \wRegOut_6_3[5] , \wRegOut_6_3[4] , \wRegOut_6_3[3] , \wRegOut_6_3[2] , 
        \wRegOut_6_3[1] , \wRegOut_6_3[0] }), .P_Out({\wRegInBot_6_3[31] , 
        \wRegInBot_6_3[30] , \wRegInBot_6_3[29] , \wRegInBot_6_3[28] , 
        \wRegInBot_6_3[27] , \wRegInBot_6_3[26] , \wRegInBot_6_3[25] , 
        \wRegInBot_6_3[24] , \wRegInBot_6_3[23] , \wRegInBot_6_3[22] , 
        \wRegInBot_6_3[21] , \wRegInBot_6_3[20] , \wRegInBot_6_3[19] , 
        \wRegInBot_6_3[18] , \wRegInBot_6_3[17] , \wRegInBot_6_3[16] , 
        \wRegInBot_6_3[15] , \wRegInBot_6_3[14] , \wRegInBot_6_3[13] , 
        \wRegInBot_6_3[12] , \wRegInBot_6_3[11] , \wRegInBot_6_3[10] , 
        \wRegInBot_6_3[9] , \wRegInBot_6_3[8] , \wRegInBot_6_3[7] , 
        \wRegInBot_6_3[6] , \wRegInBot_6_3[5] , \wRegInBot_6_3[4] , 
        \wRegInBot_6_3[3] , \wRegInBot_6_3[2] , \wRegInBot_6_3[1] , 
        \wRegInBot_6_3[0] }), .L_WR(\wRegEnTop_7_6[0] ), .L_In({
        \wRegOut_7_6[31] , \wRegOut_7_6[30] , \wRegOut_7_6[29] , 
        \wRegOut_7_6[28] , \wRegOut_7_6[27] , \wRegOut_7_6[26] , 
        \wRegOut_7_6[25] , \wRegOut_7_6[24] , \wRegOut_7_6[23] , 
        \wRegOut_7_6[22] , \wRegOut_7_6[21] , \wRegOut_7_6[20] , 
        \wRegOut_7_6[19] , \wRegOut_7_6[18] , \wRegOut_7_6[17] , 
        \wRegOut_7_6[16] , \wRegOut_7_6[15] , \wRegOut_7_6[14] , 
        \wRegOut_7_6[13] , \wRegOut_7_6[12] , \wRegOut_7_6[11] , 
        \wRegOut_7_6[10] , \wRegOut_7_6[9] , \wRegOut_7_6[8] , 
        \wRegOut_7_6[7] , \wRegOut_7_6[6] , \wRegOut_7_6[5] , \wRegOut_7_6[4] , 
        \wRegOut_7_6[3] , \wRegOut_7_6[2] , \wRegOut_7_6[1] , \wRegOut_7_6[0] 
        }), .L_Out({\wRegInTop_7_6[31] , \wRegInTop_7_6[30] , 
        \wRegInTop_7_6[29] , \wRegInTop_7_6[28] , \wRegInTop_7_6[27] , 
        \wRegInTop_7_6[26] , \wRegInTop_7_6[25] , \wRegInTop_7_6[24] , 
        \wRegInTop_7_6[23] , \wRegInTop_7_6[22] , \wRegInTop_7_6[21] , 
        \wRegInTop_7_6[20] , \wRegInTop_7_6[19] , \wRegInTop_7_6[18] , 
        \wRegInTop_7_6[17] , \wRegInTop_7_6[16] , \wRegInTop_7_6[15] , 
        \wRegInTop_7_6[14] , \wRegInTop_7_6[13] , \wRegInTop_7_6[12] , 
        \wRegInTop_7_6[11] , \wRegInTop_7_6[10] , \wRegInTop_7_6[9] , 
        \wRegInTop_7_6[8] , \wRegInTop_7_6[7] , \wRegInTop_7_6[6] , 
        \wRegInTop_7_6[5] , \wRegInTop_7_6[4] , \wRegInTop_7_6[3] , 
        \wRegInTop_7_6[2] , \wRegInTop_7_6[1] , \wRegInTop_7_6[0] }), .R_WR(
        \wRegEnTop_7_7[0] ), .R_In({\wRegOut_7_7[31] , \wRegOut_7_7[30] , 
        \wRegOut_7_7[29] , \wRegOut_7_7[28] , \wRegOut_7_7[27] , 
        \wRegOut_7_7[26] , \wRegOut_7_7[25] , \wRegOut_7_7[24] , 
        \wRegOut_7_7[23] , \wRegOut_7_7[22] , \wRegOut_7_7[21] , 
        \wRegOut_7_7[20] , \wRegOut_7_7[19] , \wRegOut_7_7[18] , 
        \wRegOut_7_7[17] , \wRegOut_7_7[16] , \wRegOut_7_7[15] , 
        \wRegOut_7_7[14] , \wRegOut_7_7[13] , \wRegOut_7_7[12] , 
        \wRegOut_7_7[11] , \wRegOut_7_7[10] , \wRegOut_7_7[9] , 
        \wRegOut_7_7[8] , \wRegOut_7_7[7] , \wRegOut_7_7[6] , \wRegOut_7_7[5] , 
        \wRegOut_7_7[4] , \wRegOut_7_7[3] , \wRegOut_7_7[2] , \wRegOut_7_7[1] , 
        \wRegOut_7_7[0] }), .R_Out({\wRegInTop_7_7[31] , \wRegInTop_7_7[30] , 
        \wRegInTop_7_7[29] , \wRegInTop_7_7[28] , \wRegInTop_7_7[27] , 
        \wRegInTop_7_7[26] , \wRegInTop_7_7[25] , \wRegInTop_7_7[24] , 
        \wRegInTop_7_7[23] , \wRegInTop_7_7[22] , \wRegInTop_7_7[21] , 
        \wRegInTop_7_7[20] , \wRegInTop_7_7[19] , \wRegInTop_7_7[18] , 
        \wRegInTop_7_7[17] , \wRegInTop_7_7[16] , \wRegInTop_7_7[15] , 
        \wRegInTop_7_7[14] , \wRegInTop_7_7[13] , \wRegInTop_7_7[12] , 
        \wRegInTop_7_7[11] , \wRegInTop_7_7[10] , \wRegInTop_7_7[9] , 
        \wRegInTop_7_7[8] , \wRegInTop_7_7[7] , \wRegInTop_7_7[6] , 
        \wRegInTop_7_7[5] , \wRegInTop_7_7[4] , \wRegInTop_7_7[3] , 
        \wRegInTop_7_7[2] , \wRegInTop_7_7[1] , \wRegInTop_7_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_47 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink175[31] , \ScanLink175[30] , \ScanLink175[29] , 
        \ScanLink175[28] , \ScanLink175[27] , \ScanLink175[26] , 
        \ScanLink175[25] , \ScanLink175[24] , \ScanLink175[23] , 
        \ScanLink175[22] , \ScanLink175[21] , \ScanLink175[20] , 
        \ScanLink175[19] , \ScanLink175[18] , \ScanLink175[17] , 
        \ScanLink175[16] , \ScanLink175[15] , \ScanLink175[14] , 
        \ScanLink175[13] , \ScanLink175[12] , \ScanLink175[11] , 
        \ScanLink175[10] , \ScanLink175[9] , \ScanLink175[8] , 
        \ScanLink175[7] , \ScanLink175[6] , \ScanLink175[5] , \ScanLink175[4] , 
        \ScanLink175[3] , \ScanLink175[2] , \ScanLink175[1] , \ScanLink175[0] 
        }), .ScanOut({\ScanLink174[31] , \ScanLink174[30] , \ScanLink174[29] , 
        \ScanLink174[28] , \ScanLink174[27] , \ScanLink174[26] , 
        \ScanLink174[25] , \ScanLink174[24] , \ScanLink174[23] , 
        \ScanLink174[22] , \ScanLink174[21] , \ScanLink174[20] , 
        \ScanLink174[19] , \ScanLink174[18] , \ScanLink174[17] , 
        \ScanLink174[16] , \ScanLink174[15] , \ScanLink174[14] , 
        \ScanLink174[13] , \ScanLink174[12] , \ScanLink174[11] , 
        \ScanLink174[10] , \ScanLink174[9] , \ScanLink174[8] , 
        \ScanLink174[7] , \ScanLink174[6] , \ScanLink174[5] , \ScanLink174[4] , 
        \ScanLink174[3] , \ScanLink174[2] , \ScanLink174[1] , \ScanLink174[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_47[31] , 
        \wRegOut_7_47[30] , \wRegOut_7_47[29] , \wRegOut_7_47[28] , 
        \wRegOut_7_47[27] , \wRegOut_7_47[26] , \wRegOut_7_47[25] , 
        \wRegOut_7_47[24] , \wRegOut_7_47[23] , \wRegOut_7_47[22] , 
        \wRegOut_7_47[21] , \wRegOut_7_47[20] , \wRegOut_7_47[19] , 
        \wRegOut_7_47[18] , \wRegOut_7_47[17] , \wRegOut_7_47[16] , 
        \wRegOut_7_47[15] , \wRegOut_7_47[14] , \wRegOut_7_47[13] , 
        \wRegOut_7_47[12] , \wRegOut_7_47[11] , \wRegOut_7_47[10] , 
        \wRegOut_7_47[9] , \wRegOut_7_47[8] , \wRegOut_7_47[7] , 
        \wRegOut_7_47[6] , \wRegOut_7_47[5] , \wRegOut_7_47[4] , 
        \wRegOut_7_47[3] , \wRegOut_7_47[2] , \wRegOut_7_47[1] , 
        \wRegOut_7_47[0] }), .Enable1(\wRegEnTop_7_47[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_47[31] , \wRegInTop_7_47[30] , \wRegInTop_7_47[29] , 
        \wRegInTop_7_47[28] , \wRegInTop_7_47[27] , \wRegInTop_7_47[26] , 
        \wRegInTop_7_47[25] , \wRegInTop_7_47[24] , \wRegInTop_7_47[23] , 
        \wRegInTop_7_47[22] , \wRegInTop_7_47[21] , \wRegInTop_7_47[20] , 
        \wRegInTop_7_47[19] , \wRegInTop_7_47[18] , \wRegInTop_7_47[17] , 
        \wRegInTop_7_47[16] , \wRegInTop_7_47[15] , \wRegInTop_7_47[14] , 
        \wRegInTop_7_47[13] , \wRegInTop_7_47[12] , \wRegInTop_7_47[11] , 
        \wRegInTop_7_47[10] , \wRegInTop_7_47[9] , \wRegInTop_7_47[8] , 
        \wRegInTop_7_47[7] , \wRegInTop_7_47[6] , \wRegInTop_7_47[5] , 
        \wRegInTop_7_47[4] , \wRegInTop_7_47[3] , \wRegInTop_7_47[2] , 
        \wRegInTop_7_47[1] , \wRegInTop_7_47[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink78[31] , \ScanLink78[30] , \ScanLink78[29] , 
        \ScanLink78[28] , \ScanLink78[27] , \ScanLink78[26] , \ScanLink78[25] , 
        \ScanLink78[24] , \ScanLink78[23] , \ScanLink78[22] , \ScanLink78[21] , 
        \ScanLink78[20] , \ScanLink78[19] , \ScanLink78[18] , \ScanLink78[17] , 
        \ScanLink78[16] , \ScanLink78[15] , \ScanLink78[14] , \ScanLink78[13] , 
        \ScanLink78[12] , \ScanLink78[11] , \ScanLink78[10] , \ScanLink78[9] , 
        \ScanLink78[8] , \ScanLink78[7] , \ScanLink78[6] , \ScanLink78[5] , 
        \ScanLink78[4] , \ScanLink78[3] , \ScanLink78[2] , \ScanLink78[1] , 
        \ScanLink78[0] }), .ScanOut({\ScanLink77[31] , \ScanLink77[30] , 
        \ScanLink77[29] , \ScanLink77[28] , \ScanLink77[27] , \ScanLink77[26] , 
        \ScanLink77[25] , \ScanLink77[24] , \ScanLink77[23] , \ScanLink77[22] , 
        \ScanLink77[21] , \ScanLink77[20] , \ScanLink77[19] , \ScanLink77[18] , 
        \ScanLink77[17] , \ScanLink77[16] , \ScanLink77[15] , \ScanLink77[14] , 
        \ScanLink77[13] , \ScanLink77[12] , \ScanLink77[11] , \ScanLink77[10] , 
        \ScanLink77[9] , \ScanLink77[8] , \ScanLink77[7] , \ScanLink77[6] , 
        \ScanLink77[5] , \ScanLink77[4] , \ScanLink77[3] , \ScanLink77[2] , 
        \ScanLink77[1] , \ScanLink77[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_14[31] , \wRegOut_6_14[30] , 
        \wRegOut_6_14[29] , \wRegOut_6_14[28] , \wRegOut_6_14[27] , 
        \wRegOut_6_14[26] , \wRegOut_6_14[25] , \wRegOut_6_14[24] , 
        \wRegOut_6_14[23] , \wRegOut_6_14[22] , \wRegOut_6_14[21] , 
        \wRegOut_6_14[20] , \wRegOut_6_14[19] , \wRegOut_6_14[18] , 
        \wRegOut_6_14[17] , \wRegOut_6_14[16] , \wRegOut_6_14[15] , 
        \wRegOut_6_14[14] , \wRegOut_6_14[13] , \wRegOut_6_14[12] , 
        \wRegOut_6_14[11] , \wRegOut_6_14[10] , \wRegOut_6_14[9] , 
        \wRegOut_6_14[8] , \wRegOut_6_14[7] , \wRegOut_6_14[6] , 
        \wRegOut_6_14[5] , \wRegOut_6_14[4] , \wRegOut_6_14[3] , 
        \wRegOut_6_14[2] , \wRegOut_6_14[1] , \wRegOut_6_14[0] }), .Enable1(
        \wRegEnTop_6_14[0] ), .Enable2(\wRegEnBot_6_14[0] ), .In1({
        \wRegInTop_6_14[31] , \wRegInTop_6_14[30] , \wRegInTop_6_14[29] , 
        \wRegInTop_6_14[28] , \wRegInTop_6_14[27] , \wRegInTop_6_14[26] , 
        \wRegInTop_6_14[25] , \wRegInTop_6_14[24] , \wRegInTop_6_14[23] , 
        \wRegInTop_6_14[22] , \wRegInTop_6_14[21] , \wRegInTop_6_14[20] , 
        \wRegInTop_6_14[19] , \wRegInTop_6_14[18] , \wRegInTop_6_14[17] , 
        \wRegInTop_6_14[16] , \wRegInTop_6_14[15] , \wRegInTop_6_14[14] , 
        \wRegInTop_6_14[13] , \wRegInTop_6_14[12] , \wRegInTop_6_14[11] , 
        \wRegInTop_6_14[10] , \wRegInTop_6_14[9] , \wRegInTop_6_14[8] , 
        \wRegInTop_6_14[7] , \wRegInTop_6_14[6] , \wRegInTop_6_14[5] , 
        \wRegInTop_6_14[4] , \wRegInTop_6_14[3] , \wRegInTop_6_14[2] , 
        \wRegInTop_6_14[1] , \wRegInTop_6_14[0] }), .In2({\wRegInBot_6_14[31] , 
        \wRegInBot_6_14[30] , \wRegInBot_6_14[29] , \wRegInBot_6_14[28] , 
        \wRegInBot_6_14[27] , \wRegInBot_6_14[26] , \wRegInBot_6_14[25] , 
        \wRegInBot_6_14[24] , \wRegInBot_6_14[23] , \wRegInBot_6_14[22] , 
        \wRegInBot_6_14[21] , \wRegInBot_6_14[20] , \wRegInBot_6_14[19] , 
        \wRegInBot_6_14[18] , \wRegInBot_6_14[17] , \wRegInBot_6_14[16] , 
        \wRegInBot_6_14[15] , \wRegInBot_6_14[14] , \wRegInBot_6_14[13] , 
        \wRegInBot_6_14[12] , \wRegInBot_6_14[11] , \wRegInBot_6_14[10] , 
        \wRegInBot_6_14[9] , \wRegInBot_6_14[8] , \wRegInBot_6_14[7] , 
        \wRegInBot_6_14[6] , \wRegInBot_6_14[5] , \wRegInBot_6_14[4] , 
        \wRegInBot_6_14[3] , \wRegInBot_6_14[2] , \wRegInBot_6_14[1] , 
        \wRegInBot_6_14[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_60 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink188[31] , \ScanLink188[30] , \ScanLink188[29] , 
        \ScanLink188[28] , \ScanLink188[27] , \ScanLink188[26] , 
        \ScanLink188[25] , \ScanLink188[24] , \ScanLink188[23] , 
        \ScanLink188[22] , \ScanLink188[21] , \ScanLink188[20] , 
        \ScanLink188[19] , \ScanLink188[18] , \ScanLink188[17] , 
        \ScanLink188[16] , \ScanLink188[15] , \ScanLink188[14] , 
        \ScanLink188[13] , \ScanLink188[12] , \ScanLink188[11] , 
        \ScanLink188[10] , \ScanLink188[9] , \ScanLink188[8] , 
        \ScanLink188[7] , \ScanLink188[6] , \ScanLink188[5] , \ScanLink188[4] , 
        \ScanLink188[3] , \ScanLink188[2] , \ScanLink188[1] , \ScanLink188[0] 
        }), .ScanOut({\ScanLink187[31] , \ScanLink187[30] , \ScanLink187[29] , 
        \ScanLink187[28] , \ScanLink187[27] , \ScanLink187[26] , 
        \ScanLink187[25] , \ScanLink187[24] , \ScanLink187[23] , 
        \ScanLink187[22] , \ScanLink187[21] , \ScanLink187[20] , 
        \ScanLink187[19] , \ScanLink187[18] , \ScanLink187[17] , 
        \ScanLink187[16] , \ScanLink187[15] , \ScanLink187[14] , 
        \ScanLink187[13] , \ScanLink187[12] , \ScanLink187[11] , 
        \ScanLink187[10] , \ScanLink187[9] , \ScanLink187[8] , 
        \ScanLink187[7] , \ScanLink187[6] , \ScanLink187[5] , \ScanLink187[4] , 
        \ScanLink187[3] , \ScanLink187[2] , \ScanLink187[1] , \ScanLink187[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_60[31] , 
        \wRegOut_7_60[30] , \wRegOut_7_60[29] , \wRegOut_7_60[28] , 
        \wRegOut_7_60[27] , \wRegOut_7_60[26] , \wRegOut_7_60[25] , 
        \wRegOut_7_60[24] , \wRegOut_7_60[23] , \wRegOut_7_60[22] , 
        \wRegOut_7_60[21] , \wRegOut_7_60[20] , \wRegOut_7_60[19] , 
        \wRegOut_7_60[18] , \wRegOut_7_60[17] , \wRegOut_7_60[16] , 
        \wRegOut_7_60[15] , \wRegOut_7_60[14] , \wRegOut_7_60[13] , 
        \wRegOut_7_60[12] , \wRegOut_7_60[11] , \wRegOut_7_60[10] , 
        \wRegOut_7_60[9] , \wRegOut_7_60[8] , \wRegOut_7_60[7] , 
        \wRegOut_7_60[6] , \wRegOut_7_60[5] , \wRegOut_7_60[4] , 
        \wRegOut_7_60[3] , \wRegOut_7_60[2] , \wRegOut_7_60[1] , 
        \wRegOut_7_60[0] }), .Enable1(\wRegEnTop_7_60[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_60[31] , \wRegInTop_7_60[30] , \wRegInTop_7_60[29] , 
        \wRegInTop_7_60[28] , \wRegInTop_7_60[27] , \wRegInTop_7_60[26] , 
        \wRegInTop_7_60[25] , \wRegInTop_7_60[24] , \wRegInTop_7_60[23] , 
        \wRegInTop_7_60[22] , \wRegInTop_7_60[21] , \wRegInTop_7_60[20] , 
        \wRegInTop_7_60[19] , \wRegInTop_7_60[18] , \wRegInTop_7_60[17] , 
        \wRegInTop_7_60[16] , \wRegInTop_7_60[15] , \wRegInTop_7_60[14] , 
        \wRegInTop_7_60[13] , \wRegInTop_7_60[12] , \wRegInTop_7_60[11] , 
        \wRegInTop_7_60[10] , \wRegInTop_7_60[9] , \wRegInTop_7_60[8] , 
        \wRegInTop_7_60[7] , \wRegInTop_7_60[6] , \wRegInTop_7_60[5] , 
        \wRegInTop_7_60[4] , \wRegInTop_7_60[3] , \wRegInTop_7_60[2] , 
        \wRegInTop_7_60[1] , \wRegInTop_7_60[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_55 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink183[31] , \ScanLink183[30] , \ScanLink183[29] , 
        \ScanLink183[28] , \ScanLink183[27] , \ScanLink183[26] , 
        \ScanLink183[25] , \ScanLink183[24] , \ScanLink183[23] , 
        \ScanLink183[22] , \ScanLink183[21] , \ScanLink183[20] , 
        \ScanLink183[19] , \ScanLink183[18] , \ScanLink183[17] , 
        \ScanLink183[16] , \ScanLink183[15] , \ScanLink183[14] , 
        \ScanLink183[13] , \ScanLink183[12] , \ScanLink183[11] , 
        \ScanLink183[10] , \ScanLink183[9] , \ScanLink183[8] , 
        \ScanLink183[7] , \ScanLink183[6] , \ScanLink183[5] , \ScanLink183[4] , 
        \ScanLink183[3] , \ScanLink183[2] , \ScanLink183[1] , \ScanLink183[0] 
        }), .ScanOut({\ScanLink182[31] , \ScanLink182[30] , \ScanLink182[29] , 
        \ScanLink182[28] , \ScanLink182[27] , \ScanLink182[26] , 
        \ScanLink182[25] , \ScanLink182[24] , \ScanLink182[23] , 
        \ScanLink182[22] , \ScanLink182[21] , \ScanLink182[20] , 
        \ScanLink182[19] , \ScanLink182[18] , \ScanLink182[17] , 
        \ScanLink182[16] , \ScanLink182[15] , \ScanLink182[14] , 
        \ScanLink182[13] , \ScanLink182[12] , \ScanLink182[11] , 
        \ScanLink182[10] , \ScanLink182[9] , \ScanLink182[8] , 
        \ScanLink182[7] , \ScanLink182[6] , \ScanLink182[5] , \ScanLink182[4] , 
        \ScanLink182[3] , \ScanLink182[2] , \ScanLink182[1] , \ScanLink182[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_55[31] , 
        \wRegOut_7_55[30] , \wRegOut_7_55[29] , \wRegOut_7_55[28] , 
        \wRegOut_7_55[27] , \wRegOut_7_55[26] , \wRegOut_7_55[25] , 
        \wRegOut_7_55[24] , \wRegOut_7_55[23] , \wRegOut_7_55[22] , 
        \wRegOut_7_55[21] , \wRegOut_7_55[20] , \wRegOut_7_55[19] , 
        \wRegOut_7_55[18] , \wRegOut_7_55[17] , \wRegOut_7_55[16] , 
        \wRegOut_7_55[15] , \wRegOut_7_55[14] , \wRegOut_7_55[13] , 
        \wRegOut_7_55[12] , \wRegOut_7_55[11] , \wRegOut_7_55[10] , 
        \wRegOut_7_55[9] , \wRegOut_7_55[8] , \wRegOut_7_55[7] , 
        \wRegOut_7_55[6] , \wRegOut_7_55[5] , \wRegOut_7_55[4] , 
        \wRegOut_7_55[3] , \wRegOut_7_55[2] , \wRegOut_7_55[1] , 
        \wRegOut_7_55[0] }), .Enable1(\wRegEnTop_7_55[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_55[31] , \wRegInTop_7_55[30] , \wRegInTop_7_55[29] , 
        \wRegInTop_7_55[28] , \wRegInTop_7_55[27] , \wRegInTop_7_55[26] , 
        \wRegInTop_7_55[25] , \wRegInTop_7_55[24] , \wRegInTop_7_55[23] , 
        \wRegInTop_7_55[22] , \wRegInTop_7_55[21] , \wRegInTop_7_55[20] , 
        \wRegInTop_7_55[19] , \wRegInTop_7_55[18] , \wRegInTop_7_55[17] , 
        \wRegInTop_7_55[16] , \wRegInTop_7_55[15] , \wRegInTop_7_55[14] , 
        \wRegInTop_7_55[13] , \wRegInTop_7_55[12] , \wRegInTop_7_55[11] , 
        \wRegInTop_7_55[10] , \wRegInTop_7_55[9] , \wRegInTop_7_55[8] , 
        \wRegInTop_7_55[7] , \wRegInTop_7_55[6] , \wRegInTop_7_55[5] , 
        \wRegInTop_7_55[4] , \wRegInTop_7_55[3] , \wRegInTop_7_55[2] , 
        \wRegInTop_7_55[1] , \wRegInTop_7_55[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_21 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink85[31] , \ScanLink85[30] , \ScanLink85[29] , 
        \ScanLink85[28] , \ScanLink85[27] , \ScanLink85[26] , \ScanLink85[25] , 
        \ScanLink85[24] , \ScanLink85[23] , \ScanLink85[22] , \ScanLink85[21] , 
        \ScanLink85[20] , \ScanLink85[19] , \ScanLink85[18] , \ScanLink85[17] , 
        \ScanLink85[16] , \ScanLink85[15] , \ScanLink85[14] , \ScanLink85[13] , 
        \ScanLink85[12] , \ScanLink85[11] , \ScanLink85[10] , \ScanLink85[9] , 
        \ScanLink85[8] , \ScanLink85[7] , \ScanLink85[6] , \ScanLink85[5] , 
        \ScanLink85[4] , \ScanLink85[3] , \ScanLink85[2] , \ScanLink85[1] , 
        \ScanLink85[0] }), .ScanOut({\ScanLink84[31] , \ScanLink84[30] , 
        \ScanLink84[29] , \ScanLink84[28] , \ScanLink84[27] , \ScanLink84[26] , 
        \ScanLink84[25] , \ScanLink84[24] , \ScanLink84[23] , \ScanLink84[22] , 
        \ScanLink84[21] , \ScanLink84[20] , \ScanLink84[19] , \ScanLink84[18] , 
        \ScanLink84[17] , \ScanLink84[16] , \ScanLink84[15] , \ScanLink84[14] , 
        \ScanLink84[13] , \ScanLink84[12] , \ScanLink84[11] , \ScanLink84[10] , 
        \ScanLink84[9] , \ScanLink84[8] , \ScanLink84[7] , \ScanLink84[6] , 
        \ScanLink84[5] , \ScanLink84[4] , \ScanLink84[3] , \ScanLink84[2] , 
        \ScanLink84[1] , \ScanLink84[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_21[31] , \wRegOut_6_21[30] , 
        \wRegOut_6_21[29] , \wRegOut_6_21[28] , \wRegOut_6_21[27] , 
        \wRegOut_6_21[26] , \wRegOut_6_21[25] , \wRegOut_6_21[24] , 
        \wRegOut_6_21[23] , \wRegOut_6_21[22] , \wRegOut_6_21[21] , 
        \wRegOut_6_21[20] , \wRegOut_6_21[19] , \wRegOut_6_21[18] , 
        \wRegOut_6_21[17] , \wRegOut_6_21[16] , \wRegOut_6_21[15] , 
        \wRegOut_6_21[14] , \wRegOut_6_21[13] , \wRegOut_6_21[12] , 
        \wRegOut_6_21[11] , \wRegOut_6_21[10] , \wRegOut_6_21[9] , 
        \wRegOut_6_21[8] , \wRegOut_6_21[7] , \wRegOut_6_21[6] , 
        \wRegOut_6_21[5] , \wRegOut_6_21[4] , \wRegOut_6_21[3] , 
        \wRegOut_6_21[2] , \wRegOut_6_21[1] , \wRegOut_6_21[0] }), .Enable1(
        \wRegEnTop_6_21[0] ), .Enable2(\wRegEnBot_6_21[0] ), .In1({
        \wRegInTop_6_21[31] , \wRegInTop_6_21[30] , \wRegInTop_6_21[29] , 
        \wRegInTop_6_21[28] , \wRegInTop_6_21[27] , \wRegInTop_6_21[26] , 
        \wRegInTop_6_21[25] , \wRegInTop_6_21[24] , \wRegInTop_6_21[23] , 
        \wRegInTop_6_21[22] , \wRegInTop_6_21[21] , \wRegInTop_6_21[20] , 
        \wRegInTop_6_21[19] , \wRegInTop_6_21[18] , \wRegInTop_6_21[17] , 
        \wRegInTop_6_21[16] , \wRegInTop_6_21[15] , \wRegInTop_6_21[14] , 
        \wRegInTop_6_21[13] , \wRegInTop_6_21[12] , \wRegInTop_6_21[11] , 
        \wRegInTop_6_21[10] , \wRegInTop_6_21[9] , \wRegInTop_6_21[8] , 
        \wRegInTop_6_21[7] , \wRegInTop_6_21[6] , \wRegInTop_6_21[5] , 
        \wRegInTop_6_21[4] , \wRegInTop_6_21[3] , \wRegInTop_6_21[2] , 
        \wRegInTop_6_21[1] , \wRegInTop_6_21[0] }), .In2({\wRegInBot_6_21[31] , 
        \wRegInBot_6_21[30] , \wRegInBot_6_21[29] , \wRegInBot_6_21[28] , 
        \wRegInBot_6_21[27] , \wRegInBot_6_21[26] , \wRegInBot_6_21[25] , 
        \wRegInBot_6_21[24] , \wRegInBot_6_21[23] , \wRegInBot_6_21[22] , 
        \wRegInBot_6_21[21] , \wRegInBot_6_21[20] , \wRegInBot_6_21[19] , 
        \wRegInBot_6_21[18] , \wRegInBot_6_21[17] , \wRegInBot_6_21[16] , 
        \wRegInBot_6_21[15] , \wRegInBot_6_21[14] , \wRegInBot_6_21[13] , 
        \wRegInBot_6_21[12] , \wRegInBot_6_21[11] , \wRegInBot_6_21[10] , 
        \wRegInBot_6_21[9] , \wRegInBot_6_21[8] , \wRegInBot_6_21[7] , 
        \wRegInBot_6_21[6] , \wRegInBot_6_21[5] , \wRegInBot_6_21[4] , 
        \wRegInBot_6_21[3] , \wRegInBot_6_21[2] , \wRegInBot_6_21[1] , 
        \wRegInBot_6_21[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_72 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink200[31] , \ScanLink200[30] , \ScanLink200[29] , 
        \ScanLink200[28] , \ScanLink200[27] , \ScanLink200[26] , 
        \ScanLink200[25] , \ScanLink200[24] , \ScanLink200[23] , 
        \ScanLink200[22] , \ScanLink200[21] , \ScanLink200[20] , 
        \ScanLink200[19] , \ScanLink200[18] , \ScanLink200[17] , 
        \ScanLink200[16] , \ScanLink200[15] , \ScanLink200[14] , 
        \ScanLink200[13] , \ScanLink200[12] , \ScanLink200[11] , 
        \ScanLink200[10] , \ScanLink200[9] , \ScanLink200[8] , 
        \ScanLink200[7] , \ScanLink200[6] , \ScanLink200[5] , \ScanLink200[4] , 
        \ScanLink200[3] , \ScanLink200[2] , \ScanLink200[1] , \ScanLink200[0] 
        }), .ScanOut({\ScanLink199[31] , \ScanLink199[30] , \ScanLink199[29] , 
        \ScanLink199[28] , \ScanLink199[27] , \ScanLink199[26] , 
        \ScanLink199[25] , \ScanLink199[24] , \ScanLink199[23] , 
        \ScanLink199[22] , \ScanLink199[21] , \ScanLink199[20] , 
        \ScanLink199[19] , \ScanLink199[18] , \ScanLink199[17] , 
        \ScanLink199[16] , \ScanLink199[15] , \ScanLink199[14] , 
        \ScanLink199[13] , \ScanLink199[12] , \ScanLink199[11] , 
        \ScanLink199[10] , \ScanLink199[9] , \ScanLink199[8] , 
        \ScanLink199[7] , \ScanLink199[6] , \ScanLink199[5] , \ScanLink199[4] , 
        \ScanLink199[3] , \ScanLink199[2] , \ScanLink199[1] , \ScanLink199[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_72[31] , 
        \wRegOut_7_72[30] , \wRegOut_7_72[29] , \wRegOut_7_72[28] , 
        \wRegOut_7_72[27] , \wRegOut_7_72[26] , \wRegOut_7_72[25] , 
        \wRegOut_7_72[24] , \wRegOut_7_72[23] , \wRegOut_7_72[22] , 
        \wRegOut_7_72[21] , \wRegOut_7_72[20] , \wRegOut_7_72[19] , 
        \wRegOut_7_72[18] , \wRegOut_7_72[17] , \wRegOut_7_72[16] , 
        \wRegOut_7_72[15] , \wRegOut_7_72[14] , \wRegOut_7_72[13] , 
        \wRegOut_7_72[12] , \wRegOut_7_72[11] , \wRegOut_7_72[10] , 
        \wRegOut_7_72[9] , \wRegOut_7_72[8] , \wRegOut_7_72[7] , 
        \wRegOut_7_72[6] , \wRegOut_7_72[5] , \wRegOut_7_72[4] , 
        \wRegOut_7_72[3] , \wRegOut_7_72[2] , \wRegOut_7_72[1] , 
        \wRegOut_7_72[0] }), .Enable1(\wRegEnTop_7_72[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_72[31] , \wRegInTop_7_72[30] , \wRegInTop_7_72[29] , 
        \wRegInTop_7_72[28] , \wRegInTop_7_72[27] , \wRegInTop_7_72[26] , 
        \wRegInTop_7_72[25] , \wRegInTop_7_72[24] , \wRegInTop_7_72[23] , 
        \wRegInTop_7_72[22] , \wRegInTop_7_72[21] , \wRegInTop_7_72[20] , 
        \wRegInTop_7_72[19] , \wRegInTop_7_72[18] , \wRegInTop_7_72[17] , 
        \wRegInTop_7_72[16] , \wRegInTop_7_72[15] , \wRegInTop_7_72[14] , 
        \wRegInTop_7_72[13] , \wRegInTop_7_72[12] , \wRegInTop_7_72[11] , 
        \wRegInTop_7_72[10] , \wRegInTop_7_72[9] , \wRegInTop_7_72[8] , 
        \wRegInTop_7_72[7] , \wRegInTop_7_72[6] , \wRegInTop_7_72[5] , 
        \wRegInTop_7_72[4] , \wRegInTop_7_72[3] , \wRegInTop_7_72[2] , 
        \wRegInTop_7_72[1] , \wRegInTop_7_72[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink26[31] , \ScanLink26[30] , \ScanLink26[29] , 
        \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , \ScanLink26[25] , 
        \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , \ScanLink26[21] , 
        \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , \ScanLink26[17] , 
        \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , \ScanLink26[13] , 
        \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , \ScanLink26[9] , 
        \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , \ScanLink26[5] , 
        \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , \ScanLink26[1] , 
        \ScanLink26[0] }), .ScanOut({\ScanLink25[31] , \ScanLink25[30] , 
        \ScanLink25[29] , \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , 
        \ScanLink25[25] , \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , 
        \ScanLink25[21] , \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , 
        \ScanLink25[17] , \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , 
        \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , 
        \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , 
        \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , 
        \ScanLink25[1] , \ScanLink25[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_10[31] , \wRegOut_4_10[30] , 
        \wRegOut_4_10[29] , \wRegOut_4_10[28] , \wRegOut_4_10[27] , 
        \wRegOut_4_10[26] , \wRegOut_4_10[25] , \wRegOut_4_10[24] , 
        \wRegOut_4_10[23] , \wRegOut_4_10[22] , \wRegOut_4_10[21] , 
        \wRegOut_4_10[20] , \wRegOut_4_10[19] , \wRegOut_4_10[18] , 
        \wRegOut_4_10[17] , \wRegOut_4_10[16] , \wRegOut_4_10[15] , 
        \wRegOut_4_10[14] , \wRegOut_4_10[13] , \wRegOut_4_10[12] , 
        \wRegOut_4_10[11] , \wRegOut_4_10[10] , \wRegOut_4_10[9] , 
        \wRegOut_4_10[8] , \wRegOut_4_10[7] , \wRegOut_4_10[6] , 
        \wRegOut_4_10[5] , \wRegOut_4_10[4] , \wRegOut_4_10[3] , 
        \wRegOut_4_10[2] , \wRegOut_4_10[1] , \wRegOut_4_10[0] }), .Enable1(
        \wRegEnTop_4_10[0] ), .Enable2(\wRegEnBot_4_10[0] ), .In1({
        \wRegInTop_4_10[31] , \wRegInTop_4_10[30] , \wRegInTop_4_10[29] , 
        \wRegInTop_4_10[28] , \wRegInTop_4_10[27] , \wRegInTop_4_10[26] , 
        \wRegInTop_4_10[25] , \wRegInTop_4_10[24] , \wRegInTop_4_10[23] , 
        \wRegInTop_4_10[22] , \wRegInTop_4_10[21] , \wRegInTop_4_10[20] , 
        \wRegInTop_4_10[19] , \wRegInTop_4_10[18] , \wRegInTop_4_10[17] , 
        \wRegInTop_4_10[16] , \wRegInTop_4_10[15] , \wRegInTop_4_10[14] , 
        \wRegInTop_4_10[13] , \wRegInTop_4_10[12] , \wRegInTop_4_10[11] , 
        \wRegInTop_4_10[10] , \wRegInTop_4_10[9] , \wRegInTop_4_10[8] , 
        \wRegInTop_4_10[7] , \wRegInTop_4_10[6] , \wRegInTop_4_10[5] , 
        \wRegInTop_4_10[4] , \wRegInTop_4_10[3] , \wRegInTop_4_10[2] , 
        \wRegInTop_4_10[1] , \wRegInTop_4_10[0] }), .In2({\wRegInBot_4_10[31] , 
        \wRegInBot_4_10[30] , \wRegInBot_4_10[29] , \wRegInBot_4_10[28] , 
        \wRegInBot_4_10[27] , \wRegInBot_4_10[26] , \wRegInBot_4_10[25] , 
        \wRegInBot_4_10[24] , \wRegInBot_4_10[23] , \wRegInBot_4_10[22] , 
        \wRegInBot_4_10[21] , \wRegInBot_4_10[20] , \wRegInBot_4_10[19] , 
        \wRegInBot_4_10[18] , \wRegInBot_4_10[17] , \wRegInBot_4_10[16] , 
        \wRegInBot_4_10[15] , \wRegInBot_4_10[14] , \wRegInBot_4_10[13] , 
        \wRegInBot_4_10[12] , \wRegInBot_4_10[11] , \wRegInBot_4_10[10] , 
        \wRegInBot_4_10[9] , \wRegInBot_4_10[8] , \wRegInBot_4_10[7] , 
        \wRegInBot_4_10[6] , \wRegInBot_4_10[5] , \wRegInBot_4_10[4] , 
        \wRegInBot_4_10[3] , \wRegInBot_4_10[2] , \wRegInBot_4_10[1] , 
        \wRegInBot_4_10[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink72[31] , \ScanLink72[30] , \ScanLink72[29] , 
        \ScanLink72[28] , \ScanLink72[27] , \ScanLink72[26] , \ScanLink72[25] , 
        \ScanLink72[24] , \ScanLink72[23] , \ScanLink72[22] , \ScanLink72[21] , 
        \ScanLink72[20] , \ScanLink72[19] , \ScanLink72[18] , \ScanLink72[17] , 
        \ScanLink72[16] , \ScanLink72[15] , \ScanLink72[14] , \ScanLink72[13] , 
        \ScanLink72[12] , \ScanLink72[11] , \ScanLink72[10] , \ScanLink72[9] , 
        \ScanLink72[8] , \ScanLink72[7] , \ScanLink72[6] , \ScanLink72[5] , 
        \ScanLink72[4] , \ScanLink72[3] , \ScanLink72[2] , \ScanLink72[1] , 
        \ScanLink72[0] }), .ScanOut({\ScanLink71[31] , \ScanLink71[30] , 
        \ScanLink71[29] , \ScanLink71[28] , \ScanLink71[27] , \ScanLink71[26] , 
        \ScanLink71[25] , \ScanLink71[24] , \ScanLink71[23] , \ScanLink71[22] , 
        \ScanLink71[21] , \ScanLink71[20] , \ScanLink71[19] , \ScanLink71[18] , 
        \ScanLink71[17] , \ScanLink71[16] , \ScanLink71[15] , \ScanLink71[14] , 
        \ScanLink71[13] , \ScanLink71[12] , \ScanLink71[11] , \ScanLink71[10] , 
        \ScanLink71[9] , \ScanLink71[8] , \ScanLink71[7] , \ScanLink71[6] , 
        \ScanLink71[5] , \ScanLink71[4] , \ScanLink71[3] , \ScanLink71[2] , 
        \ScanLink71[1] , \ScanLink71[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_6_8[31] , \wRegOut_6_8[30] , \wRegOut_6_8[29] , 
        \wRegOut_6_8[28] , \wRegOut_6_8[27] , \wRegOut_6_8[26] , 
        \wRegOut_6_8[25] , \wRegOut_6_8[24] , \wRegOut_6_8[23] , 
        \wRegOut_6_8[22] , \wRegOut_6_8[21] , \wRegOut_6_8[20] , 
        \wRegOut_6_8[19] , \wRegOut_6_8[18] , \wRegOut_6_8[17] , 
        \wRegOut_6_8[16] , \wRegOut_6_8[15] , \wRegOut_6_8[14] , 
        \wRegOut_6_8[13] , \wRegOut_6_8[12] , \wRegOut_6_8[11] , 
        \wRegOut_6_8[10] , \wRegOut_6_8[9] , \wRegOut_6_8[8] , 
        \wRegOut_6_8[7] , \wRegOut_6_8[6] , \wRegOut_6_8[5] , \wRegOut_6_8[4] , 
        \wRegOut_6_8[3] , \wRegOut_6_8[2] , \wRegOut_6_8[1] , \wRegOut_6_8[0] 
        }), .Enable1(\wRegEnTop_6_8[0] ), .Enable2(\wRegEnBot_6_8[0] ), .In1({
        \wRegInTop_6_8[31] , \wRegInTop_6_8[30] , \wRegInTop_6_8[29] , 
        \wRegInTop_6_8[28] , \wRegInTop_6_8[27] , \wRegInTop_6_8[26] , 
        \wRegInTop_6_8[25] , \wRegInTop_6_8[24] , \wRegInTop_6_8[23] , 
        \wRegInTop_6_8[22] , \wRegInTop_6_8[21] , \wRegInTop_6_8[20] , 
        \wRegInTop_6_8[19] , \wRegInTop_6_8[18] , \wRegInTop_6_8[17] , 
        \wRegInTop_6_8[16] , \wRegInTop_6_8[15] , \wRegInTop_6_8[14] , 
        \wRegInTop_6_8[13] , \wRegInTop_6_8[12] , \wRegInTop_6_8[11] , 
        \wRegInTop_6_8[10] , \wRegInTop_6_8[9] , \wRegInTop_6_8[8] , 
        \wRegInTop_6_8[7] , \wRegInTop_6_8[6] , \wRegInTop_6_8[5] , 
        \wRegInTop_6_8[4] , \wRegInTop_6_8[3] , \wRegInTop_6_8[2] , 
        \wRegInTop_6_8[1] , \wRegInTop_6_8[0] }), .In2({\wRegInBot_6_8[31] , 
        \wRegInBot_6_8[30] , \wRegInBot_6_8[29] , \wRegInBot_6_8[28] , 
        \wRegInBot_6_8[27] , \wRegInBot_6_8[26] , \wRegInBot_6_8[25] , 
        \wRegInBot_6_8[24] , \wRegInBot_6_8[23] , \wRegInBot_6_8[22] , 
        \wRegInBot_6_8[21] , \wRegInBot_6_8[20] , \wRegInBot_6_8[19] , 
        \wRegInBot_6_8[18] , \wRegInBot_6_8[17] , \wRegInBot_6_8[16] , 
        \wRegInBot_6_8[15] , \wRegInBot_6_8[14] , \wRegInBot_6_8[13] , 
        \wRegInBot_6_8[12] , \wRegInBot_6_8[11] , \wRegInBot_6_8[10] , 
        \wRegInBot_6_8[9] , \wRegInBot_6_8[8] , \wRegInBot_6_8[7] , 
        \wRegInBot_6_8[6] , \wRegInBot_6_8[5] , \wRegInBot_6_8[4] , 
        \wRegInBot_6_8[3] , \wRegInBot_6_8[2] , \wRegInBot_6_8[1] , 
        \wRegInBot_6_8[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_6_54 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink118[31] , \ScanLink118[30] , \ScanLink118[29] , 
        \ScanLink118[28] , \ScanLink118[27] , \ScanLink118[26] , 
        \ScanLink118[25] , \ScanLink118[24] , \ScanLink118[23] , 
        \ScanLink118[22] , \ScanLink118[21] , \ScanLink118[20] , 
        \ScanLink118[19] , \ScanLink118[18] , \ScanLink118[17] , 
        \ScanLink118[16] , \ScanLink118[15] , \ScanLink118[14] , 
        \ScanLink118[13] , \ScanLink118[12] , \ScanLink118[11] , 
        \ScanLink118[10] , \ScanLink118[9] , \ScanLink118[8] , 
        \ScanLink118[7] , \ScanLink118[6] , \ScanLink118[5] , \ScanLink118[4] , 
        \ScanLink118[3] , \ScanLink118[2] , \ScanLink118[1] , \ScanLink118[0] 
        }), .ScanOut({\ScanLink117[31] , \ScanLink117[30] , \ScanLink117[29] , 
        \ScanLink117[28] , \ScanLink117[27] , \ScanLink117[26] , 
        \ScanLink117[25] , \ScanLink117[24] , \ScanLink117[23] , 
        \ScanLink117[22] , \ScanLink117[21] , \ScanLink117[20] , 
        \ScanLink117[19] , \ScanLink117[18] , \ScanLink117[17] , 
        \ScanLink117[16] , \ScanLink117[15] , \ScanLink117[14] , 
        \ScanLink117[13] , \ScanLink117[12] , \ScanLink117[11] , 
        \ScanLink117[10] , \ScanLink117[9] , \ScanLink117[8] , 
        \ScanLink117[7] , \ScanLink117[6] , \ScanLink117[5] , \ScanLink117[4] , 
        \ScanLink117[3] , \ScanLink117[2] , \ScanLink117[1] , \ScanLink117[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_6_54[31] , 
        \wRegOut_6_54[30] , \wRegOut_6_54[29] , \wRegOut_6_54[28] , 
        \wRegOut_6_54[27] , \wRegOut_6_54[26] , \wRegOut_6_54[25] , 
        \wRegOut_6_54[24] , \wRegOut_6_54[23] , \wRegOut_6_54[22] , 
        \wRegOut_6_54[21] , \wRegOut_6_54[20] , \wRegOut_6_54[19] , 
        \wRegOut_6_54[18] , \wRegOut_6_54[17] , \wRegOut_6_54[16] , 
        \wRegOut_6_54[15] , \wRegOut_6_54[14] , \wRegOut_6_54[13] , 
        \wRegOut_6_54[12] , \wRegOut_6_54[11] , \wRegOut_6_54[10] , 
        \wRegOut_6_54[9] , \wRegOut_6_54[8] , \wRegOut_6_54[7] , 
        \wRegOut_6_54[6] , \wRegOut_6_54[5] , \wRegOut_6_54[4] , 
        \wRegOut_6_54[3] , \wRegOut_6_54[2] , \wRegOut_6_54[1] , 
        \wRegOut_6_54[0] }), .Enable1(\wRegEnTop_6_54[0] ), .Enable2(
        \wRegEnBot_6_54[0] ), .In1({\wRegInTop_6_54[31] , \wRegInTop_6_54[30] , 
        \wRegInTop_6_54[29] , \wRegInTop_6_54[28] , \wRegInTop_6_54[27] , 
        \wRegInTop_6_54[26] , \wRegInTop_6_54[25] , \wRegInTop_6_54[24] , 
        \wRegInTop_6_54[23] , \wRegInTop_6_54[22] , \wRegInTop_6_54[21] , 
        \wRegInTop_6_54[20] , \wRegInTop_6_54[19] , \wRegInTop_6_54[18] , 
        \wRegInTop_6_54[17] , \wRegInTop_6_54[16] , \wRegInTop_6_54[15] , 
        \wRegInTop_6_54[14] , \wRegInTop_6_54[13] , \wRegInTop_6_54[12] , 
        \wRegInTop_6_54[11] , \wRegInTop_6_54[10] , \wRegInTop_6_54[9] , 
        \wRegInTop_6_54[8] , \wRegInTop_6_54[7] , \wRegInTop_6_54[6] , 
        \wRegInTop_6_54[5] , \wRegInTop_6_54[4] , \wRegInTop_6_54[3] , 
        \wRegInTop_6_54[2] , \wRegInTop_6_54[1] , \wRegInTop_6_54[0] }), .In2(
        {\wRegInBot_6_54[31] , \wRegInBot_6_54[30] , \wRegInBot_6_54[29] , 
        \wRegInBot_6_54[28] , \wRegInBot_6_54[27] , \wRegInBot_6_54[26] , 
        \wRegInBot_6_54[25] , \wRegInBot_6_54[24] , \wRegInBot_6_54[23] , 
        \wRegInBot_6_54[22] , \wRegInBot_6_54[21] , \wRegInBot_6_54[20] , 
        \wRegInBot_6_54[19] , \wRegInBot_6_54[18] , \wRegInBot_6_54[17] , 
        \wRegInBot_6_54[16] , \wRegInBot_6_54[15] , \wRegInBot_6_54[14] , 
        \wRegInBot_6_54[13] , \wRegInBot_6_54[12] , \wRegInBot_6_54[11] , 
        \wRegInBot_6_54[10] , \wRegInBot_6_54[9] , \wRegInBot_6_54[8] , 
        \wRegInBot_6_54[7] , \wRegInBot_6_54[6] , \wRegInBot_6_54[5] , 
        \wRegInBot_6_54[4] , \wRegInBot_6_54[3] , \wRegInBot_6_54[2] , 
        \wRegInBot_6_54[1] , \wRegInBot_6_54[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_97 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink225[31] , \ScanLink225[30] , \ScanLink225[29] , 
        \ScanLink225[28] , \ScanLink225[27] , \ScanLink225[26] , 
        \ScanLink225[25] , \ScanLink225[24] , \ScanLink225[23] , 
        \ScanLink225[22] , \ScanLink225[21] , \ScanLink225[20] , 
        \ScanLink225[19] , \ScanLink225[18] , \ScanLink225[17] , 
        \ScanLink225[16] , \ScanLink225[15] , \ScanLink225[14] , 
        \ScanLink225[13] , \ScanLink225[12] , \ScanLink225[11] , 
        \ScanLink225[10] , \ScanLink225[9] , \ScanLink225[8] , 
        \ScanLink225[7] , \ScanLink225[6] , \ScanLink225[5] , \ScanLink225[4] , 
        \ScanLink225[3] , \ScanLink225[2] , \ScanLink225[1] , \ScanLink225[0] 
        }), .ScanOut({\ScanLink224[31] , \ScanLink224[30] , \ScanLink224[29] , 
        \ScanLink224[28] , \ScanLink224[27] , \ScanLink224[26] , 
        \ScanLink224[25] , \ScanLink224[24] , \ScanLink224[23] , 
        \ScanLink224[22] , \ScanLink224[21] , \ScanLink224[20] , 
        \ScanLink224[19] , \ScanLink224[18] , \ScanLink224[17] , 
        \ScanLink224[16] , \ScanLink224[15] , \ScanLink224[14] , 
        \ScanLink224[13] , \ScanLink224[12] , \ScanLink224[11] , 
        \ScanLink224[10] , \ScanLink224[9] , \ScanLink224[8] , 
        \ScanLink224[7] , \ScanLink224[6] , \ScanLink224[5] , \ScanLink224[4] , 
        \ScanLink224[3] , \ScanLink224[2] , \ScanLink224[1] , \ScanLink224[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_97[31] , 
        \wRegOut_7_97[30] , \wRegOut_7_97[29] , \wRegOut_7_97[28] , 
        \wRegOut_7_97[27] , \wRegOut_7_97[26] , \wRegOut_7_97[25] , 
        \wRegOut_7_97[24] , \wRegOut_7_97[23] , \wRegOut_7_97[22] , 
        \wRegOut_7_97[21] , \wRegOut_7_97[20] , \wRegOut_7_97[19] , 
        \wRegOut_7_97[18] , \wRegOut_7_97[17] , \wRegOut_7_97[16] , 
        \wRegOut_7_97[15] , \wRegOut_7_97[14] , \wRegOut_7_97[13] , 
        \wRegOut_7_97[12] , \wRegOut_7_97[11] , \wRegOut_7_97[10] , 
        \wRegOut_7_97[9] , \wRegOut_7_97[8] , \wRegOut_7_97[7] , 
        \wRegOut_7_97[6] , \wRegOut_7_97[5] , \wRegOut_7_97[4] , 
        \wRegOut_7_97[3] , \wRegOut_7_97[2] , \wRegOut_7_97[1] , 
        \wRegOut_7_97[0] }), .Enable1(\wRegEnTop_7_97[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_97[31] , \wRegInTop_7_97[30] , \wRegInTop_7_97[29] , 
        \wRegInTop_7_97[28] , \wRegInTop_7_97[27] , \wRegInTop_7_97[26] , 
        \wRegInTop_7_97[25] , \wRegInTop_7_97[24] , \wRegInTop_7_97[23] , 
        \wRegInTop_7_97[22] , \wRegInTop_7_97[21] , \wRegInTop_7_97[20] , 
        \wRegInTop_7_97[19] , \wRegInTop_7_97[18] , \wRegInTop_7_97[17] , 
        \wRegInTop_7_97[16] , \wRegInTop_7_97[15] , \wRegInTop_7_97[14] , 
        \wRegInTop_7_97[13] , \wRegInTop_7_97[12] , \wRegInTop_7_97[11] , 
        \wRegInTop_7_97[10] , \wRegInTop_7_97[9] , \wRegInTop_7_97[8] , 
        \wRegInTop_7_97[7] , \wRegInTop_7_97[6] , \wRegInTop_7_97[5] , 
        \wRegInTop_7_97[4] , \wRegInTop_7_97[3] , \wRegInTop_7_97[2] , 
        \wRegInTop_7_97[1] , \wRegInTop_7_97[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_108 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink236[31] , \ScanLink236[30] , \ScanLink236[29] , 
        \ScanLink236[28] , \ScanLink236[27] , \ScanLink236[26] , 
        \ScanLink236[25] , \ScanLink236[24] , \ScanLink236[23] , 
        \ScanLink236[22] , \ScanLink236[21] , \ScanLink236[20] , 
        \ScanLink236[19] , \ScanLink236[18] , \ScanLink236[17] , 
        \ScanLink236[16] , \ScanLink236[15] , \ScanLink236[14] , 
        \ScanLink236[13] , \ScanLink236[12] , \ScanLink236[11] , 
        \ScanLink236[10] , \ScanLink236[9] , \ScanLink236[8] , 
        \ScanLink236[7] , \ScanLink236[6] , \ScanLink236[5] , \ScanLink236[4] , 
        \ScanLink236[3] , \ScanLink236[2] , \ScanLink236[1] , \ScanLink236[0] 
        }), .ScanOut({\ScanLink235[31] , \ScanLink235[30] , \ScanLink235[29] , 
        \ScanLink235[28] , \ScanLink235[27] , \ScanLink235[26] , 
        \ScanLink235[25] , \ScanLink235[24] , \ScanLink235[23] , 
        \ScanLink235[22] , \ScanLink235[21] , \ScanLink235[20] , 
        \ScanLink235[19] , \ScanLink235[18] , \ScanLink235[17] , 
        \ScanLink235[16] , \ScanLink235[15] , \ScanLink235[14] , 
        \ScanLink235[13] , \ScanLink235[12] , \ScanLink235[11] , 
        \ScanLink235[10] , \ScanLink235[9] , \ScanLink235[8] , 
        \ScanLink235[7] , \ScanLink235[6] , \ScanLink235[5] , \ScanLink235[4] , 
        \ScanLink235[3] , \ScanLink235[2] , \ScanLink235[1] , \ScanLink235[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_108[31] , 
        \wRegOut_7_108[30] , \wRegOut_7_108[29] , \wRegOut_7_108[28] , 
        \wRegOut_7_108[27] , \wRegOut_7_108[26] , \wRegOut_7_108[25] , 
        \wRegOut_7_108[24] , \wRegOut_7_108[23] , \wRegOut_7_108[22] , 
        \wRegOut_7_108[21] , \wRegOut_7_108[20] , \wRegOut_7_108[19] , 
        \wRegOut_7_108[18] , \wRegOut_7_108[17] , \wRegOut_7_108[16] , 
        \wRegOut_7_108[15] , \wRegOut_7_108[14] , \wRegOut_7_108[13] , 
        \wRegOut_7_108[12] , \wRegOut_7_108[11] , \wRegOut_7_108[10] , 
        \wRegOut_7_108[9] , \wRegOut_7_108[8] , \wRegOut_7_108[7] , 
        \wRegOut_7_108[6] , \wRegOut_7_108[5] , \wRegOut_7_108[4] , 
        \wRegOut_7_108[3] , \wRegOut_7_108[2] , \wRegOut_7_108[1] , 
        \wRegOut_7_108[0] }), .Enable1(\wRegEnTop_7_108[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_108[31] , \wRegInTop_7_108[30] , 
        \wRegInTop_7_108[29] , \wRegInTop_7_108[28] , \wRegInTop_7_108[27] , 
        \wRegInTop_7_108[26] , \wRegInTop_7_108[25] , \wRegInTop_7_108[24] , 
        \wRegInTop_7_108[23] , \wRegInTop_7_108[22] , \wRegInTop_7_108[21] , 
        \wRegInTop_7_108[20] , \wRegInTop_7_108[19] , \wRegInTop_7_108[18] , 
        \wRegInTop_7_108[17] , \wRegInTop_7_108[16] , \wRegInTop_7_108[15] , 
        \wRegInTop_7_108[14] , \wRegInTop_7_108[13] , \wRegInTop_7_108[12] , 
        \wRegInTop_7_108[11] , \wRegInTop_7_108[10] , \wRegInTop_7_108[9] , 
        \wRegInTop_7_108[8] , \wRegInTop_7_108[7] , \wRegInTop_7_108[6] , 
        \wRegInTop_7_108[5] , \wRegInTop_7_108[4] , \wRegInTop_7_108[3] , 
        \wRegInTop_7_108[2] , \wRegInTop_7_108[1] , \wRegInTop_7_108[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_0_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_0[0] ), .P_WR(\wRegEnBot_0_0[0] ), .P_In({\wRegOut_0_0[31] , 
        \wRegOut_0_0[30] , \wRegOut_0_0[29] , \wRegOut_0_0[28] , 
        \wRegOut_0_0[27] , \wRegOut_0_0[26] , \wRegOut_0_0[25] , 
        \wRegOut_0_0[24] , \wRegOut_0_0[23] , \wRegOut_0_0[22] , 
        \wRegOut_0_0[21] , \wRegOut_0_0[20] , \wRegOut_0_0[19] , 
        \wRegOut_0_0[18] , \wRegOut_0_0[17] , \wRegOut_0_0[16] , 
        \wRegOut_0_0[15] , \wRegOut_0_0[14] , \wRegOut_0_0[13] , 
        \wRegOut_0_0[12] , \wRegOut_0_0[11] , \wRegOut_0_0[10] , 
        \wRegOut_0_0[9] , \wRegOut_0_0[8] , \wRegOut_0_0[7] , \wRegOut_0_0[6] , 
        \wRegOut_0_0[5] , \wRegOut_0_0[4] , \wRegOut_0_0[3] , \wRegOut_0_0[2] , 
        \wRegOut_0_0[1] , \wRegOut_0_0[0] }), .P_Out({\wRegInBot_0_0[31] , 
        \wRegInBot_0_0[30] , \wRegInBot_0_0[29] , \wRegInBot_0_0[28] , 
        \wRegInBot_0_0[27] , \wRegInBot_0_0[26] , \wRegInBot_0_0[25] , 
        \wRegInBot_0_0[24] , \wRegInBot_0_0[23] , \wRegInBot_0_0[22] , 
        \wRegInBot_0_0[21] , \wRegInBot_0_0[20] , \wRegInBot_0_0[19] , 
        \wRegInBot_0_0[18] , \wRegInBot_0_0[17] , \wRegInBot_0_0[16] , 
        \wRegInBot_0_0[15] , \wRegInBot_0_0[14] , \wRegInBot_0_0[13] , 
        \wRegInBot_0_0[12] , \wRegInBot_0_0[11] , \wRegInBot_0_0[10] , 
        \wRegInBot_0_0[9] , \wRegInBot_0_0[8] , \wRegInBot_0_0[7] , 
        \wRegInBot_0_0[6] , \wRegInBot_0_0[5] , \wRegInBot_0_0[4] , 
        \wRegInBot_0_0[3] , \wRegInBot_0_0[2] , \wRegInBot_0_0[1] , 
        \wRegInBot_0_0[0] }), .L_WR(\wRegEnTop_1_0[0] ), .L_In({
        \wRegOut_1_0[31] , \wRegOut_1_0[30] , \wRegOut_1_0[29] , 
        \wRegOut_1_0[28] , \wRegOut_1_0[27] , \wRegOut_1_0[26] , 
        \wRegOut_1_0[25] , \wRegOut_1_0[24] , \wRegOut_1_0[23] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[21] , \wRegOut_1_0[20] , 
        \wRegOut_1_0[19] , \wRegOut_1_0[18] , \wRegOut_1_0[17] , 
        \wRegOut_1_0[16] , \wRegOut_1_0[15] , \wRegOut_1_0[14] , 
        \wRegOut_1_0[13] , \wRegOut_1_0[12] , \wRegOut_1_0[11] , 
        \wRegOut_1_0[10] , \wRegOut_1_0[9] , \wRegOut_1_0[8] , 
        \wRegOut_1_0[7] , \wRegOut_1_0[6] , \wRegOut_1_0[5] , \wRegOut_1_0[4] , 
        \wRegOut_1_0[3] , \wRegOut_1_0[2] , \wRegOut_1_0[1] , \wRegOut_1_0[0] 
        }), .L_Out({\wRegInTop_1_0[31] , \wRegInTop_1_0[30] , 
        \wRegInTop_1_0[29] , \wRegInTop_1_0[28] , \wRegInTop_1_0[27] , 
        \wRegInTop_1_0[26] , \wRegInTop_1_0[25] , \wRegInTop_1_0[24] , 
        \wRegInTop_1_0[23] , \wRegInTop_1_0[22] , \wRegInTop_1_0[21] , 
        \wRegInTop_1_0[20] , \wRegInTop_1_0[19] , \wRegInTop_1_0[18] , 
        \wRegInTop_1_0[17] , \wRegInTop_1_0[16] , \wRegInTop_1_0[15] , 
        \wRegInTop_1_0[14] , \wRegInTop_1_0[13] , \wRegInTop_1_0[12] , 
        \wRegInTop_1_0[11] , \wRegInTop_1_0[10] , \wRegInTop_1_0[9] , 
        \wRegInTop_1_0[8] , \wRegInTop_1_0[7] , \wRegInTop_1_0[6] , 
        \wRegInTop_1_0[5] , \wRegInTop_1_0[4] , \wRegInTop_1_0[3] , 
        \wRegInTop_1_0[2] , \wRegInTop_1_0[1] , \wRegInTop_1_0[0] }), .R_WR(
        \wRegEnTop_1_1[0] ), .R_In({\wRegOut_1_1[31] , \wRegOut_1_1[30] , 
        \wRegOut_1_1[29] , \wRegOut_1_1[28] , \wRegOut_1_1[27] , 
        \wRegOut_1_1[26] , \wRegOut_1_1[25] , \wRegOut_1_1[24] , 
        \wRegOut_1_1[23] , \wRegOut_1_1[22] , \wRegOut_1_1[21] , 
        \wRegOut_1_1[20] , \wRegOut_1_1[19] , \wRegOut_1_1[18] , 
        \wRegOut_1_1[17] , \wRegOut_1_1[16] , \wRegOut_1_1[15] , 
        \wRegOut_1_1[14] , \wRegOut_1_1[13] , \wRegOut_1_1[12] , 
        \wRegOut_1_1[11] , \wRegOut_1_1[10] , \wRegOut_1_1[9] , 
        \wRegOut_1_1[8] , \wRegOut_1_1[7] , \wRegOut_1_1[6] , \wRegOut_1_1[5] , 
        \wRegOut_1_1[4] , \wRegOut_1_1[3] , \wRegOut_1_1[2] , \wRegOut_1_1[1] , 
        \wRegOut_1_1[0] }), .R_Out({\wRegInTop_1_1[31] , \wRegInTop_1_1[30] , 
        \wRegInTop_1_1[29] , \wRegInTop_1_1[28] , \wRegInTop_1_1[27] , 
        \wRegInTop_1_1[26] , \wRegInTop_1_1[25] , \wRegInTop_1_1[24] , 
        \wRegInTop_1_1[23] , \wRegInTop_1_1[22] , \wRegInTop_1_1[21] , 
        \wRegInTop_1_1[20] , \wRegInTop_1_1[19] , \wRegInTop_1_1[18] , 
        \wRegInTop_1_1[17] , \wRegInTop_1_1[16] , \wRegInTop_1_1[15] , 
        \wRegInTop_1_1[14] , \wRegInTop_1_1[13] , \wRegInTop_1_1[12] , 
        \wRegInTop_1_1[11] , \wRegInTop_1_1[10] , \wRegInTop_1_1[9] , 
        \wRegInTop_1_1[8] , \wRegInTop_1_1[7] , \wRegInTop_1_1[6] , 
        \wRegInTop_1_1[5] , \wRegInTop_1_1[4] , \wRegInTop_1_1[3] , 
        \wRegInTop_1_1[2] , \wRegInTop_1_1[1] , \wRegInTop_1_1[0] }) );
    BHeap_Node_WIDTH32 BHN_5_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_6[0] ), .P_In({\wRegOut_5_6[31] , 
        \wRegOut_5_6[30] , \wRegOut_5_6[29] , \wRegOut_5_6[28] , 
        \wRegOut_5_6[27] , \wRegOut_5_6[26] , \wRegOut_5_6[25] , 
        \wRegOut_5_6[24] , \wRegOut_5_6[23] , \wRegOut_5_6[22] , 
        \wRegOut_5_6[21] , \wRegOut_5_6[20] , \wRegOut_5_6[19] , 
        \wRegOut_5_6[18] , \wRegOut_5_6[17] , \wRegOut_5_6[16] , 
        \wRegOut_5_6[15] , \wRegOut_5_6[14] , \wRegOut_5_6[13] , 
        \wRegOut_5_6[12] , \wRegOut_5_6[11] , \wRegOut_5_6[10] , 
        \wRegOut_5_6[9] , \wRegOut_5_6[8] , \wRegOut_5_6[7] , \wRegOut_5_6[6] , 
        \wRegOut_5_6[5] , \wRegOut_5_6[4] , \wRegOut_5_6[3] , \wRegOut_5_6[2] , 
        \wRegOut_5_6[1] , \wRegOut_5_6[0] }), .P_Out({\wRegInBot_5_6[31] , 
        \wRegInBot_5_6[30] , \wRegInBot_5_6[29] , \wRegInBot_5_6[28] , 
        \wRegInBot_5_6[27] , \wRegInBot_5_6[26] , \wRegInBot_5_6[25] , 
        \wRegInBot_5_6[24] , \wRegInBot_5_6[23] , \wRegInBot_5_6[22] , 
        \wRegInBot_5_6[21] , \wRegInBot_5_6[20] , \wRegInBot_5_6[19] , 
        \wRegInBot_5_6[18] , \wRegInBot_5_6[17] , \wRegInBot_5_6[16] , 
        \wRegInBot_5_6[15] , \wRegInBot_5_6[14] , \wRegInBot_5_6[13] , 
        \wRegInBot_5_6[12] , \wRegInBot_5_6[11] , \wRegInBot_5_6[10] , 
        \wRegInBot_5_6[9] , \wRegInBot_5_6[8] , \wRegInBot_5_6[7] , 
        \wRegInBot_5_6[6] , \wRegInBot_5_6[5] , \wRegInBot_5_6[4] , 
        \wRegInBot_5_6[3] , \wRegInBot_5_6[2] , \wRegInBot_5_6[1] , 
        \wRegInBot_5_6[0] }), .L_WR(\wRegEnTop_6_12[0] ), .L_In({
        \wRegOut_6_12[31] , \wRegOut_6_12[30] , \wRegOut_6_12[29] , 
        \wRegOut_6_12[28] , \wRegOut_6_12[27] , \wRegOut_6_12[26] , 
        \wRegOut_6_12[25] , \wRegOut_6_12[24] , \wRegOut_6_12[23] , 
        \wRegOut_6_12[22] , \wRegOut_6_12[21] , \wRegOut_6_12[20] , 
        \wRegOut_6_12[19] , \wRegOut_6_12[18] , \wRegOut_6_12[17] , 
        \wRegOut_6_12[16] , \wRegOut_6_12[15] , \wRegOut_6_12[14] , 
        \wRegOut_6_12[13] , \wRegOut_6_12[12] , \wRegOut_6_12[11] , 
        \wRegOut_6_12[10] , \wRegOut_6_12[9] , \wRegOut_6_12[8] , 
        \wRegOut_6_12[7] , \wRegOut_6_12[6] , \wRegOut_6_12[5] , 
        \wRegOut_6_12[4] , \wRegOut_6_12[3] , \wRegOut_6_12[2] , 
        \wRegOut_6_12[1] , \wRegOut_6_12[0] }), .L_Out({\wRegInTop_6_12[31] , 
        \wRegInTop_6_12[30] , \wRegInTop_6_12[29] , \wRegInTop_6_12[28] , 
        \wRegInTop_6_12[27] , \wRegInTop_6_12[26] , \wRegInTop_6_12[25] , 
        \wRegInTop_6_12[24] , \wRegInTop_6_12[23] , \wRegInTop_6_12[22] , 
        \wRegInTop_6_12[21] , \wRegInTop_6_12[20] , \wRegInTop_6_12[19] , 
        \wRegInTop_6_12[18] , \wRegInTop_6_12[17] , \wRegInTop_6_12[16] , 
        \wRegInTop_6_12[15] , \wRegInTop_6_12[14] , \wRegInTop_6_12[13] , 
        \wRegInTop_6_12[12] , \wRegInTop_6_12[11] , \wRegInTop_6_12[10] , 
        \wRegInTop_6_12[9] , \wRegInTop_6_12[8] , \wRegInTop_6_12[7] , 
        \wRegInTop_6_12[6] , \wRegInTop_6_12[5] , \wRegInTop_6_12[4] , 
        \wRegInTop_6_12[3] , \wRegInTop_6_12[2] , \wRegInTop_6_12[1] , 
        \wRegInTop_6_12[0] }), .R_WR(\wRegEnTop_6_13[0] ), .R_In({
        \wRegOut_6_13[31] , \wRegOut_6_13[30] , \wRegOut_6_13[29] , 
        \wRegOut_6_13[28] , \wRegOut_6_13[27] , \wRegOut_6_13[26] , 
        \wRegOut_6_13[25] , \wRegOut_6_13[24] , \wRegOut_6_13[23] , 
        \wRegOut_6_13[22] , \wRegOut_6_13[21] , \wRegOut_6_13[20] , 
        \wRegOut_6_13[19] , \wRegOut_6_13[18] , \wRegOut_6_13[17] , 
        \wRegOut_6_13[16] , \wRegOut_6_13[15] , \wRegOut_6_13[14] , 
        \wRegOut_6_13[13] , \wRegOut_6_13[12] , \wRegOut_6_13[11] , 
        \wRegOut_6_13[10] , \wRegOut_6_13[9] , \wRegOut_6_13[8] , 
        \wRegOut_6_13[7] , \wRegOut_6_13[6] , \wRegOut_6_13[5] , 
        \wRegOut_6_13[4] , \wRegOut_6_13[3] , \wRegOut_6_13[2] , 
        \wRegOut_6_13[1] , \wRegOut_6_13[0] }), .R_Out({\wRegInTop_6_13[31] , 
        \wRegInTop_6_13[30] , \wRegInTop_6_13[29] , \wRegInTop_6_13[28] , 
        \wRegInTop_6_13[27] , \wRegInTop_6_13[26] , \wRegInTop_6_13[25] , 
        \wRegInTop_6_13[24] , \wRegInTop_6_13[23] , \wRegInTop_6_13[22] , 
        \wRegInTop_6_13[21] , \wRegInTop_6_13[20] , \wRegInTop_6_13[19] , 
        \wRegInTop_6_13[18] , \wRegInTop_6_13[17] , \wRegInTop_6_13[16] , 
        \wRegInTop_6_13[15] , \wRegInTop_6_13[14] , \wRegInTop_6_13[13] , 
        \wRegInTop_6_13[12] , \wRegInTop_6_13[11] , \wRegInTop_6_13[10] , 
        \wRegInTop_6_13[9] , \wRegInTop_6_13[8] , \wRegInTop_6_13[7] , 
        \wRegInTop_6_13[6] , \wRegInTop_6_13[5] , \wRegInTop_6_13[4] , 
        \wRegInTop_6_13[3] , \wRegInTop_6_13[2] , \wRegInTop_6_13[1] , 
        \wRegInTop_6_13[0] }) );
    BHeap_Control_CWIDTH4_IDWIDTH1_WIDTH32_SCAN1 BHC ( .Clk(Clk), .Reset(Reset
        ), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink0[31] , \ScanLink0[30] , \ScanLink0[29] , 
        \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , \ScanLink0[25] , 
        \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , \ScanLink0[21] , 
        \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , \ScanLink0[17] , 
        \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , \ScanLink0[13] , 
        \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , \ScanLink0[9] , 
        \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , \ScanLink0[5] , 
        \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , \ScanLink0[1] , 
        \ScanLink0[0] }), .ScanOut({\ScanLink255[31] , \ScanLink255[30] , 
        \ScanLink255[29] , \ScanLink255[28] , \ScanLink255[27] , 
        \ScanLink255[26] , \ScanLink255[25] , \ScanLink255[24] , 
        \ScanLink255[23] , \ScanLink255[22] , \ScanLink255[21] , 
        \ScanLink255[20] , \ScanLink255[19] , \ScanLink255[18] , 
        \ScanLink255[17] , \ScanLink255[16] , \ScanLink255[15] , 
        \ScanLink255[14] , \ScanLink255[13] , \ScanLink255[12] , 
        \ScanLink255[11] , \ScanLink255[10] , \ScanLink255[9] , 
        \ScanLink255[8] , \ScanLink255[7] , \ScanLink255[6] , \ScanLink255[5] , 
        \ScanLink255[4] , \ScanLink255[3] , \ScanLink255[2] , \ScanLink255[1] , 
        \ScanLink255[0] }), .ScanEnable(\ScanEnable[0] ), .ScanId(1'b0), .Id(
        1'b1), .Go(\wCtrlOut_7[0] ), .Done(\wCtrlOut_0[0] ) );
    BHeap_Node_WIDTH32 BHN_6_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_40[0] ), .P_In({\wRegOut_6_40[31] , 
        \wRegOut_6_40[30] , \wRegOut_6_40[29] , \wRegOut_6_40[28] , 
        \wRegOut_6_40[27] , \wRegOut_6_40[26] , \wRegOut_6_40[25] , 
        \wRegOut_6_40[24] , \wRegOut_6_40[23] , \wRegOut_6_40[22] , 
        \wRegOut_6_40[21] , \wRegOut_6_40[20] , \wRegOut_6_40[19] , 
        \wRegOut_6_40[18] , \wRegOut_6_40[17] , \wRegOut_6_40[16] , 
        \wRegOut_6_40[15] , \wRegOut_6_40[14] , \wRegOut_6_40[13] , 
        \wRegOut_6_40[12] , \wRegOut_6_40[11] , \wRegOut_6_40[10] , 
        \wRegOut_6_40[9] , \wRegOut_6_40[8] , \wRegOut_6_40[7] , 
        \wRegOut_6_40[6] , \wRegOut_6_40[5] , \wRegOut_6_40[4] , 
        \wRegOut_6_40[3] , \wRegOut_6_40[2] , \wRegOut_6_40[1] , 
        \wRegOut_6_40[0] }), .P_Out({\wRegInBot_6_40[31] , 
        \wRegInBot_6_40[30] , \wRegInBot_6_40[29] , \wRegInBot_6_40[28] , 
        \wRegInBot_6_40[27] , \wRegInBot_6_40[26] , \wRegInBot_6_40[25] , 
        \wRegInBot_6_40[24] , \wRegInBot_6_40[23] , \wRegInBot_6_40[22] , 
        \wRegInBot_6_40[21] , \wRegInBot_6_40[20] , \wRegInBot_6_40[19] , 
        \wRegInBot_6_40[18] , \wRegInBot_6_40[17] , \wRegInBot_6_40[16] , 
        \wRegInBot_6_40[15] , \wRegInBot_6_40[14] , \wRegInBot_6_40[13] , 
        \wRegInBot_6_40[12] , \wRegInBot_6_40[11] , \wRegInBot_6_40[10] , 
        \wRegInBot_6_40[9] , \wRegInBot_6_40[8] , \wRegInBot_6_40[7] , 
        \wRegInBot_6_40[6] , \wRegInBot_6_40[5] , \wRegInBot_6_40[4] , 
        \wRegInBot_6_40[3] , \wRegInBot_6_40[2] , \wRegInBot_6_40[1] , 
        \wRegInBot_6_40[0] }), .L_WR(\wRegEnTop_7_80[0] ), .L_In({
        \wRegOut_7_80[31] , \wRegOut_7_80[30] , \wRegOut_7_80[29] , 
        \wRegOut_7_80[28] , \wRegOut_7_80[27] , \wRegOut_7_80[26] , 
        \wRegOut_7_80[25] , \wRegOut_7_80[24] , \wRegOut_7_80[23] , 
        \wRegOut_7_80[22] , \wRegOut_7_80[21] , \wRegOut_7_80[20] , 
        \wRegOut_7_80[19] , \wRegOut_7_80[18] , \wRegOut_7_80[17] , 
        \wRegOut_7_80[16] , \wRegOut_7_80[15] , \wRegOut_7_80[14] , 
        \wRegOut_7_80[13] , \wRegOut_7_80[12] , \wRegOut_7_80[11] , 
        \wRegOut_7_80[10] , \wRegOut_7_80[9] , \wRegOut_7_80[8] , 
        \wRegOut_7_80[7] , \wRegOut_7_80[6] , \wRegOut_7_80[5] , 
        \wRegOut_7_80[4] , \wRegOut_7_80[3] , \wRegOut_7_80[2] , 
        \wRegOut_7_80[1] , \wRegOut_7_80[0] }), .L_Out({\wRegInTop_7_80[31] , 
        \wRegInTop_7_80[30] , \wRegInTop_7_80[29] , \wRegInTop_7_80[28] , 
        \wRegInTop_7_80[27] , \wRegInTop_7_80[26] , \wRegInTop_7_80[25] , 
        \wRegInTop_7_80[24] , \wRegInTop_7_80[23] , \wRegInTop_7_80[22] , 
        \wRegInTop_7_80[21] , \wRegInTop_7_80[20] , \wRegInTop_7_80[19] , 
        \wRegInTop_7_80[18] , \wRegInTop_7_80[17] , \wRegInTop_7_80[16] , 
        \wRegInTop_7_80[15] , \wRegInTop_7_80[14] , \wRegInTop_7_80[13] , 
        \wRegInTop_7_80[12] , \wRegInTop_7_80[11] , \wRegInTop_7_80[10] , 
        \wRegInTop_7_80[9] , \wRegInTop_7_80[8] , \wRegInTop_7_80[7] , 
        \wRegInTop_7_80[6] , \wRegInTop_7_80[5] , \wRegInTop_7_80[4] , 
        \wRegInTop_7_80[3] , \wRegInTop_7_80[2] , \wRegInTop_7_80[1] , 
        \wRegInTop_7_80[0] }), .R_WR(\wRegEnTop_7_81[0] ), .R_In({
        \wRegOut_7_81[31] , \wRegOut_7_81[30] , \wRegOut_7_81[29] , 
        \wRegOut_7_81[28] , \wRegOut_7_81[27] , \wRegOut_7_81[26] , 
        \wRegOut_7_81[25] , \wRegOut_7_81[24] , \wRegOut_7_81[23] , 
        \wRegOut_7_81[22] , \wRegOut_7_81[21] , \wRegOut_7_81[20] , 
        \wRegOut_7_81[19] , \wRegOut_7_81[18] , \wRegOut_7_81[17] , 
        \wRegOut_7_81[16] , \wRegOut_7_81[15] , \wRegOut_7_81[14] , 
        \wRegOut_7_81[13] , \wRegOut_7_81[12] , \wRegOut_7_81[11] , 
        \wRegOut_7_81[10] , \wRegOut_7_81[9] , \wRegOut_7_81[8] , 
        \wRegOut_7_81[7] , \wRegOut_7_81[6] , \wRegOut_7_81[5] , 
        \wRegOut_7_81[4] , \wRegOut_7_81[3] , \wRegOut_7_81[2] , 
        \wRegOut_7_81[1] , \wRegOut_7_81[0] }), .R_Out({\wRegInTop_7_81[31] , 
        \wRegInTop_7_81[30] , \wRegInTop_7_81[29] , \wRegInTop_7_81[28] , 
        \wRegInTop_7_81[27] , \wRegInTop_7_81[26] , \wRegInTop_7_81[25] , 
        \wRegInTop_7_81[24] , \wRegInTop_7_81[23] , \wRegInTop_7_81[22] , 
        \wRegInTop_7_81[21] , \wRegInTop_7_81[20] , \wRegInTop_7_81[19] , 
        \wRegInTop_7_81[18] , \wRegInTop_7_81[17] , \wRegInTop_7_81[16] , 
        \wRegInTop_7_81[15] , \wRegInTop_7_81[14] , \wRegInTop_7_81[13] , 
        \wRegInTop_7_81[12] , \wRegInTop_7_81[11] , \wRegInTop_7_81[10] , 
        \wRegInTop_7_81[9] , \wRegInTop_7_81[8] , \wRegInTop_7_81[7] , 
        \wRegInTop_7_81[6] , \wRegInTop_7_81[5] , \wRegInTop_7_81[4] , 
        \wRegInTop_7_81[3] , \wRegInTop_7_81[2] , \wRegInTop_7_81[1] , 
        \wRegInTop_7_81[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink36[31] , \ScanLink36[30] , \ScanLink36[29] , 
        \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , \ScanLink36[25] , 
        \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , \ScanLink36[21] , 
        \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , \ScanLink36[17] , 
        \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , \ScanLink36[13] , 
        \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , \ScanLink36[9] , 
        \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , \ScanLink36[5] , 
        \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , \ScanLink36[1] , 
        \ScanLink36[0] }), .ScanOut({\ScanLink35[31] , \ScanLink35[30] , 
        \ScanLink35[29] , \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , 
        \ScanLink35[25] , \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , 
        \ScanLink35[21] , \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , 
        \ScanLink35[17] , \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , 
        \ScanLink35[13] , \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , 
        \ScanLink35[9] , \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , 
        \ScanLink35[5] , \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , 
        \ScanLink35[1] , \ScanLink35[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_4[31] , \wRegOut_5_4[30] , \wRegOut_5_4[29] , 
        \wRegOut_5_4[28] , \wRegOut_5_4[27] , \wRegOut_5_4[26] , 
        \wRegOut_5_4[25] , \wRegOut_5_4[24] , \wRegOut_5_4[23] , 
        \wRegOut_5_4[22] , \wRegOut_5_4[21] , \wRegOut_5_4[20] , 
        \wRegOut_5_4[19] , \wRegOut_5_4[18] , \wRegOut_5_4[17] , 
        \wRegOut_5_4[16] , \wRegOut_5_4[15] , \wRegOut_5_4[14] , 
        \wRegOut_5_4[13] , \wRegOut_5_4[12] , \wRegOut_5_4[11] , 
        \wRegOut_5_4[10] , \wRegOut_5_4[9] , \wRegOut_5_4[8] , 
        \wRegOut_5_4[7] , \wRegOut_5_4[6] , \wRegOut_5_4[5] , \wRegOut_5_4[4] , 
        \wRegOut_5_4[3] , \wRegOut_5_4[2] , \wRegOut_5_4[1] , \wRegOut_5_4[0] 
        }), .Enable1(\wRegEnTop_5_4[0] ), .Enable2(\wRegEnBot_5_4[0] ), .In1({
        \wRegInTop_5_4[31] , \wRegInTop_5_4[30] , \wRegInTop_5_4[29] , 
        \wRegInTop_5_4[28] , \wRegInTop_5_4[27] , \wRegInTop_5_4[26] , 
        \wRegInTop_5_4[25] , \wRegInTop_5_4[24] , \wRegInTop_5_4[23] , 
        \wRegInTop_5_4[22] , \wRegInTop_5_4[21] , \wRegInTop_5_4[20] , 
        \wRegInTop_5_4[19] , \wRegInTop_5_4[18] , \wRegInTop_5_4[17] , 
        \wRegInTop_5_4[16] , \wRegInTop_5_4[15] , \wRegInTop_5_4[14] , 
        \wRegInTop_5_4[13] , \wRegInTop_5_4[12] , \wRegInTop_5_4[11] , 
        \wRegInTop_5_4[10] , \wRegInTop_5_4[9] , \wRegInTop_5_4[8] , 
        \wRegInTop_5_4[7] , \wRegInTop_5_4[6] , \wRegInTop_5_4[5] , 
        \wRegInTop_5_4[4] , \wRegInTop_5_4[3] , \wRegInTop_5_4[2] , 
        \wRegInTop_5_4[1] , \wRegInTop_5_4[0] }), .In2({\wRegInBot_5_4[31] , 
        \wRegInBot_5_4[30] , \wRegInBot_5_4[29] , \wRegInBot_5_4[28] , 
        \wRegInBot_5_4[27] , \wRegInBot_5_4[26] , \wRegInBot_5_4[25] , 
        \wRegInBot_5_4[24] , \wRegInBot_5_4[23] , \wRegInBot_5_4[22] , 
        \wRegInBot_5_4[21] , \wRegInBot_5_4[20] , \wRegInBot_5_4[19] , 
        \wRegInBot_5_4[18] , \wRegInBot_5_4[17] , \wRegInBot_5_4[16] , 
        \wRegInBot_5_4[15] , \wRegInBot_5_4[14] , \wRegInBot_5_4[13] , 
        \wRegInBot_5_4[12] , \wRegInBot_5_4[11] , \wRegInBot_5_4[10] , 
        \wRegInBot_5_4[9] , \wRegInBot_5_4[8] , \wRegInBot_5_4[7] , 
        \wRegInBot_5_4[6] , \wRegInBot_5_4[5] , \wRegInBot_5_4[4] , 
        \wRegInBot_5_4[3] , \wRegInBot_5_4[2] , \wRegInBot_5_4[1] , 
        \wRegInBot_5_4[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_20 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink148[31] , \ScanLink148[30] , \ScanLink148[29] , 
        \ScanLink148[28] , \ScanLink148[27] , \ScanLink148[26] , 
        \ScanLink148[25] , \ScanLink148[24] , \ScanLink148[23] , 
        \ScanLink148[22] , \ScanLink148[21] , \ScanLink148[20] , 
        \ScanLink148[19] , \ScanLink148[18] , \ScanLink148[17] , 
        \ScanLink148[16] , \ScanLink148[15] , \ScanLink148[14] , 
        \ScanLink148[13] , \ScanLink148[12] , \ScanLink148[11] , 
        \ScanLink148[10] , \ScanLink148[9] , \ScanLink148[8] , 
        \ScanLink148[7] , \ScanLink148[6] , \ScanLink148[5] , \ScanLink148[4] , 
        \ScanLink148[3] , \ScanLink148[2] , \ScanLink148[1] , \ScanLink148[0] 
        }), .ScanOut({\ScanLink147[31] , \ScanLink147[30] , \ScanLink147[29] , 
        \ScanLink147[28] , \ScanLink147[27] , \ScanLink147[26] , 
        \ScanLink147[25] , \ScanLink147[24] , \ScanLink147[23] , 
        \ScanLink147[22] , \ScanLink147[21] , \ScanLink147[20] , 
        \ScanLink147[19] , \ScanLink147[18] , \ScanLink147[17] , 
        \ScanLink147[16] , \ScanLink147[15] , \ScanLink147[14] , 
        \ScanLink147[13] , \ScanLink147[12] , \ScanLink147[11] , 
        \ScanLink147[10] , \ScanLink147[9] , \ScanLink147[8] , 
        \ScanLink147[7] , \ScanLink147[6] , \ScanLink147[5] , \ScanLink147[4] , 
        \ScanLink147[3] , \ScanLink147[2] , \ScanLink147[1] , \ScanLink147[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_20[31] , 
        \wRegOut_7_20[30] , \wRegOut_7_20[29] , \wRegOut_7_20[28] , 
        \wRegOut_7_20[27] , \wRegOut_7_20[26] , \wRegOut_7_20[25] , 
        \wRegOut_7_20[24] , \wRegOut_7_20[23] , \wRegOut_7_20[22] , 
        \wRegOut_7_20[21] , \wRegOut_7_20[20] , \wRegOut_7_20[19] , 
        \wRegOut_7_20[18] , \wRegOut_7_20[17] , \wRegOut_7_20[16] , 
        \wRegOut_7_20[15] , \wRegOut_7_20[14] , \wRegOut_7_20[13] , 
        \wRegOut_7_20[12] , \wRegOut_7_20[11] , \wRegOut_7_20[10] , 
        \wRegOut_7_20[9] , \wRegOut_7_20[8] , \wRegOut_7_20[7] , 
        \wRegOut_7_20[6] , \wRegOut_7_20[5] , \wRegOut_7_20[4] , 
        \wRegOut_7_20[3] , \wRegOut_7_20[2] , \wRegOut_7_20[1] , 
        \wRegOut_7_20[0] }), .Enable1(\wRegEnTop_7_20[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_20[31] , \wRegInTop_7_20[30] , \wRegInTop_7_20[29] , 
        \wRegInTop_7_20[28] , \wRegInTop_7_20[27] , \wRegInTop_7_20[26] , 
        \wRegInTop_7_20[25] , \wRegInTop_7_20[24] , \wRegInTop_7_20[23] , 
        \wRegInTop_7_20[22] , \wRegInTop_7_20[21] , \wRegInTop_7_20[20] , 
        \wRegInTop_7_20[19] , \wRegInTop_7_20[18] , \wRegInTop_7_20[17] , 
        \wRegInTop_7_20[16] , \wRegInTop_7_20[15] , \wRegInTop_7_20[14] , 
        \wRegInTop_7_20[13] , \wRegInTop_7_20[12] , \wRegInTop_7_20[11] , 
        \wRegInTop_7_20[10] , \wRegInTop_7_20[9] , \wRegInTop_7_20[8] , 
        \wRegInTop_7_20[7] , \wRegInTop_7_20[6] , \wRegInTop_7_20[5] , 
        \wRegInTop_7_20[4] , \wRegInTop_7_20[3] , \wRegInTop_7_20[2] , 
        \wRegInTop_7_20[1] , \wRegInTop_7_20[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_113 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink241[31] , \ScanLink241[30] , \ScanLink241[29] , 
        \ScanLink241[28] , \ScanLink241[27] , \ScanLink241[26] , 
        \ScanLink241[25] , \ScanLink241[24] , \ScanLink241[23] , 
        \ScanLink241[22] , \ScanLink241[21] , \ScanLink241[20] , 
        \ScanLink241[19] , \ScanLink241[18] , \ScanLink241[17] , 
        \ScanLink241[16] , \ScanLink241[15] , \ScanLink241[14] , 
        \ScanLink241[13] , \ScanLink241[12] , \ScanLink241[11] , 
        \ScanLink241[10] , \ScanLink241[9] , \ScanLink241[8] , 
        \ScanLink241[7] , \ScanLink241[6] , \ScanLink241[5] , \ScanLink241[4] , 
        \ScanLink241[3] , \ScanLink241[2] , \ScanLink241[1] , \ScanLink241[0] 
        }), .ScanOut({\ScanLink240[31] , \ScanLink240[30] , \ScanLink240[29] , 
        \ScanLink240[28] , \ScanLink240[27] , \ScanLink240[26] , 
        \ScanLink240[25] , \ScanLink240[24] , \ScanLink240[23] , 
        \ScanLink240[22] , \ScanLink240[21] , \ScanLink240[20] , 
        \ScanLink240[19] , \ScanLink240[18] , \ScanLink240[17] , 
        \ScanLink240[16] , \ScanLink240[15] , \ScanLink240[14] , 
        \ScanLink240[13] , \ScanLink240[12] , \ScanLink240[11] , 
        \ScanLink240[10] , \ScanLink240[9] , \ScanLink240[8] , 
        \ScanLink240[7] , \ScanLink240[6] , \ScanLink240[5] , \ScanLink240[4] , 
        \ScanLink240[3] , \ScanLink240[2] , \ScanLink240[1] , \ScanLink240[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_113[31] , 
        \wRegOut_7_113[30] , \wRegOut_7_113[29] , \wRegOut_7_113[28] , 
        \wRegOut_7_113[27] , \wRegOut_7_113[26] , \wRegOut_7_113[25] , 
        \wRegOut_7_113[24] , \wRegOut_7_113[23] , \wRegOut_7_113[22] , 
        \wRegOut_7_113[21] , \wRegOut_7_113[20] , \wRegOut_7_113[19] , 
        \wRegOut_7_113[18] , \wRegOut_7_113[17] , \wRegOut_7_113[16] , 
        \wRegOut_7_113[15] , \wRegOut_7_113[14] , \wRegOut_7_113[13] , 
        \wRegOut_7_113[12] , \wRegOut_7_113[11] , \wRegOut_7_113[10] , 
        \wRegOut_7_113[9] , \wRegOut_7_113[8] , \wRegOut_7_113[7] , 
        \wRegOut_7_113[6] , \wRegOut_7_113[5] , \wRegOut_7_113[4] , 
        \wRegOut_7_113[3] , \wRegOut_7_113[2] , \wRegOut_7_113[1] , 
        \wRegOut_7_113[0] }), .Enable1(\wRegEnTop_7_113[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_113[31] , \wRegInTop_7_113[30] , 
        \wRegInTop_7_113[29] , \wRegInTop_7_113[28] , \wRegInTop_7_113[27] , 
        \wRegInTop_7_113[26] , \wRegInTop_7_113[25] , \wRegInTop_7_113[24] , 
        \wRegInTop_7_113[23] , \wRegInTop_7_113[22] , \wRegInTop_7_113[21] , 
        \wRegInTop_7_113[20] , \wRegInTop_7_113[19] , \wRegInTop_7_113[18] , 
        \wRegInTop_7_113[17] , \wRegInTop_7_113[16] , \wRegInTop_7_113[15] , 
        \wRegInTop_7_113[14] , \wRegInTop_7_113[13] , \wRegInTop_7_113[12] , 
        \wRegInTop_7_113[11] , \wRegInTop_7_113[10] , \wRegInTop_7_113[9] , 
        \wRegInTop_7_113[8] , \wRegInTop_7_113[7] , \wRegInTop_7_113[6] , 
        \wRegInTop_7_113[5] , \wRegInTop_7_113[4] , \wRegInTop_7_113[3] , 
        \wRegInTop_7_113[2] , \wRegInTop_7_113[1] , \wRegInTop_7_113[0] }), 
        .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_1[0] ), .P_WR(\wRegEnBot_1_0[0] ), .P_In({\wRegOut_1_0[31] , 
        \wRegOut_1_0[30] , \wRegOut_1_0[29] , \wRegOut_1_0[28] , 
        \wRegOut_1_0[27] , \wRegOut_1_0[26] , \wRegOut_1_0[25] , 
        \wRegOut_1_0[24] , \wRegOut_1_0[23] , \wRegOut_1_0[22] , 
        \wRegOut_1_0[21] , \wRegOut_1_0[20] , \wRegOut_1_0[19] , 
        \wRegOut_1_0[18] , \wRegOut_1_0[17] , \wRegOut_1_0[16] , 
        \wRegOut_1_0[15] , \wRegOut_1_0[14] , \wRegOut_1_0[13] , 
        \wRegOut_1_0[12] , \wRegOut_1_0[11] , \wRegOut_1_0[10] , 
        \wRegOut_1_0[9] , \wRegOut_1_0[8] , \wRegOut_1_0[7] , \wRegOut_1_0[6] , 
        \wRegOut_1_0[5] , \wRegOut_1_0[4] , \wRegOut_1_0[3] , \wRegOut_1_0[2] , 
        \wRegOut_1_0[1] , \wRegOut_1_0[0] }), .P_Out({\wRegInBot_1_0[31] , 
        \wRegInBot_1_0[30] , \wRegInBot_1_0[29] , \wRegInBot_1_0[28] , 
        \wRegInBot_1_0[27] , \wRegInBot_1_0[26] , \wRegInBot_1_0[25] , 
        \wRegInBot_1_0[24] , \wRegInBot_1_0[23] , \wRegInBot_1_0[22] , 
        \wRegInBot_1_0[21] , \wRegInBot_1_0[20] , \wRegInBot_1_0[19] , 
        \wRegInBot_1_0[18] , \wRegInBot_1_0[17] , \wRegInBot_1_0[16] , 
        \wRegInBot_1_0[15] , \wRegInBot_1_0[14] , \wRegInBot_1_0[13] , 
        \wRegInBot_1_0[12] , \wRegInBot_1_0[11] , \wRegInBot_1_0[10] , 
        \wRegInBot_1_0[9] , \wRegInBot_1_0[8] , \wRegInBot_1_0[7] , 
        \wRegInBot_1_0[6] , \wRegInBot_1_0[5] , \wRegInBot_1_0[4] , 
        \wRegInBot_1_0[3] , \wRegInBot_1_0[2] , \wRegInBot_1_0[1] , 
        \wRegInBot_1_0[0] }), .L_WR(\wRegEnTop_2_0[0] ), .L_In({
        \wRegOut_2_0[31] , \wRegOut_2_0[30] , \wRegOut_2_0[29] , 
        \wRegOut_2_0[28] , \wRegOut_2_0[27] , \wRegOut_2_0[26] , 
        \wRegOut_2_0[25] , \wRegOut_2_0[24] , \wRegOut_2_0[23] , 
        \wRegOut_2_0[22] , \wRegOut_2_0[21] , \wRegOut_2_0[20] , 
        \wRegOut_2_0[19] , \wRegOut_2_0[18] , \wRegOut_2_0[17] , 
        \wRegOut_2_0[16] , \wRegOut_2_0[15] , \wRegOut_2_0[14] , 
        \wRegOut_2_0[13] , \wRegOut_2_0[12] , \wRegOut_2_0[11] , 
        \wRegOut_2_0[10] , \wRegOut_2_0[9] , \wRegOut_2_0[8] , 
        \wRegOut_2_0[7] , \wRegOut_2_0[6] , \wRegOut_2_0[5] , \wRegOut_2_0[4] , 
        \wRegOut_2_0[3] , \wRegOut_2_0[2] , \wRegOut_2_0[1] , \wRegOut_2_0[0] 
        }), .L_Out({\wRegInTop_2_0[31] , \wRegInTop_2_0[30] , 
        \wRegInTop_2_0[29] , \wRegInTop_2_0[28] , \wRegInTop_2_0[27] , 
        \wRegInTop_2_0[26] , \wRegInTop_2_0[25] , \wRegInTop_2_0[24] , 
        \wRegInTop_2_0[23] , \wRegInTop_2_0[22] , \wRegInTop_2_0[21] , 
        \wRegInTop_2_0[20] , \wRegInTop_2_0[19] , \wRegInTop_2_0[18] , 
        \wRegInTop_2_0[17] , \wRegInTop_2_0[16] , \wRegInTop_2_0[15] , 
        \wRegInTop_2_0[14] , \wRegInTop_2_0[13] , \wRegInTop_2_0[12] , 
        \wRegInTop_2_0[11] , \wRegInTop_2_0[10] , \wRegInTop_2_0[9] , 
        \wRegInTop_2_0[8] , \wRegInTop_2_0[7] , \wRegInTop_2_0[6] , 
        \wRegInTop_2_0[5] , \wRegInTop_2_0[4] , \wRegInTop_2_0[3] , 
        \wRegInTop_2_0[2] , \wRegInTop_2_0[1] , \wRegInTop_2_0[0] }), .R_WR(
        \wRegEnTop_2_1[0] ), .R_In({\wRegOut_2_1[31] , \wRegOut_2_1[30] , 
        \wRegOut_2_1[29] , \wRegOut_2_1[28] , \wRegOut_2_1[27] , 
        \wRegOut_2_1[26] , \wRegOut_2_1[25] , \wRegOut_2_1[24] , 
        \wRegOut_2_1[23] , \wRegOut_2_1[22] , \wRegOut_2_1[21] , 
        \wRegOut_2_1[20] , \wRegOut_2_1[19] , \wRegOut_2_1[18] , 
        \wRegOut_2_1[17] , \wRegOut_2_1[16] , \wRegOut_2_1[15] , 
        \wRegOut_2_1[14] , \wRegOut_2_1[13] , \wRegOut_2_1[12] , 
        \wRegOut_2_1[11] , \wRegOut_2_1[10] , \wRegOut_2_1[9] , 
        \wRegOut_2_1[8] , \wRegOut_2_1[7] , \wRegOut_2_1[6] , \wRegOut_2_1[5] , 
        \wRegOut_2_1[4] , \wRegOut_2_1[3] , \wRegOut_2_1[2] , \wRegOut_2_1[1] , 
        \wRegOut_2_1[0] }), .R_Out({\wRegInTop_2_1[31] , \wRegInTop_2_1[30] , 
        \wRegInTop_2_1[29] , \wRegInTop_2_1[28] , \wRegInTop_2_1[27] , 
        \wRegInTop_2_1[26] , \wRegInTop_2_1[25] , \wRegInTop_2_1[24] , 
        \wRegInTop_2_1[23] , \wRegInTop_2_1[22] , \wRegInTop_2_1[21] , 
        \wRegInTop_2_1[20] , \wRegInTop_2_1[19] , \wRegInTop_2_1[18] , 
        \wRegInTop_2_1[17] , \wRegInTop_2_1[16] , \wRegInTop_2_1[15] , 
        \wRegInTop_2_1[14] , \wRegInTop_2_1[13] , \wRegInTop_2_1[12] , 
        \wRegInTop_2_1[11] , \wRegInTop_2_1[10] , \wRegInTop_2_1[9] , 
        \wRegInTop_2_1[8] , \wRegInTop_2_1[7] , \wRegInTop_2_1[6] , 
        \wRegInTop_2_1[5] , \wRegInTop_2_1[4] , \wRegInTop_2_1[3] , 
        \wRegInTop_2_1[2] , \wRegInTop_2_1[1] , \wRegInTop_2_1[0] }) );
    BHeap_Node_WIDTH32 BHN_4_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_6[0] ), .P_In({\wRegOut_4_6[31] , 
        \wRegOut_4_6[30] , \wRegOut_4_6[29] , \wRegOut_4_6[28] , 
        \wRegOut_4_6[27] , \wRegOut_4_6[26] , \wRegOut_4_6[25] , 
        \wRegOut_4_6[24] , \wRegOut_4_6[23] , \wRegOut_4_6[22] , 
        \wRegOut_4_6[21] , \wRegOut_4_6[20] , \wRegOut_4_6[19] , 
        \wRegOut_4_6[18] , \wRegOut_4_6[17] , \wRegOut_4_6[16] , 
        \wRegOut_4_6[15] , \wRegOut_4_6[14] , \wRegOut_4_6[13] , 
        \wRegOut_4_6[12] , \wRegOut_4_6[11] , \wRegOut_4_6[10] , 
        \wRegOut_4_6[9] , \wRegOut_4_6[8] , \wRegOut_4_6[7] , \wRegOut_4_6[6] , 
        \wRegOut_4_6[5] , \wRegOut_4_6[4] , \wRegOut_4_6[3] , \wRegOut_4_6[2] , 
        \wRegOut_4_6[1] , \wRegOut_4_6[0] }), .P_Out({\wRegInBot_4_6[31] , 
        \wRegInBot_4_6[30] , \wRegInBot_4_6[29] , \wRegInBot_4_6[28] , 
        \wRegInBot_4_6[27] , \wRegInBot_4_6[26] , \wRegInBot_4_6[25] , 
        \wRegInBot_4_6[24] , \wRegInBot_4_6[23] , \wRegInBot_4_6[22] , 
        \wRegInBot_4_6[21] , \wRegInBot_4_6[20] , \wRegInBot_4_6[19] , 
        \wRegInBot_4_6[18] , \wRegInBot_4_6[17] , \wRegInBot_4_6[16] , 
        \wRegInBot_4_6[15] , \wRegInBot_4_6[14] , \wRegInBot_4_6[13] , 
        \wRegInBot_4_6[12] , \wRegInBot_4_6[11] , \wRegInBot_4_6[10] , 
        \wRegInBot_4_6[9] , \wRegInBot_4_6[8] , \wRegInBot_4_6[7] , 
        \wRegInBot_4_6[6] , \wRegInBot_4_6[5] , \wRegInBot_4_6[4] , 
        \wRegInBot_4_6[3] , \wRegInBot_4_6[2] , \wRegInBot_4_6[1] , 
        \wRegInBot_4_6[0] }), .L_WR(\wRegEnTop_5_12[0] ), .L_In({
        \wRegOut_5_12[31] , \wRegOut_5_12[30] , \wRegOut_5_12[29] , 
        \wRegOut_5_12[28] , \wRegOut_5_12[27] , \wRegOut_5_12[26] , 
        \wRegOut_5_12[25] , \wRegOut_5_12[24] , \wRegOut_5_12[23] , 
        \wRegOut_5_12[22] , \wRegOut_5_12[21] , \wRegOut_5_12[20] , 
        \wRegOut_5_12[19] , \wRegOut_5_12[18] , \wRegOut_5_12[17] , 
        \wRegOut_5_12[16] , \wRegOut_5_12[15] , \wRegOut_5_12[14] , 
        \wRegOut_5_12[13] , \wRegOut_5_12[12] , \wRegOut_5_12[11] , 
        \wRegOut_5_12[10] , \wRegOut_5_12[9] , \wRegOut_5_12[8] , 
        \wRegOut_5_12[7] , \wRegOut_5_12[6] , \wRegOut_5_12[5] , 
        \wRegOut_5_12[4] , \wRegOut_5_12[3] , \wRegOut_5_12[2] , 
        \wRegOut_5_12[1] , \wRegOut_5_12[0] }), .L_Out({\wRegInTop_5_12[31] , 
        \wRegInTop_5_12[30] , \wRegInTop_5_12[29] , \wRegInTop_5_12[28] , 
        \wRegInTop_5_12[27] , \wRegInTop_5_12[26] , \wRegInTop_5_12[25] , 
        \wRegInTop_5_12[24] , \wRegInTop_5_12[23] , \wRegInTop_5_12[22] , 
        \wRegInTop_5_12[21] , \wRegInTop_5_12[20] , \wRegInTop_5_12[19] , 
        \wRegInTop_5_12[18] , \wRegInTop_5_12[17] , \wRegInTop_5_12[16] , 
        \wRegInTop_5_12[15] , \wRegInTop_5_12[14] , \wRegInTop_5_12[13] , 
        \wRegInTop_5_12[12] , \wRegInTop_5_12[11] , \wRegInTop_5_12[10] , 
        \wRegInTop_5_12[9] , \wRegInTop_5_12[8] , \wRegInTop_5_12[7] , 
        \wRegInTop_5_12[6] , \wRegInTop_5_12[5] , \wRegInTop_5_12[4] , 
        \wRegInTop_5_12[3] , \wRegInTop_5_12[2] , \wRegInTop_5_12[1] , 
        \wRegInTop_5_12[0] }), .R_WR(\wRegEnTop_5_13[0] ), .R_In({
        \wRegOut_5_13[31] , \wRegOut_5_13[30] , \wRegOut_5_13[29] , 
        \wRegOut_5_13[28] , \wRegOut_5_13[27] , \wRegOut_5_13[26] , 
        \wRegOut_5_13[25] , \wRegOut_5_13[24] , \wRegOut_5_13[23] , 
        \wRegOut_5_13[22] , \wRegOut_5_13[21] , \wRegOut_5_13[20] , 
        \wRegOut_5_13[19] , \wRegOut_5_13[18] , \wRegOut_5_13[17] , 
        \wRegOut_5_13[16] , \wRegOut_5_13[15] , \wRegOut_5_13[14] , 
        \wRegOut_5_13[13] , \wRegOut_5_13[12] , \wRegOut_5_13[11] , 
        \wRegOut_5_13[10] , \wRegOut_5_13[9] , \wRegOut_5_13[8] , 
        \wRegOut_5_13[7] , \wRegOut_5_13[6] , \wRegOut_5_13[5] , 
        \wRegOut_5_13[4] , \wRegOut_5_13[3] , \wRegOut_5_13[2] , 
        \wRegOut_5_13[1] , \wRegOut_5_13[0] }), .R_Out({\wRegInTop_5_13[31] , 
        \wRegInTop_5_13[30] , \wRegInTop_5_13[29] , \wRegInTop_5_13[28] , 
        \wRegInTop_5_13[27] , \wRegInTop_5_13[26] , \wRegInTop_5_13[25] , 
        \wRegInTop_5_13[24] , \wRegInTop_5_13[23] , \wRegInTop_5_13[22] , 
        \wRegInTop_5_13[21] , \wRegInTop_5_13[20] , \wRegInTop_5_13[19] , 
        \wRegInTop_5_13[18] , \wRegInTop_5_13[17] , \wRegInTop_5_13[16] , 
        \wRegInTop_5_13[15] , \wRegInTop_5_13[14] , \wRegInTop_5_13[13] , 
        \wRegInTop_5_13[12] , \wRegInTop_5_13[11] , \wRegInTop_5_13[10] , 
        \wRegInTop_5_13[9] , \wRegInTop_5_13[8] , \wRegInTop_5_13[7] , 
        \wRegInTop_5_13[6] , \wRegInTop_5_13[5] , \wRegInTop_5_13[4] , 
        \wRegInTop_5_13[3] , \wRegInTop_5_13[2] , \wRegInTop_5_13[1] , 
        \wRegInTop_5_13[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink136[31] , \ScanLink136[30] , \ScanLink136[29] , 
        \ScanLink136[28] , \ScanLink136[27] , \ScanLink136[26] , 
        \ScanLink136[25] , \ScanLink136[24] , \ScanLink136[23] , 
        \ScanLink136[22] , \ScanLink136[21] , \ScanLink136[20] , 
        \ScanLink136[19] , \ScanLink136[18] , \ScanLink136[17] , 
        \ScanLink136[16] , \ScanLink136[15] , \ScanLink136[14] , 
        \ScanLink136[13] , \ScanLink136[12] , \ScanLink136[11] , 
        \ScanLink136[10] , \ScanLink136[9] , \ScanLink136[8] , 
        \ScanLink136[7] , \ScanLink136[6] , \ScanLink136[5] , \ScanLink136[4] , 
        \ScanLink136[3] , \ScanLink136[2] , \ScanLink136[1] , \ScanLink136[0] 
        }), .ScanOut({\ScanLink135[31] , \ScanLink135[30] , \ScanLink135[29] , 
        \ScanLink135[28] , \ScanLink135[27] , \ScanLink135[26] , 
        \ScanLink135[25] , \ScanLink135[24] , \ScanLink135[23] , 
        \ScanLink135[22] , \ScanLink135[21] , \ScanLink135[20] , 
        \ScanLink135[19] , \ScanLink135[18] , \ScanLink135[17] , 
        \ScanLink135[16] , \ScanLink135[15] , \ScanLink135[14] , 
        \ScanLink135[13] , \ScanLink135[12] , \ScanLink135[11] , 
        \ScanLink135[10] , \ScanLink135[9] , \ScanLink135[8] , 
        \ScanLink135[7] , \ScanLink135[6] , \ScanLink135[5] , \ScanLink135[4] , 
        \ScanLink135[3] , \ScanLink135[2] , \ScanLink135[1] , \ScanLink135[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_8[31] , 
        \wRegOut_7_8[30] , \wRegOut_7_8[29] , \wRegOut_7_8[28] , 
        \wRegOut_7_8[27] , \wRegOut_7_8[26] , \wRegOut_7_8[25] , 
        \wRegOut_7_8[24] , \wRegOut_7_8[23] , \wRegOut_7_8[22] , 
        \wRegOut_7_8[21] , \wRegOut_7_8[20] , \wRegOut_7_8[19] , 
        \wRegOut_7_8[18] , \wRegOut_7_8[17] , \wRegOut_7_8[16] , 
        \wRegOut_7_8[15] , \wRegOut_7_8[14] , \wRegOut_7_8[13] , 
        \wRegOut_7_8[12] , \wRegOut_7_8[11] , \wRegOut_7_8[10] , 
        \wRegOut_7_8[9] , \wRegOut_7_8[8] , \wRegOut_7_8[7] , \wRegOut_7_8[6] , 
        \wRegOut_7_8[5] , \wRegOut_7_8[4] , \wRegOut_7_8[3] , \wRegOut_7_8[2] , 
        \wRegOut_7_8[1] , \wRegOut_7_8[0] }), .Enable1(\wRegEnTop_7_8[0] ), 
        .Enable2(1'b0), .In1({\wRegInTop_7_8[31] , \wRegInTop_7_8[30] , 
        \wRegInTop_7_8[29] , \wRegInTop_7_8[28] , \wRegInTop_7_8[27] , 
        \wRegInTop_7_8[26] , \wRegInTop_7_8[25] , \wRegInTop_7_8[24] , 
        \wRegInTop_7_8[23] , \wRegInTop_7_8[22] , \wRegInTop_7_8[21] , 
        \wRegInTop_7_8[20] , \wRegInTop_7_8[19] , \wRegInTop_7_8[18] , 
        \wRegInTop_7_8[17] , \wRegInTop_7_8[16] , \wRegInTop_7_8[15] , 
        \wRegInTop_7_8[14] , \wRegInTop_7_8[13] , \wRegInTop_7_8[12] , 
        \wRegInTop_7_8[11] , \wRegInTop_7_8[10] , \wRegInTop_7_8[9] , 
        \wRegInTop_7_8[8] , \wRegInTop_7_8[7] , \wRegInTop_7_8[6] , 
        \wRegInTop_7_8[5] , \wRegInTop_7_8[4] , \wRegInTop_7_8[3] , 
        \wRegInTop_7_8[2] , \wRegInTop_7_8[1] , \wRegInTop_7_8[0] }), .In2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_7_69 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink197[31] , \ScanLink197[30] , \ScanLink197[29] , 
        \ScanLink197[28] , \ScanLink197[27] , \ScanLink197[26] , 
        \ScanLink197[25] , \ScanLink197[24] , \ScanLink197[23] , 
        \ScanLink197[22] , \ScanLink197[21] , \ScanLink197[20] , 
        \ScanLink197[19] , \ScanLink197[18] , \ScanLink197[17] , 
        \ScanLink197[16] , \ScanLink197[15] , \ScanLink197[14] , 
        \ScanLink197[13] , \ScanLink197[12] , \ScanLink197[11] , 
        \ScanLink197[10] , \ScanLink197[9] , \ScanLink197[8] , 
        \ScanLink197[7] , \ScanLink197[6] , \ScanLink197[5] , \ScanLink197[4] , 
        \ScanLink197[3] , \ScanLink197[2] , \ScanLink197[1] , \ScanLink197[0] 
        }), .ScanOut({\ScanLink196[31] , \ScanLink196[30] , \ScanLink196[29] , 
        \ScanLink196[28] , \ScanLink196[27] , \ScanLink196[26] , 
        \ScanLink196[25] , \ScanLink196[24] , \ScanLink196[23] , 
        \ScanLink196[22] , \ScanLink196[21] , \ScanLink196[20] , 
        \ScanLink196[19] , \ScanLink196[18] , \ScanLink196[17] , 
        \ScanLink196[16] , \ScanLink196[15] , \ScanLink196[14] , 
        \ScanLink196[13] , \ScanLink196[12] , \ScanLink196[11] , 
        \ScanLink196[10] , \ScanLink196[9] , \ScanLink196[8] , 
        \ScanLink196[7] , \ScanLink196[6] , \ScanLink196[5] , \ScanLink196[4] , 
        \ScanLink196[3] , \ScanLink196[2] , \ScanLink196[1] , \ScanLink196[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Out({\wRegOut_7_69[31] , 
        \wRegOut_7_69[30] , \wRegOut_7_69[29] , \wRegOut_7_69[28] , 
        \wRegOut_7_69[27] , \wRegOut_7_69[26] , \wRegOut_7_69[25] , 
        \wRegOut_7_69[24] , \wRegOut_7_69[23] , \wRegOut_7_69[22] , 
        \wRegOut_7_69[21] , \wRegOut_7_69[20] , \wRegOut_7_69[19] , 
        \wRegOut_7_69[18] , \wRegOut_7_69[17] , \wRegOut_7_69[16] , 
        \wRegOut_7_69[15] , \wRegOut_7_69[14] , \wRegOut_7_69[13] , 
        \wRegOut_7_69[12] , \wRegOut_7_69[11] , \wRegOut_7_69[10] , 
        \wRegOut_7_69[9] , \wRegOut_7_69[8] , \wRegOut_7_69[7] , 
        \wRegOut_7_69[6] , \wRegOut_7_69[5] , \wRegOut_7_69[4] , 
        \wRegOut_7_69[3] , \wRegOut_7_69[2] , \wRegOut_7_69[1] , 
        \wRegOut_7_69[0] }), .Enable1(\wRegEnTop_7_69[0] ), .Enable2(1'b0), 
        .In1({\wRegInTop_7_69[31] , \wRegInTop_7_69[30] , \wRegInTop_7_69[29] , 
        \wRegInTop_7_69[28] , \wRegInTop_7_69[27] , \wRegInTop_7_69[26] , 
        \wRegInTop_7_69[25] , \wRegInTop_7_69[24] , \wRegInTop_7_69[23] , 
        \wRegInTop_7_69[22] , \wRegInTop_7_69[21] , \wRegInTop_7_69[20] , 
        \wRegInTop_7_69[19] , \wRegInTop_7_69[18] , \wRegInTop_7_69[17] , 
        \wRegInTop_7_69[16] , \wRegInTop_7_69[15] , \wRegInTop_7_69[14] , 
        \wRegInTop_7_69[13] , \wRegInTop_7_69[12] , \wRegInTop_7_69[11] , 
        \wRegInTop_7_69[10] , \wRegInTop_7_69[9] , \wRegInTop_7_69[8] , 
        \wRegInTop_7_69[7] , \wRegInTop_7_69[6] , \wRegInTop_7_69[5] , 
        \wRegInTop_7_69[4] , \wRegInTop_7_69[3] , \wRegInTop_7_69[2] , 
        \wRegInTop_7_69[1] , \wRegInTop_7_69[0] }), .In2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_6_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_35[0] ), .P_In({\wRegOut_6_35[31] , 
        \wRegOut_6_35[30] , \wRegOut_6_35[29] , \wRegOut_6_35[28] , 
        \wRegOut_6_35[27] , \wRegOut_6_35[26] , \wRegOut_6_35[25] , 
        \wRegOut_6_35[24] , \wRegOut_6_35[23] , \wRegOut_6_35[22] , 
        \wRegOut_6_35[21] , \wRegOut_6_35[20] , \wRegOut_6_35[19] , 
        \wRegOut_6_35[18] , \wRegOut_6_35[17] , \wRegOut_6_35[16] , 
        \wRegOut_6_35[15] , \wRegOut_6_35[14] , \wRegOut_6_35[13] , 
        \wRegOut_6_35[12] , \wRegOut_6_35[11] , \wRegOut_6_35[10] , 
        \wRegOut_6_35[9] , \wRegOut_6_35[8] , \wRegOut_6_35[7] , 
        \wRegOut_6_35[6] , \wRegOut_6_35[5] , \wRegOut_6_35[4] , 
        \wRegOut_6_35[3] , \wRegOut_6_35[2] , \wRegOut_6_35[1] , 
        \wRegOut_6_35[0] }), .P_Out({\wRegInBot_6_35[31] , 
        \wRegInBot_6_35[30] , \wRegInBot_6_35[29] , \wRegInBot_6_35[28] , 
        \wRegInBot_6_35[27] , \wRegInBot_6_35[26] , \wRegInBot_6_35[25] , 
        \wRegInBot_6_35[24] , \wRegInBot_6_35[23] , \wRegInBot_6_35[22] , 
        \wRegInBot_6_35[21] , \wRegInBot_6_35[20] , \wRegInBot_6_35[19] , 
        \wRegInBot_6_35[18] , \wRegInBot_6_35[17] , \wRegInBot_6_35[16] , 
        \wRegInBot_6_35[15] , \wRegInBot_6_35[14] , \wRegInBot_6_35[13] , 
        \wRegInBot_6_35[12] , \wRegInBot_6_35[11] , \wRegInBot_6_35[10] , 
        \wRegInBot_6_35[9] , \wRegInBot_6_35[8] , \wRegInBot_6_35[7] , 
        \wRegInBot_6_35[6] , \wRegInBot_6_35[5] , \wRegInBot_6_35[4] , 
        \wRegInBot_6_35[3] , \wRegInBot_6_35[2] , \wRegInBot_6_35[1] , 
        \wRegInBot_6_35[0] }), .L_WR(\wRegEnTop_7_70[0] ), .L_In({
        \wRegOut_7_70[31] , \wRegOut_7_70[30] , \wRegOut_7_70[29] , 
        \wRegOut_7_70[28] , \wRegOut_7_70[27] , \wRegOut_7_70[26] , 
        \wRegOut_7_70[25] , \wRegOut_7_70[24] , \wRegOut_7_70[23] , 
        \wRegOut_7_70[22] , \wRegOut_7_70[21] , \wRegOut_7_70[20] , 
        \wRegOut_7_70[19] , \wRegOut_7_70[18] , \wRegOut_7_70[17] , 
        \wRegOut_7_70[16] , \wRegOut_7_70[15] , \wRegOut_7_70[14] , 
        \wRegOut_7_70[13] , \wRegOut_7_70[12] , \wRegOut_7_70[11] , 
        \wRegOut_7_70[10] , \wRegOut_7_70[9] , \wRegOut_7_70[8] , 
        \wRegOut_7_70[7] , \wRegOut_7_70[6] , \wRegOut_7_70[5] , 
        \wRegOut_7_70[4] , \wRegOut_7_70[3] , \wRegOut_7_70[2] , 
        \wRegOut_7_70[1] , \wRegOut_7_70[0] }), .L_Out({\wRegInTop_7_70[31] , 
        \wRegInTop_7_70[30] , \wRegInTop_7_70[29] , \wRegInTop_7_70[28] , 
        \wRegInTop_7_70[27] , \wRegInTop_7_70[26] , \wRegInTop_7_70[25] , 
        \wRegInTop_7_70[24] , \wRegInTop_7_70[23] , \wRegInTop_7_70[22] , 
        \wRegInTop_7_70[21] , \wRegInTop_7_70[20] , \wRegInTop_7_70[19] , 
        \wRegInTop_7_70[18] , \wRegInTop_7_70[17] , \wRegInTop_7_70[16] , 
        \wRegInTop_7_70[15] , \wRegInTop_7_70[14] , \wRegInTop_7_70[13] , 
        \wRegInTop_7_70[12] , \wRegInTop_7_70[11] , \wRegInTop_7_70[10] , 
        \wRegInTop_7_70[9] , \wRegInTop_7_70[8] , \wRegInTop_7_70[7] , 
        \wRegInTop_7_70[6] , \wRegInTop_7_70[5] , \wRegInTop_7_70[4] , 
        \wRegInTop_7_70[3] , \wRegInTop_7_70[2] , \wRegInTop_7_70[1] , 
        \wRegInTop_7_70[0] }), .R_WR(\wRegEnTop_7_71[0] ), .R_In({
        \wRegOut_7_71[31] , \wRegOut_7_71[30] , \wRegOut_7_71[29] , 
        \wRegOut_7_71[28] , \wRegOut_7_71[27] , \wRegOut_7_71[26] , 
        \wRegOut_7_71[25] , \wRegOut_7_71[24] , \wRegOut_7_71[23] , 
        \wRegOut_7_71[22] , \wRegOut_7_71[21] , \wRegOut_7_71[20] , 
        \wRegOut_7_71[19] , \wRegOut_7_71[18] , \wRegOut_7_71[17] , 
        \wRegOut_7_71[16] , \wRegOut_7_71[15] , \wRegOut_7_71[14] , 
        \wRegOut_7_71[13] , \wRegOut_7_71[12] , \wRegOut_7_71[11] , 
        \wRegOut_7_71[10] , \wRegOut_7_71[9] , \wRegOut_7_71[8] , 
        \wRegOut_7_71[7] , \wRegOut_7_71[6] , \wRegOut_7_71[5] , 
        \wRegOut_7_71[4] , \wRegOut_7_71[3] , \wRegOut_7_71[2] , 
        \wRegOut_7_71[1] , \wRegOut_7_71[0] }), .R_Out({\wRegInTop_7_71[31] , 
        \wRegInTop_7_71[30] , \wRegInTop_7_71[29] , \wRegInTop_7_71[28] , 
        \wRegInTop_7_71[27] , \wRegInTop_7_71[26] , \wRegInTop_7_71[25] , 
        \wRegInTop_7_71[24] , \wRegInTop_7_71[23] , \wRegInTop_7_71[22] , 
        \wRegInTop_7_71[21] , \wRegInTop_7_71[20] , \wRegInTop_7_71[19] , 
        \wRegInTop_7_71[18] , \wRegInTop_7_71[17] , \wRegInTop_7_71[16] , 
        \wRegInTop_7_71[15] , \wRegInTop_7_71[14] , \wRegInTop_7_71[13] , 
        \wRegInTop_7_71[12] , \wRegInTop_7_71[11] , \wRegInTop_7_71[10] , 
        \wRegInTop_7_71[9] , \wRegInTop_7_71[8] , \wRegInTop_7_71[7] , 
        \wRegInTop_7_71[6] , \wRegInTop_7_71[5] , \wRegInTop_7_71[4] , 
        \wRegInTop_7_71[3] , \wRegInTop_7_71[2] , \wRegInTop_7_71[1] , 
        \wRegInTop_7_71[0] }) );
    BHeap_Node_WIDTH32 BHN_5_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_5[0] ), .P_WR(\wRegEnBot_5_22[0] ), .P_In({\wRegOut_5_22[31] , 
        \wRegOut_5_22[30] , \wRegOut_5_22[29] , \wRegOut_5_22[28] , 
        \wRegOut_5_22[27] , \wRegOut_5_22[26] , \wRegOut_5_22[25] , 
        \wRegOut_5_22[24] , \wRegOut_5_22[23] , \wRegOut_5_22[22] , 
        \wRegOut_5_22[21] , \wRegOut_5_22[20] , \wRegOut_5_22[19] , 
        \wRegOut_5_22[18] , \wRegOut_5_22[17] , \wRegOut_5_22[16] , 
        \wRegOut_5_22[15] , \wRegOut_5_22[14] , \wRegOut_5_22[13] , 
        \wRegOut_5_22[12] , \wRegOut_5_22[11] , \wRegOut_5_22[10] , 
        \wRegOut_5_22[9] , \wRegOut_5_22[8] , \wRegOut_5_22[7] , 
        \wRegOut_5_22[6] , \wRegOut_5_22[5] , \wRegOut_5_22[4] , 
        \wRegOut_5_22[3] , \wRegOut_5_22[2] , \wRegOut_5_22[1] , 
        \wRegOut_5_22[0] }), .P_Out({\wRegInBot_5_22[31] , 
        \wRegInBot_5_22[30] , \wRegInBot_5_22[29] , \wRegInBot_5_22[28] , 
        \wRegInBot_5_22[27] , \wRegInBot_5_22[26] , \wRegInBot_5_22[25] , 
        \wRegInBot_5_22[24] , \wRegInBot_5_22[23] , \wRegInBot_5_22[22] , 
        \wRegInBot_5_22[21] , \wRegInBot_5_22[20] , \wRegInBot_5_22[19] , 
        \wRegInBot_5_22[18] , \wRegInBot_5_22[17] , \wRegInBot_5_22[16] , 
        \wRegInBot_5_22[15] , \wRegInBot_5_22[14] , \wRegInBot_5_22[13] , 
        \wRegInBot_5_22[12] , \wRegInBot_5_22[11] , \wRegInBot_5_22[10] , 
        \wRegInBot_5_22[9] , \wRegInBot_5_22[8] , \wRegInBot_5_22[7] , 
        \wRegInBot_5_22[6] , \wRegInBot_5_22[5] , \wRegInBot_5_22[4] , 
        \wRegInBot_5_22[3] , \wRegInBot_5_22[2] , \wRegInBot_5_22[1] , 
        \wRegInBot_5_22[0] }), .L_WR(\wRegEnTop_6_44[0] ), .L_In({
        \wRegOut_6_44[31] , \wRegOut_6_44[30] , \wRegOut_6_44[29] , 
        \wRegOut_6_44[28] , \wRegOut_6_44[27] , \wRegOut_6_44[26] , 
        \wRegOut_6_44[25] , \wRegOut_6_44[24] , \wRegOut_6_44[23] , 
        \wRegOut_6_44[22] , \wRegOut_6_44[21] , \wRegOut_6_44[20] , 
        \wRegOut_6_44[19] , \wRegOut_6_44[18] , \wRegOut_6_44[17] , 
        \wRegOut_6_44[16] , \wRegOut_6_44[15] , \wRegOut_6_44[14] , 
        \wRegOut_6_44[13] , \wRegOut_6_44[12] , \wRegOut_6_44[11] , 
        \wRegOut_6_44[10] , \wRegOut_6_44[9] , \wRegOut_6_44[8] , 
        \wRegOut_6_44[7] , \wRegOut_6_44[6] , \wRegOut_6_44[5] , 
        \wRegOut_6_44[4] , \wRegOut_6_44[3] , \wRegOut_6_44[2] , 
        \wRegOut_6_44[1] , \wRegOut_6_44[0] }), .L_Out({\wRegInTop_6_44[31] , 
        \wRegInTop_6_44[30] , \wRegInTop_6_44[29] , \wRegInTop_6_44[28] , 
        \wRegInTop_6_44[27] , \wRegInTop_6_44[26] , \wRegInTop_6_44[25] , 
        \wRegInTop_6_44[24] , \wRegInTop_6_44[23] , \wRegInTop_6_44[22] , 
        \wRegInTop_6_44[21] , \wRegInTop_6_44[20] , \wRegInTop_6_44[19] , 
        \wRegInTop_6_44[18] , \wRegInTop_6_44[17] , \wRegInTop_6_44[16] , 
        \wRegInTop_6_44[15] , \wRegInTop_6_44[14] , \wRegInTop_6_44[13] , 
        \wRegInTop_6_44[12] , \wRegInTop_6_44[11] , \wRegInTop_6_44[10] , 
        \wRegInTop_6_44[9] , \wRegInTop_6_44[8] , \wRegInTop_6_44[7] , 
        \wRegInTop_6_44[6] , \wRegInTop_6_44[5] , \wRegInTop_6_44[4] , 
        \wRegInTop_6_44[3] , \wRegInTop_6_44[2] , \wRegInTop_6_44[1] , 
        \wRegInTop_6_44[0] }), .R_WR(\wRegEnTop_6_45[0] ), .R_In({
        \wRegOut_6_45[31] , \wRegOut_6_45[30] , \wRegOut_6_45[29] , 
        \wRegOut_6_45[28] , \wRegOut_6_45[27] , \wRegOut_6_45[26] , 
        \wRegOut_6_45[25] , \wRegOut_6_45[24] , \wRegOut_6_45[23] , 
        \wRegOut_6_45[22] , \wRegOut_6_45[21] , \wRegOut_6_45[20] , 
        \wRegOut_6_45[19] , \wRegOut_6_45[18] , \wRegOut_6_45[17] , 
        \wRegOut_6_45[16] , \wRegOut_6_45[15] , \wRegOut_6_45[14] , 
        \wRegOut_6_45[13] , \wRegOut_6_45[12] , \wRegOut_6_45[11] , 
        \wRegOut_6_45[10] , \wRegOut_6_45[9] , \wRegOut_6_45[8] , 
        \wRegOut_6_45[7] , \wRegOut_6_45[6] , \wRegOut_6_45[5] , 
        \wRegOut_6_45[4] , \wRegOut_6_45[3] , \wRegOut_6_45[2] , 
        \wRegOut_6_45[1] , \wRegOut_6_45[0] }), .R_Out({\wRegInTop_6_45[31] , 
        \wRegInTop_6_45[30] , \wRegInTop_6_45[29] , \wRegInTop_6_45[28] , 
        \wRegInTop_6_45[27] , \wRegInTop_6_45[26] , \wRegInTop_6_45[25] , 
        \wRegInTop_6_45[24] , \wRegInTop_6_45[23] , \wRegInTop_6_45[22] , 
        \wRegInTop_6_45[21] , \wRegInTop_6_45[20] , \wRegInTop_6_45[19] , 
        \wRegInTop_6_45[18] , \wRegInTop_6_45[17] , \wRegInTop_6_45[16] , 
        \wRegInTop_6_45[15] , \wRegInTop_6_45[14] , \wRegInTop_6_45[13] , 
        \wRegInTop_6_45[12] , \wRegInTop_6_45[11] , \wRegInTop_6_45[10] , 
        \wRegInTop_6_45[9] , \wRegInTop_6_45[8] , \wRegInTop_6_45[7] , 
        \wRegInTop_6_45[6] , \wRegInTop_6_45[5] , \wRegInTop_6_45[4] , 
        \wRegInTop_6_45[3] , \wRegInTop_6_45[2] , \wRegInTop_6_45[1] , 
        \wRegInTop_6_45[0] }) );
    BHeap_Node_WIDTH32 BHN_6_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_6[0] ), .P_WR(\wRegEnBot_6_12[0] ), .P_In({\wRegOut_6_12[31] , 
        \wRegOut_6_12[30] , \wRegOut_6_12[29] , \wRegOut_6_12[28] , 
        \wRegOut_6_12[27] , \wRegOut_6_12[26] , \wRegOut_6_12[25] , 
        \wRegOut_6_12[24] , \wRegOut_6_12[23] , \wRegOut_6_12[22] , 
        \wRegOut_6_12[21] , \wRegOut_6_12[20] , \wRegOut_6_12[19] , 
        \wRegOut_6_12[18] , \wRegOut_6_12[17] , \wRegOut_6_12[16] , 
        \wRegOut_6_12[15] , \wRegOut_6_12[14] , \wRegOut_6_12[13] , 
        \wRegOut_6_12[12] , \wRegOut_6_12[11] , \wRegOut_6_12[10] , 
        \wRegOut_6_12[9] , \wRegOut_6_12[8] , \wRegOut_6_12[7] , 
        \wRegOut_6_12[6] , \wRegOut_6_12[5] , \wRegOut_6_12[4] , 
        \wRegOut_6_12[3] , \wRegOut_6_12[2] , \wRegOut_6_12[1] , 
        \wRegOut_6_12[0] }), .P_Out({\wRegInBot_6_12[31] , 
        \wRegInBot_6_12[30] , \wRegInBot_6_12[29] , \wRegInBot_6_12[28] , 
        \wRegInBot_6_12[27] , \wRegInBot_6_12[26] , \wRegInBot_6_12[25] , 
        \wRegInBot_6_12[24] , \wRegInBot_6_12[23] , \wRegInBot_6_12[22] , 
        \wRegInBot_6_12[21] , \wRegInBot_6_12[20] , \wRegInBot_6_12[19] , 
        \wRegInBot_6_12[18] , \wRegInBot_6_12[17] , \wRegInBot_6_12[16] , 
        \wRegInBot_6_12[15] , \wRegInBot_6_12[14] , \wRegInBot_6_12[13] , 
        \wRegInBot_6_12[12] , \wRegInBot_6_12[11] , \wRegInBot_6_12[10] , 
        \wRegInBot_6_12[9] , \wRegInBot_6_12[8] , \wRegInBot_6_12[7] , 
        \wRegInBot_6_12[6] , \wRegInBot_6_12[5] , \wRegInBot_6_12[4] , 
        \wRegInBot_6_12[3] , \wRegInBot_6_12[2] , \wRegInBot_6_12[1] , 
        \wRegInBot_6_12[0] }), .L_WR(\wRegEnTop_7_24[0] ), .L_In({
        \wRegOut_7_24[31] , \wRegOut_7_24[30] , \wRegOut_7_24[29] , 
        \wRegOut_7_24[28] , \wRegOut_7_24[27] , \wRegOut_7_24[26] , 
        \wRegOut_7_24[25] , \wRegOut_7_24[24] , \wRegOut_7_24[23] , 
        \wRegOut_7_24[22] , \wRegOut_7_24[21] , \wRegOut_7_24[20] , 
        \wRegOut_7_24[19] , \wRegOut_7_24[18] , \wRegOut_7_24[17] , 
        \wRegOut_7_24[16] , \wRegOut_7_24[15] , \wRegOut_7_24[14] , 
        \wRegOut_7_24[13] , \wRegOut_7_24[12] , \wRegOut_7_24[11] , 
        \wRegOut_7_24[10] , \wRegOut_7_24[9] , \wRegOut_7_24[8] , 
        \wRegOut_7_24[7] , \wRegOut_7_24[6] , \wRegOut_7_24[5] , 
        \wRegOut_7_24[4] , \wRegOut_7_24[3] , \wRegOut_7_24[2] , 
        \wRegOut_7_24[1] , \wRegOut_7_24[0] }), .L_Out({\wRegInTop_7_24[31] , 
        \wRegInTop_7_24[30] , \wRegInTop_7_24[29] , \wRegInTop_7_24[28] , 
        \wRegInTop_7_24[27] , \wRegInTop_7_24[26] , \wRegInTop_7_24[25] , 
        \wRegInTop_7_24[24] , \wRegInTop_7_24[23] , \wRegInTop_7_24[22] , 
        \wRegInTop_7_24[21] , \wRegInTop_7_24[20] , \wRegInTop_7_24[19] , 
        \wRegInTop_7_24[18] , \wRegInTop_7_24[17] , \wRegInTop_7_24[16] , 
        \wRegInTop_7_24[15] , \wRegInTop_7_24[14] , \wRegInTop_7_24[13] , 
        \wRegInTop_7_24[12] , \wRegInTop_7_24[11] , \wRegInTop_7_24[10] , 
        \wRegInTop_7_24[9] , \wRegInTop_7_24[8] , \wRegInTop_7_24[7] , 
        \wRegInTop_7_24[6] , \wRegInTop_7_24[5] , \wRegInTop_7_24[4] , 
        \wRegInTop_7_24[3] , \wRegInTop_7_24[2] , \wRegInTop_7_24[1] , 
        \wRegInTop_7_24[0] }), .R_WR(\wRegEnTop_7_25[0] ), .R_In({
        \wRegOut_7_25[31] , \wRegOut_7_25[30] , \wRegOut_7_25[29] , 
        \wRegOut_7_25[28] , \wRegOut_7_25[27] , \wRegOut_7_25[26] , 
        \wRegOut_7_25[25] , \wRegOut_7_25[24] , \wRegOut_7_25[23] , 
        \wRegOut_7_25[22] , \wRegOut_7_25[21] , \wRegOut_7_25[20] , 
        \wRegOut_7_25[19] , \wRegOut_7_25[18] , \wRegOut_7_25[17] , 
        \wRegOut_7_25[16] , \wRegOut_7_25[15] , \wRegOut_7_25[14] , 
        \wRegOut_7_25[13] , \wRegOut_7_25[12] , \wRegOut_7_25[11] , 
        \wRegOut_7_25[10] , \wRegOut_7_25[9] , \wRegOut_7_25[8] , 
        \wRegOut_7_25[7] , \wRegOut_7_25[6] , \wRegOut_7_25[5] , 
        \wRegOut_7_25[4] , \wRegOut_7_25[3] , \wRegOut_7_25[2] , 
        \wRegOut_7_25[1] , \wRegOut_7_25[0] }), .R_Out({\wRegInTop_7_25[31] , 
        \wRegInTop_7_25[30] , \wRegInTop_7_25[29] , \wRegInTop_7_25[28] , 
        \wRegInTop_7_25[27] , \wRegInTop_7_25[26] , \wRegInTop_7_25[25] , 
        \wRegInTop_7_25[24] , \wRegInTop_7_25[23] , \wRegInTop_7_25[22] , 
        \wRegInTop_7_25[21] , \wRegInTop_7_25[20] , \wRegInTop_7_25[19] , 
        \wRegInTop_7_25[18] , \wRegInTop_7_25[17] , \wRegInTop_7_25[16] , 
        \wRegInTop_7_25[15] , \wRegInTop_7_25[14] , \wRegInTop_7_25[13] , 
        \wRegInTop_7_25[12] , \wRegInTop_7_25[11] , \wRegInTop_7_25[10] , 
        \wRegInTop_7_25[9] , \wRegInTop_7_25[8] , \wRegInTop_7_25[7] , 
        \wRegInTop_7_25[6] , \wRegInTop_7_25[5] , \wRegInTop_7_25[4] , 
        \wRegInTop_7_25[3] , \wRegInTop_7_25[2] , \wRegInTop_7_25[1] , 
        \wRegInTop_7_25[0] }) );
endmodule

