
module EdgeAux_DW01_add_16_0 ( A, B, CI, SUM, CO );
input  [15:0] A;
input  [15:0] B;
output [15:0] SUM;
input  CI;
output CO;
    wire \carry[15] , \carry[13] , \carry[9] , \carry[4] , \carry[6] , 
        \carry[2] , \carry[14] , \carry[11] , \carry[10] , \carry[12] , 
        \carry[8] , \carry[7] , \carry[3] , \carry[5] , \carry[1] , n1;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_8 ( .CI(\carry[8] ), .A(A[8]), .B(B[8]), .S(SUM[8]), .CO(
        \carry[9] ) );
    VMW_FADD U1_11 ( .CI(\carry[11] ), .A(A[11]), .B(B[11]), .S(SUM[11]), .CO(
        \carry[12] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]), .CO(
        \carry[8] ) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_9 ( .CI(\carry[9] ), .A(A[9]), .B(B[9]), .S(SUM[9]), .CO(
        \carry[10] ) );
    VMW_FADD U1_10 ( .CI(\carry[10] ), .A(A[10]), .B(B[10]), .S(SUM[10]), .CO(
        \carry[11] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
    VMW_FADD U1_12 ( .CI(\carry[12] ), .A(A[12]), .B(B[12]), .S(SUM[12]), .CO(
        \carry[13] ) );
    VMW_FADD U1_15 ( .CI(\carry[15] ), .A(A[15]), .B(B[15]), .S(SUM[15]) );
    VMW_FADD U1_14 ( .CI(\carry[14] ), .A(A[14]), .B(B[14]), .S(SUM[14]), .CO(
        \carry[15] ) );
    VMW_FADD U1_13 ( .CI(\carry[13] ), .A(A[13]), .B(B[13]), .S(SUM[13]), .CO(
        \carry[14] ) );
endmodule


module EdgeAux ( Eid, InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [10:0] Eid;
input  [10:0] WeightAddr;
input  [15:0] InEdge;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire \Weight[11] , \Weight[6] , \Weight[15] , \Weight[2] , \Weight[0] , 
        \Weight[9] , \Weight[13] , \Weight[4] , \Weight[12] , \Weight[5] , 
        \Weight[1] , \Weight[8] , \Weight[14] , \Weight[3] , \Weight[10] , 
        \Weight[7] , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
        n101, n102, n103, n104, n105, n106, n107, n108;
    VMW_PULLDOWN U15 ( .Z(n108) );
    VMW_AO22 U16 ( .A(\Weight[9] ), .B(n76), .C(WeightData[9]), .D(n77), .Z(
        n98) );
    VMW_AO22 U17 ( .A(\Weight[8] ), .B(n76), .C(WeightData[8]), .D(n77), .Z(
        n99) );
    VMW_AO22 U18 ( .A(\Weight[7] ), .B(n76), .C(WeightData[7]), .D(n77), .Z(
        n100) );
    VMW_AO22 U19 ( .A(\Weight[6] ), .B(n76), .C(WeightData[6]), .D(n77), .Z(
        n101) );
    VMW_AO22 U20 ( .A(\Weight[5] ), .B(n76), .C(WeightData[5]), .D(n77), .Z(
        n102) );
    VMW_AO22 U21 ( .A(\Weight[4] ), .B(n76), .C(WeightData[4]), .D(n77), .Z(
        n103) );
    VMW_AO22 U22 ( .A(\Weight[3] ), .B(n76), .C(WeightData[3]), .D(n77), .Z(
        n104) );
    VMW_AO22 U23 ( .A(\Weight[2] ), .B(n76), .C(WeightData[2]), .D(n77), .Z(
        n105) );
    VMW_AO22 U24 ( .A(\Weight[1] ), .B(n76), .C(WeightData[1]), .D(n77), .Z(
        n106) );
    VMW_AO22 U25 ( .A(\Weight[15] ), .B(n76), .C(WeightData[15]), .D(n77), .Z(
        n92) );
    VMW_AO22 U26 ( .A(\Weight[14] ), .B(n76), .C(WeightData[14]), .D(n77), .Z(
        n93) );
    VMW_AO22 U27 ( .A(\Weight[13] ), .B(n76), .C(WeightData[13]), .D(n77), .Z(
        n94) );
    VMW_AO22 U28 ( .A(\Weight[12] ), .B(n76), .C(WeightData[12]), .D(n77), .Z(
        n95) );
    VMW_AO22 U29 ( .A(\Weight[11] ), .B(n76), .C(WeightData[11]), .D(n77), .Z(
        n96) );
    VMW_AO22 U30 ( .A(\Weight[10] ), .B(n76), .C(WeightData[10]), .D(n77), .Z(
        n97) );
    VMW_AO22 U31 ( .A(\Weight[0] ), .B(n76), .C(WeightData[0]), .D(n77), .Z(
        n107) );
    VMW_AND3 U32 ( .A(n79), .B(n80), .C(n81), .Z(n78) );
    VMW_AND4 U33 ( .A(n83), .B(n84), .C(n85), .D(n78), .Z(n82) );
    VMW_AND3 U34 ( .A(n87), .B(n88), .C(n89), .Z(n86) );
    VMW_AND4 U35 ( .A(n90), .B(n91), .C(n86), .D(n82), .Z(n77) );
    VMW_XNOR2 U36 ( .A(WeightAddr[4]), .B(Eid[4]), .Z(n80) );
    VMW_XNOR2 U37 ( .A(WeightAddr[0]), .B(Eid[0]), .Z(n79) );
    VMW_XNOR2 U38 ( .A(WeightAddr[3]), .B(Eid[3]), .Z(n81) );
    VMW_XNOR2 U39 ( .A(WeightAddr[7]), .B(Eid[7]), .Z(n84) );
    VMW_XNOR2 U40 ( .A(WeightAddr[5]), .B(Eid[5]), .Z(n83) );
    VMW_XNOR2 U41 ( .A(WeightAddr[6]), .B(Eid[6]), .Z(n85) );
    VMW_XNOR2 U42 ( .A(WeightAddr[10]), .B(Eid[10]), .Z(n88) );
    VMW_XNOR2 U43 ( .A(WeightAddr[8]), .B(Eid[8]), .Z(n87) );
    VMW_XNOR2 U44 ( .A(WeightAddr[9]), .B(Eid[9]), .Z(n89) );
    VMW_XNOR2 U45 ( .A(WeightAddr[2]), .B(Eid[2]), .Z(n91) );
    VMW_XNOR2 U46 ( .A(WeightAddr[1]), .B(Eid[1]), .Z(n90) );
    VMW_INV U47 ( .A(n77), .Z(n76) );
    VMW_FD \Weight_reg[15]  ( .D(n92), .CP(Clk), .Q(\Weight[15] ) );
    VMW_FD \Weight_reg[14]  ( .D(n93), .CP(Clk), .Q(\Weight[14] ) );
    VMW_FD \Weight_reg[13]  ( .D(n94), .CP(Clk), .Q(\Weight[13] ) );
    VMW_FD \Weight_reg[12]  ( .D(n95), .CP(Clk), .Q(\Weight[12] ) );
    VMW_FD \Weight_reg[11]  ( .D(n96), .CP(Clk), .Q(\Weight[11] ) );
    VMW_FD \Weight_reg[10]  ( .D(n97), .CP(Clk), .Q(\Weight[10] ) );
    VMW_FD \Weight_reg[9]  ( .D(n98), .CP(Clk), .Q(\Weight[9] ) );
    VMW_FD \Weight_reg[8]  ( .D(n99), .CP(Clk), .Q(\Weight[8] ) );
    VMW_FD \Weight_reg[7]  ( .D(n100), .CP(Clk), .Q(\Weight[7] ) );
    VMW_FD \Weight_reg[6]  ( .D(n101), .CP(Clk), .Q(\Weight[6] ) );
    VMW_FD \Weight_reg[5]  ( .D(n102), .CP(Clk), .Q(\Weight[5] ) );
    VMW_FD \Weight_reg[4]  ( .D(n103), .CP(Clk), .Q(\Weight[4] ) );
    VMW_FD \Weight_reg[3]  ( .D(n104), .CP(Clk), .Q(\Weight[3] ) );
    VMW_FD \Weight_reg[2]  ( .D(n105), .CP(Clk), .Q(\Weight[2] ) );
    VMW_FD \Weight_reg[1]  ( .D(n106), .CP(Clk), .Q(\Weight[1] ) );
    VMW_FD \Weight_reg[0]  ( .D(n107), .CP(Clk), .Q(\Weight[0] ) );
    EdgeAux_DW01_add_16_0 add_92 ( .A({\Weight[15] , \Weight[14] , 
        \Weight[13] , \Weight[12] , \Weight[11] , \Weight[10] , \Weight[9] , 
        \Weight[8] , \Weight[7] , \Weight[6] , \Weight[5] , \Weight[4] , 
        \Weight[3] , \Weight[2] , \Weight[1] , \Weight[0] }), .B(InEdge), .CI(
        n108), .SUM(OutEdge) );
endmodule


module NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_7 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_6 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n92, n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n105, n106, 
        n107, n108, n109, n110, n111, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n93), .C(n91), .D(n89), .Z(n92) );
    VMW_NAND2 U20 ( .A(n95), .B(B[10]), .Z(n94) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n92), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n95), .C(n99), .D(n97), .Z(n100) );
    VMW_NAND2 U24 ( .A(n102), .B(B[12]), .Z(n101) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n100), .D(n94), .Z(n103) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n102), .C(n106), .D(n103), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n101), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n113), .D(n110), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n102) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n93) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n95) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n118, n119, n121, n122, n123, n124, n125, n126, n127, 
        n129, n130, n131, n132, n133, n134, n135, n137, n138, n139, n140, n141, 
        n142, n143, n145, n146, n147, n148, n149, n150, n151, n153, n154, n155, 
        n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
        n168, n169;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n119), .B(B[2]), .Z(n118) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n119), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n127), .B(B[4]), .Z(n126) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n125), .D(n118), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n127), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n135), .B(B[6]), .Z(n134) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n132), .D(n126), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n135), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n146), .C(n140), .D(n134), .Z(n145) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n147) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n149), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U20 ( .A(n151), .B(B[10]), .Z(n150) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n154), .C(n148), .D(n142), .Z(n153) );
    VMW_NAND2 U22 ( .A(n154), .B(A[9]), .Z(n155) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n151), .C(n155), .D(n153), .Z(n156) );
    VMW_NAND2 U24 ( .A(n158), .B(B[12]), .Z(n157) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n160), .C(n156), .D(n150), .Z(n159) );
    VMW_NAND2 U26 ( .A(n160), .B(A[11]), .Z(n161) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n158), .C(n161), .D(n159), .Z(n162) );
    VMW_NAND2 U28 ( .A(n164), .B(B[14]), .Z(n163) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n166), .C(n162), .D(n157), .Z(n165) );
    VMW_NAND2 U30 ( .A(n166), .B(A[13]), .Z(n167) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n164), .C(n167), .D(n165), .Z(n168) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n169), .C(n168), .D(n163), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n158) );
    VMW_INV U34 ( .A(B[7]), .Z(n146) );
    VMW_INV U35 ( .A(A[7]), .Z(n149) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n151) );
    VMW_INV U39 ( .A(B[9]), .Z(n154) );
    VMW_INV U40 ( .A(A[4]), .Z(n127) );
    VMW_INV U41 ( .A(A[8]), .Z(n143) );
    VMW_INV U42 ( .A(A[14]), .Z(n164) );
    VMW_INV U43 ( .A(B[11]), .Z(n160) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n169) );
    VMW_INV U48 ( .A(B[13]), .Z(n166) );
    VMW_INV U49 ( .A(A[6]), .Z(n135) );
    VMW_INV U50 ( .A(A[2]), .Z(n119) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
        n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
        n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
        n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
        n217, n218;
    VMW_OAI21 U3 ( .A(B[15]), .B(n170), .C(n171), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n173), .B(B[2]), .Z(n172) );
    VMW_AO22 U5 ( .A(n175), .B(B[0]), .C(n176), .D(B[1]), .Z(n174) );
    VMW_OR2 U6 ( .A(B[2]), .B(n173), .Z(n177) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n176), .C(n177), .D(n174), .Z(n178) );
    VMW_NAND2 U8 ( .A(n180), .B(B[4]), .Z(n179) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n182), .C(n178), .D(n172), .Z(n181) );
    VMW_OR2 U10 ( .A(B[4]), .B(n180), .Z(n183) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n185), .C(n183), .D(n181), .Z(n184) );
    VMW_NAND2 U12 ( .A(n187), .B(B[6]), .Z(n186) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n189), .C(n184), .D(n179), .Z(n188) );
    VMW_OR2 U14 ( .A(B[6]), .B(n187), .Z(n190) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n192), .C(n190), .D(n188), .Z(n191) );
    VMW_NAND2 U16 ( .A(n194), .B(B[8]), .Z(n193) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n196), .C(n191), .D(n186), .Z(n195) );
    VMW_OR2 U18 ( .A(B[8]), .B(n194), .Z(n197) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n199), .C(n197), .D(n195), .Z(n198) );
    VMW_NAND2 U20 ( .A(n201), .B(B[10]), .Z(n200) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n203), .C(n198), .D(n193), .Z(n202) );
    VMW_NAND2 U22 ( .A(n203), .B(A[9]), .Z(n204) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n201), .C(n204), .D(n202), .Z(n205) );
    VMW_NAND2 U24 ( .A(n207), .B(B[12]), .Z(n206) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n209), .C(n205), .D(n200), .Z(n208) );
    VMW_NAND2 U26 ( .A(n209), .B(A[11]), .Z(n210) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n207), .C(n210), .D(n208), .Z(n211) );
    VMW_NAND2 U28 ( .A(n213), .B(B[14]), .Z(n212) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n215), .C(n211), .D(n206), .Z(n214) );
    VMW_NAND2 U30 ( .A(n215), .B(A[13]), .Z(n216) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n213), .C(n216), .D(n214), .Z(n217) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n218), .C(n217), .D(n212), .Z(n171) );
    VMW_INV U33 ( .A(A[12]), .Z(n207) );
    VMW_INV U34 ( .A(B[7]), .Z(n196) );
    VMW_INV U35 ( .A(A[7]), .Z(n199) );
    VMW_INV U36 ( .A(A[3]), .Z(n185) );
    VMW_INV U37 ( .A(B[3]), .Z(n182) );
    VMW_INV U38 ( .A(A[10]), .Z(n201) );
    VMW_INV U39 ( .A(B[9]), .Z(n203) );
    VMW_INV U40 ( .A(A[4]), .Z(n180) );
    VMW_INV U41 ( .A(A[8]), .Z(n194) );
    VMW_INV U42 ( .A(A[14]), .Z(n213) );
    VMW_INV U43 ( .A(B[11]), .Z(n209) );
    VMW_INV U44 ( .A(A[5]), .Z(n192) );
    VMW_INV U45 ( .A(B[5]), .Z(n189) );
    VMW_INV U46 ( .A(A[1]), .Z(n176) );
    VMW_INV U47 ( .A(B[15]), .Z(n218) );
    VMW_INV U48 ( .A(B[13]), .Z(n215) );
    VMW_INV U49 ( .A(A[6]), .Z(n187) );
    VMW_INV U50 ( .A(A[2]), .Z(n173) );
    VMW_INV U51 ( .A(A[0]), .Z(n175) );
    VMW_INV U52 ( .A(A[15]), .Z(n170) );
endmodule


module NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267;
    VMW_OAI21 U3 ( .A(B[15]), .B(n219), .C(n220), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n222), .B(B[2]), .Z(n221) );
    VMW_AO22 U5 ( .A(n224), .B(B[0]), .C(n225), .D(B[1]), .Z(n223) );
    VMW_OR2 U6 ( .A(B[2]), .B(n222), .Z(n226) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n225), .C(n226), .D(n223), .Z(n227) );
    VMW_NAND2 U8 ( .A(n229), .B(B[4]), .Z(n228) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n231), .C(n227), .D(n221), .Z(n230) );
    VMW_OR2 U10 ( .A(B[4]), .B(n229), .Z(n232) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n234), .C(n232), .D(n230), .Z(n233) );
    VMW_NAND2 U12 ( .A(n236), .B(B[6]), .Z(n235) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n238), .C(n233), .D(n228), .Z(n237) );
    VMW_OR2 U14 ( .A(B[6]), .B(n236), .Z(n239) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n241), .C(n239), .D(n237), .Z(n240) );
    VMW_NAND2 U16 ( .A(n243), .B(B[8]), .Z(n242) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n245), .C(n240), .D(n235), .Z(n244) );
    VMW_OR2 U18 ( .A(B[8]), .B(n243), .Z(n246) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n248), .C(n246), .D(n244), .Z(n247) );
    VMW_NAND2 U20 ( .A(n250), .B(B[10]), .Z(n249) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n252), .C(n247), .D(n242), .Z(n251) );
    VMW_NAND2 U22 ( .A(n252), .B(A[9]), .Z(n253) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n250), .C(n253), .D(n251), .Z(n254) );
    VMW_NAND2 U24 ( .A(n256), .B(B[12]), .Z(n255) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n258), .C(n254), .D(n249), .Z(n257) );
    VMW_NAND2 U26 ( .A(n258), .B(A[11]), .Z(n259) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n256), .C(n259), .D(n257), .Z(n260) );
    VMW_NAND2 U28 ( .A(n262), .B(B[14]), .Z(n261) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n264), .C(n260), .D(n255), .Z(n263) );
    VMW_NAND2 U30 ( .A(n264), .B(A[13]), .Z(n265) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n262), .C(n265), .D(n263), .Z(n266) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n267), .C(n266), .D(n261), .Z(n220) );
    VMW_INV U33 ( .A(A[12]), .Z(n256) );
    VMW_INV U34 ( .A(B[7]), .Z(n245) );
    VMW_INV U35 ( .A(A[7]), .Z(n248) );
    VMW_INV U36 ( .A(A[3]), .Z(n234) );
    VMW_INV U37 ( .A(B[3]), .Z(n231) );
    VMW_INV U38 ( .A(A[10]), .Z(n250) );
    VMW_INV U39 ( .A(B[9]), .Z(n252) );
    VMW_INV U40 ( .A(A[4]), .Z(n229) );
    VMW_INV U41 ( .A(A[8]), .Z(n243) );
    VMW_INV U42 ( .A(A[14]), .Z(n262) );
    VMW_INV U43 ( .A(B[11]), .Z(n258) );
    VMW_INV U44 ( .A(A[5]), .Z(n241) );
    VMW_INV U45 ( .A(B[5]), .Z(n238) );
    VMW_INV U46 ( .A(A[1]), .Z(n225) );
    VMW_INV U47 ( .A(B[15]), .Z(n267) );
    VMW_INV U48 ( .A(B[13]), .Z(n264) );
    VMW_INV U49 ( .A(A[6]), .Z(n236) );
    VMW_INV U50 ( .A(A[2]), .Z(n222) );
    VMW_INV U51 ( .A(A[0]), .Z(n224) );
    VMW_INV U52 ( .A(A[15]), .Z(n219) );
endmodule


module NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
        n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
        n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
        n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
        n315, n316;
    VMW_OAI21 U3 ( .A(B[15]), .B(n268), .C(n269), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n271), .B(B[2]), .Z(n270) );
    VMW_AO22 U5 ( .A(n273), .B(B[0]), .C(n274), .D(B[1]), .Z(n272) );
    VMW_OR2 U6 ( .A(B[2]), .B(n271), .Z(n275) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n274), .C(n275), .D(n272), .Z(n276) );
    VMW_NAND2 U8 ( .A(n278), .B(B[4]), .Z(n277) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n280), .C(n276), .D(n270), .Z(n279) );
    VMW_OR2 U10 ( .A(B[4]), .B(n278), .Z(n281) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n283), .C(n281), .D(n279), .Z(n282) );
    VMW_NAND2 U12 ( .A(n285), .B(B[6]), .Z(n284) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n287), .C(n282), .D(n277), .Z(n286) );
    VMW_OR2 U14 ( .A(B[6]), .B(n285), .Z(n288) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n290), .C(n288), .D(n286), .Z(n289) );
    VMW_NAND2 U16 ( .A(n292), .B(B[8]), .Z(n291) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n294), .C(n289), .D(n284), .Z(n293) );
    VMW_OR2 U18 ( .A(B[8]), .B(n292), .Z(n295) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n297), .C(n295), .D(n293), .Z(n296) );
    VMW_NAND2 U20 ( .A(n299), .B(B[10]), .Z(n298) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n301), .C(n296), .D(n291), .Z(n300) );
    VMW_NAND2 U22 ( .A(n301), .B(A[9]), .Z(n302) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n299), .C(n302), .D(n300), .Z(n303) );
    VMW_NAND2 U24 ( .A(n305), .B(B[12]), .Z(n304) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n307), .C(n303), .D(n298), .Z(n306) );
    VMW_NAND2 U26 ( .A(n307), .B(A[11]), .Z(n308) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n305), .C(n308), .D(n306), .Z(n309) );
    VMW_NAND2 U28 ( .A(n311), .B(B[14]), .Z(n310) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n313), .C(n309), .D(n304), .Z(n312) );
    VMW_NAND2 U30 ( .A(n313), .B(A[13]), .Z(n314) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n311), .C(n314), .D(n312), .Z(n315) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n316), .C(n315), .D(n310), .Z(n269) );
    VMW_INV U33 ( .A(A[12]), .Z(n305) );
    VMW_INV U34 ( .A(B[7]), .Z(n294) );
    VMW_INV U35 ( .A(A[7]), .Z(n297) );
    VMW_INV U36 ( .A(A[3]), .Z(n283) );
    VMW_INV U37 ( .A(B[3]), .Z(n280) );
    VMW_INV U38 ( .A(A[10]), .Z(n299) );
    VMW_INV U39 ( .A(B[9]), .Z(n301) );
    VMW_INV U40 ( .A(A[4]), .Z(n278) );
    VMW_INV U41 ( .A(A[8]), .Z(n292) );
    VMW_INV U42 ( .A(A[14]), .Z(n311) );
    VMW_INV U43 ( .A(B[11]), .Z(n307) );
    VMW_INV U44 ( .A(A[5]), .Z(n290) );
    VMW_INV U45 ( .A(B[5]), .Z(n287) );
    VMW_INV U46 ( .A(A[1]), .Z(n274) );
    VMW_INV U47 ( .A(B[15]), .Z(n316) );
    VMW_INV U48 ( .A(B[13]), .Z(n313) );
    VMW_INV U49 ( .A(A[6]), .Z(n285) );
    VMW_INV U50 ( .A(A[2]), .Z(n271) );
    VMW_INV U51 ( .A(A[0]), .Z(n273) );
    VMW_INV U52 ( .A(A[15]), .Z(n268) );
endmodule


module NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
        n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
        n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
        n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
        n364, n365;
    VMW_OAI21 U3 ( .A(B[15]), .B(n317), .C(n318), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n320), .B(B[2]), .Z(n319) );
    VMW_AO22 U5 ( .A(n322), .B(B[0]), .C(n323), .D(B[1]), .Z(n321) );
    VMW_OR2 U6 ( .A(B[2]), .B(n320), .Z(n324) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n323), .C(n324), .D(n321), .Z(n325) );
    VMW_NAND2 U8 ( .A(n327), .B(B[4]), .Z(n326) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n329), .C(n325), .D(n319), .Z(n328) );
    VMW_OR2 U10 ( .A(B[4]), .B(n327), .Z(n330) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n332), .C(n330), .D(n328), .Z(n331) );
    VMW_NAND2 U12 ( .A(n334), .B(B[6]), .Z(n333) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n336), .C(n331), .D(n326), .Z(n335) );
    VMW_OR2 U14 ( .A(B[6]), .B(n334), .Z(n337) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n339), .C(n337), .D(n335), .Z(n338) );
    VMW_NAND2 U16 ( .A(n341), .B(B[8]), .Z(n340) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n343), .C(n338), .D(n333), .Z(n342) );
    VMW_OR2 U18 ( .A(B[8]), .B(n341), .Z(n344) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n346), .C(n344), .D(n342), .Z(n345) );
    VMW_NAND2 U20 ( .A(n348), .B(B[10]), .Z(n347) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n350), .C(n345), .D(n340), .Z(n349) );
    VMW_NAND2 U22 ( .A(n350), .B(A[9]), .Z(n351) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n348), .C(n351), .D(n349), .Z(n352) );
    VMW_NAND2 U24 ( .A(n354), .B(B[12]), .Z(n353) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n356), .C(n352), .D(n347), .Z(n355) );
    VMW_NAND2 U26 ( .A(n356), .B(A[11]), .Z(n357) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n354), .C(n357), .D(n355), .Z(n358) );
    VMW_NAND2 U28 ( .A(n360), .B(B[14]), .Z(n359) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n362), .C(n358), .D(n353), .Z(n361) );
    VMW_NAND2 U30 ( .A(n362), .B(A[13]), .Z(n363) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n360), .C(n363), .D(n361), .Z(n364) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n365), .C(n364), .D(n359), .Z(n318) );
    VMW_INV U33 ( .A(A[12]), .Z(n354) );
    VMW_INV U34 ( .A(B[7]), .Z(n343) );
    VMW_INV U35 ( .A(A[7]), .Z(n346) );
    VMW_INV U36 ( .A(A[3]), .Z(n332) );
    VMW_INV U37 ( .A(B[3]), .Z(n329) );
    VMW_INV U38 ( .A(A[10]), .Z(n348) );
    VMW_INV U39 ( .A(B[9]), .Z(n350) );
    VMW_INV U40 ( .A(A[4]), .Z(n327) );
    VMW_INV U41 ( .A(A[8]), .Z(n341) );
    VMW_INV U42 ( .A(A[14]), .Z(n360) );
    VMW_INV U43 ( .A(B[11]), .Z(n356) );
    VMW_INV U44 ( .A(A[5]), .Z(n339) );
    VMW_INV U45 ( .A(B[5]), .Z(n336) );
    VMW_INV U46 ( .A(A[1]), .Z(n323) );
    VMW_INV U47 ( .A(B[15]), .Z(n365) );
    VMW_INV U48 ( .A(B[13]), .Z(n362) );
    VMW_INV U49 ( .A(A[6]), .Z(n334) );
    VMW_INV U50 ( .A(A[2]), .Z(n320) );
    VMW_INV U51 ( .A(A[0]), .Z(n322) );
    VMW_INV U52 ( .A(A[15]), .Z(n317) );
endmodule


module NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
        n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
        n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
        n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
        n413, n414;
    VMW_OAI21 U3 ( .A(B[15]), .B(n366), .C(n367), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n369), .B(B[2]), .Z(n368) );
    VMW_AO22 U5 ( .A(n371), .B(B[0]), .C(n372), .D(B[1]), .Z(n370) );
    VMW_OR2 U6 ( .A(B[2]), .B(n369), .Z(n373) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n372), .C(n373), .D(n370), .Z(n374) );
    VMW_NAND2 U8 ( .A(n376), .B(B[4]), .Z(n375) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n378), .C(n374), .D(n368), .Z(n377) );
    VMW_OR2 U10 ( .A(B[4]), .B(n376), .Z(n379) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n381), .C(n379), .D(n377), .Z(n380) );
    VMW_NAND2 U12 ( .A(n383), .B(B[6]), .Z(n382) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n385), .C(n380), .D(n375), .Z(n384) );
    VMW_OR2 U14 ( .A(B[6]), .B(n383), .Z(n386) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n388), .C(n386), .D(n384), .Z(n387) );
    VMW_NAND2 U16 ( .A(n390), .B(B[8]), .Z(n389) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n392), .C(n387), .D(n382), .Z(n391) );
    VMW_OR2 U18 ( .A(B[8]), .B(n390), .Z(n393) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n395), .C(n393), .D(n391), .Z(n394) );
    VMW_NAND2 U20 ( .A(n397), .B(B[10]), .Z(n396) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n399), .C(n394), .D(n389), .Z(n398) );
    VMW_NAND2 U22 ( .A(n399), .B(A[9]), .Z(n400) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n397), .C(n400), .D(n398), .Z(n401) );
    VMW_NAND2 U24 ( .A(n403), .B(B[12]), .Z(n402) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n405), .C(n401), .D(n396), .Z(n404) );
    VMW_NAND2 U26 ( .A(n405), .B(A[11]), .Z(n406) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n403), .C(n406), .D(n404), .Z(n407) );
    VMW_NAND2 U28 ( .A(n409), .B(B[14]), .Z(n408) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n411), .C(n407), .D(n402), .Z(n410) );
    VMW_NAND2 U30 ( .A(n411), .B(A[13]), .Z(n412) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n409), .C(n412), .D(n410), .Z(n413) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n414), .C(n413), .D(n408), .Z(n367) );
    VMW_INV U33 ( .A(A[12]), .Z(n403) );
    VMW_INV U34 ( .A(B[7]), .Z(n392) );
    VMW_INV U35 ( .A(A[7]), .Z(n395) );
    VMW_INV U36 ( .A(A[3]), .Z(n381) );
    VMW_INV U37 ( .A(B[3]), .Z(n378) );
    VMW_INV U38 ( .A(A[10]), .Z(n397) );
    VMW_INV U39 ( .A(B[9]), .Z(n399) );
    VMW_INV U40 ( .A(A[4]), .Z(n376) );
    VMW_INV U41 ( .A(A[8]), .Z(n390) );
    VMW_INV U42 ( .A(A[14]), .Z(n409) );
    VMW_INV U43 ( .A(B[11]), .Z(n405) );
    VMW_INV U44 ( .A(A[5]), .Z(n388) );
    VMW_INV U45 ( .A(B[5]), .Z(n385) );
    VMW_INV U46 ( .A(A[1]), .Z(n372) );
    VMW_INV U47 ( .A(B[15]), .Z(n414) );
    VMW_INV U48 ( .A(B[13]), .Z(n411) );
    VMW_INV U49 ( .A(A[6]), .Z(n383) );
    VMW_INV U50 ( .A(A[2]), .Z(n369) );
    VMW_INV U51 ( .A(A[0]), .Z(n371) );
    VMW_INV U52 ( .A(A[15]), .Z(n366) );
endmodule


module NodeAux_INDEGREE8_SOURCE1 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp240[2] , \temp334[3] , \temp424[2] , \temp604[10] , 
        \temp424[14] , n152, \temp694[10] , \temp604[3] , \temp784[12] , n112, 
        \temp424[10] , \temp604[14] , \temp424[6] , \temp240[6] , \temp334[7] , 
        \path[2] , \temp604[7] , \temp694[14] , \path[0] , \temp604[5] , 
        \temp784[14] , \temp424[4] , \temp240[4] , \temp334[5] , \temp424[12] , 
        \temp334[8] , n120, \temp784[10] , \temp240[9] , \temp424[9] , 
        \temp694[12] , \temp604[1] , \temp604[8] , \temp604[12] , \temp334[1] , 
        \temp424[0] , \temp240[0] , \temp240[14] , \temp514[3] , \temp334[10] , 
        \temp694[2] , \temp784[7] , \temp514[13] , \OutEdge166[13] , 
        \OutEdge166[3] , n128, \temp694[6] , \temp784[3] , \temp334[14] , 
        \temp514[7] , \OutEdge166[7] , \temp240[10] , \temp784[8] , 
        \temp514[15] , \OutEdge166[15] , \OutEdge166[5] , n96, \temp514[5] , 
        \temp240[12] , \temp784[1] , \temp694[4] , \temp514[8] , 
        \OutEdge166[11] , \OutEdge166[1] , \temp694[9] , \temp514[11] , 
        \temp334[12] , \temp694[0] , \temp784[5] , \temp514[1] , 
        \OutEdge166[8] , \temp514[9] , \OutEdge166[10] , \OutEdge166[0] , 
        \temp694[8] , \temp514[10] , \temp694[1] , \temp334[13] , \temp514[0] , 
        \temp784[4] , \OutEdge166[9] , \temp514[14] , \temp784[9] , n136, 
        \OutEdge166[14] , \OutEdge166[4] , \temp240[13] , \temp514[4] , 
        \temp784[0] , \temp694[5] , \temp784[2] , \temp334[15] , \temp694[7] , 
        \temp240[11] , \temp514[6] , n144, \OutEdge166[6] , \temp514[2] , n104, 
        \temp240[15] , \temp694[3] , \temp334[11] , \temp784[6] , 
        \temp514[12] , \OutEdge166[12] , \OutEdge166[2] , \temp334[9] , 
        \temp240[8] , \temp424[8] , \temp784[11] , \temp694[13] , \temp604[0] , 
        \temp604[13] , \temp604[9] , \temp334[0] , \temp240[1] , \temp424[1] , 
        \path[1] , \temp604[4] , \temp784[15] , \temp424[5] , \temp240[5] , 
        \temp334[4] , \temp424[13] , \temp424[11] , \temp604[15] , 
        \temp424[7] , \temp240[7] , \temp334[6] , \path[3] , \temp694[15] , 
        \temp604[6] , \temp334[2] , \temp424[3] , \temp240[3] , \temp604[11] , 
        \temp424[15] , \temp604[2] , \temp694[11] , \temp784[13] , n967, n968, 
        n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
        n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
        n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
        n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U109 ( .Z(n1006) );
    VMW_PULLDOWN U110 ( .Z(n1005) );
    VMW_PULLDOWN U111 ( .Z(n1008) );
    VMW_PULLDOWN U112 ( .Z(n1009) );
    VMW_PULLDOWN U113 ( .Z(n1004) );
    VMW_PULLDOWN U114 ( .Z(n1011) );
    VMW_PULLDOWN U115 ( .Z(n1007) );
    VMW_PULLDOWN U116 ( .Z(n1010) );
    VMW_AO22 U117 ( .A(InEdges[127]), .B(n967), .C(n968), .D(\temp784[15] ), 
        .Z(\OutEdge166[15] ) );
    VMW_AO22 U118 ( .A(InEdges[126]), .B(n967), .C(n968), .D(\temp784[14] ), 
        .Z(\OutEdge166[14] ) );
    VMW_AO22 U119 ( .A(InEdges[125]), .B(n967), .C(n968), .D(\temp784[13] ), 
        .Z(\OutEdge166[13] ) );
    VMW_AO22 U120 ( .A(InEdges[124]), .B(n967), .C(n968), .D(\temp784[12] ), 
        .Z(\OutEdge166[12] ) );
    VMW_AO22 U121 ( .A(InEdges[123]), .B(n967), .C(n968), .D(\temp784[11] ), 
        .Z(\OutEdge166[11] ) );
    VMW_AO22 U122 ( .A(InEdges[122]), .B(n967), .C(n968), .D(\temp784[10] ), 
        .Z(\OutEdge166[10] ) );
    VMW_AO22 U123 ( .A(InEdges[121]), .B(n967), .C(n968), .D(\temp784[9] ), 
        .Z(\OutEdge166[9] ) );
    VMW_AO22 U124 ( .A(InEdges[120]), .B(n967), .C(n968), .D(\temp784[8] ), 
        .Z(\OutEdge166[8] ) );
    VMW_AO22 U125 ( .A(InEdges[119]), .B(n967), .C(n968), .D(\temp784[7] ), 
        .Z(\OutEdge166[7] ) );
    VMW_AO22 U126 ( .A(InEdges[118]), .B(n967), .C(n968), .D(\temp784[6] ), 
        .Z(\OutEdge166[6] ) );
    VMW_AO22 U127 ( .A(InEdges[117]), .B(n967), .C(n968), .D(\temp784[5] ), 
        .Z(\OutEdge166[5] ) );
    VMW_AO22 U128 ( .A(InEdges[116]), .B(n967), .C(n968), .D(\temp784[4] ), 
        .Z(\OutEdge166[4] ) );
    VMW_AO22 U129 ( .A(InEdges[115]), .B(n967), .C(n968), .D(\temp784[3] ), 
        .Z(\OutEdge166[3] ) );
    VMW_AO22 U130 ( .A(InEdges[114]), .B(n967), .C(n968), .D(\temp784[2] ), 
        .Z(\OutEdge166[2] ) );
    VMW_AO22 U131 ( .A(InEdges[113]), .B(n967), .C(n968), .D(\temp784[1] ), 
        .Z(\OutEdge166[1] ) );
    VMW_AO22 U132 ( .A(InEdges[112]), .B(n967), .C(n968), .D(\temp784[0] ), 
        .Z(\OutEdge166[0] ) );
    VMW_OR2 U133 ( .A(n969), .B(n967), .Z(n1003) );
    VMW_AO21 U134 ( .A(Start), .B(\path[3] ), .C(n970), .Z(n1002) );
    VMW_NAND2 U135 ( .A(n971), .B(n972), .Z(n1001) );
    VMW_NAND2 U136 ( .A(n971), .B(n973), .Z(n1000) );
    VMW_AND5 U137 ( .A(n974), .B(n968), .C(n975), .D(n976), .E(n977), .Z(n970)
         );
    VMW_OR4 U138 ( .A(n144), .B(n136), .C(n128), .D(n974), .Z(n978) );
    VMW_AO22 U139 ( .A(\temp694[9] ), .B(n976), .C(InEdges[105]), .D(n144), 
        .Z(\temp784[9] ) );
    VMW_AO22 U140 ( .A(\temp694[8] ), .B(n976), .C(InEdges[104]), .D(n144), 
        .Z(\temp784[8] ) );
    VMW_AO22 U141 ( .A(\temp694[7] ), .B(n976), .C(InEdges[103]), .D(n144), 
        .Z(\temp784[7] ) );
    VMW_AO22 U142 ( .A(\temp694[6] ), .B(n976), .C(InEdges[102]), .D(n144), 
        .Z(\temp784[6] ) );
    VMW_AO22 U143 ( .A(\temp694[5] ), .B(n976), .C(InEdges[101]), .D(n144), 
        .Z(\temp784[5] ) );
    VMW_AO22 U144 ( .A(\temp694[4] ), .B(n976), .C(InEdges[100]), .D(n144), 
        .Z(\temp784[4] ) );
    VMW_AO22 U145 ( .A(\temp694[3] ), .B(n976), .C(InEdges[99]), .D(n144), .Z(
        \temp784[3] ) );
    VMW_AO22 U146 ( .A(\temp694[2] ), .B(n976), .C(InEdges[98]), .D(n144), .Z(
        \temp784[2] ) );
    VMW_AO22 U147 ( .A(\temp694[1] ), .B(n976), .C(InEdges[97]), .D(n144), .Z(
        \temp784[1] ) );
    VMW_AO22 U148 ( .A(\temp694[15] ), .B(n976), .C(InEdges[111]), .D(n144), 
        .Z(\temp784[15] ) );
    VMW_AO22 U149 ( .A(\temp694[14] ), .B(n976), .C(InEdges[110]), .D(n144), 
        .Z(\temp784[14] ) );
    VMW_AO22 U150 ( .A(\temp694[13] ), .B(n976), .C(InEdges[109]), .D(n144), 
        .Z(\temp784[13] ) );
    VMW_AO22 U151 ( .A(\temp694[12] ), .B(n976), .C(InEdges[108]), .D(n144), 
        .Z(\temp784[12] ) );
    VMW_AO22 U152 ( .A(\temp694[11] ), .B(n976), .C(InEdges[107]), .D(n144), 
        .Z(\temp784[11] ) );
    VMW_AO22 U153 ( .A(\temp694[10] ), .B(n976), .C(InEdges[106]), .D(n144), 
        .Z(\temp784[10] ) );
    VMW_AO22 U154 ( .A(\temp694[0] ), .B(n976), .C(InEdges[96]), .D(n144), .Z(
        \temp784[0] ) );
    VMW_AND4 U155 ( .A(n979), .B(n980), .C(n981), .D(n982), .Z(n974) );
    VMW_NOR2 U156 ( .A(Start), .B(n152), .Z(n968) );
    VMW_AND2 U157 ( .A(n152), .B(n983), .Z(n967) );
    VMW_OAI22 U158 ( .A(n978), .B(Start), .C(\path[2] ), .D(n983), .Z(n972) );
    VMW_AO21 U159 ( .A(n985), .B(n986), .C(n144), .Z(n984) );
    VMW_OAI22 U160 ( .A(n987), .B(Start), .C(\path[0] ), .D(n983), .Z(n973) );
    VMW_AND2 U161 ( .A(n977), .B(n975), .Z(n985) );
    VMW_AND4 U162 ( .A(n989), .B(n990), .C(n991), .D(n992), .Z(n988) );
    VMW_INV U163 ( .A(n120), .Z(n982) );
    VMW_INV U164 ( .A(n136), .Z(n977) );
    VMW_INV U165 ( .A(n112), .Z(n980) );
    VMW_OAI211 U166 ( .A(n96), .B(n104), .C(n980), .D(n982), .Z(n986) );
    VMW_AO21 U167 ( .A(n979), .B(n96), .C(n112), .Z(n993) );
    VMW_AO21 U168 ( .A(n982), .B(n993), .C(n128), .Z(n994) );
    VMW_AND5 U169 ( .A(n995), .B(n996), .C(n997), .D(n998), .E(n988), .Z(n999)
         );
    VMW_XNOR2 U170 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n992) );
    VMW_XNOR2 U171 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n991) );
    VMW_XNOR2 U172 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n990) );
    VMW_XNOR2 U173 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n989) );
    VMW_XNOR2 U174 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n998) );
    VMW_XNOR2 U175 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n997) );
    VMW_XNOR2 U176 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n996) );
    VMW_XNOR2 U177 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n995) );
    VMW_AO22 U178 ( .A(InEdges[9]), .B(n96), .C(OutEdge[9]), .D(n981), .Z(
        \temp240[9] ) );
    VMW_AO22 U179 ( .A(\temp240[9] ), .B(n979), .C(InEdges[25]), .D(n104), .Z(
        \temp334[9] ) );
    VMW_AO22 U180 ( .A(InEdges[41]), .B(n112), .C(\temp334[9] ), .D(n980), .Z(
        \temp424[9] ) );
    VMW_AO22 U181 ( .A(InEdges[57]), .B(n120), .C(\temp424[9] ), .D(n982), .Z(
        \temp514[9] ) );
    VMW_AO22 U182 ( .A(\temp514[9] ), .B(n975), .C(InEdges[73]), .D(n128), .Z(
        \temp604[9] ) );
    VMW_AO22 U183 ( .A(InEdges[89]), .B(n136), .C(\temp604[9] ), .D(n977), .Z(
        \temp694[9] ) );
    VMW_AO22 U184 ( .A(InEdges[8]), .B(n96), .C(OutEdge[8]), .D(n981), .Z(
        \temp240[8] ) );
    VMW_AO22 U185 ( .A(\temp240[8] ), .B(n979), .C(InEdges[24]), .D(n104), .Z(
        \temp334[8] ) );
    VMW_AO22 U186 ( .A(InEdges[40]), .B(n112), .C(\temp334[8] ), .D(n980), .Z(
        \temp424[8] ) );
    VMW_AO22 U187 ( .A(InEdges[56]), .B(n120), .C(\temp424[8] ), .D(n982), .Z(
        \temp514[8] ) );
    VMW_AO22 U188 ( .A(\temp514[8] ), .B(n975), .C(InEdges[72]), .D(n128), .Z(
        \temp604[8] ) );
    VMW_AO22 U189 ( .A(InEdges[88]), .B(n136), .C(\temp604[8] ), .D(n977), .Z(
        \temp694[8] ) );
    VMW_AO22 U190 ( .A(InEdges[7]), .B(n96), .C(OutEdge[7]), .D(n981), .Z(
        \temp240[7] ) );
    VMW_AO22 U191 ( .A(\temp240[7] ), .B(n979), .C(InEdges[23]), .D(n104), .Z(
        \temp334[7] ) );
    VMW_AO22 U192 ( .A(InEdges[39]), .B(n112), .C(\temp334[7] ), .D(n980), .Z(
        \temp424[7] ) );
    VMW_AO22 U193 ( .A(InEdges[55]), .B(n120), .C(\temp424[7] ), .D(n982), .Z(
        \temp514[7] ) );
    VMW_AO22 U194 ( .A(\temp514[7] ), .B(n975), .C(InEdges[71]), .D(n128), .Z(
        \temp604[7] ) );
    VMW_AO22 U195 ( .A(InEdges[87]), .B(n136), .C(\temp604[7] ), .D(n977), .Z(
        \temp694[7] ) );
    VMW_AO22 U196 ( .A(InEdges[6]), .B(n96), .C(OutEdge[6]), .D(n981), .Z(
        \temp240[6] ) );
    VMW_AO22 U197 ( .A(\temp240[6] ), .B(n979), .C(InEdges[22]), .D(n104), .Z(
        \temp334[6] ) );
    VMW_AO22 U198 ( .A(InEdges[38]), .B(n112), .C(\temp334[6] ), .D(n980), .Z(
        \temp424[6] ) );
    VMW_AO22 U199 ( .A(InEdges[54]), .B(n120), .C(\temp424[6] ), .D(n982), .Z(
        \temp514[6] ) );
    VMW_AO22 U200 ( .A(\temp514[6] ), .B(n975), .C(InEdges[70]), .D(n128), .Z(
        \temp604[6] ) );
    VMW_AO22 U201 ( .A(InEdges[86]), .B(n136), .C(\temp604[6] ), .D(n977), .Z(
        \temp694[6] ) );
    VMW_AO22 U202 ( .A(InEdges[5]), .B(n96), .C(OutEdge[5]), .D(n981), .Z(
        \temp240[5] ) );
    VMW_AO22 U203 ( .A(\temp240[5] ), .B(n979), .C(InEdges[21]), .D(n104), .Z(
        \temp334[5] ) );
    VMW_AO22 U204 ( .A(InEdges[37]), .B(n112), .C(\temp334[5] ), .D(n980), .Z(
        \temp424[5] ) );
    VMW_AO22 U205 ( .A(InEdges[53]), .B(n120), .C(\temp424[5] ), .D(n982), .Z(
        \temp514[5] ) );
    VMW_AO22 U206 ( .A(\temp514[5] ), .B(n975), .C(InEdges[69]), .D(n128), .Z(
        \temp604[5] ) );
    VMW_AO22 U207 ( .A(InEdges[85]), .B(n136), .C(\temp604[5] ), .D(n977), .Z(
        \temp694[5] ) );
    VMW_AO22 U208 ( .A(InEdges[4]), .B(n96), .C(OutEdge[4]), .D(n981), .Z(
        \temp240[4] ) );
    VMW_AO22 U209 ( .A(\temp240[4] ), .B(n979), .C(InEdges[20]), .D(n104), .Z(
        \temp334[4] ) );
    VMW_AO22 U210 ( .A(InEdges[36]), .B(n112), .C(\temp334[4] ), .D(n980), .Z(
        \temp424[4] ) );
    VMW_AO22 U211 ( .A(InEdges[52]), .B(n120), .C(\temp424[4] ), .D(n982), .Z(
        \temp514[4] ) );
    VMW_AO22 U212 ( .A(\temp514[4] ), .B(n975), .C(InEdges[68]), .D(n128), .Z(
        \temp604[4] ) );
    VMW_AO22 U213 ( .A(InEdges[84]), .B(n136), .C(\temp604[4] ), .D(n977), .Z(
        \temp694[4] ) );
    VMW_AO22 U214 ( .A(InEdges[3]), .B(n96), .C(OutEdge[3]), .D(n981), .Z(
        \temp240[3] ) );
    VMW_AO22 U215 ( .A(\temp240[3] ), .B(n979), .C(InEdges[19]), .D(n104), .Z(
        \temp334[3] ) );
    VMW_AO22 U216 ( .A(InEdges[35]), .B(n112), .C(\temp334[3] ), .D(n980), .Z(
        \temp424[3] ) );
    VMW_AO22 U217 ( .A(InEdges[51]), .B(n120), .C(\temp424[3] ), .D(n982), .Z(
        \temp514[3] ) );
    VMW_AO22 U218 ( .A(\temp514[3] ), .B(n975), .C(InEdges[67]), .D(n128), .Z(
        \temp604[3] ) );
    VMW_AO22 U219 ( .A(InEdges[83]), .B(n136), .C(\temp604[3] ), .D(n977), .Z(
        \temp694[3] ) );
    VMW_AO22 U220 ( .A(InEdges[2]), .B(n96), .C(OutEdge[2]), .D(n981), .Z(
        \temp240[2] ) );
    VMW_AO22 U221 ( .A(\temp240[2] ), .B(n979), .C(InEdges[18]), .D(n104), .Z(
        \temp334[2] ) );
    VMW_AO22 U222 ( .A(InEdges[34]), .B(n112), .C(\temp334[2] ), .D(n980), .Z(
        \temp424[2] ) );
    VMW_AO22 U223 ( .A(InEdges[50]), .B(n120), .C(\temp424[2] ), .D(n982), .Z(
        \temp514[2] ) );
    VMW_AO22 U224 ( .A(\temp514[2] ), .B(n975), .C(InEdges[66]), .D(n128), .Z(
        \temp604[2] ) );
    VMW_AO22 U225 ( .A(InEdges[82]), .B(n136), .C(\temp604[2] ), .D(n977), .Z(
        \temp694[2] ) );
    VMW_AO22 U226 ( .A(InEdges[1]), .B(n96), .C(OutEdge[1]), .D(n981), .Z(
        \temp240[1] ) );
    VMW_AO22 U227 ( .A(\temp240[1] ), .B(n979), .C(InEdges[17]), .D(n104), .Z(
        \temp334[1] ) );
    VMW_AO22 U228 ( .A(InEdges[33]), .B(n112), .C(\temp334[1] ), .D(n980), .Z(
        \temp424[1] ) );
    VMW_AO22 U229 ( .A(InEdges[49]), .B(n120), .C(\temp424[1] ), .D(n982), .Z(
        \temp514[1] ) );
    VMW_AO22 U230 ( .A(\temp514[1] ), .B(n975), .C(InEdges[65]), .D(n128), .Z(
        \temp604[1] ) );
    VMW_AO22 U231 ( .A(InEdges[81]), .B(n136), .C(\temp604[1] ), .D(n977), .Z(
        \temp694[1] ) );
    VMW_AO22 U232 ( .A(InEdges[15]), .B(n96), .C(OutEdge[15]), .D(n981), .Z(
        \temp240[15] ) );
    VMW_AO22 U233 ( .A(\temp240[15] ), .B(n979), .C(InEdges[31]), .D(n104), 
        .Z(\temp334[15] ) );
    VMW_AO22 U234 ( .A(InEdges[47]), .B(n112), .C(\temp334[15] ), .D(n980), 
        .Z(\temp424[15] ) );
    VMW_AO22 U235 ( .A(InEdges[63]), .B(n120), .C(\temp424[15] ), .D(n982), 
        .Z(\temp514[15] ) );
    VMW_AO22 U236 ( .A(\temp514[15] ), .B(n975), .C(InEdges[79]), .D(n128), 
        .Z(\temp604[15] ) );
    VMW_AO22 U237 ( .A(InEdges[95]), .B(n136), .C(\temp604[15] ), .D(n977), 
        .Z(\temp694[15] ) );
    VMW_AO22 U238 ( .A(InEdges[14]), .B(n96), .C(OutEdge[14]), .D(n981), .Z(
        \temp240[14] ) );
    VMW_AO22 U239 ( .A(\temp240[14] ), .B(n979), .C(InEdges[30]), .D(n104), 
        .Z(\temp334[14] ) );
    VMW_AO22 U240 ( .A(InEdges[46]), .B(n112), .C(\temp334[14] ), .D(n980), 
        .Z(\temp424[14] ) );
    VMW_AO22 U241 ( .A(InEdges[62]), .B(n120), .C(\temp424[14] ), .D(n982), 
        .Z(\temp514[14] ) );
    VMW_AO22 U242 ( .A(\temp514[14] ), .B(n975), .C(InEdges[78]), .D(n128), 
        .Z(\temp604[14] ) );
    VMW_AO22 U243 ( .A(InEdges[94]), .B(n136), .C(\temp604[14] ), .D(n977), 
        .Z(\temp694[14] ) );
    VMW_AO22 U244 ( .A(InEdges[13]), .B(n96), .C(OutEdge[13]), .D(n981), .Z(
        \temp240[13] ) );
    VMW_AO22 U245 ( .A(\temp240[13] ), .B(n979), .C(InEdges[29]), .D(n104), 
        .Z(\temp334[13] ) );
    VMW_AO22 U246 ( .A(InEdges[45]), .B(n112), .C(\temp334[13] ), .D(n980), 
        .Z(\temp424[13] ) );
    VMW_AO22 U247 ( .A(InEdges[61]), .B(n120), .C(\temp424[13] ), .D(n982), 
        .Z(\temp514[13] ) );
    VMW_AO22 U248 ( .A(\temp514[13] ), .B(n975), .C(InEdges[77]), .D(n128), 
        .Z(\temp604[13] ) );
    VMW_AO22 U249 ( .A(InEdges[93]), .B(n136), .C(\temp604[13] ), .D(n977), 
        .Z(\temp694[13] ) );
    VMW_AO22 U250 ( .A(InEdges[12]), .B(n96), .C(OutEdge[12]), .D(n981), .Z(
        \temp240[12] ) );
    VMW_AO22 U251 ( .A(\temp240[12] ), .B(n979), .C(InEdges[28]), .D(n104), 
        .Z(\temp334[12] ) );
    VMW_AO22 U252 ( .A(InEdges[44]), .B(n112), .C(\temp334[12] ), .D(n980), 
        .Z(\temp424[12] ) );
    VMW_AO22 U253 ( .A(InEdges[60]), .B(n120), .C(\temp424[12] ), .D(n982), 
        .Z(\temp514[12] ) );
    VMW_AO22 U254 ( .A(\temp514[12] ), .B(n975), .C(InEdges[76]), .D(n128), 
        .Z(\temp604[12] ) );
    VMW_AO22 U255 ( .A(InEdges[92]), .B(n136), .C(\temp604[12] ), .D(n977), 
        .Z(\temp694[12] ) );
    VMW_AO22 U256 ( .A(InEdges[11]), .B(n96), .C(OutEdge[11]), .D(n981), .Z(
        \temp240[11] ) );
    VMW_AO22 U257 ( .A(\temp240[11] ), .B(n979), .C(InEdges[27]), .D(n104), 
        .Z(\temp334[11] ) );
    VMW_AO22 U258 ( .A(InEdges[43]), .B(n112), .C(\temp334[11] ), .D(n980), 
        .Z(\temp424[11] ) );
    VMW_AO22 U259 ( .A(InEdges[59]), .B(n120), .C(\temp424[11] ), .D(n982), 
        .Z(\temp514[11] ) );
    VMW_AO22 U260 ( .A(\temp514[11] ), .B(n975), .C(InEdges[75]), .D(n128), 
        .Z(\temp604[11] ) );
    VMW_AO22 U261 ( .A(InEdges[91]), .B(n136), .C(\temp604[11] ), .D(n977), 
        .Z(\temp694[11] ) );
    VMW_AO22 U262 ( .A(InEdges[10]), .B(n96), .C(OutEdge[10]), .D(n981), .Z(
        \temp240[10] ) );
    VMW_AO22 U263 ( .A(\temp240[10] ), .B(n979), .C(InEdges[26]), .D(n104), 
        .Z(\temp334[10] ) );
    VMW_AO22 U264 ( .A(InEdges[42]), .B(n112), .C(\temp334[10] ), .D(n980), 
        .Z(\temp424[10] ) );
    VMW_AO22 U265 ( .A(InEdges[58]), .B(n120), .C(\temp424[10] ), .D(n982), 
        .Z(\temp514[10] ) );
    VMW_AO22 U266 ( .A(\temp514[10] ), .B(n975), .C(InEdges[74]), .D(n128), 
        .Z(\temp604[10] ) );
    VMW_AO22 U267 ( .A(InEdges[90]), .B(n136), .C(\temp604[10] ), .D(n977), 
        .Z(\temp694[10] ) );
    VMW_AO22 U268 ( .A(InEdges[0]), .B(n96), .C(OutEdge[0]), .D(n981), .Z(
        \temp240[0] ) );
    VMW_AO22 U269 ( .A(\temp240[0] ), .B(n979), .C(InEdges[16]), .D(n104), .Z(
        \temp334[0] ) );
    VMW_AO22 U270 ( .A(InEdges[32]), .B(n112), .C(\temp334[0] ), .D(n980), .Z(
        \temp424[0] ) );
    VMW_AO22 U271 ( .A(InEdges[48]), .B(n120), .C(\temp424[0] ), .D(n982), .Z(
        \temp514[0] ) );
    VMW_AO22 U272 ( .A(\temp514[0] ), .B(n975), .C(InEdges[64]), .D(n128), .Z(
        \temp604[0] ) );
    VMW_AO22 U273 ( .A(InEdges[80]), .B(n136), .C(\temp604[0] ), .D(n977), .Z(
        \temp694[0] ) );
    VMW_AO22 U274 ( .A(n984), .B(n983), .C(\path[1] ), .D(Start), .Z(n969) );
    VMW_AOI21 U275 ( .A(n977), .B(n994), .C(n144), .Z(n987) );
    VMW_INV U276 ( .A(n128), .Z(n975) );
    VMW_INV U277 ( .A(n144), .Z(n976) );
    VMW_INV U278 ( .A(n96), .Z(n981) );
    VMW_INV U279 ( .A(n104), .Z(n979) );
    VMW_INV U280 ( .A(Start), .Z(n983) );
    VMW_INV U281 ( .A(n967), .Z(n971) );
    VMW_BUFIZ U282 ( .A(\path[3] ), .E(n999), .Z(\PathData[3] ) );
    VMW_BUFIZ U283 ( .A(\path[1] ), .E(n999), .Z(\PathData[1] ) );
    VMW_BUFIZ U284 ( .A(\path[0] ), .E(n999), .Z(\PathData[0] ) );
    VMW_BUFIZ U285 ( .A(\path[2] ), .E(n999), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n1000), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n1001), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n1002), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n1003), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge166[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge166[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge166[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge166[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge166[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge166[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge166[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge166[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge166[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge166[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge166[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge166[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge166[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge166[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge166[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge166[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_7 lte_55_2 ( .A({\temp334[15] , 
        \temp334[14] , \temp334[13] , \temp334[12] , \temp334[11] , 
        \temp334[10] , \temp334[9] , \temp334[8] , \temp334[7] , \temp334[6] , 
        \temp334[5] , \temp334[4] , \temp334[3] , \temp334[2] , \temp334[1] , 
        \temp334[0] }), .B(InEdges[47:32]), .LEQ(n1011), .TC(n1011), .GE_GT(
        n112) );
    NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_6 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n1010), .TC(n1010), .GE_GT(n96) );
    NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_5 lte_55_4 ( .A({\temp514[15] , 
        \temp514[14] , \temp514[13] , \temp514[12] , \temp514[11] , 
        \temp514[10] , \temp514[9] , \temp514[8] , \temp514[7] , \temp514[6] , 
        \temp514[5] , \temp514[4] , \temp514[3] , \temp514[2] , \temp514[1] , 
        \temp514[0] }), .B(InEdges[79:64]), .LEQ(n1009), .TC(n1009), .GE_GT(
        n128) );
    NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_4 lte_55_5 ( .A({\temp604[15] , 
        \temp604[14] , \temp604[13] , \temp604[12] , \temp604[11] , 
        \temp604[10] , \temp604[9] , \temp604[8] , \temp604[7] , \temp604[6] , 
        \temp604[5] , \temp604[4] , \temp604[3] , \temp604[2] , \temp604[1] , 
        \temp604[0] }), .B(InEdges[95:80]), .LEQ(n1008), .TC(n1008), .GE_GT(
        n136) );
    NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_3 lte_55_1 ( .A({\temp240[15] , 
        \temp240[14] , \temp240[13] , \temp240[12] , \temp240[11] , 
        \temp240[10] , \temp240[9] , \temp240[8] , \temp240[7] , \temp240[6] , 
        \temp240[5] , \temp240[4] , \temp240[3] , \temp240[2] , \temp240[1] , 
        \temp240[0] }), .B(InEdges[31:16]), .LEQ(n1007), .TC(n1007), .GE_GT(
        n104) );
    NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_2 lte_55_7 ( .A({\temp784[15] , 
        \temp784[14] , \temp784[13] , \temp784[12] , \temp784[11] , 
        \temp784[10] , \temp784[9] , \temp784[8] , \temp784[7] , \temp784[6] , 
        \temp784[5] , \temp784[4] , \temp784[3] , \temp784[2] , \temp784[1] , 
        \temp784[0] }), .B(InEdges[127:112]), .LEQ(n1006), .TC(n1006), .GE_GT(
        n152) );
    NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_1 lte_55_6 ( .A({\temp694[15] , 
        \temp694[14] , \temp694[13] , \temp694[12] , \temp694[11] , 
        \temp694[10] , \temp694[9] , \temp694[8] , \temp694[7] , \temp694[6] , 
        \temp694[5] , \temp694[4] , \temp694[3] , \temp694[2] , \temp694[1] , 
        \temp694[0] }), .B(InEdges[111:96]), .LEQ(n1005), .TC(n1005), .GE_GT(
        n144) );
    NodeAux_INDEGREE8_SOURCE1_DW01_cmp2_16_0 lte_55_3 ( .A({\temp424[15] , 
        \temp424[14] , \temp424[13] , \temp424[12] , \temp424[11] , 
        \temp424[10] , \temp424[9] , \temp424[8] , \temp424[7] , \temp424[6] , 
        \temp424[5] , \temp424[4] , \temp424[3] , \temp424[2] , \temp424[1] , 
        \temp424[0] }), .B(InEdges[63:48]), .LEQ(n1004), .TC(n1004), .GE_GT(
        n120) );
endmodule


module NodeAux_INDEGREE1_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE1_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , n82, \OutEdge96[11] , \OutEdge96[5] , 
        \OutEdge96[15] , \OutEdge96[8] , \OutEdge96[1] , \OutEdge96[3] , 
        \OutEdge96[7] , \OutEdge96[13] , \OutEdge96[6] , \OutEdge96[12] , 
        \OutEdge96[2] , \OutEdge96[9] , \OutEdge96[14] , \OutEdge96[0] , 
        \OutEdge96[10] , \OutEdge96[4] , \path[1] , \path[3] , n267, n268, 
        n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
        n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
        n293, n294, n295, n296, n297, n298, n299;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U46 ( .Z(n299) );
    VMW_AO22 U47 ( .A(OutEdge[15]), .B(n267), .C(n268), .D(InEdges[15]), .Z(
        \OutEdge96[15] ) );
    VMW_OR2 U48 ( .A(n269), .B(Start), .Z(\OutEdge96[14] ) );
    VMW_OR2 U49 ( .A(n270), .B(Start), .Z(\OutEdge96[13] ) );
    VMW_OR2 U50 ( .A(n271), .B(Start), .Z(\OutEdge96[12] ) );
    VMW_OR2 U51 ( .A(n272), .B(Start), .Z(\OutEdge96[11] ) );
    VMW_OR2 U52 ( .A(n273), .B(Start), .Z(\OutEdge96[10] ) );
    VMW_OR2 U53 ( .A(n274), .B(Start), .Z(\OutEdge96[9] ) );
    VMW_OR2 U54 ( .A(n275), .B(Start), .Z(\OutEdge96[8] ) );
    VMW_OR2 U55 ( .A(n276), .B(Start), .Z(\OutEdge96[7] ) );
    VMW_OR2 U56 ( .A(n277), .B(Start), .Z(\OutEdge96[6] ) );
    VMW_OR2 U57 ( .A(n278), .B(Start), .Z(\OutEdge96[5] ) );
    VMW_OR2 U58 ( .A(n279), .B(Start), .Z(\OutEdge96[4] ) );
    VMW_OR2 U59 ( .A(n280), .B(Start), .Z(\OutEdge96[3] ) );
    VMW_OR2 U60 ( .A(n281), .B(Start), .Z(\OutEdge96[2] ) );
    VMW_OR2 U61 ( .A(n282), .B(Start), .Z(\OutEdge96[1] ) );
    VMW_OR2 U62 ( .A(n283), .B(Start), .Z(\OutEdge96[0] ) );
    VMW_AO21 U63 ( .A(\path[1] ), .B(Start), .C(n267), .Z(n298) );
    VMW_AO21 U64 ( .A(Start), .B(\path[3] ), .C(n267), .Z(n297) );
    VMW_AO21 U65 ( .A(\path[2] ), .B(Start), .C(n267), .Z(n296) );
    VMW_AO21 U66 ( .A(\path[0] ), .B(Start), .C(n267), .Z(n295) );
    VMW_INV U67 ( .A(n82), .Z(n284) );
    VMW_NOR2 U68 ( .A(Start), .B(n82), .Z(n267) );
    VMW_AND4 U69 ( .A(n286), .B(n287), .C(n288), .D(n289), .Z(n285) );
    VMW_NOR2 U70 ( .A(Start), .B(n284), .Z(n268) );
    VMW_AND5 U71 ( .A(n290), .B(n291), .C(n292), .D(n293), .E(n285), .Z(n294)
         );
    VMW_XNOR2 U72 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n289) );
    VMW_XNOR2 U73 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n288) );
    VMW_XNOR2 U74 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n287) );
    VMW_XNOR2 U75 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n286) );
    VMW_XNOR2 U76 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n293) );
    VMW_XNOR2 U77 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n292) );
    VMW_XNOR2 U78 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n291) );
    VMW_XNOR2 U79 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n290) );
    VMW_AO22 U80 ( .A(InEdges[9]), .B(n82), .C(OutEdge[9]), .D(n284), .Z(n274)
         );
    VMW_AO22 U81 ( .A(InEdges[8]), .B(n82), .C(OutEdge[8]), .D(n284), .Z(n275)
         );
    VMW_AO22 U82 ( .A(InEdges[7]), .B(n82), .C(OutEdge[7]), .D(n284), .Z(n276)
         );
    VMW_AO22 U83 ( .A(InEdges[6]), .B(n82), .C(OutEdge[6]), .D(n284), .Z(n277)
         );
    VMW_AO22 U84 ( .A(InEdges[5]), .B(n82), .C(OutEdge[5]), .D(n284), .Z(n278)
         );
    VMW_AO22 U85 ( .A(InEdges[4]), .B(n82), .C(OutEdge[4]), .D(n284), .Z(n279)
         );
    VMW_AO22 U86 ( .A(InEdges[3]), .B(n82), .C(OutEdge[3]), .D(n284), .Z(n280)
         );
    VMW_AO22 U87 ( .A(InEdges[2]), .B(n82), .C(OutEdge[2]), .D(n284), .Z(n281)
         );
    VMW_AO22 U88 ( .A(InEdges[1]), .B(n82), .C(OutEdge[1]), .D(n284), .Z(n282)
         );
    VMW_AO22 U89 ( .A(InEdges[14]), .B(n82), .C(OutEdge[14]), .D(n284), .Z(
        n269) );
    VMW_AO22 U90 ( .A(InEdges[13]), .B(n82), .C(OutEdge[13]), .D(n284), .Z(
        n270) );
    VMW_AO22 U91 ( .A(InEdges[12]), .B(n82), .C(OutEdge[12]), .D(n284), .Z(
        n271) );
    VMW_AO22 U92 ( .A(InEdges[11]), .B(n82), .C(OutEdge[11]), .D(n284), .Z(
        n272) );
    VMW_AO22 U93 ( .A(InEdges[10]), .B(n82), .C(OutEdge[10]), .D(n284), .Z(
        n273) );
    VMW_AO22 U94 ( .A(InEdges[0]), .B(n82), .C(OutEdge[0]), .D(n284), .Z(n283)
         );
    VMW_BUFIZ U95 ( .A(\path[3] ), .E(n294), .Z(\PathData[3] ) );
    VMW_BUFIZ U96 ( .A(\path[1] ), .E(n294), .Z(\PathData[1] ) );
    VMW_BUFIZ U97 ( .A(\path[0] ), .E(n294), .Z(\PathData[0] ) );
    VMW_BUFIZ U98 ( .A(\path[2] ), .E(n294), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n295), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n296), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n297), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n298), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge96[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge96[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge96[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge96[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge96[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge96[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge96[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge96[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge96[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge96[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge96[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge96[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge96[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge96[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge96[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge96[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE1_SOURCE0_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges), 
        .LEQ(n299), .TC(n299), .GE_GT(n82) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n85) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n85), .D(n82), .Z(n86) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n86), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n93) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n93), .D(n90), .Z(n94) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n94), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n96), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n102), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n112) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n112), .D(n110), .Z(n113) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n114), .C(n113), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n114) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE2_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp180[1] , \temp180[8] , \OutEdge106[5] , \temp180[5] , 
        \OutEdge106[8] , \OutEdge106[1] , \path[2] , \path[0] , 
        \OutEdge106[3] , \temp180[7] , \OutEdge106[7] , \temp180[3] , 
        \OutEdge106[13] , \temp180[12] , \temp180[10] , \OutEdge106[11] , 
        \OutEdge106[15] , \temp180[14] , n84, \OutEdge106[14] , \temp180[15] , 
        \temp180[11] , \OutEdge106[10] , \OutEdge106[12] , \temp180[13] , 
        \OutEdge106[6] , \temp180[2] , \path[1] , n92, \OutEdge106[2] , 
        \temp180[6] , \temp180[4] , \OutEdge106[9] , \OutEdge106[0] , 
        \path[3] , \temp180[0] , \temp180[9] , \OutEdge106[4] , n367, n368, 
        n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
        n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
        n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U55 ( .Z(n402) );
    VMW_PULLDOWN U56 ( .Z(n403) );
    VMW_NOR2 U57 ( .A(Start), .B(n367), .Z(\OutEdge106[15] ) );
    VMW_NAND2 U58 ( .A(n368), .B(n369), .Z(\OutEdge106[14] ) );
    VMW_NAND2 U59 ( .A(n370), .B(n369), .Z(\OutEdge106[13] ) );
    VMW_NAND2 U60 ( .A(n371), .B(n369), .Z(\OutEdge106[12] ) );
    VMW_NAND2 U61 ( .A(n372), .B(n369), .Z(\OutEdge106[11] ) );
    VMW_NAND2 U62 ( .A(n373), .B(n369), .Z(\OutEdge106[10] ) );
    VMW_NAND2 U63 ( .A(n374), .B(n369), .Z(\OutEdge106[9] ) );
    VMW_NAND2 U64 ( .A(n375), .B(n369), .Z(\OutEdge106[8] ) );
    VMW_NAND2 U65 ( .A(n376), .B(n369), .Z(\OutEdge106[7] ) );
    VMW_NAND2 U66 ( .A(n377), .B(n369), .Z(\OutEdge106[6] ) );
    VMW_NAND2 U67 ( .A(n378), .B(n369), .Z(\OutEdge106[5] ) );
    VMW_NAND2 U68 ( .A(n379), .B(n369), .Z(\OutEdge106[4] ) );
    VMW_NAND2 U69 ( .A(n380), .B(n369), .Z(\OutEdge106[3] ) );
    VMW_NAND2 U70 ( .A(n381), .B(n369), .Z(\OutEdge106[2] ) );
    VMW_NAND2 U71 ( .A(n382), .B(n369), .Z(\OutEdge106[1] ) );
    VMW_NAND2 U72 ( .A(n383), .B(n369), .Z(\OutEdge106[0] ) );
    VMW_AO21 U73 ( .A(Start), .B(\path[1] ), .C(n384), .Z(n401) );
    VMW_AO21 U74 ( .A(\path[3] ), .B(Start), .C(n384), .Z(n400) );
    VMW_AO21 U75 ( .A(Start), .B(\path[2] ), .C(n384), .Z(n399) );
    VMW_OR2 U76 ( .A(n386), .B(n92), .Z(n385) );
    VMW_AO22 U77 ( .A(OutEdge[15]), .B(n386), .C(InEdges[15]), .D(n84), .Z(
        \temp180[15] ) );
    VMW_OAI22 U78 ( .A(\path[0] ), .B(n369), .C(n385), .D(Start), .Z(n387) );
    VMW_MUX2I U79 ( .A(\temp180[15] ), .B(InEdges[31]), .S(n92), .Z(n367) );
    VMW_AND4 U80 ( .A(n389), .B(n390), .C(n391), .D(n392), .Z(n388) );
    VMW_NOR3 U81 ( .A(Start), .B(n84), .C(n92), .Z(n384) );
    VMW_AND5 U82 ( .A(n393), .B(n394), .C(n395), .D(n396), .E(n388), .Z(n397)
         );
    VMW_XNOR2 U83 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n392) );
    VMW_XNOR2 U84 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n391) );
    VMW_XNOR2 U85 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n390) );
    VMW_XNOR2 U86 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n389) );
    VMW_XNOR2 U87 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n396) );
    VMW_XNOR2 U88 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n395) );
    VMW_XNOR2 U89 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n394) );
    VMW_XNOR2 U90 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n393) );
    VMW_AO22 U91 ( .A(OutEdge[9]), .B(n386), .C(InEdges[9]), .D(n84), .Z(
        \temp180[9] ) );
    VMW_AO22 U92 ( .A(OutEdge[8]), .B(n386), .C(InEdges[8]), .D(n84), .Z(
        \temp180[8] ) );
    VMW_AO22 U93 ( .A(OutEdge[7]), .B(n386), .C(InEdges[7]), .D(n84), .Z(
        \temp180[7] ) );
    VMW_AO22 U94 ( .A(OutEdge[6]), .B(n386), .C(InEdges[6]), .D(n84), .Z(
        \temp180[6] ) );
    VMW_AO22 U95 ( .A(OutEdge[5]), .B(n386), .C(InEdges[5]), .D(n84), .Z(
        \temp180[5] ) );
    VMW_AO22 U96 ( .A(OutEdge[4]), .B(n386), .C(InEdges[4]), .D(n84), .Z(
        \temp180[4] ) );
    VMW_AO22 U97 ( .A(OutEdge[3]), .B(n386), .C(InEdges[3]), .D(n84), .Z(
        \temp180[3] ) );
    VMW_AO22 U98 ( .A(OutEdge[2]), .B(n386), .C(InEdges[2]), .D(n84), .Z(
        \temp180[2] ) );
    VMW_AO22 U99 ( .A(OutEdge[1]), .B(n386), .C(InEdges[1]), .D(n84), .Z(
        \temp180[1] ) );
    VMW_AO22 U100 ( .A(OutEdge[14]), .B(n386), .C(InEdges[14]), .D(n84), .Z(
        \temp180[14] ) );
    VMW_AO22 U101 ( .A(OutEdge[13]), .B(n386), .C(InEdges[13]), .D(n84), .Z(
        \temp180[13] ) );
    VMW_AO22 U102 ( .A(OutEdge[12]), .B(n386), .C(InEdges[12]), .D(n84), .Z(
        \temp180[12] ) );
    VMW_AO22 U103 ( .A(OutEdge[11]), .B(n386), .C(InEdges[11]), .D(n84), .Z(
        \temp180[11] ) );
    VMW_AO22 U104 ( .A(OutEdge[10]), .B(n386), .C(InEdges[10]), .D(n84), .Z(
        \temp180[10] ) );
    VMW_AO22 U105 ( .A(OutEdge[0]), .B(n386), .C(InEdges[0]), .D(n84), .Z(
        \temp180[0] ) );
    VMW_MUX2I U106 ( .A(\temp180[9] ), .B(InEdges[25]), .S(n92), .Z(n374) );
    VMW_MUX2I U107 ( .A(\temp180[8] ), .B(InEdges[24]), .S(n92), .Z(n375) );
    VMW_MUX2I U108 ( .A(\temp180[7] ), .B(InEdges[23]), .S(n92), .Z(n376) );
    VMW_MUX2I U109 ( .A(\temp180[6] ), .B(InEdges[22]), .S(n92), .Z(n377) );
    VMW_MUX2I U110 ( .A(\temp180[5] ), .B(InEdges[21]), .S(n92), .Z(n378) );
    VMW_MUX2I U111 ( .A(\temp180[4] ), .B(InEdges[20]), .S(n92), .Z(n379) );
    VMW_MUX2I U112 ( .A(\temp180[3] ), .B(InEdges[19]), .S(n92), .Z(n380) );
    VMW_MUX2I U113 ( .A(\temp180[2] ), .B(InEdges[18]), .S(n92), .Z(n381) );
    VMW_MUX2I U114 ( .A(\temp180[1] ), .B(InEdges[17]), .S(n92), .Z(n382) );
    VMW_MUX2I U115 ( .A(\temp180[14] ), .B(InEdges[30]), .S(n92), .Z(n368) );
    VMW_MUX2I U116 ( .A(\temp180[13] ), .B(InEdges[29]), .S(n92), .Z(n370) );
    VMW_MUX2I U117 ( .A(\temp180[12] ), .B(InEdges[28]), .S(n92), .Z(n371) );
    VMW_MUX2I U118 ( .A(\temp180[11] ), .B(InEdges[27]), .S(n92), .Z(n372) );
    VMW_MUX2I U119 ( .A(\temp180[10] ), .B(InEdges[26]), .S(n92), .Z(n373) );
    VMW_MUX2I U120 ( .A(\temp180[0] ), .B(InEdges[16]), .S(n92), .Z(n383) );
    VMW_INV U121 ( .A(n84), .Z(n386) );
    VMW_INV U122 ( .A(Start), .Z(n369) );
    VMW_INV U123 ( .A(n387), .Z(n398) );
    VMW_BUFIZ U124 ( .A(\path[3] ), .E(n397), .Z(\PathData[3] ) );
    VMW_BUFIZ U125 ( .A(\path[1] ), .E(n397), .Z(\PathData[1] ) );
    VMW_BUFIZ U126 ( .A(\path[0] ), .E(n397), .Z(\PathData[0] ) );
    VMW_BUFIZ U127 ( .A(\path[2] ), .E(n397), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n398), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n399), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n400), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n401), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge106[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge106[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge106[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge106[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge106[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge106[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge106[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge106[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge106[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge106[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge106[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge106[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge106[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge106[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge106[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge106[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n403), .TC(n403), .GE_GT(n84) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 lte_55_1 ( .A({\temp180[15] , 
        \temp180[14] , \temp180[13] , \temp180[12] , \temp180[11] , 
        \temp180[10] , \temp180[9] , \temp180[8] , \temp180[7] , \temp180[6] , 
        \temp180[5] , \temp180[4] , \temp180[3] , \temp180[2] , \temp180[1] , 
        \temp180[0] }), .B(InEdges[31:16]), .LEQ(n402), .TC(n402), .GE_GT(n92)
         );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, 
        n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, n107, 
        n108, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n104), .B(B[12]), .Z(n103) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n96), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n104), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n103), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n104) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
        n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
        n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
        n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
        n163, n164;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n119), .B(B[2]), .Z(n118) );
    VMW_AO22 U5 ( .A(n121), .B(B[0]), .C(n122), .D(B[1]), .Z(n120) );
    VMW_OR2 U6 ( .A(B[2]), .B(n119), .Z(n123) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n122), .C(n123), .D(n120), .Z(n124) );
    VMW_NAND2 U8 ( .A(n126), .B(B[4]), .Z(n125) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n128), .C(n124), .D(n118), .Z(n127) );
    VMW_OR2 U10 ( .A(B[4]), .B(n126), .Z(n129) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n131), .C(n129), .D(n127), .Z(n130) );
    VMW_NAND2 U12 ( .A(n133), .B(B[6]), .Z(n132) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n135), .C(n130), .D(n125), .Z(n134) );
    VMW_OR2 U14 ( .A(B[6]), .B(n133), .Z(n136) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n138), .C(n136), .D(n134), .Z(n137) );
    VMW_NAND2 U16 ( .A(n140), .B(B[8]), .Z(n139) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n142), .C(n137), .D(n132), .Z(n141) );
    VMW_OR2 U18 ( .A(B[8]), .B(n140), .Z(n143) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n145), .C(n143), .D(n141), .Z(n144) );
    VMW_NAND2 U20 ( .A(n147), .B(B[10]), .Z(n146) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n149), .C(n144), .D(n139), .Z(n148) );
    VMW_NAND2 U22 ( .A(n149), .B(A[9]), .Z(n150) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n147), .C(n150), .D(n148), .Z(n151) );
    VMW_NAND2 U24 ( .A(n153), .B(B[12]), .Z(n152) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n155), .C(n151), .D(n146), .Z(n154) );
    VMW_NAND2 U26 ( .A(n155), .B(A[11]), .Z(n156) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n153), .C(n156), .D(n154), .Z(n157) );
    VMW_NAND2 U28 ( .A(n159), .B(B[14]), .Z(n158) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n161), .C(n157), .D(n152), .Z(n160) );
    VMW_NAND2 U30 ( .A(n161), .B(A[13]), .Z(n162) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n159), .C(n162), .D(n160), .Z(n163) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n164), .C(n163), .D(n158), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n153) );
    VMW_INV U34 ( .A(B[7]), .Z(n142) );
    VMW_INV U35 ( .A(A[7]), .Z(n145) );
    VMW_INV U36 ( .A(A[3]), .Z(n131) );
    VMW_INV U37 ( .A(B[3]), .Z(n128) );
    VMW_INV U38 ( .A(A[10]), .Z(n147) );
    VMW_INV U39 ( .A(B[9]), .Z(n149) );
    VMW_INV U40 ( .A(A[4]), .Z(n126) );
    VMW_INV U41 ( .A(A[8]), .Z(n140) );
    VMW_INV U42 ( .A(A[14]), .Z(n159) );
    VMW_INV U43 ( .A(B[11]), .Z(n155) );
    VMW_INV U44 ( .A(A[5]), .Z(n138) );
    VMW_INV U45 ( .A(B[5]), .Z(n135) );
    VMW_INV U46 ( .A(A[1]), .Z(n122) );
    VMW_INV U47 ( .A(B[15]), .Z(n164) );
    VMW_INV U48 ( .A(B[13]), .Z(n161) );
    VMW_INV U49 ( .A(A[6]), .Z(n133) );
    VMW_INV U50 ( .A(A[2]), .Z(n119) );
    VMW_INV U51 ( .A(A[0]), .Z(n121) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE3_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp284[0] , \OutEdge116[6] , \temp284[9] , \temp284[11] , 
        \temp190[2] , \OutEdge116[2] , \temp284[4] , \temp190[6] , 
        \temp284[15] , \path[2] , \OutEdge116[9] , \path[0] , \temp190[4] , 
        \OutEdge116[0] , \temp284[6] , \temp284[13] , \temp190[0] , 
        \temp284[2] , \OutEdge116[4] , \temp190[9] , \temp190[10] , 
        \OutEdge116[11] , \OutEdge116[15] , \temp190[14] , \OutEdge116[13] , 
        \temp190[12] , n94, \OutEdge116[12] , \temp190[13] , n86, 
        \OutEdge116[14] , \temp190[15] , \temp190[11] , \OutEdge116[10] , 
        \temp284[12] , \temp190[1] , \temp284[3] , \OutEdge116[5] , 
        \temp190[8] , \path[1] , \OutEdge116[8] , \temp190[5] , 
        \OutEdge116[1] , \temp284[7] , n102, \OutEdge116[3] , \temp284[5] , 
        \temp190[7] , \temp284[14] , \path[3] , \temp284[1] , \OutEdge116[7] , 
        \temp284[8] , \temp284[10] , \temp190[3] , n467, n468, n469, n470, 
        n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
        n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
        n507, n508;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U64 ( .Z(n506) );
    VMW_PULLDOWN U65 ( .Z(n508) );
    VMW_PULLDOWN U66 ( .Z(n507) );
    VMW_NOR2 U67 ( .A(Start), .B(n467), .Z(\OutEdge116[15] ) );
    VMW_NAND2 U68 ( .A(n468), .B(n469), .Z(\OutEdge116[14] ) );
    VMW_NAND2 U69 ( .A(n470), .B(n469), .Z(\OutEdge116[13] ) );
    VMW_NAND2 U70 ( .A(n471), .B(n469), .Z(\OutEdge116[12] ) );
    VMW_NAND2 U71 ( .A(n472), .B(n469), .Z(\OutEdge116[11] ) );
    VMW_NAND2 U72 ( .A(n473), .B(n469), .Z(\OutEdge116[10] ) );
    VMW_NAND2 U73 ( .A(n474), .B(n469), .Z(\OutEdge116[9] ) );
    VMW_NAND2 U74 ( .A(n475), .B(n469), .Z(\OutEdge116[8] ) );
    VMW_NAND2 U75 ( .A(n476), .B(n469), .Z(\OutEdge116[7] ) );
    VMW_NAND2 U76 ( .A(n477), .B(n469), .Z(\OutEdge116[6] ) );
    VMW_NAND2 U77 ( .A(n478), .B(n469), .Z(\OutEdge116[5] ) );
    VMW_NAND2 U78 ( .A(n479), .B(n469), .Z(\OutEdge116[4] ) );
    VMW_NAND2 U79 ( .A(n480), .B(n469), .Z(\OutEdge116[3] ) );
    VMW_NAND2 U80 ( .A(n481), .B(n469), .Z(\OutEdge116[2] ) );
    VMW_NAND2 U81 ( .A(n482), .B(n469), .Z(\OutEdge116[1] ) );
    VMW_NAND2 U82 ( .A(n483), .B(n469), .Z(\OutEdge116[0] ) );
    VMW_OR2 U83 ( .A(n484), .B(n485), .Z(n505) );
    VMW_AO21 U84 ( .A(\path[3] ), .B(Start), .C(n486), .Z(n504) );
    VMW_AO21 U85 ( .A(Start), .B(\path[2] ), .C(n486), .Z(n503) );
    VMW_AO22 U86 ( .A(InEdges[31]), .B(n94), .C(\temp190[15] ), .D(n487), .Z(
        \temp284[15] ) );
    VMW_INV U87 ( .A(Start), .Z(n469) );
    VMW_AND3 U88 ( .A(n469), .B(n488), .C(n487), .Z(n485) );
    VMW_OAI22 U89 ( .A(\path[0] ), .B(n469), .C(n490), .D(Start), .Z(n489) );
    VMW_MUX2I U90 ( .A(\temp284[15] ), .B(InEdges[47]), .S(n102), .Z(n467) );
    VMW_AND4 U91 ( .A(n492), .B(n493), .C(n494), .D(n495), .Z(n491) );
    VMW_NOR2 U92 ( .A(n102), .B(n496), .Z(n486) );
    VMW_AND5 U93 ( .A(n497), .B(n498), .C(n499), .D(n500), .E(n491), .Z(n501)
         );
    VMW_XNOR2 U94 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n495) );
    VMW_XNOR2 U95 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n494) );
    VMW_XNOR2 U96 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n493) );
    VMW_XNOR2 U97 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n492) );
    VMW_XNOR2 U98 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n500) );
    VMW_XNOR2 U99 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n499) );
    VMW_XNOR2 U100 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n498) );
    VMW_XNOR2 U101 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n497) );
    VMW_AO22 U102 ( .A(OutEdge[9]), .B(n488), .C(InEdges[9]), .D(n86), .Z(
        \temp190[9] ) );
    VMW_AO22 U103 ( .A(InEdges[25]), .B(n94), .C(\temp190[9] ), .D(n487), .Z(
        \temp284[9] ) );
    VMW_AO22 U104 ( .A(OutEdge[8]), .B(n488), .C(InEdges[8]), .D(n86), .Z(
        \temp190[8] ) );
    VMW_AO22 U105 ( .A(InEdges[24]), .B(n94), .C(\temp190[8] ), .D(n487), .Z(
        \temp284[8] ) );
    VMW_AO22 U106 ( .A(OutEdge[7]), .B(n488), .C(InEdges[7]), .D(n86), .Z(
        \temp190[7] ) );
    VMW_AO22 U107 ( .A(InEdges[23]), .B(n94), .C(\temp190[7] ), .D(n487), .Z(
        \temp284[7] ) );
    VMW_AO22 U108 ( .A(OutEdge[6]), .B(n488), .C(InEdges[6]), .D(n86), .Z(
        \temp190[6] ) );
    VMW_AO22 U109 ( .A(InEdges[22]), .B(n94), .C(\temp190[6] ), .D(n487), .Z(
        \temp284[6] ) );
    VMW_AO22 U110 ( .A(OutEdge[5]), .B(n488), .C(InEdges[5]), .D(n86), .Z(
        \temp190[5] ) );
    VMW_AO22 U111 ( .A(InEdges[21]), .B(n94), .C(\temp190[5] ), .D(n487), .Z(
        \temp284[5] ) );
    VMW_AO22 U112 ( .A(OutEdge[4]), .B(n488), .C(InEdges[4]), .D(n86), .Z(
        \temp190[4] ) );
    VMW_AO22 U113 ( .A(InEdges[20]), .B(n94), .C(\temp190[4] ), .D(n487), .Z(
        \temp284[4] ) );
    VMW_AO22 U114 ( .A(OutEdge[3]), .B(n488), .C(InEdges[3]), .D(n86), .Z(
        \temp190[3] ) );
    VMW_AO22 U115 ( .A(InEdges[19]), .B(n94), .C(\temp190[3] ), .D(n487), .Z(
        \temp284[3] ) );
    VMW_AO22 U116 ( .A(OutEdge[2]), .B(n488), .C(InEdges[2]), .D(n86), .Z(
        \temp190[2] ) );
    VMW_AO22 U117 ( .A(InEdges[18]), .B(n94), .C(\temp190[2] ), .D(n487), .Z(
        \temp284[2] ) );
    VMW_AO22 U118 ( .A(OutEdge[1]), .B(n488), .C(InEdges[1]), .D(n86), .Z(
        \temp190[1] ) );
    VMW_AO22 U119 ( .A(InEdges[17]), .B(n94), .C(\temp190[1] ), .D(n487), .Z(
        \temp284[1] ) );
    VMW_AO22 U120 ( .A(OutEdge[15]), .B(n488), .C(InEdges[15]), .D(n86), .Z(
        \temp190[15] ) );
    VMW_AO22 U121 ( .A(OutEdge[14]), .B(n488), .C(InEdges[14]), .D(n86), .Z(
        \temp190[14] ) );
    VMW_AO22 U122 ( .A(InEdges[30]), .B(n94), .C(\temp190[14] ), .D(n487), .Z(
        \temp284[14] ) );
    VMW_AO22 U123 ( .A(OutEdge[13]), .B(n488), .C(InEdges[13]), .D(n86), .Z(
        \temp190[13] ) );
    VMW_AO22 U124 ( .A(InEdges[29]), .B(n94), .C(\temp190[13] ), .D(n487), .Z(
        \temp284[13] ) );
    VMW_AO22 U125 ( .A(OutEdge[12]), .B(n488), .C(InEdges[12]), .D(n86), .Z(
        \temp190[12] ) );
    VMW_AO22 U126 ( .A(InEdges[28]), .B(n94), .C(\temp190[12] ), .D(n487), .Z(
        \temp284[12] ) );
    VMW_AO22 U127 ( .A(OutEdge[11]), .B(n488), .C(InEdges[11]), .D(n86), .Z(
        \temp190[11] ) );
    VMW_AO22 U128 ( .A(InEdges[27]), .B(n94), .C(\temp190[11] ), .D(n487), .Z(
        \temp284[11] ) );
    VMW_AO22 U129 ( .A(OutEdge[10]), .B(n488), .C(InEdges[10]), .D(n86), .Z(
        \temp190[10] ) );
    VMW_AO22 U130 ( .A(InEdges[26]), .B(n94), .C(\temp190[10] ), .D(n487), .Z(
        \temp284[10] ) );
    VMW_AO22 U131 ( .A(OutEdge[0]), .B(n488), .C(InEdges[0]), .D(n86), .Z(
        \temp190[0] ) );
    VMW_AO22 U132 ( .A(InEdges[16]), .B(n94), .C(\temp190[0] ), .D(n487), .Z(
        \temp284[0] ) );
    VMW_AO22 U133 ( .A(\path[1] ), .B(Start), .C(n102), .D(n469), .Z(n484) );
    VMW_AOI21 U134 ( .A(n487), .B(n86), .C(n102), .Z(n490) );
    VMW_MUX2I U135 ( .A(\temp284[9] ), .B(InEdges[41]), .S(n102), .Z(n474) );
    VMW_MUX2I U136 ( .A(\temp284[8] ), .B(InEdges[40]), .S(n102), .Z(n475) );
    VMW_MUX2I U137 ( .A(\temp284[7] ), .B(InEdges[39]), .S(n102), .Z(n476) );
    VMW_MUX2I U138 ( .A(\temp284[6] ), .B(InEdges[38]), .S(n102), .Z(n477) );
    VMW_MUX2I U139 ( .A(\temp284[5] ), .B(InEdges[37]), .S(n102), .Z(n478) );
    VMW_MUX2I U140 ( .A(\temp284[4] ), .B(InEdges[36]), .S(n102), .Z(n479) );
    VMW_MUX2I U141 ( .A(\temp284[3] ), .B(InEdges[35]), .S(n102), .Z(n480) );
    VMW_MUX2I U142 ( .A(\temp284[2] ), .B(InEdges[34]), .S(n102), .Z(n481) );
    VMW_MUX2I U143 ( .A(\temp284[1] ), .B(InEdges[33]), .S(n102), .Z(n482) );
    VMW_MUX2I U144 ( .A(\temp284[14] ), .B(InEdges[46]), .S(n102), .Z(n468) );
    VMW_MUX2I U145 ( .A(\temp284[13] ), .B(InEdges[45]), .S(n102), .Z(n470) );
    VMW_MUX2I U146 ( .A(\temp284[12] ), .B(InEdges[44]), .S(n102), .Z(n471) );
    VMW_MUX2I U147 ( .A(\temp284[11] ), .B(InEdges[43]), .S(n102), .Z(n472) );
    VMW_MUX2I U148 ( .A(\temp284[10] ), .B(InEdges[42]), .S(n102), .Z(n473) );
    VMW_MUX2I U149 ( .A(\temp284[0] ), .B(InEdges[32]), .S(n102), .Z(n483) );
    VMW_INV U150 ( .A(n94), .Z(n487) );
    VMW_INV U151 ( .A(n86), .Z(n488) );
    VMW_INV U152 ( .A(n485), .Z(n496) );
    VMW_INV U153 ( .A(n489), .Z(n502) );
    VMW_BUFIZ U154 ( .A(\path[3] ), .E(n501), .Z(\PathData[3] ) );
    VMW_BUFIZ U155 ( .A(\path[1] ), .E(n501), .Z(\PathData[1] ) );
    VMW_BUFIZ U156 ( .A(\path[0] ), .E(n501), .Z(\PathData[0] ) );
    VMW_BUFIZ U157 ( .A(\path[2] ), .E(n501), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n502), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n503), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n504), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n505), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge116[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge116[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge116[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge116[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge116[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge116[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge116[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge116[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge116[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge116[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge116[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge116[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge116[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge116[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge116[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge116[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp190[15] , 
        \temp190[14] , \temp190[13] , \temp190[12] , \temp190[11] , 
        \temp190[10] , \temp190[9] , \temp190[8] , \temp190[7] , \temp190[6] , 
        \temp190[5] , \temp190[4] , \temp190[3] , \temp190[2] , \temp190[1] , 
        \temp190[0] }), .B(InEdges[31:16]), .LEQ(n508), .TC(n508), .GE_GT(n94)
         );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n507), .TC(n507), .GE_GT(n86) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 lte_55_2 ( .A({\temp284[15] , 
        \temp284[14] , \temp284[13] , \temp284[12] , \temp284[11] , 
        \temp284[10] , \temp284[9] , \temp284[8] , \temp284[7] , \temp284[6] , 
        \temp284[5] , \temp284[4] , \temp284[3] , \temp284[2] , \temp284[1] , 
        \temp284[0] }), .B(InEdges[47:32]), .LEQ(n506), .TC(n506), .GE_GT(n102
        ) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, 
        n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, 
        n108, n109, n110, n111, n113, n114, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n95), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n113), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n113), .B(A[13]), .Z(n114) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n114), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n113) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
        n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
        n164, n165;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n127), .B(B[4]), .Z(n126) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n129), .C(n125), .D(n119), .Z(n128) );
    VMW_OR2 U10 ( .A(B[4]), .B(n127), .Z(n130) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n132), .C(n130), .D(n128), .Z(n131) );
    VMW_NAND2 U12 ( .A(n134), .B(B[6]), .Z(n133) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n136), .C(n131), .D(n126), .Z(n135) );
    VMW_OR2 U14 ( .A(B[6]), .B(n134), .Z(n137) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n139), .C(n137), .D(n135), .Z(n138) );
    VMW_NAND2 U16 ( .A(n141), .B(B[8]), .Z(n140) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n143), .C(n138), .D(n133), .Z(n142) );
    VMW_OR2 U18 ( .A(B[8]), .B(n141), .Z(n144) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n146), .C(n144), .D(n142), .Z(n145) );
    VMW_NAND2 U20 ( .A(n148), .B(B[10]), .Z(n147) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n150), .C(n145), .D(n140), .Z(n149) );
    VMW_NAND2 U22 ( .A(n150), .B(A[9]), .Z(n151) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n148), .C(n151), .D(n149), .Z(n152) );
    VMW_NAND2 U24 ( .A(n154), .B(B[12]), .Z(n153) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n156), .C(n152), .D(n147), .Z(n155) );
    VMW_NAND2 U26 ( .A(n156), .B(A[11]), .Z(n157) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n154), .C(n157), .D(n155), .Z(n158) );
    VMW_NAND2 U28 ( .A(n160), .B(B[14]), .Z(n159) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n162), .C(n158), .D(n153), .Z(n161) );
    VMW_NAND2 U30 ( .A(n162), .B(A[13]), .Z(n163) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n160), .C(n163), .D(n161), .Z(n164) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n165), .C(n164), .D(n159), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n154) );
    VMW_INV U34 ( .A(B[7]), .Z(n143) );
    VMW_INV U35 ( .A(A[7]), .Z(n146) );
    VMW_INV U36 ( .A(A[3]), .Z(n132) );
    VMW_INV U37 ( .A(B[3]), .Z(n129) );
    VMW_INV U38 ( .A(A[10]), .Z(n148) );
    VMW_INV U39 ( .A(B[9]), .Z(n150) );
    VMW_INV U40 ( .A(A[4]), .Z(n127) );
    VMW_INV U41 ( .A(A[8]), .Z(n141) );
    VMW_INV U42 ( .A(A[14]), .Z(n160) );
    VMW_INV U43 ( .A(B[11]), .Z(n156) );
    VMW_INV U44 ( .A(A[5]), .Z(n139) );
    VMW_INV U45 ( .A(B[5]), .Z(n136) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n165) );
    VMW_INV U48 ( .A(B[13]), .Z(n162) );
    VMW_INV U49 ( .A(A[6]), .Z(n134) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
        n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
        n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
        n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
        n213, n214;
    VMW_OAI21 U3 ( .A(B[15]), .B(n166), .C(n167), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n169), .B(B[2]), .Z(n168) );
    VMW_AO22 U5 ( .A(n171), .B(B[0]), .C(n172), .D(B[1]), .Z(n170) );
    VMW_OR2 U6 ( .A(B[2]), .B(n169), .Z(n173) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n172), .C(n173), .D(n170), .Z(n174) );
    VMW_NAND2 U8 ( .A(n176), .B(B[4]), .Z(n175) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n178), .C(n174), .D(n168), .Z(n177) );
    VMW_OR2 U10 ( .A(B[4]), .B(n176), .Z(n179) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n181), .C(n179), .D(n177), .Z(n180) );
    VMW_NAND2 U12 ( .A(n183), .B(B[6]), .Z(n182) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n185), .C(n180), .D(n175), .Z(n184) );
    VMW_OR2 U14 ( .A(B[6]), .B(n183), .Z(n186) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n188), .C(n186), .D(n184), .Z(n187) );
    VMW_NAND2 U16 ( .A(n190), .B(B[8]), .Z(n189) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n192), .C(n187), .D(n182), .Z(n191) );
    VMW_OR2 U18 ( .A(B[8]), .B(n190), .Z(n193) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n195), .C(n193), .D(n191), .Z(n194) );
    VMW_NAND2 U20 ( .A(n197), .B(B[10]), .Z(n196) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n199), .C(n194), .D(n189), .Z(n198) );
    VMW_NAND2 U22 ( .A(n199), .B(A[9]), .Z(n200) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n197), .C(n200), .D(n198), .Z(n201) );
    VMW_NAND2 U24 ( .A(n203), .B(B[12]), .Z(n202) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n205), .C(n201), .D(n196), .Z(n204) );
    VMW_NAND2 U26 ( .A(n205), .B(A[11]), .Z(n206) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n203), .C(n206), .D(n204), .Z(n207) );
    VMW_NAND2 U28 ( .A(n209), .B(B[14]), .Z(n208) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n211), .C(n207), .D(n202), .Z(n210) );
    VMW_NAND2 U30 ( .A(n211), .B(A[13]), .Z(n212) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n209), .C(n212), .D(n210), .Z(n213) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n214), .C(n213), .D(n208), .Z(n167) );
    VMW_INV U33 ( .A(A[12]), .Z(n203) );
    VMW_INV U34 ( .A(B[7]), .Z(n192) );
    VMW_INV U35 ( .A(A[7]), .Z(n195) );
    VMW_INV U36 ( .A(A[3]), .Z(n181) );
    VMW_INV U37 ( .A(B[3]), .Z(n178) );
    VMW_INV U38 ( .A(A[10]), .Z(n197) );
    VMW_INV U39 ( .A(B[9]), .Z(n199) );
    VMW_INV U40 ( .A(A[4]), .Z(n176) );
    VMW_INV U41 ( .A(A[8]), .Z(n190) );
    VMW_INV U42 ( .A(A[14]), .Z(n209) );
    VMW_INV U43 ( .A(B[11]), .Z(n205) );
    VMW_INV U44 ( .A(A[5]), .Z(n188) );
    VMW_INV U45 ( .A(B[5]), .Z(n185) );
    VMW_INV U46 ( .A(A[1]), .Z(n172) );
    VMW_INV U47 ( .A(B[15]), .Z(n214) );
    VMW_INV U48 ( .A(B[13]), .Z(n211) );
    VMW_INV U49 ( .A(A[6]), .Z(n183) );
    VMW_INV U50 ( .A(A[2]), .Z(n169) );
    VMW_INV U51 ( .A(A[0]), .Z(n171) );
    VMW_INV U52 ( .A(A[15]), .Z(n166) );
endmodule


module NodeAux_INDEGREE4_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp200[0] , \temp384[15] , \OutEdge126[12] , \temp200[15] , 
        \temp200[9] , \temp384[6] , \temp294[3] , n112, \temp294[13] , 
        \temp384[11] , \temp200[4] , \temp294[7] , \temp384[2] , \path[2] , 
        \temp200[11] , \temp200[13] , \path[0] , \temp294[5] , \temp384[0] , 
        \temp384[13] , \temp200[6] , \temp384[9] , \OutEdge126[14] , 
        \temp294[11] , \temp384[4] , \temp294[1] , \OutEdge126[10] , 
        \temp294[15] , \temp200[2] , \temp294[8] , \OutEdge126[8] , 
        \OutEdge126[1] , \OutEdge126[5] , n96, \OutEdge126[7] , 
        \OutEdge126[3] , \OutEdge126[2] , \OutEdge126[6] , \OutEdge126[4] , 
        n104, \OutEdge126[9] , n88, \OutEdge126[0] , \temp384[5] , 
        \temp294[0] , \OutEdge126[11] , \temp294[14] , \temp200[3] , 
        \temp294[9] , \path[1] , \temp200[12] , \temp294[4] , \temp384[1] , 
        \temp384[12] , \temp384[8] , \temp200[7] , \OutEdge126[15] , 
        \temp294[10] , \temp294[12] , \temp384[10] , \temp200[5] , 
        \temp294[6] , \temp384[3] , \path[3] , \temp200[10] , \temp200[1] , 
        \temp384[14] , \OutEdge126[13] , \temp200[14] , \temp384[7] , 
        \temp200[8] , \temp294[2] , n567, n568, n569, n570, n571, n572, n573, 
        n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
        n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, 
        n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
        n610, n611;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U73 ( .Z(n608) );
    VMW_PULLDOWN U74 ( .Z(n609) );
    VMW_PULLDOWN U75 ( .Z(n610) );
    VMW_PULLDOWN U76 ( .Z(n611) );
    VMW_NOR2 U77 ( .A(Start), .B(n567), .Z(\OutEdge126[15] ) );
    VMW_NAND2 U78 ( .A(n568), .B(n569), .Z(\OutEdge126[14] ) );
    VMW_NAND2 U79 ( .A(n570), .B(n569), .Z(\OutEdge126[13] ) );
    VMW_NAND2 U80 ( .A(n571), .B(n569), .Z(\OutEdge126[12] ) );
    VMW_NAND2 U81 ( .A(n572), .B(n569), .Z(\OutEdge126[11] ) );
    VMW_NAND2 U82 ( .A(n573), .B(n569), .Z(\OutEdge126[10] ) );
    VMW_NAND2 U83 ( .A(n574), .B(n569), .Z(\OutEdge126[9] ) );
    VMW_NAND2 U84 ( .A(n575), .B(n569), .Z(\OutEdge126[8] ) );
    VMW_NAND2 U85 ( .A(n576), .B(n569), .Z(\OutEdge126[7] ) );
    VMW_NAND2 U86 ( .A(n577), .B(n569), .Z(\OutEdge126[6] ) );
    VMW_NAND2 U87 ( .A(n578), .B(n569), .Z(\OutEdge126[5] ) );
    VMW_NAND2 U88 ( .A(n579), .B(n569), .Z(\OutEdge126[4] ) );
    VMW_NAND2 U89 ( .A(n580), .B(n569), .Z(\OutEdge126[3] ) );
    VMW_NAND2 U90 ( .A(n581), .B(n569), .Z(\OutEdge126[2] ) );
    VMW_NAND2 U91 ( .A(n582), .B(n569), .Z(\OutEdge126[1] ) );
    VMW_NAND2 U92 ( .A(n583), .B(n569), .Z(\OutEdge126[0] ) );
    VMW_AO21 U93 ( .A(Start), .B(\path[3] ), .C(n584), .Z(n606) );
    VMW_AO21 U94 ( .A(\path[2] ), .B(Start), .C(n584), .Z(n605) );
    VMW_OAI211 U95 ( .A(n96), .B(n88), .C(n586), .D(n587), .Z(n585) );
    VMW_NAND2 U96 ( .A(n586), .B(n589), .Z(n588) );
    VMW_AO22 U97 ( .A(\temp294[15] ), .B(n587), .C(InEdges[47]), .D(n104), .Z(
        \temp384[15] ) );
    VMW_INV U98 ( .A(n88), .Z(n590) );
    VMW_INV U99 ( .A(Start), .Z(n569) );
    VMW_OAI22 U100 ( .A(n585), .B(Start), .C(\path[1] ), .D(n569), .Z(n591) );
    VMW_OAI22 U101 ( .A(n588), .B(Start), .C(\path[0] ), .D(n569), .Z(n592) );
    VMW_MUX2I U102 ( .A(\temp384[15] ), .B(InEdges[63]), .S(n112), .Z(n567) );
    VMW_AND4 U103 ( .A(n594), .B(n595), .C(n596), .D(n597), .Z(n593) );
    VMW_INV U104 ( .A(n96), .Z(n598) );
    VMW_AND5 U105 ( .A(n590), .B(n569), .C(n586), .D(n587), .E(n598), .Z(n584)
         );
    VMW_OAI21 U106 ( .A(n96), .B(n590), .C(n587), .Z(n589) );
    VMW_AND5 U107 ( .A(n599), .B(n600), .C(n601), .D(n602), .E(n593), .Z(n603)
         );
    VMW_XNOR2 U108 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n597) );
    VMW_XNOR2 U109 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n596) );
    VMW_XNOR2 U110 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n595) );
    VMW_XNOR2 U111 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n594) );
    VMW_XNOR2 U112 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n602) );
    VMW_XNOR2 U113 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n601) );
    VMW_XNOR2 U114 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n600) );
    VMW_XNOR2 U115 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n599) );
    VMW_AO22 U116 ( .A(InEdges[9]), .B(n88), .C(OutEdge[9]), .D(n590), .Z(
        \temp200[9] ) );
    VMW_AO22 U117 ( .A(InEdges[25]), .B(n96), .C(\temp200[9] ), .D(n598), .Z(
        \temp294[9] ) );
    VMW_AO22 U118 ( .A(\temp294[9] ), .B(n587), .C(InEdges[41]), .D(n104), .Z(
        \temp384[9] ) );
    VMW_AO22 U119 ( .A(InEdges[8]), .B(n88), .C(OutEdge[8]), .D(n590), .Z(
        \temp200[8] ) );
    VMW_AO22 U120 ( .A(InEdges[24]), .B(n96), .C(\temp200[8] ), .D(n598), .Z(
        \temp294[8] ) );
    VMW_AO22 U121 ( .A(\temp294[8] ), .B(n587), .C(InEdges[40]), .D(n104), .Z(
        \temp384[8] ) );
    VMW_AO22 U122 ( .A(InEdges[7]), .B(n88), .C(OutEdge[7]), .D(n590), .Z(
        \temp200[7] ) );
    VMW_AO22 U123 ( .A(InEdges[23]), .B(n96), .C(\temp200[7] ), .D(n598), .Z(
        \temp294[7] ) );
    VMW_AO22 U124 ( .A(\temp294[7] ), .B(n587), .C(InEdges[39]), .D(n104), .Z(
        \temp384[7] ) );
    VMW_AO22 U125 ( .A(InEdges[6]), .B(n88), .C(OutEdge[6]), .D(n590), .Z(
        \temp200[6] ) );
    VMW_AO22 U126 ( .A(InEdges[22]), .B(n96), .C(\temp200[6] ), .D(n598), .Z(
        \temp294[6] ) );
    VMW_AO22 U127 ( .A(\temp294[6] ), .B(n587), .C(InEdges[38]), .D(n104), .Z(
        \temp384[6] ) );
    VMW_AO22 U128 ( .A(InEdges[5]), .B(n88), .C(OutEdge[5]), .D(n590), .Z(
        \temp200[5] ) );
    VMW_AO22 U129 ( .A(InEdges[21]), .B(n96), .C(\temp200[5] ), .D(n598), .Z(
        \temp294[5] ) );
    VMW_AO22 U130 ( .A(\temp294[5] ), .B(n587), .C(InEdges[37]), .D(n104), .Z(
        \temp384[5] ) );
    VMW_AO22 U131 ( .A(InEdges[4]), .B(n88), .C(OutEdge[4]), .D(n590), .Z(
        \temp200[4] ) );
    VMW_AO22 U132 ( .A(InEdges[20]), .B(n96), .C(\temp200[4] ), .D(n598), .Z(
        \temp294[4] ) );
    VMW_AO22 U133 ( .A(\temp294[4] ), .B(n587), .C(InEdges[36]), .D(n104), .Z(
        \temp384[4] ) );
    VMW_AO22 U134 ( .A(InEdges[3]), .B(n88), .C(OutEdge[3]), .D(n590), .Z(
        \temp200[3] ) );
    VMW_AO22 U135 ( .A(InEdges[19]), .B(n96), .C(\temp200[3] ), .D(n598), .Z(
        \temp294[3] ) );
    VMW_AO22 U136 ( .A(\temp294[3] ), .B(n587), .C(InEdges[35]), .D(n104), .Z(
        \temp384[3] ) );
    VMW_AO22 U137 ( .A(InEdges[2]), .B(n88), .C(OutEdge[2]), .D(n590), .Z(
        \temp200[2] ) );
    VMW_AO22 U138 ( .A(InEdges[18]), .B(n96), .C(\temp200[2] ), .D(n598), .Z(
        \temp294[2] ) );
    VMW_AO22 U139 ( .A(\temp294[2] ), .B(n587), .C(InEdges[34]), .D(n104), .Z(
        \temp384[2] ) );
    VMW_AO22 U140 ( .A(InEdges[1]), .B(n88), .C(OutEdge[1]), .D(n590), .Z(
        \temp200[1] ) );
    VMW_AO22 U141 ( .A(InEdges[17]), .B(n96), .C(\temp200[1] ), .D(n598), .Z(
        \temp294[1] ) );
    VMW_AO22 U142 ( .A(\temp294[1] ), .B(n587), .C(InEdges[33]), .D(n104), .Z(
        \temp384[1] ) );
    VMW_AO22 U143 ( .A(InEdges[15]), .B(n88), .C(OutEdge[15]), .D(n590), .Z(
        \temp200[15] ) );
    VMW_AO22 U144 ( .A(InEdges[31]), .B(n96), .C(\temp200[15] ), .D(n598), .Z(
        \temp294[15] ) );
    VMW_AO22 U145 ( .A(InEdges[14]), .B(n88), .C(OutEdge[14]), .D(n590), .Z(
        \temp200[14] ) );
    VMW_AO22 U146 ( .A(InEdges[30]), .B(n96), .C(\temp200[14] ), .D(n598), .Z(
        \temp294[14] ) );
    VMW_AO22 U147 ( .A(\temp294[14] ), .B(n587), .C(InEdges[46]), .D(n104), 
        .Z(\temp384[14] ) );
    VMW_AO22 U148 ( .A(InEdges[13]), .B(n88), .C(OutEdge[13]), .D(n590), .Z(
        \temp200[13] ) );
    VMW_AO22 U149 ( .A(InEdges[29]), .B(n96), .C(\temp200[13] ), .D(n598), .Z(
        \temp294[13] ) );
    VMW_AO22 U150 ( .A(\temp294[13] ), .B(n587), .C(InEdges[45]), .D(n104), 
        .Z(\temp384[13] ) );
    VMW_AO22 U151 ( .A(InEdges[12]), .B(n88), .C(OutEdge[12]), .D(n590), .Z(
        \temp200[12] ) );
    VMW_AO22 U152 ( .A(InEdges[28]), .B(n96), .C(\temp200[12] ), .D(n598), .Z(
        \temp294[12] ) );
    VMW_AO22 U153 ( .A(\temp294[12] ), .B(n587), .C(InEdges[44]), .D(n104), 
        .Z(\temp384[12] ) );
    VMW_AO22 U154 ( .A(InEdges[11]), .B(n88), .C(OutEdge[11]), .D(n590), .Z(
        \temp200[11] ) );
    VMW_AO22 U155 ( .A(InEdges[27]), .B(n96), .C(\temp200[11] ), .D(n598), .Z(
        \temp294[11] ) );
    VMW_AO22 U156 ( .A(\temp294[11] ), .B(n587), .C(InEdges[43]), .D(n104), 
        .Z(\temp384[11] ) );
    VMW_AO22 U157 ( .A(InEdges[10]), .B(n88), .C(OutEdge[10]), .D(n590), .Z(
        \temp200[10] ) );
    VMW_AO22 U158 ( .A(InEdges[26]), .B(n96), .C(\temp200[10] ), .D(n598), .Z(
        \temp294[10] ) );
    VMW_AO22 U159 ( .A(\temp294[10] ), .B(n587), .C(InEdges[42]), .D(n104), 
        .Z(\temp384[10] ) );
    VMW_AO22 U160 ( .A(InEdges[0]), .B(n88), .C(OutEdge[0]), .D(n590), .Z(
        \temp200[0] ) );
    VMW_AO22 U161 ( .A(InEdges[16]), .B(n96), .C(\temp200[0] ), .D(n598), .Z(
        \temp294[0] ) );
    VMW_AO22 U162 ( .A(\temp294[0] ), .B(n587), .C(InEdges[32]), .D(n104), .Z(
        \temp384[0] ) );
    VMW_MUX2I U163 ( .A(\temp384[9] ), .B(InEdges[57]), .S(n112), .Z(n574) );
    VMW_MUX2I U164 ( .A(\temp384[8] ), .B(InEdges[56]), .S(n112), .Z(n575) );
    VMW_MUX2I U165 ( .A(\temp384[7] ), .B(InEdges[55]), .S(n112), .Z(n576) );
    VMW_MUX2I U166 ( .A(\temp384[6] ), .B(InEdges[54]), .S(n112), .Z(n577) );
    VMW_MUX2I U167 ( .A(\temp384[5] ), .B(InEdges[53]), .S(n112), .Z(n578) );
    VMW_MUX2I U168 ( .A(\temp384[4] ), .B(InEdges[52]), .S(n112), .Z(n579) );
    VMW_MUX2I U169 ( .A(\temp384[3] ), .B(InEdges[51]), .S(n112), .Z(n580) );
    VMW_MUX2I U170 ( .A(\temp384[2] ), .B(InEdges[50]), .S(n112), .Z(n581) );
    VMW_MUX2I U171 ( .A(\temp384[1] ), .B(InEdges[49]), .S(n112), .Z(n582) );
    VMW_MUX2I U172 ( .A(\temp384[14] ), .B(InEdges[62]), .S(n112), .Z(n568) );
    VMW_MUX2I U173 ( .A(\temp384[13] ), .B(InEdges[61]), .S(n112), .Z(n570) );
    VMW_MUX2I U174 ( .A(\temp384[12] ), .B(InEdges[60]), .S(n112), .Z(n571) );
    VMW_MUX2I U175 ( .A(\temp384[11] ), .B(InEdges[59]), .S(n112), .Z(n572) );
    VMW_MUX2I U176 ( .A(\temp384[10] ), .B(InEdges[58]), .S(n112), .Z(n573) );
    VMW_MUX2I U177 ( .A(\temp384[0] ), .B(InEdges[48]), .S(n112), .Z(n583) );
    VMW_INV U178 ( .A(n104), .Z(n587) );
    VMW_INV U179 ( .A(n112), .Z(n586) );
    VMW_INV U180 ( .A(n591), .Z(n607) );
    VMW_INV U181 ( .A(n592), .Z(n604) );
    VMW_BUFIZ U182 ( .A(\path[3] ), .E(n603), .Z(\PathData[3] ) );
    VMW_BUFIZ U183 ( .A(\path[1] ), .E(n603), .Z(\PathData[1] ) );
    VMW_BUFIZ U184 ( .A(\path[0] ), .E(n603), .Z(\PathData[0] ) );
    VMW_BUFIZ U185 ( .A(\path[2] ), .E(n603), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n604), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n605), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n606), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n607), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge126[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge126[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge126[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge126[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge126[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge126[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge126[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge126[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge126[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge126[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge126[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge126[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge126[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge126[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge126[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge126[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n611), .TC(n611), .GE_GT(n88) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp200[15] , 
        \temp200[14] , \temp200[13] , \temp200[12] , \temp200[11] , 
        \temp200[10] , \temp200[9] , \temp200[8] , \temp200[7] , \temp200[6] , 
        \temp200[5] , \temp200[4] , \temp200[3] , \temp200[2] , \temp200[1] , 
        \temp200[0] }), .B(InEdges[31:16]), .LEQ(n610), .TC(n610), .GE_GT(n96)
         );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp294[15] , 
        \temp294[14] , \temp294[13] , \temp294[12] , \temp294[11] , 
        \temp294[10] , \temp294[9] , \temp294[8] , \temp294[7] , \temp294[6] , 
        \temp294[5] , \temp294[4] , \temp294[3] , \temp294[2] , \temp294[1] , 
        \temp294[0] }), .B(InEdges[47:32]), .LEQ(n609), .TC(n609), .GE_GT(n104
        ) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp384[15] , 
        \temp384[14] , \temp384[13] , \temp384[12] , \temp384[11] , 
        \temp384[10] , \temp384[9] , \temp384[8] , \temp384[7] , \temp384[6] , 
        \temp384[5] , \temp384[4] , \temp384[3] , \temp384[2] , \temp384[1] , 
        \temp384[0] }), .B(InEdges[63:48]), .LEQ(n608), .TC(n608), .GE_GT(n112
        ) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n91, n92, 
        n93, n94, n95, n96, n97, n99, n100, n101, n102, n103, n104, n105, n107, 
        n108, n109, n110, n111, n112, n113, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n100), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n104), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, 
        n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
        n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
        n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
        n165, n166;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n123), .B(B[0]), .C(n124), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n124), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n135), .B(B[6]), .Z(n134) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n137), .C(n132), .D(n127), .Z(n136) );
    VMW_OR2 U14 ( .A(B[6]), .B(n135), .Z(n138) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n140), .C(n138), .D(n136), .Z(n139) );
    VMW_NAND2 U16 ( .A(n142), .B(B[8]), .Z(n141) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n144), .C(n139), .D(n134), .Z(n143) );
    VMW_OR2 U18 ( .A(B[8]), .B(n142), .Z(n145) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n147), .C(n145), .D(n143), .Z(n146) );
    VMW_NAND2 U20 ( .A(n149), .B(B[10]), .Z(n148) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n151), .C(n146), .D(n141), .Z(n150) );
    VMW_NAND2 U22 ( .A(n151), .B(A[9]), .Z(n152) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n149), .C(n152), .D(n150), .Z(n153) );
    VMW_NAND2 U24 ( .A(n155), .B(B[12]), .Z(n154) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n157), .C(n153), .D(n148), .Z(n156) );
    VMW_NAND2 U26 ( .A(n157), .B(A[11]), .Z(n158) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n155), .C(n158), .D(n156), .Z(n159) );
    VMW_NAND2 U28 ( .A(n161), .B(B[14]), .Z(n160) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n163), .C(n159), .D(n154), .Z(n162) );
    VMW_NAND2 U30 ( .A(n163), .B(A[13]), .Z(n164) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n161), .C(n164), .D(n162), .Z(n165) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n166), .C(n165), .D(n160), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n155) );
    VMW_INV U34 ( .A(B[7]), .Z(n144) );
    VMW_INV U35 ( .A(A[7]), .Z(n147) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n149) );
    VMW_INV U39 ( .A(B[9]), .Z(n151) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n142) );
    VMW_INV U42 ( .A(A[14]), .Z(n161) );
    VMW_INV U43 ( .A(B[11]), .Z(n157) );
    VMW_INV U44 ( .A(A[5]), .Z(n140) );
    VMW_INV U45 ( .A(B[5]), .Z(n137) );
    VMW_INV U46 ( .A(A[1]), .Z(n124) );
    VMW_INV U47 ( .A(B[15]), .Z(n166) );
    VMW_INV U48 ( .A(B[13]), .Z(n163) );
    VMW_INV U49 ( .A(A[6]), .Z(n135) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n123) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
        n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
        n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
        n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
        n214, n215;
    VMW_OAI21 U3 ( .A(B[15]), .B(n167), .C(n168), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n170), .B(B[2]), .Z(n169) );
    VMW_AO22 U5 ( .A(n172), .B(B[0]), .C(n173), .D(B[1]), .Z(n171) );
    VMW_OR2 U6 ( .A(B[2]), .B(n170), .Z(n174) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n173), .C(n174), .D(n171), .Z(n175) );
    VMW_NAND2 U8 ( .A(n177), .B(B[4]), .Z(n176) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n179), .C(n175), .D(n169), .Z(n178) );
    VMW_OR2 U10 ( .A(B[4]), .B(n177), .Z(n180) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n182), .C(n180), .D(n178), .Z(n181) );
    VMW_NAND2 U12 ( .A(n184), .B(B[6]), .Z(n183) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n186), .C(n181), .D(n176), .Z(n185) );
    VMW_OR2 U14 ( .A(B[6]), .B(n184), .Z(n187) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n189), .C(n187), .D(n185), .Z(n188) );
    VMW_NAND2 U16 ( .A(n191), .B(B[8]), .Z(n190) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n193), .C(n188), .D(n183), .Z(n192) );
    VMW_OR2 U18 ( .A(B[8]), .B(n191), .Z(n194) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n196), .C(n194), .D(n192), .Z(n195) );
    VMW_NAND2 U20 ( .A(n198), .B(B[10]), .Z(n197) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n200), .C(n195), .D(n190), .Z(n199) );
    VMW_NAND2 U22 ( .A(n200), .B(A[9]), .Z(n201) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n198), .C(n201), .D(n199), .Z(n202) );
    VMW_NAND2 U24 ( .A(n204), .B(B[12]), .Z(n203) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n206), .C(n202), .D(n197), .Z(n205) );
    VMW_NAND2 U26 ( .A(n206), .B(A[11]), .Z(n207) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n204), .C(n207), .D(n205), .Z(n208) );
    VMW_NAND2 U28 ( .A(n210), .B(B[14]), .Z(n209) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n212), .C(n208), .D(n203), .Z(n211) );
    VMW_NAND2 U30 ( .A(n212), .B(A[13]), .Z(n213) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n210), .C(n213), .D(n211), .Z(n214) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n215), .C(n214), .D(n209), .Z(n168) );
    VMW_INV U33 ( .A(A[12]), .Z(n204) );
    VMW_INV U34 ( .A(B[7]), .Z(n193) );
    VMW_INV U35 ( .A(A[7]), .Z(n196) );
    VMW_INV U36 ( .A(A[3]), .Z(n182) );
    VMW_INV U37 ( .A(B[3]), .Z(n179) );
    VMW_INV U38 ( .A(A[10]), .Z(n198) );
    VMW_INV U39 ( .A(B[9]), .Z(n200) );
    VMW_INV U40 ( .A(A[4]), .Z(n177) );
    VMW_INV U41 ( .A(A[8]), .Z(n191) );
    VMW_INV U42 ( .A(A[14]), .Z(n210) );
    VMW_INV U43 ( .A(B[11]), .Z(n206) );
    VMW_INV U44 ( .A(A[5]), .Z(n189) );
    VMW_INV U45 ( .A(B[5]), .Z(n186) );
    VMW_INV U46 ( .A(A[1]), .Z(n173) );
    VMW_INV U47 ( .A(B[15]), .Z(n215) );
    VMW_INV U48 ( .A(B[13]), .Z(n212) );
    VMW_INV U49 ( .A(A[6]), .Z(n184) );
    VMW_INV U50 ( .A(A[2]), .Z(n170) );
    VMW_INV U51 ( .A(A[0]), .Z(n172) );
    VMW_INV U52 ( .A(A[15]), .Z(n167) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
        n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
        n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
        n263, n264;
    VMW_OAI21 U3 ( .A(B[15]), .B(n216), .C(n217), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n219), .B(B[2]), .Z(n218) );
    VMW_AO22 U5 ( .A(n221), .B(B[0]), .C(n222), .D(B[1]), .Z(n220) );
    VMW_OR2 U6 ( .A(B[2]), .B(n219), .Z(n223) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n222), .C(n223), .D(n220), .Z(n224) );
    VMW_NAND2 U8 ( .A(n226), .B(B[4]), .Z(n225) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n228), .C(n224), .D(n218), .Z(n227) );
    VMW_OR2 U10 ( .A(B[4]), .B(n226), .Z(n229) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n231), .C(n229), .D(n227), .Z(n230) );
    VMW_NAND2 U12 ( .A(n233), .B(B[6]), .Z(n232) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n235), .C(n230), .D(n225), .Z(n234) );
    VMW_OR2 U14 ( .A(B[6]), .B(n233), .Z(n236) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n238), .C(n236), .D(n234), .Z(n237) );
    VMW_NAND2 U16 ( .A(n240), .B(B[8]), .Z(n239) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n242), .C(n237), .D(n232), .Z(n241) );
    VMW_OR2 U18 ( .A(B[8]), .B(n240), .Z(n243) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n245), .C(n243), .D(n241), .Z(n244) );
    VMW_NAND2 U20 ( .A(n247), .B(B[10]), .Z(n246) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n249), .C(n244), .D(n239), .Z(n248) );
    VMW_NAND2 U22 ( .A(n249), .B(A[9]), .Z(n250) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n247), .C(n250), .D(n248), .Z(n251) );
    VMW_NAND2 U24 ( .A(n253), .B(B[12]), .Z(n252) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n255), .C(n251), .D(n246), .Z(n254) );
    VMW_NAND2 U26 ( .A(n255), .B(A[11]), .Z(n256) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n253), .C(n256), .D(n254), .Z(n257) );
    VMW_NAND2 U28 ( .A(n259), .B(B[14]), .Z(n258) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n261), .C(n257), .D(n252), .Z(n260) );
    VMW_NAND2 U30 ( .A(n261), .B(A[13]), .Z(n262) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n259), .C(n262), .D(n260), .Z(n263) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n264), .C(n263), .D(n258), .Z(n217) );
    VMW_INV U33 ( .A(A[12]), .Z(n253) );
    VMW_INV U34 ( .A(B[7]), .Z(n242) );
    VMW_INV U35 ( .A(A[7]), .Z(n245) );
    VMW_INV U36 ( .A(A[3]), .Z(n231) );
    VMW_INV U37 ( .A(B[3]), .Z(n228) );
    VMW_INV U38 ( .A(A[10]), .Z(n247) );
    VMW_INV U39 ( .A(B[9]), .Z(n249) );
    VMW_INV U40 ( .A(A[4]), .Z(n226) );
    VMW_INV U41 ( .A(A[8]), .Z(n240) );
    VMW_INV U42 ( .A(A[14]), .Z(n259) );
    VMW_INV U43 ( .A(B[11]), .Z(n255) );
    VMW_INV U44 ( .A(A[5]), .Z(n238) );
    VMW_INV U45 ( .A(B[5]), .Z(n235) );
    VMW_INV U46 ( .A(A[1]), .Z(n222) );
    VMW_INV U47 ( .A(B[15]), .Z(n264) );
    VMW_INV U48 ( .A(B[13]), .Z(n261) );
    VMW_INV U49 ( .A(A[6]), .Z(n233) );
    VMW_INV U50 ( .A(A[2]), .Z(n219) );
    VMW_INV U51 ( .A(A[0]), .Z(n221) );
    VMW_INV U52 ( .A(A[15]), .Z(n216) );
endmodule


module NodeAux_INDEGREE5_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp210[13] , \temp484[4] , \temp394[5] , \temp304[13] , 
        \temp210[3] , \temp394[13] , \OutEdge136[14] , \temp394[1] , 
        \temp484[0] , \OutEdge136[10] , \path[2] , \temp394[8] , \temp210[7] , 
        \temp484[9] , \temp394[15] , \path[0] , \temp210[5] , \OutEdge136[12] , 
        \temp210[15] , \temp304[15] , \temp394[3] , \temp484[2] , \temp210[1] , 
        n90, \temp394[11] , \temp484[6] , \temp394[7] , \temp210[8] , 
        \temp304[11] , \temp210[11] , n98, n114, \OutEdge136[2] , \temp304[4] , 
        \OutEdge136[6] , \temp304[9] , \temp304[0] , \temp484[13] , n106, 
        \temp304[2] , \temp484[11] , \OutEdge136[4] , \temp484[15] , 
        \temp304[6] , \OutEdge136[9] , \OutEdge136[0] , \temp484[14] , 
        \OutEdge136[8] , \temp304[7] , \OutEdge136[1] , \temp304[3] , 
        \temp484[10] , \OutEdge136[5] , \OutEdge136[7] , \temp304[8] , 
        \temp304[1] , \temp484[12] , \OutEdge136[3] , \temp304[5] , 
        \temp394[10] , \temp210[0] , \temp484[7] , \temp210[9] , \temp304[10] , 
        \temp394[6] , \temp210[10] , \temp210[4] , \path[1] , \temp394[14] , 
        \OutEdge136[13] , \temp210[14] , \temp394[2] , n122, \temp304[14] , 
        \temp484[3] , \temp394[0] , \temp484[1] , \OutEdge136[11] , 
        \temp210[6] , \path[3] , \temp394[9] , \temp484[8] , \temp210[12] , 
        \temp484[5] , \temp304[12] , \temp394[4] , \OutEdge136[15] , 
        \temp394[12] , \temp210[2] , n667, n668, n669, n670, n671, n672, n673, 
        n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
        n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
        n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
        n710, n711, n712, n713, n714;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U82 ( .Z(n713) );
    VMW_PULLDOWN U83 ( .Z(n710) );
    VMW_PULLDOWN U84 ( .Z(n712) );
    VMW_PULLDOWN U85 ( .Z(n711) );
    VMW_PULLDOWN U86 ( .Z(n714) );
    VMW_AO21 U87 ( .A(\temp484[15] ), .B(n667), .C(n668), .Z(\OutEdge136[15] )
         );
    VMW_OR2 U88 ( .A(n669), .B(Start), .Z(\OutEdge136[14] ) );
    VMW_OR2 U89 ( .A(n670), .B(Start), .Z(\OutEdge136[13] ) );
    VMW_OR2 U90 ( .A(n671), .B(Start), .Z(\OutEdge136[12] ) );
    VMW_OR2 U91 ( .A(n672), .B(Start), .Z(\OutEdge136[11] ) );
    VMW_OR2 U92 ( .A(n673), .B(Start), .Z(\OutEdge136[10] ) );
    VMW_OR2 U93 ( .A(n674), .B(Start), .Z(\OutEdge136[9] ) );
    VMW_OR2 U94 ( .A(n675), .B(Start), .Z(\OutEdge136[8] ) );
    VMW_OR2 U95 ( .A(n676), .B(Start), .Z(\OutEdge136[7] ) );
    VMW_OR2 U96 ( .A(n677), .B(Start), .Z(\OutEdge136[6] ) );
    VMW_OR2 U97 ( .A(n678), .B(Start), .Z(\OutEdge136[5] ) );
    VMW_OR2 U98 ( .A(n679), .B(Start), .Z(\OutEdge136[4] ) );
    VMW_OR2 U99 ( .A(n680), .B(Start), .Z(\OutEdge136[3] ) );
    VMW_OR2 U100 ( .A(n681), .B(Start), .Z(\OutEdge136[2] ) );
    VMW_OR2 U101 ( .A(n682), .B(Start), .Z(\OutEdge136[1] ) );
    VMW_OR2 U102 ( .A(n683), .B(Start), .Z(\OutEdge136[0] ) );
    VMW_AO22 U103 ( .A(\path[1] ), .B(Start), .C(n667), .D(n684), .Z(n709) );
    VMW_AO22 U104 ( .A(Start), .B(\path[3] ), .C(n685), .D(n686), .Z(n708) );
    VMW_OR2 U105 ( .A(n685), .B(n687), .Z(n707) );
    VMW_AO21 U106 ( .A(Start), .B(\path[0] ), .C(n688), .Z(n706) );
    VMW_AO22 U107 ( .A(\temp394[15] ), .B(n689), .C(InEdges[63]), .D(n114), 
        .Z(\temp484[15] ) );
    VMW_NOR5 U108 ( .A(n90), .B(Start), .C(n114), .D(n106), .E(n98), .Z(n685)
         );
    VMW_INV U109 ( .A(Start), .Z(n690) );
    VMW_INV U110 ( .A(n122), .Z(n686) );
    VMW_AND2 U111 ( .A(n690), .B(n686), .Z(n667) );
    VMW_AO22 U112 ( .A(\path[2] ), .B(Start), .C(n122), .D(n690), .Z(n687) );
    VMW_AND4 U113 ( .A(n692), .B(n693), .C(n694), .D(n695), .Z(n691) );
    VMW_INV U114 ( .A(n114), .Z(n689) );
    VMW_INV U115 ( .A(n106), .Z(n696) );
    VMW_OAI211 U116 ( .A(n90), .B(n98), .C(n696), .D(n689), .Z(n684) );
    VMW_OAI21 U117 ( .A(n98), .B(n698), .C(n696), .Z(n697) );
    VMW_AOI21 U118 ( .A(n689), .B(n697), .C(n699), .Z(n688) );
    VMW_AND5 U119 ( .A(n700), .B(n701), .C(n702), .D(n703), .E(n691), .Z(n705)
         );
    VMW_AND3 U120 ( .A(n122), .B(n690), .C(InEdges[79]), .Z(n668) );
    VMW_XNOR2 U121 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n695) );
    VMW_XNOR2 U122 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n694) );
    VMW_XNOR2 U123 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n693) );
    VMW_XNOR2 U124 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n692) );
    VMW_XNOR2 U125 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n703) );
    VMW_XNOR2 U126 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n702) );
    VMW_XNOR2 U127 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n701) );
    VMW_XNOR2 U128 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n700) );
    VMW_AO22 U129 ( .A(OutEdge[9]), .B(n698), .C(InEdges[9]), .D(n90), .Z(
        \temp210[9] ) );
    VMW_AO22 U130 ( .A(\temp210[9] ), .B(n704), .C(InEdges[25]), .D(n98), .Z(
        \temp304[9] ) );
    VMW_AO22 U131 ( .A(InEdges[41]), .B(n106), .C(\temp304[9] ), .D(n696), .Z(
        \temp394[9] ) );
    VMW_AO22 U132 ( .A(InEdges[57]), .B(n114), .C(\temp394[9] ), .D(n689), .Z(
        \temp484[9] ) );
    VMW_AO22 U133 ( .A(OutEdge[8]), .B(n698), .C(InEdges[8]), .D(n90), .Z(
        \temp210[8] ) );
    VMW_AO22 U134 ( .A(\temp210[8] ), .B(n704), .C(InEdges[24]), .D(n98), .Z(
        \temp304[8] ) );
    VMW_AO22 U135 ( .A(InEdges[40]), .B(n106), .C(\temp304[8] ), .D(n696), .Z(
        \temp394[8] ) );
    VMW_AO22 U136 ( .A(InEdges[56]), .B(n114), .C(\temp394[8] ), .D(n689), .Z(
        \temp484[8] ) );
    VMW_AO22 U137 ( .A(OutEdge[7]), .B(n698), .C(InEdges[7]), .D(n90), .Z(
        \temp210[7] ) );
    VMW_AO22 U138 ( .A(\temp210[7] ), .B(n704), .C(InEdges[23]), .D(n98), .Z(
        \temp304[7] ) );
    VMW_AO22 U139 ( .A(InEdges[39]), .B(n106), .C(\temp304[7] ), .D(n696), .Z(
        \temp394[7] ) );
    VMW_AO22 U140 ( .A(InEdges[55]), .B(n114), .C(\temp394[7] ), .D(n689), .Z(
        \temp484[7] ) );
    VMW_AO22 U141 ( .A(OutEdge[6]), .B(n698), .C(InEdges[6]), .D(n90), .Z(
        \temp210[6] ) );
    VMW_AO22 U142 ( .A(\temp210[6] ), .B(n704), .C(InEdges[22]), .D(n98), .Z(
        \temp304[6] ) );
    VMW_AO22 U143 ( .A(InEdges[38]), .B(n106), .C(\temp304[6] ), .D(n696), .Z(
        \temp394[6] ) );
    VMW_AO22 U144 ( .A(InEdges[54]), .B(n114), .C(\temp394[6] ), .D(n689), .Z(
        \temp484[6] ) );
    VMW_AO22 U145 ( .A(OutEdge[5]), .B(n698), .C(InEdges[5]), .D(n90), .Z(
        \temp210[5] ) );
    VMW_AO22 U146 ( .A(\temp210[5] ), .B(n704), .C(InEdges[21]), .D(n98), .Z(
        \temp304[5] ) );
    VMW_AO22 U147 ( .A(InEdges[37]), .B(n106), .C(\temp304[5] ), .D(n696), .Z(
        \temp394[5] ) );
    VMW_AO22 U148 ( .A(InEdges[53]), .B(n114), .C(\temp394[5] ), .D(n689), .Z(
        \temp484[5] ) );
    VMW_AO22 U149 ( .A(OutEdge[4]), .B(n698), .C(InEdges[4]), .D(n90), .Z(
        \temp210[4] ) );
    VMW_AO22 U150 ( .A(\temp210[4] ), .B(n704), .C(InEdges[20]), .D(n98), .Z(
        \temp304[4] ) );
    VMW_AO22 U151 ( .A(InEdges[36]), .B(n106), .C(\temp304[4] ), .D(n696), .Z(
        \temp394[4] ) );
    VMW_AO22 U152 ( .A(InEdges[52]), .B(n114), .C(\temp394[4] ), .D(n689), .Z(
        \temp484[4] ) );
    VMW_AO22 U153 ( .A(OutEdge[3]), .B(n698), .C(InEdges[3]), .D(n90), .Z(
        \temp210[3] ) );
    VMW_AO22 U154 ( .A(\temp210[3] ), .B(n704), .C(InEdges[19]), .D(n98), .Z(
        \temp304[3] ) );
    VMW_AO22 U155 ( .A(InEdges[35]), .B(n106), .C(\temp304[3] ), .D(n696), .Z(
        \temp394[3] ) );
    VMW_AO22 U156 ( .A(InEdges[51]), .B(n114), .C(\temp394[3] ), .D(n689), .Z(
        \temp484[3] ) );
    VMW_AO22 U157 ( .A(OutEdge[2]), .B(n698), .C(InEdges[2]), .D(n90), .Z(
        \temp210[2] ) );
    VMW_AO22 U158 ( .A(\temp210[2] ), .B(n704), .C(InEdges[18]), .D(n98), .Z(
        \temp304[2] ) );
    VMW_AO22 U159 ( .A(InEdges[34]), .B(n106), .C(\temp304[2] ), .D(n696), .Z(
        \temp394[2] ) );
    VMW_AO22 U160 ( .A(InEdges[50]), .B(n114), .C(\temp394[2] ), .D(n689), .Z(
        \temp484[2] ) );
    VMW_AO22 U161 ( .A(OutEdge[1]), .B(n698), .C(InEdges[1]), .D(n90), .Z(
        \temp210[1] ) );
    VMW_AO22 U162 ( .A(\temp210[1] ), .B(n704), .C(InEdges[17]), .D(n98), .Z(
        \temp304[1] ) );
    VMW_AO22 U163 ( .A(InEdges[33]), .B(n106), .C(\temp304[1] ), .D(n696), .Z(
        \temp394[1] ) );
    VMW_AO22 U164 ( .A(InEdges[49]), .B(n114), .C(\temp394[1] ), .D(n689), .Z(
        \temp484[1] ) );
    VMW_AO22 U165 ( .A(OutEdge[15]), .B(n698), .C(InEdges[15]), .D(n90), .Z(
        \temp210[15] ) );
    VMW_AO22 U166 ( .A(\temp210[15] ), .B(n704), .C(InEdges[31]), .D(n98), .Z(
        \temp304[15] ) );
    VMW_AO22 U167 ( .A(InEdges[47]), .B(n106), .C(\temp304[15] ), .D(n696), 
        .Z(\temp394[15] ) );
    VMW_AO22 U168 ( .A(OutEdge[14]), .B(n698), .C(InEdges[14]), .D(n90), .Z(
        \temp210[14] ) );
    VMW_AO22 U169 ( .A(\temp210[14] ), .B(n704), .C(InEdges[30]), .D(n98), .Z(
        \temp304[14] ) );
    VMW_AO22 U170 ( .A(InEdges[46]), .B(n106), .C(\temp304[14] ), .D(n696), 
        .Z(\temp394[14] ) );
    VMW_AO22 U171 ( .A(InEdges[62]), .B(n114), .C(\temp394[14] ), .D(n689), 
        .Z(\temp484[14] ) );
    VMW_AO22 U172 ( .A(OutEdge[13]), .B(n698), .C(InEdges[13]), .D(n90), .Z(
        \temp210[13] ) );
    VMW_AO22 U173 ( .A(\temp210[13] ), .B(n704), .C(InEdges[29]), .D(n98), .Z(
        \temp304[13] ) );
    VMW_AO22 U174 ( .A(InEdges[45]), .B(n106), .C(\temp304[13] ), .D(n696), 
        .Z(\temp394[13] ) );
    VMW_AO22 U175 ( .A(InEdges[61]), .B(n114), .C(\temp394[13] ), .D(n689), 
        .Z(\temp484[13] ) );
    VMW_AO22 U176 ( .A(OutEdge[12]), .B(n698), .C(InEdges[12]), .D(n90), .Z(
        \temp210[12] ) );
    VMW_AO22 U177 ( .A(\temp210[12] ), .B(n704), .C(InEdges[28]), .D(n98), .Z(
        \temp304[12] ) );
    VMW_AO22 U178 ( .A(InEdges[44]), .B(n106), .C(\temp304[12] ), .D(n696), 
        .Z(\temp394[12] ) );
    VMW_AO22 U179 ( .A(InEdges[60]), .B(n114), .C(\temp394[12] ), .D(n689), 
        .Z(\temp484[12] ) );
    VMW_AO22 U180 ( .A(OutEdge[11]), .B(n698), .C(InEdges[11]), .D(n90), .Z(
        \temp210[11] ) );
    VMW_AO22 U181 ( .A(\temp210[11] ), .B(n704), .C(InEdges[27]), .D(n98), .Z(
        \temp304[11] ) );
    VMW_AO22 U182 ( .A(InEdges[43]), .B(n106), .C(\temp304[11] ), .D(n696), 
        .Z(\temp394[11] ) );
    VMW_AO22 U183 ( .A(InEdges[59]), .B(n114), .C(\temp394[11] ), .D(n689), 
        .Z(\temp484[11] ) );
    VMW_AO22 U184 ( .A(OutEdge[10]), .B(n698), .C(InEdges[10]), .D(n90), .Z(
        \temp210[10] ) );
    VMW_AO22 U185 ( .A(\temp210[10] ), .B(n704), .C(InEdges[26]), .D(n98), .Z(
        \temp304[10] ) );
    VMW_AO22 U186 ( .A(InEdges[42]), .B(n106), .C(\temp304[10] ), .D(n696), 
        .Z(\temp394[10] ) );
    VMW_AO22 U187 ( .A(InEdges[58]), .B(n114), .C(\temp394[10] ), .D(n689), 
        .Z(\temp484[10] ) );
    VMW_AO22 U188 ( .A(OutEdge[0]), .B(n698), .C(InEdges[0]), .D(n90), .Z(
        \temp210[0] ) );
    VMW_AO22 U189 ( .A(\temp210[0] ), .B(n704), .C(InEdges[16]), .D(n98), .Z(
        \temp304[0] ) );
    VMW_AO22 U190 ( .A(InEdges[32]), .B(n106), .C(\temp304[0] ), .D(n696), .Z(
        \temp394[0] ) );
    VMW_AO22 U191 ( .A(InEdges[48]), .B(n114), .C(\temp394[0] ), .D(n689), .Z(
        \temp484[0] ) );
    VMW_AO22 U192 ( .A(\temp484[9] ), .B(n686), .C(InEdges[73]), .D(n122), .Z(
        n674) );
    VMW_AO22 U193 ( .A(\temp484[8] ), .B(n686), .C(InEdges[72]), .D(n122), .Z(
        n675) );
    VMW_AO22 U194 ( .A(\temp484[7] ), .B(n686), .C(InEdges[71]), .D(n122), .Z(
        n676) );
    VMW_AO22 U195 ( .A(\temp484[6] ), .B(n686), .C(InEdges[70]), .D(n122), .Z(
        n677) );
    VMW_AO22 U196 ( .A(\temp484[5] ), .B(n686), .C(InEdges[69]), .D(n122), .Z(
        n678) );
    VMW_AO22 U197 ( .A(\temp484[4] ), .B(n686), .C(InEdges[68]), .D(n122), .Z(
        n679) );
    VMW_AO22 U198 ( .A(\temp484[3] ), .B(n686), .C(InEdges[67]), .D(n122), .Z(
        n680) );
    VMW_AO22 U199 ( .A(\temp484[2] ), .B(n686), .C(InEdges[66]), .D(n122), .Z(
        n681) );
    VMW_AO22 U200 ( .A(\temp484[1] ), .B(n686), .C(InEdges[65]), .D(n122), .Z(
        n682) );
    VMW_AO22 U201 ( .A(\temp484[14] ), .B(n686), .C(InEdges[78]), .D(n122), 
        .Z(n669) );
    VMW_AO22 U202 ( .A(\temp484[13] ), .B(n686), .C(InEdges[77]), .D(n122), 
        .Z(n670) );
    VMW_AO22 U203 ( .A(\temp484[12] ), .B(n686), .C(InEdges[76]), .D(n122), 
        .Z(n671) );
    VMW_AO22 U204 ( .A(\temp484[11] ), .B(n686), .C(InEdges[75]), .D(n122), 
        .Z(n672) );
    VMW_AO22 U205 ( .A(\temp484[10] ), .B(n686), .C(InEdges[74]), .D(n122), 
        .Z(n673) );
    VMW_AO22 U206 ( .A(\temp484[0] ), .B(n686), .C(InEdges[64]), .D(n122), .Z(
        n683) );
    VMW_INV U207 ( .A(n90), .Z(n698) );
    VMW_INV U208 ( .A(n98), .Z(n704) );
    VMW_INV U209 ( .A(n667), .Z(n699) );
    VMW_BUFIZ U210 ( .A(\path[3] ), .E(n705), .Z(\PathData[3] ) );
    VMW_BUFIZ U211 ( .A(\path[1] ), .E(n705), .Z(\PathData[1] ) );
    VMW_BUFIZ U212 ( .A(\path[0] ), .E(n705), .Z(\PathData[0] ) );
    VMW_BUFIZ U213 ( .A(\path[2] ), .E(n705), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n706), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n707), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n708), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n709), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge136[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge136[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge136[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge136[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge136[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge136[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge136[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge136[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge136[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge136[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge136[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge136[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge136[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge136[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge136[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge136[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_4 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n714), .TC(n714), .GE_GT(n90) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_3 lte_55_4 ( .A({\temp484[15] , 
        \temp484[14] , \temp484[13] , \temp484[12] , \temp484[11] , 
        \temp484[10] , \temp484[9] , \temp484[8] , \temp484[7] , \temp484[6] , 
        \temp484[5] , \temp484[4] , \temp484[3] , \temp484[2] , \temp484[1] , 
        \temp484[0] }), .B(InEdges[79:64]), .LEQ(n713), .TC(n713), .GE_GT(n122
        ) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_2 lte_55_2 ( .A({\temp304[15] , 
        \temp304[14] , \temp304[13] , \temp304[12] , \temp304[11] , 
        \temp304[10] , \temp304[9] , \temp304[8] , \temp304[7] , \temp304[6] , 
        \temp304[5] , \temp304[4] , \temp304[3] , \temp304[2] , \temp304[1] , 
        \temp304[0] }), .B(InEdges[47:32]), .LEQ(n712), .TC(n712), .GE_GT(n106
        ) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_1 lte_55_1 ( .A({\temp210[15] , 
        \temp210[14] , \temp210[13] , \temp210[12] , \temp210[11] , 
        \temp210[10] , \temp210[9] , \temp210[8] , \temp210[7] , \temp210[6] , 
        \temp210[5] , \temp210[4] , \temp210[3] , \temp210[2] , \temp210[1] , 
        \temp210[0] }), .B(InEdges[31:16]), .LEQ(n711), .TC(n711), .GE_GT(n98)
         );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp394[15] , 
        \temp394[14] , \temp394[13] , \temp394[12] , \temp394[11] , 
        \temp394[10] , \temp394[9] , \temp394[8] , \temp394[7] , \temp394[6] , 
        \temp394[5] , \temp394[4] , \temp394[3] , \temp394[2] , \temp394[1] , 
        \temp394[0] }), .B(InEdges[63:48]), .LEQ(n710), .TC(n710), .GE_GT(n114
        ) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n93, n94, n95, n96, n97, n98, n99, n101, n102, n103, n104, n105, n106, 
        n107, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n91), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n99), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n107), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n125, n126, n127, n128, 
        n129, n130, n131, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
        n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
        n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
        n166, n167;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n134), .C(n131), .D(n129), .Z(n133) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n133), .D(n127), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n145), .C(n140), .D(n135), .Z(n144) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n146) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n148), .C(n146), .D(n144), .Z(n147) );
    VMW_NAND2 U20 ( .A(n150), .B(B[10]), .Z(n149) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n152), .C(n147), .D(n142), .Z(n151) );
    VMW_NAND2 U22 ( .A(n152), .B(A[9]), .Z(n153) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U24 ( .A(n156), .B(B[12]), .Z(n155) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_NAND2 U26 ( .A(n158), .B(A[11]), .Z(n159) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_NAND2 U28 ( .A(n162), .B(B[14]), .Z(n161) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_NAND2 U30 ( .A(n164), .B(A[13]), .Z(n165) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n162), .C(n165), .D(n163), .Z(n166) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n167), .C(n166), .D(n161), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n156) );
    VMW_INV U34 ( .A(B[7]), .Z(n145) );
    VMW_INV U35 ( .A(A[7]), .Z(n148) );
    VMW_INV U36 ( .A(A[3]), .Z(n134) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n150) );
    VMW_INV U39 ( .A(B[9]), .Z(n152) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n143) );
    VMW_INV U42 ( .A(A[14]), .Z(n162) );
    VMW_INV U43 ( .A(B[11]), .Z(n158) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n167) );
    VMW_INV U48 ( .A(B[13]), .Z(n164) );
    VMW_INV U49 ( .A(A[6]), .Z(n136) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
        n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216;
    VMW_OAI21 U3 ( .A(B[15]), .B(n168), .C(n169), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n171), .B(B[2]), .Z(n170) );
    VMW_AO22 U5 ( .A(n173), .B(B[0]), .C(n174), .D(B[1]), .Z(n172) );
    VMW_OR2 U6 ( .A(B[2]), .B(n171), .Z(n175) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n174), .C(n175), .D(n172), .Z(n176) );
    VMW_NAND2 U8 ( .A(n178), .B(B[4]), .Z(n177) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n180), .C(n176), .D(n170), .Z(n179) );
    VMW_OR2 U10 ( .A(B[4]), .B(n178), .Z(n181) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n183), .C(n181), .D(n179), .Z(n182) );
    VMW_NAND2 U12 ( .A(n185), .B(B[6]), .Z(n184) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n187), .C(n182), .D(n177), .Z(n186) );
    VMW_OR2 U14 ( .A(B[6]), .B(n185), .Z(n188) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n190), .C(n188), .D(n186), .Z(n189) );
    VMW_NAND2 U16 ( .A(n192), .B(B[8]), .Z(n191) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n194), .C(n189), .D(n184), .Z(n193) );
    VMW_OR2 U18 ( .A(B[8]), .B(n192), .Z(n195) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n197), .C(n195), .D(n193), .Z(n196) );
    VMW_NAND2 U20 ( .A(n199), .B(B[10]), .Z(n198) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n201), .C(n196), .D(n191), .Z(n200) );
    VMW_NAND2 U22 ( .A(n201), .B(A[9]), .Z(n202) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n199), .C(n202), .D(n200), .Z(n203) );
    VMW_NAND2 U24 ( .A(n205), .B(B[12]), .Z(n204) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n207), .C(n203), .D(n198), .Z(n206) );
    VMW_NAND2 U26 ( .A(n207), .B(A[11]), .Z(n208) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n205), .C(n208), .D(n206), .Z(n209) );
    VMW_NAND2 U28 ( .A(n211), .B(B[14]), .Z(n210) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n213), .C(n209), .D(n204), .Z(n212) );
    VMW_NAND2 U30 ( .A(n213), .B(A[13]), .Z(n214) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n211), .C(n214), .D(n212), .Z(n215) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n216), .C(n215), .D(n210), .Z(n169) );
    VMW_INV U33 ( .A(A[12]), .Z(n205) );
    VMW_INV U34 ( .A(B[7]), .Z(n194) );
    VMW_INV U35 ( .A(A[7]), .Z(n197) );
    VMW_INV U36 ( .A(A[3]), .Z(n183) );
    VMW_INV U37 ( .A(B[3]), .Z(n180) );
    VMW_INV U38 ( .A(A[10]), .Z(n199) );
    VMW_INV U39 ( .A(B[9]), .Z(n201) );
    VMW_INV U40 ( .A(A[4]), .Z(n178) );
    VMW_INV U41 ( .A(A[8]), .Z(n192) );
    VMW_INV U42 ( .A(A[14]), .Z(n211) );
    VMW_INV U43 ( .A(B[11]), .Z(n207) );
    VMW_INV U44 ( .A(A[5]), .Z(n190) );
    VMW_INV U45 ( .A(B[5]), .Z(n187) );
    VMW_INV U46 ( .A(A[1]), .Z(n174) );
    VMW_INV U47 ( .A(B[15]), .Z(n216) );
    VMW_INV U48 ( .A(B[13]), .Z(n213) );
    VMW_INV U49 ( .A(A[6]), .Z(n185) );
    VMW_INV U50 ( .A(A[2]), .Z(n171) );
    VMW_INV U51 ( .A(A[0]), .Z(n173) );
    VMW_INV U52 ( .A(A[15]), .Z(n168) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
        n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265;
    VMW_OAI21 U3 ( .A(B[15]), .B(n217), .C(n218), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n220), .B(B[2]), .Z(n219) );
    VMW_AO22 U5 ( .A(n222), .B(B[0]), .C(n223), .D(B[1]), .Z(n221) );
    VMW_OR2 U6 ( .A(B[2]), .B(n220), .Z(n224) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n223), .C(n224), .D(n221), .Z(n225) );
    VMW_NAND2 U8 ( .A(n227), .B(B[4]), .Z(n226) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n229), .C(n225), .D(n219), .Z(n228) );
    VMW_OR2 U10 ( .A(B[4]), .B(n227), .Z(n230) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n232), .C(n230), .D(n228), .Z(n231) );
    VMW_NAND2 U12 ( .A(n234), .B(B[6]), .Z(n233) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n236), .C(n231), .D(n226), .Z(n235) );
    VMW_OR2 U14 ( .A(B[6]), .B(n234), .Z(n237) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n239), .C(n237), .D(n235), .Z(n238) );
    VMW_NAND2 U16 ( .A(n241), .B(B[8]), .Z(n240) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n243), .C(n238), .D(n233), .Z(n242) );
    VMW_OR2 U18 ( .A(B[8]), .B(n241), .Z(n244) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n246), .C(n244), .D(n242), .Z(n245) );
    VMW_NAND2 U20 ( .A(n248), .B(B[10]), .Z(n247) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n250), .C(n245), .D(n240), .Z(n249) );
    VMW_NAND2 U22 ( .A(n250), .B(A[9]), .Z(n251) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n248), .C(n251), .D(n249), .Z(n252) );
    VMW_NAND2 U24 ( .A(n254), .B(B[12]), .Z(n253) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n256), .C(n252), .D(n247), .Z(n255) );
    VMW_NAND2 U26 ( .A(n256), .B(A[11]), .Z(n257) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n254), .C(n257), .D(n255), .Z(n258) );
    VMW_NAND2 U28 ( .A(n260), .B(B[14]), .Z(n259) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n262), .C(n258), .D(n253), .Z(n261) );
    VMW_NAND2 U30 ( .A(n262), .B(A[13]), .Z(n263) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n260), .C(n263), .D(n261), .Z(n264) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n265), .C(n264), .D(n259), .Z(n218) );
    VMW_INV U33 ( .A(A[12]), .Z(n254) );
    VMW_INV U34 ( .A(B[7]), .Z(n243) );
    VMW_INV U35 ( .A(A[7]), .Z(n246) );
    VMW_INV U36 ( .A(A[3]), .Z(n232) );
    VMW_INV U37 ( .A(B[3]), .Z(n229) );
    VMW_INV U38 ( .A(A[10]), .Z(n248) );
    VMW_INV U39 ( .A(B[9]), .Z(n250) );
    VMW_INV U40 ( .A(A[4]), .Z(n227) );
    VMW_INV U41 ( .A(A[8]), .Z(n241) );
    VMW_INV U42 ( .A(A[14]), .Z(n260) );
    VMW_INV U43 ( .A(B[11]), .Z(n256) );
    VMW_INV U44 ( .A(A[5]), .Z(n239) );
    VMW_INV U45 ( .A(B[5]), .Z(n236) );
    VMW_INV U46 ( .A(A[1]), .Z(n223) );
    VMW_INV U47 ( .A(B[15]), .Z(n265) );
    VMW_INV U48 ( .A(B[13]), .Z(n262) );
    VMW_INV U49 ( .A(A[6]), .Z(n234) );
    VMW_INV U50 ( .A(A[2]), .Z(n220) );
    VMW_INV U51 ( .A(A[0]), .Z(n222) );
    VMW_INV U52 ( .A(A[15]), .Z(n217) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
        n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
        n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
        n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
        n313, n314;
    VMW_OAI21 U3 ( .A(B[15]), .B(n266), .C(n267), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n269), .B(B[2]), .Z(n268) );
    VMW_AO22 U5 ( .A(n271), .B(B[0]), .C(n272), .D(B[1]), .Z(n270) );
    VMW_OR2 U6 ( .A(B[2]), .B(n269), .Z(n273) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n272), .C(n273), .D(n270), .Z(n274) );
    VMW_NAND2 U8 ( .A(n276), .B(B[4]), .Z(n275) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n278), .C(n274), .D(n268), .Z(n277) );
    VMW_OR2 U10 ( .A(B[4]), .B(n276), .Z(n279) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n281), .C(n279), .D(n277), .Z(n280) );
    VMW_NAND2 U12 ( .A(n283), .B(B[6]), .Z(n282) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n285), .C(n280), .D(n275), .Z(n284) );
    VMW_OR2 U14 ( .A(B[6]), .B(n283), .Z(n286) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n288), .C(n286), .D(n284), .Z(n287) );
    VMW_NAND2 U16 ( .A(n290), .B(B[8]), .Z(n289) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n292), .C(n287), .D(n282), .Z(n291) );
    VMW_OR2 U18 ( .A(B[8]), .B(n290), .Z(n293) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n295), .C(n293), .D(n291), .Z(n294) );
    VMW_NAND2 U20 ( .A(n297), .B(B[10]), .Z(n296) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n299), .C(n294), .D(n289), .Z(n298) );
    VMW_NAND2 U22 ( .A(n299), .B(A[9]), .Z(n300) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n297), .C(n300), .D(n298), .Z(n301) );
    VMW_NAND2 U24 ( .A(n303), .B(B[12]), .Z(n302) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n305), .C(n301), .D(n296), .Z(n304) );
    VMW_NAND2 U26 ( .A(n305), .B(A[11]), .Z(n306) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n303), .C(n306), .D(n304), .Z(n307) );
    VMW_NAND2 U28 ( .A(n309), .B(B[14]), .Z(n308) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n311), .C(n307), .D(n302), .Z(n310) );
    VMW_NAND2 U30 ( .A(n311), .B(A[13]), .Z(n312) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n309), .C(n312), .D(n310), .Z(n313) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n314), .C(n313), .D(n308), .Z(n267) );
    VMW_INV U33 ( .A(A[12]), .Z(n303) );
    VMW_INV U34 ( .A(B[7]), .Z(n292) );
    VMW_INV U35 ( .A(A[7]), .Z(n295) );
    VMW_INV U36 ( .A(A[3]), .Z(n281) );
    VMW_INV U37 ( .A(B[3]), .Z(n278) );
    VMW_INV U38 ( .A(A[10]), .Z(n297) );
    VMW_INV U39 ( .A(B[9]), .Z(n299) );
    VMW_INV U40 ( .A(A[4]), .Z(n276) );
    VMW_INV U41 ( .A(A[8]), .Z(n290) );
    VMW_INV U42 ( .A(A[14]), .Z(n309) );
    VMW_INV U43 ( .A(B[11]), .Z(n305) );
    VMW_INV U44 ( .A(A[5]), .Z(n288) );
    VMW_INV U45 ( .A(B[5]), .Z(n285) );
    VMW_INV U46 ( .A(A[1]), .Z(n272) );
    VMW_INV U47 ( .A(B[15]), .Z(n314) );
    VMW_INV U48 ( .A(B[13]), .Z(n311) );
    VMW_INV U49 ( .A(A[6]), .Z(n283) );
    VMW_INV U50 ( .A(A[2]), .Z(n269) );
    VMW_INV U51 ( .A(A[0]), .Z(n271) );
    VMW_INV U52 ( .A(A[15]), .Z(n266) );
endmodule


module NodeAux_INDEGREE6_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp494[7] , \temp584[2] , n100, \OutEdge146[7] , \temp314[15] , 
        \OutEdge146[12] , \temp314[11] , \OutEdge146[3] , \temp494[3] , 
        \temp584[6] , \path[2] , \path[0] , \temp314[13] , \temp494[1] , 
        \OutEdge146[1] , \temp584[4] , \OutEdge146[8] , \temp494[8] , n132, 
        \OutEdge146[10] , \temp584[0] , \OutEdge146[5] , \temp494[5] , 
        \OutEdge146[14] , \temp584[9] , \temp220[10] , \temp220[4] , 
        \temp314[7] , \temp494[11] , \temp404[6] , \temp584[13] , 
        \temp404[11] , \temp404[2] , \temp220[0] , \temp314[3] , \temp494[15] , 
        \temp220[14] , \temp404[15] , \temp220[9] , \temp404[9] , \temp314[8] , 
        \temp220[2] , \temp404[0] , \temp314[1] , \temp584[15] , n108, 
        \temp404[13] , \temp584[11] , \temp220[12] , \temp220[6] , 
        \temp314[5] , \temp404[4] , \temp494[13] , \temp404[12] , 
        \temp584[10] , \temp220[7] , \temp314[4] , n124, \temp494[12] , 
        \temp220[13] , \temp404[5] , \temp404[8] , \temp314[9] , \temp404[1] , 
        \temp220[3] , \temp314[0] , \temp584[14] , \temp404[3] , \temp220[15] , 
        \temp220[1] , \temp314[2] , \temp494[14] , \temp220[8] , \temp404[14] , 
        n116, \temp220[5] , \temp314[6] , \temp494[10] , \temp220[11] , 
        \temp404[7] , \temp584[12] , \temp404[10] , \temp584[1] , \temp494[4] , 
        \OutEdge146[4] , \OutEdge146[15] , \temp584[8] , \path[1] , 
        \temp494[0] , \OutEdge146[0] , \temp314[12] , n92, \temp584[5] , 
        \OutEdge146[9] , \temp494[9] , \OutEdge146[11] , \OutEdge146[13] , 
        \temp494[2] , \OutEdge146[2] , \temp314[10] , \temp584[7] , \path[3] , 
        \temp584[3] , \temp314[14] , \temp494[6] , \OutEdge146[6] , n767, n768, 
        n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
        n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
        n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
        n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
        n817, n818;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U91 ( .Z(n817) );
    VMW_PULLDOWN U92 ( .Z(n816) );
    VMW_PULLDOWN U93 ( .Z(n815) );
    VMW_PULLDOWN U94 ( .Z(n814) );
    VMW_PULLDOWN U95 ( .Z(n818) );
    VMW_PULLDOWN U96 ( .Z(n813) );
    VMW_NOR2 U97 ( .A(Start), .B(n767), .Z(\OutEdge146[15] ) );
    VMW_NAND2 U98 ( .A(n768), .B(n769), .Z(\OutEdge146[14] ) );
    VMW_NAND2 U99 ( .A(n770), .B(n769), .Z(\OutEdge146[13] ) );
    VMW_NAND2 U100 ( .A(n771), .B(n769), .Z(\OutEdge146[12] ) );
    VMW_NAND2 U101 ( .A(n772), .B(n769), .Z(\OutEdge146[11] ) );
    VMW_NAND2 U102 ( .A(n773), .B(n769), .Z(\OutEdge146[10] ) );
    VMW_NAND2 U103 ( .A(n774), .B(n769), .Z(\OutEdge146[9] ) );
    VMW_NAND2 U104 ( .A(n775), .B(n769), .Z(\OutEdge146[8] ) );
    VMW_NAND2 U105 ( .A(n776), .B(n769), .Z(\OutEdge146[7] ) );
    VMW_NAND2 U106 ( .A(n777), .B(n769), .Z(\OutEdge146[6] ) );
    VMW_NAND2 U107 ( .A(n778), .B(n769), .Z(\OutEdge146[5] ) );
    VMW_NAND2 U108 ( .A(n779), .B(n769), .Z(\OutEdge146[4] ) );
    VMW_NAND2 U109 ( .A(n780), .B(n769), .Z(\OutEdge146[3] ) );
    VMW_NAND2 U110 ( .A(n781), .B(n769), .Z(\OutEdge146[2] ) );
    VMW_NAND2 U111 ( .A(n782), .B(n769), .Z(\OutEdge146[1] ) );
    VMW_NAND2 U112 ( .A(n783), .B(n769), .Z(\OutEdge146[0] ) );
    VMW_AO21 U113 ( .A(Start), .B(\path[1] ), .C(n784), .Z(n812) );
    VMW_AO22 U114 ( .A(\path[3] ), .B(Start), .C(n785), .D(n786), .Z(n811) );
    VMW_OR2 U115 ( .A(n787), .B(n788), .Z(n809) );
    VMW_OR3 U116 ( .A(n785), .B(n124), .C(n132), .Z(n789) );
    VMW_AO22 U117 ( .A(\temp494[15] ), .B(n790), .C(InEdges[79]), .D(n124), 
        .Z(\temp584[15] ) );
    VMW_NAND2 U118 ( .A(n769), .B(n790), .Z(n791) );
    VMW_AND4 U119 ( .A(n792), .B(n793), .C(n794), .D(n795), .Z(n785) );
    VMW_INV U120 ( .A(Start), .Z(n769) );
    VMW_OAI22 U121 ( .A(n789), .B(Start), .C(\path[2] ), .D(n769), .Z(n796) );
    VMW_MUX2I U122 ( .A(\temp584[15] ), .B(InEdges[95]), .S(n132), .Z(n767) );
    VMW_NOR2 U123 ( .A(n132), .B(n791), .Z(n786) );
    VMW_AND4 U124 ( .A(n798), .B(n799), .C(n800), .D(n801), .Z(n797) );
    VMW_INV U125 ( .A(n116), .Z(n795) );
    VMW_AOI211 U126 ( .A(n794), .B(n792), .C(n108), .D(n116), .Z(n802) );
    VMW_NOR3 U127 ( .A(n802), .B(n132), .C(n791), .Z(n784) );
    VMW_OAI21 U128 ( .A(n100), .B(n794), .C(n793), .Z(n803) );
    VMW_AOI21 U129 ( .A(n795), .B(n803), .C(n791), .Z(n788) );
    VMW_AND5 U130 ( .A(n804), .B(n805), .C(n806), .D(n807), .E(n797), .Z(n808)
         );
    VMW_XNOR2 U131 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n801) );
    VMW_XNOR2 U132 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n800) );
    VMW_XNOR2 U133 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n799) );
    VMW_XNOR2 U134 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n798) );
    VMW_XNOR2 U135 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n807) );
    VMW_XNOR2 U136 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n806) );
    VMW_XNOR2 U137 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n805) );
    VMW_XNOR2 U138 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n804) );
    VMW_AO22 U139 ( .A(InEdges[9]), .B(n92), .C(OutEdge[9]), .D(n794), .Z(
        \temp220[9] ) );
    VMW_AO22 U140 ( .A(InEdges[25]), .B(n100), .C(\temp220[9] ), .D(n792), .Z(
        \temp314[9] ) );
    VMW_AO22 U141 ( .A(\temp314[9] ), .B(n793), .C(InEdges[41]), .D(n108), .Z(
        \temp404[9] ) );
    VMW_AO22 U142 ( .A(InEdges[57]), .B(n116), .C(\temp404[9] ), .D(n795), .Z(
        \temp494[9] ) );
    VMW_AO22 U143 ( .A(\temp494[9] ), .B(n790), .C(InEdges[73]), .D(n124), .Z(
        \temp584[9] ) );
    VMW_AO22 U144 ( .A(InEdges[8]), .B(n92), .C(OutEdge[8]), .D(n794), .Z(
        \temp220[8] ) );
    VMW_AO22 U145 ( .A(InEdges[24]), .B(n100), .C(\temp220[8] ), .D(n792), .Z(
        \temp314[8] ) );
    VMW_AO22 U146 ( .A(\temp314[8] ), .B(n793), .C(InEdges[40]), .D(n108), .Z(
        \temp404[8] ) );
    VMW_AO22 U147 ( .A(InEdges[56]), .B(n116), .C(\temp404[8] ), .D(n795), .Z(
        \temp494[8] ) );
    VMW_AO22 U148 ( .A(\temp494[8] ), .B(n790), .C(InEdges[72]), .D(n124), .Z(
        \temp584[8] ) );
    VMW_AO22 U149 ( .A(InEdges[7]), .B(n92), .C(OutEdge[7]), .D(n794), .Z(
        \temp220[7] ) );
    VMW_AO22 U150 ( .A(InEdges[23]), .B(n100), .C(\temp220[7] ), .D(n792), .Z(
        \temp314[7] ) );
    VMW_AO22 U151 ( .A(\temp314[7] ), .B(n793), .C(InEdges[39]), .D(n108), .Z(
        \temp404[7] ) );
    VMW_AO22 U152 ( .A(InEdges[55]), .B(n116), .C(\temp404[7] ), .D(n795), .Z(
        \temp494[7] ) );
    VMW_AO22 U153 ( .A(\temp494[7] ), .B(n790), .C(InEdges[71]), .D(n124), .Z(
        \temp584[7] ) );
    VMW_AO22 U154 ( .A(InEdges[6]), .B(n92), .C(OutEdge[6]), .D(n794), .Z(
        \temp220[6] ) );
    VMW_AO22 U155 ( .A(InEdges[22]), .B(n100), .C(\temp220[6] ), .D(n792), .Z(
        \temp314[6] ) );
    VMW_AO22 U156 ( .A(\temp314[6] ), .B(n793), .C(InEdges[38]), .D(n108), .Z(
        \temp404[6] ) );
    VMW_AO22 U157 ( .A(InEdges[54]), .B(n116), .C(\temp404[6] ), .D(n795), .Z(
        \temp494[6] ) );
    VMW_AO22 U158 ( .A(\temp494[6] ), .B(n790), .C(InEdges[70]), .D(n124), .Z(
        \temp584[6] ) );
    VMW_AO22 U159 ( .A(InEdges[5]), .B(n92), .C(OutEdge[5]), .D(n794), .Z(
        \temp220[5] ) );
    VMW_AO22 U160 ( .A(InEdges[21]), .B(n100), .C(\temp220[5] ), .D(n792), .Z(
        \temp314[5] ) );
    VMW_AO22 U161 ( .A(\temp314[5] ), .B(n793), .C(InEdges[37]), .D(n108), .Z(
        \temp404[5] ) );
    VMW_AO22 U162 ( .A(InEdges[53]), .B(n116), .C(\temp404[5] ), .D(n795), .Z(
        \temp494[5] ) );
    VMW_AO22 U163 ( .A(\temp494[5] ), .B(n790), .C(InEdges[69]), .D(n124), .Z(
        \temp584[5] ) );
    VMW_AO22 U164 ( .A(InEdges[4]), .B(n92), .C(OutEdge[4]), .D(n794), .Z(
        \temp220[4] ) );
    VMW_AO22 U165 ( .A(InEdges[20]), .B(n100), .C(\temp220[4] ), .D(n792), .Z(
        \temp314[4] ) );
    VMW_AO22 U166 ( .A(\temp314[4] ), .B(n793), .C(InEdges[36]), .D(n108), .Z(
        \temp404[4] ) );
    VMW_AO22 U167 ( .A(InEdges[52]), .B(n116), .C(\temp404[4] ), .D(n795), .Z(
        \temp494[4] ) );
    VMW_AO22 U168 ( .A(\temp494[4] ), .B(n790), .C(InEdges[68]), .D(n124), .Z(
        \temp584[4] ) );
    VMW_AO22 U169 ( .A(InEdges[3]), .B(n92), .C(OutEdge[3]), .D(n794), .Z(
        \temp220[3] ) );
    VMW_AO22 U170 ( .A(InEdges[19]), .B(n100), .C(\temp220[3] ), .D(n792), .Z(
        \temp314[3] ) );
    VMW_AO22 U171 ( .A(\temp314[3] ), .B(n793), .C(InEdges[35]), .D(n108), .Z(
        \temp404[3] ) );
    VMW_AO22 U172 ( .A(InEdges[51]), .B(n116), .C(\temp404[3] ), .D(n795), .Z(
        \temp494[3] ) );
    VMW_AO22 U173 ( .A(\temp494[3] ), .B(n790), .C(InEdges[67]), .D(n124), .Z(
        \temp584[3] ) );
    VMW_AO22 U174 ( .A(InEdges[2]), .B(n92), .C(OutEdge[2]), .D(n794), .Z(
        \temp220[2] ) );
    VMW_AO22 U175 ( .A(InEdges[18]), .B(n100), .C(\temp220[2] ), .D(n792), .Z(
        \temp314[2] ) );
    VMW_AO22 U176 ( .A(\temp314[2] ), .B(n793), .C(InEdges[34]), .D(n108), .Z(
        \temp404[2] ) );
    VMW_AO22 U177 ( .A(InEdges[50]), .B(n116), .C(\temp404[2] ), .D(n795), .Z(
        \temp494[2] ) );
    VMW_AO22 U178 ( .A(\temp494[2] ), .B(n790), .C(InEdges[66]), .D(n124), .Z(
        \temp584[2] ) );
    VMW_AO22 U179 ( .A(InEdges[1]), .B(n92), .C(OutEdge[1]), .D(n794), .Z(
        \temp220[1] ) );
    VMW_AO22 U180 ( .A(InEdges[17]), .B(n100), .C(\temp220[1] ), .D(n792), .Z(
        \temp314[1] ) );
    VMW_AO22 U181 ( .A(\temp314[1] ), .B(n793), .C(InEdges[33]), .D(n108), .Z(
        \temp404[1] ) );
    VMW_AO22 U182 ( .A(InEdges[49]), .B(n116), .C(\temp404[1] ), .D(n795), .Z(
        \temp494[1] ) );
    VMW_AO22 U183 ( .A(\temp494[1] ), .B(n790), .C(InEdges[65]), .D(n124), .Z(
        \temp584[1] ) );
    VMW_AO22 U184 ( .A(InEdges[15]), .B(n92), .C(OutEdge[15]), .D(n794), .Z(
        \temp220[15] ) );
    VMW_AO22 U185 ( .A(InEdges[31]), .B(n100), .C(\temp220[15] ), .D(n792), 
        .Z(\temp314[15] ) );
    VMW_AO22 U186 ( .A(\temp314[15] ), .B(n793), .C(InEdges[47]), .D(n108), 
        .Z(\temp404[15] ) );
    VMW_AO22 U187 ( .A(InEdges[63]), .B(n116), .C(\temp404[15] ), .D(n795), 
        .Z(\temp494[15] ) );
    VMW_AO22 U188 ( .A(InEdges[14]), .B(n92), .C(OutEdge[14]), .D(n794), .Z(
        \temp220[14] ) );
    VMW_AO22 U189 ( .A(InEdges[30]), .B(n100), .C(\temp220[14] ), .D(n792), 
        .Z(\temp314[14] ) );
    VMW_AO22 U190 ( .A(\temp314[14] ), .B(n793), .C(InEdges[46]), .D(n108), 
        .Z(\temp404[14] ) );
    VMW_AO22 U191 ( .A(InEdges[62]), .B(n116), .C(\temp404[14] ), .D(n795), 
        .Z(\temp494[14] ) );
    VMW_AO22 U192 ( .A(\temp494[14] ), .B(n790), .C(InEdges[78]), .D(n124), 
        .Z(\temp584[14] ) );
    VMW_AO22 U193 ( .A(InEdges[13]), .B(n92), .C(OutEdge[13]), .D(n794), .Z(
        \temp220[13] ) );
    VMW_AO22 U194 ( .A(InEdges[29]), .B(n100), .C(\temp220[13] ), .D(n792), 
        .Z(\temp314[13] ) );
    VMW_AO22 U195 ( .A(\temp314[13] ), .B(n793), .C(InEdges[45]), .D(n108), 
        .Z(\temp404[13] ) );
    VMW_AO22 U196 ( .A(InEdges[61]), .B(n116), .C(\temp404[13] ), .D(n795), 
        .Z(\temp494[13] ) );
    VMW_AO22 U197 ( .A(\temp494[13] ), .B(n790), .C(InEdges[77]), .D(n124), 
        .Z(\temp584[13] ) );
    VMW_AO22 U198 ( .A(InEdges[12]), .B(n92), .C(OutEdge[12]), .D(n794), .Z(
        \temp220[12] ) );
    VMW_AO22 U199 ( .A(InEdges[28]), .B(n100), .C(\temp220[12] ), .D(n792), 
        .Z(\temp314[12] ) );
    VMW_AO22 U200 ( .A(\temp314[12] ), .B(n793), .C(InEdges[44]), .D(n108), 
        .Z(\temp404[12] ) );
    VMW_AO22 U201 ( .A(InEdges[60]), .B(n116), .C(\temp404[12] ), .D(n795), 
        .Z(\temp494[12] ) );
    VMW_AO22 U202 ( .A(\temp494[12] ), .B(n790), .C(InEdges[76]), .D(n124), 
        .Z(\temp584[12] ) );
    VMW_AO22 U203 ( .A(InEdges[11]), .B(n92), .C(OutEdge[11]), .D(n794), .Z(
        \temp220[11] ) );
    VMW_AO22 U204 ( .A(InEdges[27]), .B(n100), .C(\temp220[11] ), .D(n792), 
        .Z(\temp314[11] ) );
    VMW_AO22 U205 ( .A(\temp314[11] ), .B(n793), .C(InEdges[43]), .D(n108), 
        .Z(\temp404[11] ) );
    VMW_AO22 U206 ( .A(InEdges[59]), .B(n116), .C(\temp404[11] ), .D(n795), 
        .Z(\temp494[11] ) );
    VMW_AO22 U207 ( .A(\temp494[11] ), .B(n790), .C(InEdges[75]), .D(n124), 
        .Z(\temp584[11] ) );
    VMW_AO22 U208 ( .A(InEdges[10]), .B(n92), .C(OutEdge[10]), .D(n794), .Z(
        \temp220[10] ) );
    VMW_AO22 U209 ( .A(InEdges[26]), .B(n100), .C(\temp220[10] ), .D(n792), 
        .Z(\temp314[10] ) );
    VMW_AO22 U210 ( .A(\temp314[10] ), .B(n793), .C(InEdges[42]), .D(n108), 
        .Z(\temp404[10] ) );
    VMW_AO22 U211 ( .A(InEdges[58]), .B(n116), .C(\temp404[10] ), .D(n795), 
        .Z(\temp494[10] ) );
    VMW_AO22 U212 ( .A(\temp494[10] ), .B(n790), .C(InEdges[74]), .D(n124), 
        .Z(\temp584[10] ) );
    VMW_AO22 U213 ( .A(InEdges[0]), .B(n92), .C(OutEdge[0]), .D(n794), .Z(
        \temp220[0] ) );
    VMW_AO22 U214 ( .A(InEdges[16]), .B(n100), .C(\temp220[0] ), .D(n792), .Z(
        \temp314[0] ) );
    VMW_AO22 U215 ( .A(\temp314[0] ), .B(n793), .C(InEdges[32]), .D(n108), .Z(
        \temp404[0] ) );
    VMW_AO22 U216 ( .A(InEdges[48]), .B(n116), .C(\temp404[0] ), .D(n795), .Z(
        \temp494[0] ) );
    VMW_AO22 U217 ( .A(\temp494[0] ), .B(n790), .C(InEdges[64]), .D(n124), .Z(
        \temp584[0] ) );
    VMW_AO22 U218 ( .A(n132), .B(n769), .C(\path[0] ), .D(Start), .Z(n787) );
    VMW_MUX2I U219 ( .A(\temp584[9] ), .B(InEdges[89]), .S(n132), .Z(n774) );
    VMW_MUX2I U220 ( .A(\temp584[8] ), .B(InEdges[88]), .S(n132), .Z(n775) );
    VMW_MUX2I U221 ( .A(\temp584[7] ), .B(InEdges[87]), .S(n132), .Z(n776) );
    VMW_MUX2I U222 ( .A(\temp584[6] ), .B(InEdges[86]), .S(n132), .Z(n777) );
    VMW_MUX2I U223 ( .A(\temp584[5] ), .B(InEdges[85]), .S(n132), .Z(n778) );
    VMW_MUX2I U224 ( .A(\temp584[4] ), .B(InEdges[84]), .S(n132), .Z(n779) );
    VMW_MUX2I U225 ( .A(\temp584[3] ), .B(InEdges[83]), .S(n132), .Z(n780) );
    VMW_MUX2I U226 ( .A(\temp584[2] ), .B(InEdges[82]), .S(n132), .Z(n781) );
    VMW_MUX2I U227 ( .A(\temp584[1] ), .B(InEdges[81]), .S(n132), .Z(n782) );
    VMW_MUX2I U228 ( .A(\temp584[14] ), .B(InEdges[94]), .S(n132), .Z(n768) );
    VMW_MUX2I U229 ( .A(\temp584[13] ), .B(InEdges[93]), .S(n132), .Z(n770) );
    VMW_MUX2I U230 ( .A(\temp584[12] ), .B(InEdges[92]), .S(n132), .Z(n771) );
    VMW_MUX2I U231 ( .A(\temp584[11] ), .B(InEdges[91]), .S(n132), .Z(n772) );
    VMW_MUX2I U232 ( .A(\temp584[10] ), .B(InEdges[90]), .S(n132), .Z(n773) );
    VMW_MUX2I U233 ( .A(\temp584[0] ), .B(InEdges[80]), .S(n132), .Z(n783) );
    VMW_INV U234 ( .A(n100), .Z(n792) );
    VMW_INV U235 ( .A(n92), .Z(n794) );
    VMW_INV U236 ( .A(n108), .Z(n793) );
    VMW_INV U237 ( .A(n124), .Z(n790) );
    VMW_INV U238 ( .A(n796), .Z(n810) );
    VMW_BUFIZ U239 ( .A(\path[3] ), .E(n808), .Z(\PathData[3] ) );
    VMW_BUFIZ U240 ( .A(\path[1] ), .E(n808), .Z(\PathData[1] ) );
    VMW_BUFIZ U241 ( .A(\path[0] ), .E(n808), .Z(\PathData[0] ) );
    VMW_BUFIZ U242 ( .A(\path[2] ), .E(n808), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n809), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n810), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n811), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n812), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge146[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge146[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge146[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge146[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge146[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge146[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge146[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge146[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge146[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge146[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge146[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge146[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge146[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge146[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge146[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge146[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_5 lte_55_1 ( .A({\temp220[15] , 
        \temp220[14] , \temp220[13] , \temp220[12] , \temp220[11] , 
        \temp220[10] , \temp220[9] , \temp220[8] , \temp220[7] , \temp220[6] , 
        \temp220[5] , \temp220[4] , \temp220[3] , \temp220[2] , \temp220[1] , 
        \temp220[0] }), .B(InEdges[31:16]), .LEQ(n818), .TC(n818), .GE_GT(n100
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_4 lte_55_5 ( .A({\temp584[15] , 
        \temp584[14] , \temp584[13] , \temp584[12] , \temp584[11] , 
        \temp584[10] , \temp584[9] , \temp584[8] , \temp584[7] , \temp584[6] , 
        \temp584[5] , \temp584[4] , \temp584[3] , \temp584[2] , \temp584[1] , 
        \temp584[0] }), .B(InEdges[95:80]), .LEQ(n817), .TC(n817), .GE_GT(n132
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_3 lte_55_4 ( .A({\temp494[15] , 
        \temp494[14] , \temp494[13] , \temp494[12] , \temp494[11] , 
        \temp494[10] , \temp494[9] , \temp494[8] , \temp494[7] , \temp494[6] , 
        \temp494[5] , \temp494[4] , \temp494[3] , \temp494[2] , \temp494[1] , 
        \temp494[0] }), .B(InEdges[79:64]), .LEQ(n816), .TC(n816), .GE_GT(n124
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_2 lte_55_3 ( .A({\temp404[15] , 
        \temp404[14] , \temp404[13] , \temp404[12] , \temp404[11] , 
        \temp404[10] , \temp404[9] , \temp404[8] , \temp404[7] , \temp404[6] , 
        \temp404[5] , \temp404[4] , \temp404[3] , \temp404[2] , \temp404[1] , 
        \temp404[0] }), .B(InEdges[63:48]), .LEQ(n815), .TC(n815), .GE_GT(n116
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp314[15] , 
        \temp314[14] , \temp314[13] , \temp314[12] , \temp314[11] , 
        \temp314[10] , \temp314[9] , \temp314[8] , \temp314[7] , \temp314[6] , 
        \temp314[5] , \temp314[4] , \temp314[3] , \temp314[2] , \temp314[1] , 
        \temp314[0] }), .B(InEdges[47:32]), .LEQ(n814), .TC(n814), .GE_GT(n108
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n813), .TC(n813), .GE_GT(n92) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_6 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n92, n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, 
        n107, n108, n109, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n93), .C(n91), .D(n89), .Z(n92) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n92), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n99), .D(n97), .Z(n100) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n101) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n107), .D(n101), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n93) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n119, n120, n121, n122, n123, n124, n125, n127, n128, 
        n129, n130, n131, n132, n133, n135, n136, n137, n138, n139, n140, n141, 
        n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
        n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
        n167, n168;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n125), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n132), .D(n127), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n144), .B(B[8]), .Z(n143) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n146), .C(n140), .D(n135), .Z(n145) );
    VMW_OR2 U18 ( .A(B[8]), .B(n144), .Z(n147) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n149), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U20 ( .A(n151), .B(B[10]), .Z(n150) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n153), .C(n148), .D(n143), .Z(n152) );
    VMW_NAND2 U22 ( .A(n153), .B(A[9]), .Z(n154) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n151), .C(n154), .D(n152), .Z(n155) );
    VMW_NAND2 U24 ( .A(n157), .B(B[12]), .Z(n156) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n159), .C(n155), .D(n150), .Z(n158) );
    VMW_NAND2 U26 ( .A(n159), .B(A[11]), .Z(n160) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n157), .C(n160), .D(n158), .Z(n161) );
    VMW_NAND2 U28 ( .A(n163), .B(B[14]), .Z(n162) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n165), .C(n161), .D(n156), .Z(n164) );
    VMW_NAND2 U30 ( .A(n165), .B(A[13]), .Z(n166) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n163), .C(n166), .D(n164), .Z(n167) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n168), .C(n167), .D(n162), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n157) );
    VMW_INV U34 ( .A(B[7]), .Z(n146) );
    VMW_INV U35 ( .A(A[7]), .Z(n149) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n151) );
    VMW_INV U39 ( .A(B[9]), .Z(n153) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n144) );
    VMW_INV U42 ( .A(A[14]), .Z(n163) );
    VMW_INV U43 ( .A(B[11]), .Z(n159) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n168) );
    VMW_INV U48 ( .A(B[13]), .Z(n165) );
    VMW_INV U49 ( .A(A[6]), .Z(n136) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
        n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
        n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
        n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
        n216, n217;
    VMW_OAI21 U3 ( .A(B[15]), .B(n169), .C(n170), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n172), .B(B[2]), .Z(n171) );
    VMW_AO22 U5 ( .A(n174), .B(B[0]), .C(n175), .D(B[1]), .Z(n173) );
    VMW_OR2 U6 ( .A(B[2]), .B(n172), .Z(n176) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n175), .C(n176), .D(n173), .Z(n177) );
    VMW_NAND2 U8 ( .A(n179), .B(B[4]), .Z(n178) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n181), .C(n177), .D(n171), .Z(n180) );
    VMW_OR2 U10 ( .A(B[4]), .B(n179), .Z(n182) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n184), .C(n182), .D(n180), .Z(n183) );
    VMW_NAND2 U12 ( .A(n186), .B(B[6]), .Z(n185) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n188), .C(n183), .D(n178), .Z(n187) );
    VMW_OR2 U14 ( .A(B[6]), .B(n186), .Z(n189) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n191), .C(n189), .D(n187), .Z(n190) );
    VMW_NAND2 U16 ( .A(n193), .B(B[8]), .Z(n192) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n195), .C(n190), .D(n185), .Z(n194) );
    VMW_OR2 U18 ( .A(B[8]), .B(n193), .Z(n196) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n198), .C(n196), .D(n194), .Z(n197) );
    VMW_NAND2 U20 ( .A(n200), .B(B[10]), .Z(n199) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n202), .C(n197), .D(n192), .Z(n201) );
    VMW_NAND2 U22 ( .A(n202), .B(A[9]), .Z(n203) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n200), .C(n203), .D(n201), .Z(n204) );
    VMW_NAND2 U24 ( .A(n206), .B(B[12]), .Z(n205) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n208), .C(n204), .D(n199), .Z(n207) );
    VMW_NAND2 U26 ( .A(n208), .B(A[11]), .Z(n209) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n206), .C(n209), .D(n207), .Z(n210) );
    VMW_NAND2 U28 ( .A(n212), .B(B[14]), .Z(n211) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n214), .C(n210), .D(n205), .Z(n213) );
    VMW_NAND2 U30 ( .A(n214), .B(A[13]), .Z(n215) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n212), .C(n215), .D(n213), .Z(n216) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n217), .C(n216), .D(n211), .Z(n170) );
    VMW_INV U33 ( .A(A[12]), .Z(n206) );
    VMW_INV U34 ( .A(B[7]), .Z(n195) );
    VMW_INV U35 ( .A(A[7]), .Z(n198) );
    VMW_INV U36 ( .A(A[3]), .Z(n184) );
    VMW_INV U37 ( .A(B[3]), .Z(n181) );
    VMW_INV U38 ( .A(A[10]), .Z(n200) );
    VMW_INV U39 ( .A(B[9]), .Z(n202) );
    VMW_INV U40 ( .A(A[4]), .Z(n179) );
    VMW_INV U41 ( .A(A[8]), .Z(n193) );
    VMW_INV U42 ( .A(A[14]), .Z(n212) );
    VMW_INV U43 ( .A(B[11]), .Z(n208) );
    VMW_INV U44 ( .A(A[5]), .Z(n191) );
    VMW_INV U45 ( .A(B[5]), .Z(n188) );
    VMW_INV U46 ( .A(A[1]), .Z(n175) );
    VMW_INV U47 ( .A(B[15]), .Z(n217) );
    VMW_INV U48 ( .A(B[13]), .Z(n214) );
    VMW_INV U49 ( .A(A[6]), .Z(n186) );
    VMW_INV U50 ( .A(A[2]), .Z(n172) );
    VMW_INV U51 ( .A(A[0]), .Z(n174) );
    VMW_INV U52 ( .A(A[15]), .Z(n169) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
        n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
        n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
        n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
        n265, n266;
    VMW_OAI21 U3 ( .A(B[15]), .B(n218), .C(n219), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n221), .B(B[2]), .Z(n220) );
    VMW_AO22 U5 ( .A(n223), .B(B[0]), .C(n224), .D(B[1]), .Z(n222) );
    VMW_OR2 U6 ( .A(B[2]), .B(n221), .Z(n225) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n224), .C(n225), .D(n222), .Z(n226) );
    VMW_NAND2 U8 ( .A(n228), .B(B[4]), .Z(n227) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n230), .C(n226), .D(n220), .Z(n229) );
    VMW_OR2 U10 ( .A(B[4]), .B(n228), .Z(n231) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n233), .C(n231), .D(n229), .Z(n232) );
    VMW_NAND2 U12 ( .A(n235), .B(B[6]), .Z(n234) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n237), .C(n232), .D(n227), .Z(n236) );
    VMW_OR2 U14 ( .A(B[6]), .B(n235), .Z(n238) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n240), .C(n238), .D(n236), .Z(n239) );
    VMW_NAND2 U16 ( .A(n242), .B(B[8]), .Z(n241) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n244), .C(n239), .D(n234), .Z(n243) );
    VMW_OR2 U18 ( .A(B[8]), .B(n242), .Z(n245) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n247), .C(n245), .D(n243), .Z(n246) );
    VMW_NAND2 U20 ( .A(n249), .B(B[10]), .Z(n248) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n251), .C(n246), .D(n241), .Z(n250) );
    VMW_NAND2 U22 ( .A(n251), .B(A[9]), .Z(n252) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n249), .C(n252), .D(n250), .Z(n253) );
    VMW_NAND2 U24 ( .A(n255), .B(B[12]), .Z(n254) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n257), .C(n253), .D(n248), .Z(n256) );
    VMW_NAND2 U26 ( .A(n257), .B(A[11]), .Z(n258) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n255), .C(n258), .D(n256), .Z(n259) );
    VMW_NAND2 U28 ( .A(n261), .B(B[14]), .Z(n260) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n263), .C(n259), .D(n254), .Z(n262) );
    VMW_NAND2 U30 ( .A(n263), .B(A[13]), .Z(n264) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n261), .C(n264), .D(n262), .Z(n265) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n266), .C(n265), .D(n260), .Z(n219) );
    VMW_INV U33 ( .A(A[12]), .Z(n255) );
    VMW_INV U34 ( .A(B[7]), .Z(n244) );
    VMW_INV U35 ( .A(A[7]), .Z(n247) );
    VMW_INV U36 ( .A(A[3]), .Z(n233) );
    VMW_INV U37 ( .A(B[3]), .Z(n230) );
    VMW_INV U38 ( .A(A[10]), .Z(n249) );
    VMW_INV U39 ( .A(B[9]), .Z(n251) );
    VMW_INV U40 ( .A(A[4]), .Z(n228) );
    VMW_INV U41 ( .A(A[8]), .Z(n242) );
    VMW_INV U42 ( .A(A[14]), .Z(n261) );
    VMW_INV U43 ( .A(B[11]), .Z(n257) );
    VMW_INV U44 ( .A(A[5]), .Z(n240) );
    VMW_INV U45 ( .A(B[5]), .Z(n237) );
    VMW_INV U46 ( .A(A[1]), .Z(n224) );
    VMW_INV U47 ( .A(B[15]), .Z(n266) );
    VMW_INV U48 ( .A(B[13]), .Z(n263) );
    VMW_INV U49 ( .A(A[6]), .Z(n235) );
    VMW_INV U50 ( .A(A[2]), .Z(n221) );
    VMW_INV U51 ( .A(A[0]), .Z(n223) );
    VMW_INV U52 ( .A(A[15]), .Z(n218) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315;
    VMW_OAI21 U3 ( .A(B[15]), .B(n267), .C(n268), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n270), .B(B[2]), .Z(n269) );
    VMW_AO22 U5 ( .A(n272), .B(B[0]), .C(n273), .D(B[1]), .Z(n271) );
    VMW_OR2 U6 ( .A(B[2]), .B(n270), .Z(n274) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n273), .C(n274), .D(n271), .Z(n275) );
    VMW_NAND2 U8 ( .A(n277), .B(B[4]), .Z(n276) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n279), .C(n275), .D(n269), .Z(n278) );
    VMW_OR2 U10 ( .A(B[4]), .B(n277), .Z(n280) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n282), .C(n280), .D(n278), .Z(n281) );
    VMW_NAND2 U12 ( .A(n284), .B(B[6]), .Z(n283) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n286), .C(n281), .D(n276), .Z(n285) );
    VMW_OR2 U14 ( .A(B[6]), .B(n284), .Z(n287) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n289), .C(n287), .D(n285), .Z(n288) );
    VMW_NAND2 U16 ( .A(n291), .B(B[8]), .Z(n290) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n293), .C(n288), .D(n283), .Z(n292) );
    VMW_OR2 U18 ( .A(B[8]), .B(n291), .Z(n294) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n296), .C(n294), .D(n292), .Z(n295) );
    VMW_NAND2 U20 ( .A(n298), .B(B[10]), .Z(n297) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n300), .C(n295), .D(n290), .Z(n299) );
    VMW_NAND2 U22 ( .A(n300), .B(A[9]), .Z(n301) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n298), .C(n301), .D(n299), .Z(n302) );
    VMW_NAND2 U24 ( .A(n304), .B(B[12]), .Z(n303) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n306), .C(n302), .D(n297), .Z(n305) );
    VMW_NAND2 U26 ( .A(n306), .B(A[11]), .Z(n307) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n304), .C(n307), .D(n305), .Z(n308) );
    VMW_NAND2 U28 ( .A(n310), .B(B[14]), .Z(n309) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n312), .C(n308), .D(n303), .Z(n311) );
    VMW_NAND2 U30 ( .A(n312), .B(A[13]), .Z(n313) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n310), .C(n313), .D(n311), .Z(n314) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n315), .C(n314), .D(n309), .Z(n268) );
    VMW_INV U33 ( .A(A[12]), .Z(n304) );
    VMW_INV U34 ( .A(B[7]), .Z(n293) );
    VMW_INV U35 ( .A(A[7]), .Z(n296) );
    VMW_INV U36 ( .A(A[3]), .Z(n282) );
    VMW_INV U37 ( .A(B[3]), .Z(n279) );
    VMW_INV U38 ( .A(A[10]), .Z(n298) );
    VMW_INV U39 ( .A(B[9]), .Z(n300) );
    VMW_INV U40 ( .A(A[4]), .Z(n277) );
    VMW_INV U41 ( .A(A[8]), .Z(n291) );
    VMW_INV U42 ( .A(A[14]), .Z(n310) );
    VMW_INV U43 ( .A(B[11]), .Z(n306) );
    VMW_INV U44 ( .A(A[5]), .Z(n289) );
    VMW_INV U45 ( .A(B[5]), .Z(n286) );
    VMW_INV U46 ( .A(A[1]), .Z(n273) );
    VMW_INV U47 ( .A(B[15]), .Z(n315) );
    VMW_INV U48 ( .A(B[13]), .Z(n312) );
    VMW_INV U49 ( .A(A[6]), .Z(n284) );
    VMW_INV U50 ( .A(A[2]), .Z(n270) );
    VMW_INV U51 ( .A(A[0]), .Z(n272) );
    VMW_INV U52 ( .A(A[15]), .Z(n267) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
        n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, 
        n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
        n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
        n363, n364;
    VMW_OAI21 U3 ( .A(B[15]), .B(n316), .C(n317), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n319), .B(B[2]), .Z(n318) );
    VMW_AO22 U5 ( .A(n321), .B(B[0]), .C(n322), .D(B[1]), .Z(n320) );
    VMW_OR2 U6 ( .A(B[2]), .B(n319), .Z(n323) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n322), .C(n323), .D(n320), .Z(n324) );
    VMW_NAND2 U8 ( .A(n326), .B(B[4]), .Z(n325) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n328), .C(n324), .D(n318), .Z(n327) );
    VMW_OR2 U10 ( .A(B[4]), .B(n326), .Z(n329) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n331), .C(n329), .D(n327), .Z(n330) );
    VMW_NAND2 U12 ( .A(n333), .B(B[6]), .Z(n332) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n335), .C(n330), .D(n325), .Z(n334) );
    VMW_OR2 U14 ( .A(B[6]), .B(n333), .Z(n336) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n338), .C(n336), .D(n334), .Z(n337) );
    VMW_NAND2 U16 ( .A(n340), .B(B[8]), .Z(n339) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n342), .C(n337), .D(n332), .Z(n341) );
    VMW_OR2 U18 ( .A(B[8]), .B(n340), .Z(n343) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n345), .C(n343), .D(n341), .Z(n344) );
    VMW_NAND2 U20 ( .A(n347), .B(B[10]), .Z(n346) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n349), .C(n344), .D(n339), .Z(n348) );
    VMW_NAND2 U22 ( .A(n349), .B(A[9]), .Z(n350) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n347), .C(n350), .D(n348), .Z(n351) );
    VMW_NAND2 U24 ( .A(n353), .B(B[12]), .Z(n352) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n355), .C(n351), .D(n346), .Z(n354) );
    VMW_NAND2 U26 ( .A(n355), .B(A[11]), .Z(n356) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n353), .C(n356), .D(n354), .Z(n357) );
    VMW_NAND2 U28 ( .A(n359), .B(B[14]), .Z(n358) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n361), .C(n357), .D(n352), .Z(n360) );
    VMW_NAND2 U30 ( .A(n361), .B(A[13]), .Z(n362) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n359), .C(n362), .D(n360), .Z(n363) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n364), .C(n363), .D(n358), .Z(n317) );
    VMW_INV U33 ( .A(A[12]), .Z(n353) );
    VMW_INV U34 ( .A(B[7]), .Z(n342) );
    VMW_INV U35 ( .A(A[7]), .Z(n345) );
    VMW_INV U36 ( .A(A[3]), .Z(n331) );
    VMW_INV U37 ( .A(B[3]), .Z(n328) );
    VMW_INV U38 ( .A(A[10]), .Z(n347) );
    VMW_INV U39 ( .A(B[9]), .Z(n349) );
    VMW_INV U40 ( .A(A[4]), .Z(n326) );
    VMW_INV U41 ( .A(A[8]), .Z(n340) );
    VMW_INV U42 ( .A(A[14]), .Z(n359) );
    VMW_INV U43 ( .A(B[11]), .Z(n355) );
    VMW_INV U44 ( .A(A[5]), .Z(n338) );
    VMW_INV U45 ( .A(B[5]), .Z(n335) );
    VMW_INV U46 ( .A(A[1]), .Z(n322) );
    VMW_INV U47 ( .A(B[15]), .Z(n364) );
    VMW_INV U48 ( .A(B[13]), .Z(n361) );
    VMW_INV U49 ( .A(A[6]), .Z(n333) );
    VMW_INV U50 ( .A(A[2]), .Z(n319) );
    VMW_INV U51 ( .A(A[0]), .Z(n321) );
    VMW_INV U52 ( .A(A[15]), .Z(n316) );
endmodule


module NodeAux_INDEGREE7_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \OutEdge156[4] , \temp324[9] , \temp594[1] , \temp324[0] , 
        \temp594[8] , \OutEdge156[10] , \OutEdge156[0] , \temp594[5] , 
        \temp684[12] , \OutEdge156[14] , \path[2] , \OutEdge156[9] , 
        \temp324[4] , \path[0] , \temp324[6] , \temp684[10] , \temp594[7] , 
        \OutEdge156[2] , \OutEdge156[12] , \temp324[2] , \OutEdge156[6] , 
        \temp594[3] , \temp684[14] , \temp504[15] , \temp684[8] , \temp504[9] , 
        \temp414[5] , \temp230[7] , \temp504[0] , \temp594[15] , \temp684[1] , 
        \temp414[13] , \temp414[8] , \temp504[11] , \temp684[5] , 
        \temp594[11] , \temp324[12] , \temp230[3] , \temp504[4] , \temp414[1] , 
        \temp230[12] , \temp230[1] , \temp504[6] , \temp414[3] , \temp230[10] , 
        n126, \temp594[13] , \temp684[7] , \temp324[10] , \temp504[13] , 
        \temp230[8] , \temp414[11] , \temp324[14] , \temp684[3] , 
        \temp230[14] , \temp414[7] , \temp230[5] , \temp504[2] , \temp414[15] , 
        n134, \temp324[15] , n118, \temp684[2] , \temp414[6] , \temp230[15] , 
        n94, \temp504[3] , \temp230[4] , \temp414[14] , \temp230[0] , 
        \temp504[7] , \temp230[11] , \temp414[2] , \temp684[6] , \temp594[12] , 
        \temp324[11] , \temp504[12] , \temp230[9] , \temp414[10] , 
        \temp414[9] , \temp414[12] , \temp504[10] , \temp684[4] , 
        \temp594[10] , \temp324[13] , \temp230[2] , \temp504[5] , 
        \temp230[13] , \temp414[0] , \temp504[14] , \temp684[9] , \temp504[8] , 
        \temp414[4] , \temp230[6] , \temp504[1] , \temp684[0] , \temp594[14] , 
        \OutEdge156[13] , \temp324[3] , \OutEdge156[7] , \temp594[2] , 
        \temp684[15] , \temp324[7] , \path[1] , \temp684[11] , \temp594[6] , 
        \OutEdge156[3] , n102, \temp594[4] , \OutEdge156[1] , \temp684[13] , 
        \OutEdge156[15] , \temp324[5] , \path[3] , \OutEdge156[8] , 
        \OutEdge156[5] , n142, \temp324[8] , \temp594[0] , \OutEdge156[11] , 
        \temp594[9] , \temp324[1] , n110, n867, n868, n869, n870, n871, n872, 
        n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
        n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
        n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
        n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
        n921, n922;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U100 ( .Z(n918) );
    VMW_PULLDOWN U101 ( .Z(n922) );
    VMW_PULLDOWN U102 ( .Z(n920) );
    VMW_PULLDOWN U103 ( .Z(n921) );
    VMW_PULLDOWN U104 ( .Z(n917) );
    VMW_PULLDOWN U105 ( .Z(n916) );
    VMW_PULLDOWN U106 ( .Z(n919) );
    VMW_AO21 U107 ( .A(\temp684[15] ), .B(n867), .C(n868), .Z(\OutEdge156[15] 
        ) );
    VMW_NAND2 U108 ( .A(n869), .B(n870), .Z(\OutEdge156[14] ) );
    VMW_NAND2 U109 ( .A(n871), .B(n870), .Z(\OutEdge156[13] ) );
    VMW_NAND2 U110 ( .A(n872), .B(n870), .Z(\OutEdge156[12] ) );
    VMW_NAND2 U111 ( .A(n873), .B(n870), .Z(\OutEdge156[11] ) );
    VMW_NAND2 U112 ( .A(n874), .B(n870), .Z(\OutEdge156[10] ) );
    VMW_NAND2 U113 ( .A(n875), .B(n870), .Z(\OutEdge156[9] ) );
    VMW_NAND2 U114 ( .A(n876), .B(n870), .Z(\OutEdge156[8] ) );
    VMW_NAND2 U115 ( .A(n877), .B(n870), .Z(\OutEdge156[7] ) );
    VMW_NAND2 U116 ( .A(n878), .B(n870), .Z(\OutEdge156[6] ) );
    VMW_NAND2 U117 ( .A(n879), .B(n870), .Z(\OutEdge156[5] ) );
    VMW_NAND2 U118 ( .A(n880), .B(n870), .Z(\OutEdge156[4] ) );
    VMW_NAND2 U119 ( .A(n881), .B(n870), .Z(\OutEdge156[3] ) );
    VMW_NAND2 U120 ( .A(n882), .B(n870), .Z(\OutEdge156[2] ) );
    VMW_NAND2 U121 ( .A(n883), .B(n870), .Z(\OutEdge156[1] ) );
    VMW_NAND2 U122 ( .A(n884), .B(n870), .Z(\OutEdge156[0] ) );
    VMW_AO21 U123 ( .A(Start), .B(\path[3] ), .C(n885), .Z(n914) );
    VMW_AO22 U124 ( .A(\path[0] ), .B(Start), .C(n867), .D(n886), .Z(n912) );
    VMW_AND4 U125 ( .A(n887), .B(n888), .C(n867), .D(n889), .Z(n885) );
    VMW_OR4 U126 ( .A(n142), .B(n126), .C(n134), .D(n889), .Z(n890) );
    VMW_AND3 U127 ( .A(n888), .B(n887), .C(n892), .Z(n891) );
    VMW_OR2 U128 ( .A(n891), .B(n142), .Z(n893) );
    VMW_AO22 U129 ( .A(\temp594[15] ), .B(n888), .C(InEdges[95]), .D(n134), 
        .Z(\temp684[15] ) );
    VMW_NOR2 U130 ( .A(Start), .B(n142), .Z(n867) );
    VMW_AND4 U131 ( .A(n894), .B(n895), .C(n896), .D(n897), .Z(n889) );
    VMW_INV U132 ( .A(Start), .Z(n870) );
    VMW_OAI22 U133 ( .A(\path[2] ), .B(n870), .C(n890), .D(Start), .Z(n898) );
    VMW_OAI22 U134 ( .A(\path[1] ), .B(n870), .C(n893), .D(Start), .Z(n899) );
    VMW_AND4 U135 ( .A(n901), .B(n902), .C(n903), .D(n904), .Z(n900) );
    VMW_INV U136 ( .A(n118), .Z(n897) );
    VMW_INV U137 ( .A(n110), .Z(n895) );
    VMW_INV U138 ( .A(n126), .Z(n887) );
    VMW_INV U139 ( .A(n134), .Z(n888) );
    VMW_OAI211 U140 ( .A(n94), .B(n102), .C(n895), .D(n897), .Z(n892) );
    VMW_AO21 U141 ( .A(n894), .B(n94), .C(n110), .Z(n905) );
    VMW_AO21 U142 ( .A(n897), .B(n905), .C(n126), .Z(n906) );
    VMW_NAND2 U143 ( .A(n888), .B(n906), .Z(n886) );
    VMW_AND5 U144 ( .A(n907), .B(n908), .C(n909), .D(n910), .E(n900), .Z(n911)
         );
    VMW_AND3 U145 ( .A(n142), .B(n870), .C(InEdges[111]), .Z(n868) );
    VMW_XNOR2 U146 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n904) );
    VMW_XNOR2 U147 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n903) );
    VMW_XNOR2 U148 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n902) );
    VMW_XNOR2 U149 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n901) );
    VMW_XNOR2 U150 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n910) );
    VMW_XNOR2 U151 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n909) );
    VMW_XNOR2 U152 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n908) );
    VMW_XNOR2 U153 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n907) );
    VMW_AO22 U154 ( .A(OutEdge[9]), .B(n896), .C(InEdges[9]), .D(n94), .Z(
        \temp230[9] ) );
    VMW_AO22 U155 ( .A(\temp230[9] ), .B(n894), .C(InEdges[25]), .D(n102), .Z(
        \temp324[9] ) );
    VMW_AO22 U156 ( .A(\temp324[9] ), .B(n895), .C(InEdges[41]), .D(n110), .Z(
        \temp414[9] ) );
    VMW_AO22 U157 ( .A(\temp414[9] ), .B(n897), .C(InEdges[57]), .D(n118), .Z(
        \temp504[9] ) );
    VMW_AO22 U158 ( .A(\temp504[9] ), .B(n887), .C(InEdges[73]), .D(n126), .Z(
        \temp594[9] ) );
    VMW_AO22 U159 ( .A(\temp594[9] ), .B(n888), .C(InEdges[89]), .D(n134), .Z(
        \temp684[9] ) );
    VMW_AO22 U160 ( .A(OutEdge[8]), .B(n896), .C(InEdges[8]), .D(n94), .Z(
        \temp230[8] ) );
    VMW_AO22 U161 ( .A(\temp230[8] ), .B(n894), .C(InEdges[24]), .D(n102), .Z(
        \temp324[8] ) );
    VMW_AO22 U162 ( .A(\temp324[8] ), .B(n895), .C(InEdges[40]), .D(n110), .Z(
        \temp414[8] ) );
    VMW_AO22 U163 ( .A(\temp414[8] ), .B(n897), .C(InEdges[56]), .D(n118), .Z(
        \temp504[8] ) );
    VMW_AO22 U164 ( .A(\temp504[8] ), .B(n887), .C(InEdges[72]), .D(n126), .Z(
        \temp594[8] ) );
    VMW_AO22 U165 ( .A(\temp594[8] ), .B(n888), .C(InEdges[88]), .D(n134), .Z(
        \temp684[8] ) );
    VMW_AO22 U166 ( .A(OutEdge[7]), .B(n896), .C(InEdges[7]), .D(n94), .Z(
        \temp230[7] ) );
    VMW_AO22 U167 ( .A(\temp230[7] ), .B(n894), .C(InEdges[23]), .D(n102), .Z(
        \temp324[7] ) );
    VMW_AO22 U168 ( .A(\temp324[7] ), .B(n895), .C(InEdges[39]), .D(n110), .Z(
        \temp414[7] ) );
    VMW_AO22 U169 ( .A(\temp414[7] ), .B(n897), .C(InEdges[55]), .D(n118), .Z(
        \temp504[7] ) );
    VMW_AO22 U170 ( .A(\temp504[7] ), .B(n887), .C(InEdges[71]), .D(n126), .Z(
        \temp594[7] ) );
    VMW_AO22 U171 ( .A(\temp594[7] ), .B(n888), .C(InEdges[87]), .D(n134), .Z(
        \temp684[7] ) );
    VMW_AO22 U172 ( .A(OutEdge[6]), .B(n896), .C(InEdges[6]), .D(n94), .Z(
        \temp230[6] ) );
    VMW_AO22 U173 ( .A(\temp230[6] ), .B(n894), .C(InEdges[22]), .D(n102), .Z(
        \temp324[6] ) );
    VMW_AO22 U174 ( .A(\temp324[6] ), .B(n895), .C(InEdges[38]), .D(n110), .Z(
        \temp414[6] ) );
    VMW_AO22 U175 ( .A(\temp414[6] ), .B(n897), .C(InEdges[54]), .D(n118), .Z(
        \temp504[6] ) );
    VMW_AO22 U176 ( .A(\temp504[6] ), .B(n887), .C(InEdges[70]), .D(n126), .Z(
        \temp594[6] ) );
    VMW_AO22 U177 ( .A(\temp594[6] ), .B(n888), .C(InEdges[86]), .D(n134), .Z(
        \temp684[6] ) );
    VMW_AO22 U178 ( .A(OutEdge[5]), .B(n896), .C(InEdges[5]), .D(n94), .Z(
        \temp230[5] ) );
    VMW_AO22 U179 ( .A(\temp230[5] ), .B(n894), .C(InEdges[21]), .D(n102), .Z(
        \temp324[5] ) );
    VMW_AO22 U180 ( .A(\temp324[5] ), .B(n895), .C(InEdges[37]), .D(n110), .Z(
        \temp414[5] ) );
    VMW_AO22 U181 ( .A(\temp414[5] ), .B(n897), .C(InEdges[53]), .D(n118), .Z(
        \temp504[5] ) );
    VMW_AO22 U182 ( .A(\temp504[5] ), .B(n887), .C(InEdges[69]), .D(n126), .Z(
        \temp594[5] ) );
    VMW_AO22 U183 ( .A(\temp594[5] ), .B(n888), .C(InEdges[85]), .D(n134), .Z(
        \temp684[5] ) );
    VMW_AO22 U184 ( .A(OutEdge[4]), .B(n896), .C(InEdges[4]), .D(n94), .Z(
        \temp230[4] ) );
    VMW_AO22 U185 ( .A(\temp230[4] ), .B(n894), .C(InEdges[20]), .D(n102), .Z(
        \temp324[4] ) );
    VMW_AO22 U186 ( .A(\temp324[4] ), .B(n895), .C(InEdges[36]), .D(n110), .Z(
        \temp414[4] ) );
    VMW_AO22 U187 ( .A(\temp414[4] ), .B(n897), .C(InEdges[52]), .D(n118), .Z(
        \temp504[4] ) );
    VMW_AO22 U188 ( .A(\temp504[4] ), .B(n887), .C(InEdges[68]), .D(n126), .Z(
        \temp594[4] ) );
    VMW_AO22 U189 ( .A(\temp594[4] ), .B(n888), .C(InEdges[84]), .D(n134), .Z(
        \temp684[4] ) );
    VMW_AO22 U190 ( .A(OutEdge[3]), .B(n896), .C(InEdges[3]), .D(n94), .Z(
        \temp230[3] ) );
    VMW_AO22 U191 ( .A(\temp230[3] ), .B(n894), .C(InEdges[19]), .D(n102), .Z(
        \temp324[3] ) );
    VMW_AO22 U192 ( .A(\temp324[3] ), .B(n895), .C(InEdges[35]), .D(n110), .Z(
        \temp414[3] ) );
    VMW_AO22 U193 ( .A(\temp414[3] ), .B(n897), .C(InEdges[51]), .D(n118), .Z(
        \temp504[3] ) );
    VMW_AO22 U194 ( .A(\temp504[3] ), .B(n887), .C(InEdges[67]), .D(n126), .Z(
        \temp594[3] ) );
    VMW_AO22 U195 ( .A(\temp594[3] ), .B(n888), .C(InEdges[83]), .D(n134), .Z(
        \temp684[3] ) );
    VMW_AO22 U196 ( .A(OutEdge[2]), .B(n896), .C(InEdges[2]), .D(n94), .Z(
        \temp230[2] ) );
    VMW_AO22 U197 ( .A(\temp230[2] ), .B(n894), .C(InEdges[18]), .D(n102), .Z(
        \temp324[2] ) );
    VMW_AO22 U198 ( .A(\temp324[2] ), .B(n895), .C(InEdges[34]), .D(n110), .Z(
        \temp414[2] ) );
    VMW_AO22 U199 ( .A(\temp414[2] ), .B(n897), .C(InEdges[50]), .D(n118), .Z(
        \temp504[2] ) );
    VMW_AO22 U200 ( .A(\temp504[2] ), .B(n887), .C(InEdges[66]), .D(n126), .Z(
        \temp594[2] ) );
    VMW_AO22 U201 ( .A(\temp594[2] ), .B(n888), .C(InEdges[82]), .D(n134), .Z(
        \temp684[2] ) );
    VMW_AO22 U202 ( .A(OutEdge[1]), .B(n896), .C(InEdges[1]), .D(n94), .Z(
        \temp230[1] ) );
    VMW_AO22 U203 ( .A(\temp230[1] ), .B(n894), .C(InEdges[17]), .D(n102), .Z(
        \temp324[1] ) );
    VMW_AO22 U204 ( .A(\temp324[1] ), .B(n895), .C(InEdges[33]), .D(n110), .Z(
        \temp414[1] ) );
    VMW_AO22 U205 ( .A(\temp414[1] ), .B(n897), .C(InEdges[49]), .D(n118), .Z(
        \temp504[1] ) );
    VMW_AO22 U206 ( .A(\temp504[1] ), .B(n887), .C(InEdges[65]), .D(n126), .Z(
        \temp594[1] ) );
    VMW_AO22 U207 ( .A(\temp594[1] ), .B(n888), .C(InEdges[81]), .D(n134), .Z(
        \temp684[1] ) );
    VMW_AO22 U208 ( .A(OutEdge[15]), .B(n896), .C(InEdges[15]), .D(n94), .Z(
        \temp230[15] ) );
    VMW_AO22 U209 ( .A(\temp230[15] ), .B(n894), .C(InEdges[31]), .D(n102), 
        .Z(\temp324[15] ) );
    VMW_AO22 U210 ( .A(\temp324[15] ), .B(n895), .C(InEdges[47]), .D(n110), 
        .Z(\temp414[15] ) );
    VMW_AO22 U211 ( .A(\temp414[15] ), .B(n897), .C(InEdges[63]), .D(n118), 
        .Z(\temp504[15] ) );
    VMW_AO22 U212 ( .A(\temp504[15] ), .B(n887), .C(InEdges[79]), .D(n126), 
        .Z(\temp594[15] ) );
    VMW_AO22 U213 ( .A(OutEdge[14]), .B(n896), .C(InEdges[14]), .D(n94), .Z(
        \temp230[14] ) );
    VMW_AO22 U214 ( .A(\temp230[14] ), .B(n894), .C(InEdges[30]), .D(n102), 
        .Z(\temp324[14] ) );
    VMW_AO22 U215 ( .A(\temp324[14] ), .B(n895), .C(InEdges[46]), .D(n110), 
        .Z(\temp414[14] ) );
    VMW_AO22 U216 ( .A(\temp414[14] ), .B(n897), .C(InEdges[62]), .D(n118), 
        .Z(\temp504[14] ) );
    VMW_AO22 U217 ( .A(\temp504[14] ), .B(n887), .C(InEdges[78]), .D(n126), 
        .Z(\temp594[14] ) );
    VMW_AO22 U218 ( .A(\temp594[14] ), .B(n888), .C(InEdges[94]), .D(n134), 
        .Z(\temp684[14] ) );
    VMW_AO22 U219 ( .A(OutEdge[13]), .B(n896), .C(InEdges[13]), .D(n94), .Z(
        \temp230[13] ) );
    VMW_AO22 U220 ( .A(\temp230[13] ), .B(n894), .C(InEdges[29]), .D(n102), 
        .Z(\temp324[13] ) );
    VMW_AO22 U221 ( .A(\temp324[13] ), .B(n895), .C(InEdges[45]), .D(n110), 
        .Z(\temp414[13] ) );
    VMW_AO22 U222 ( .A(\temp414[13] ), .B(n897), .C(InEdges[61]), .D(n118), 
        .Z(\temp504[13] ) );
    VMW_AO22 U223 ( .A(\temp504[13] ), .B(n887), .C(InEdges[77]), .D(n126), 
        .Z(\temp594[13] ) );
    VMW_AO22 U224 ( .A(\temp594[13] ), .B(n888), .C(InEdges[93]), .D(n134), 
        .Z(\temp684[13] ) );
    VMW_AO22 U225 ( .A(OutEdge[12]), .B(n896), .C(InEdges[12]), .D(n94), .Z(
        \temp230[12] ) );
    VMW_AO22 U226 ( .A(\temp230[12] ), .B(n894), .C(InEdges[28]), .D(n102), 
        .Z(\temp324[12] ) );
    VMW_AO22 U227 ( .A(\temp324[12] ), .B(n895), .C(InEdges[44]), .D(n110), 
        .Z(\temp414[12] ) );
    VMW_AO22 U228 ( .A(\temp414[12] ), .B(n897), .C(InEdges[60]), .D(n118), 
        .Z(\temp504[12] ) );
    VMW_AO22 U229 ( .A(\temp504[12] ), .B(n887), .C(InEdges[76]), .D(n126), 
        .Z(\temp594[12] ) );
    VMW_AO22 U230 ( .A(\temp594[12] ), .B(n888), .C(InEdges[92]), .D(n134), 
        .Z(\temp684[12] ) );
    VMW_AO22 U231 ( .A(OutEdge[11]), .B(n896), .C(InEdges[11]), .D(n94), .Z(
        \temp230[11] ) );
    VMW_AO22 U232 ( .A(\temp230[11] ), .B(n894), .C(InEdges[27]), .D(n102), 
        .Z(\temp324[11] ) );
    VMW_AO22 U233 ( .A(\temp324[11] ), .B(n895), .C(InEdges[43]), .D(n110), 
        .Z(\temp414[11] ) );
    VMW_AO22 U234 ( .A(\temp414[11] ), .B(n897), .C(InEdges[59]), .D(n118), 
        .Z(\temp504[11] ) );
    VMW_AO22 U235 ( .A(\temp504[11] ), .B(n887), .C(InEdges[75]), .D(n126), 
        .Z(\temp594[11] ) );
    VMW_AO22 U236 ( .A(\temp594[11] ), .B(n888), .C(InEdges[91]), .D(n134), 
        .Z(\temp684[11] ) );
    VMW_AO22 U237 ( .A(OutEdge[10]), .B(n896), .C(InEdges[10]), .D(n94), .Z(
        \temp230[10] ) );
    VMW_AO22 U238 ( .A(\temp230[10] ), .B(n894), .C(InEdges[26]), .D(n102), 
        .Z(\temp324[10] ) );
    VMW_AO22 U239 ( .A(\temp324[10] ), .B(n895), .C(InEdges[42]), .D(n110), 
        .Z(\temp414[10] ) );
    VMW_AO22 U240 ( .A(\temp414[10] ), .B(n897), .C(InEdges[58]), .D(n118), 
        .Z(\temp504[10] ) );
    VMW_AO22 U241 ( .A(\temp504[10] ), .B(n887), .C(InEdges[74]), .D(n126), 
        .Z(\temp594[10] ) );
    VMW_AO22 U242 ( .A(\temp594[10] ), .B(n888), .C(InEdges[90]), .D(n134), 
        .Z(\temp684[10] ) );
    VMW_AO22 U243 ( .A(OutEdge[0]), .B(n896), .C(InEdges[0]), .D(n94), .Z(
        \temp230[0] ) );
    VMW_AO22 U244 ( .A(\temp230[0] ), .B(n894), .C(InEdges[16]), .D(n102), .Z(
        \temp324[0] ) );
    VMW_AO22 U245 ( .A(\temp324[0] ), .B(n895), .C(InEdges[32]), .D(n110), .Z(
        \temp414[0] ) );
    VMW_AO22 U246 ( .A(\temp414[0] ), .B(n897), .C(InEdges[48]), .D(n118), .Z(
        \temp504[0] ) );
    VMW_AO22 U247 ( .A(\temp504[0] ), .B(n887), .C(InEdges[64]), .D(n126), .Z(
        \temp594[0] ) );
    VMW_AO22 U248 ( .A(\temp594[0] ), .B(n888), .C(InEdges[80]), .D(n134), .Z(
        \temp684[0] ) );
    VMW_MUX2I U249 ( .A(\temp684[9] ), .B(InEdges[105]), .S(n142), .Z(n875) );
    VMW_MUX2I U250 ( .A(\temp684[8] ), .B(InEdges[104]), .S(n142), .Z(n876) );
    VMW_MUX2I U251 ( .A(\temp684[7] ), .B(InEdges[103]), .S(n142), .Z(n877) );
    VMW_MUX2I U252 ( .A(\temp684[6] ), .B(InEdges[102]), .S(n142), .Z(n878) );
    VMW_MUX2I U253 ( .A(\temp684[5] ), .B(InEdges[101]), .S(n142), .Z(n879) );
    VMW_MUX2I U254 ( .A(\temp684[4] ), .B(InEdges[100]), .S(n142), .Z(n880) );
    VMW_MUX2I U255 ( .A(\temp684[3] ), .B(InEdges[99]), .S(n142), .Z(n881) );
    VMW_MUX2I U256 ( .A(\temp684[2] ), .B(InEdges[98]), .S(n142), .Z(n882) );
    VMW_MUX2I U257 ( .A(\temp684[1] ), .B(InEdges[97]), .S(n142), .Z(n883) );
    VMW_MUX2I U258 ( .A(\temp684[14] ), .B(InEdges[110]), .S(n142), .Z(n869)
         );
    VMW_MUX2I U259 ( .A(\temp684[13] ), .B(InEdges[109]), .S(n142), .Z(n871)
         );
    VMW_MUX2I U260 ( .A(\temp684[12] ), .B(InEdges[108]), .S(n142), .Z(n872)
         );
    VMW_MUX2I U261 ( .A(\temp684[11] ), .B(InEdges[107]), .S(n142), .Z(n873)
         );
    VMW_MUX2I U262 ( .A(\temp684[10] ), .B(InEdges[106]), .S(n142), .Z(n874)
         );
    VMW_MUX2I U263 ( .A(\temp684[0] ), .B(InEdges[96]), .S(n142), .Z(n884) );
    VMW_INV U264 ( .A(n94), .Z(n896) );
    VMW_INV U265 ( .A(n102), .Z(n894) );
    VMW_INV U266 ( .A(n898), .Z(n913) );
    VMW_INV U267 ( .A(n899), .Z(n915) );
    VMW_BUFIZ U268 ( .A(\path[3] ), .E(n911), .Z(\PathData[3] ) );
    VMW_BUFIZ U269 ( .A(\path[1] ), .E(n911), .Z(\PathData[1] ) );
    VMW_BUFIZ U270 ( .A(\path[0] ), .E(n911), .Z(\PathData[0] ) );
    VMW_BUFIZ U271 ( .A(\path[2] ), .E(n911), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n912), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n913), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n914), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n915), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge156[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge156[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge156[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge156[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge156[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge156[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge156[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge156[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge156[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge156[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge156[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge156[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge156[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge156[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge156[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge156[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_6 lte_55_5 ( .A({\temp594[15] , 
        \temp594[14] , \temp594[13] , \temp594[12] , \temp594[11] , 
        \temp594[10] , \temp594[9] , \temp594[8] , \temp594[7] , \temp594[6] , 
        \temp594[5] , \temp594[4] , \temp594[3] , \temp594[2] , \temp594[1] , 
        \temp594[0] }), .B(InEdges[95:80]), .LEQ(n922), .TC(n922), .GE_GT(n134
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_5 lte_55_3 ( .A({\temp414[15] , 
        \temp414[14] , \temp414[13] , \temp414[12] , \temp414[11] , 
        \temp414[10] , \temp414[9] , \temp414[8] , \temp414[7] , \temp414[6] , 
        \temp414[5] , \temp414[4] , \temp414[3] , \temp414[2] , \temp414[1] , 
        \temp414[0] }), .B(InEdges[63:48]), .LEQ(n921), .TC(n921), .GE_GT(n118
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_4 lte_55_4 ( .A({\temp504[15] , 
        \temp504[14] , \temp504[13] , \temp504[12] , \temp504[11] , 
        \temp504[10] , \temp504[9] , \temp504[8] , \temp504[7] , \temp504[6] , 
        \temp504[5] , \temp504[4] , \temp504[3] , \temp504[2] , \temp504[1] , 
        \temp504[0] }), .B(InEdges[79:64]), .LEQ(n920), .TC(n920), .GE_GT(n126
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_3 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n919), .TC(n919), .GE_GT(n94) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_2 lte_55_6 ( .A({\temp684[15] , 
        \temp684[14] , \temp684[13] , \temp684[12] , \temp684[11] , 
        \temp684[10] , \temp684[9] , \temp684[8] , \temp684[7] , \temp684[6] , 
        \temp684[5] , \temp684[4] , \temp684[3] , \temp684[2] , \temp684[1] , 
        \temp684[0] }), .B(InEdges[111:96]), .LEQ(n918), .TC(n918), .GE_GT(
        n142) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp324[15] , 
        \temp324[14] , \temp324[13] , \temp324[12] , \temp324[11] , 
        \temp324[10] , \temp324[9] , \temp324[8] , \temp324[7] , \temp324[6] , 
        \temp324[5] , \temp324[4] , \temp324[3] , \temp324[2] , \temp324[1] , 
        \temp324[0] }), .B(InEdges[47:32]), .LEQ(n917), .TC(n917), .GE_GT(n110
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_0 lte_55_1 ( .A({\temp230[15] , 
        \temp230[14] , \temp230[13] , \temp230[12] , \temp230[11] , 
        \temp230[10] , \temp230[9] , \temp230[8] , \temp230[7] , \temp230[6] , 
        \temp230[5] , \temp230[4] , \temp230[3] , \temp230[2] , \temp230[1] , 
        \temp230[0] }), .B(InEdges[31:16]), .LEQ(n916), .TC(n916), .GE_GT(n102
        ) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_7 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_6 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n92, n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n105, n106, 
        n107, n108, n109, n110, n111, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n93), .C(n91), .D(n89), .Z(n92) );
    VMW_NAND2 U20 ( .A(n95), .B(B[10]), .Z(n94) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n92), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n95), .C(n99), .D(n97), .Z(n100) );
    VMW_NAND2 U24 ( .A(n102), .B(B[12]), .Z(n101) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n100), .D(n94), .Z(n103) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n102), .C(n106), .D(n103), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n101), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n113), .D(n110), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n102) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n93) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n95) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n118, n119, n121, n122, n123, n124, n125, n126, n127, 
        n129, n130, n131, n132, n133, n134, n135, n137, n138, n139, n140, n141, 
        n142, n143, n145, n146, n147, n148, n149, n150, n151, n153, n154, n155, 
        n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
        n168, n169;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n119), .B(B[2]), .Z(n118) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n119), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n127), .B(B[4]), .Z(n126) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n125), .D(n118), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n127), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n135), .B(B[6]), .Z(n134) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n132), .D(n126), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n135), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n146), .C(n140), .D(n134), .Z(n145) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n147) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n149), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U20 ( .A(n151), .B(B[10]), .Z(n150) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n154), .C(n148), .D(n142), .Z(n153) );
    VMW_NAND2 U22 ( .A(n154), .B(A[9]), .Z(n155) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n151), .C(n155), .D(n153), .Z(n156) );
    VMW_NAND2 U24 ( .A(n158), .B(B[12]), .Z(n157) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n160), .C(n156), .D(n150), .Z(n159) );
    VMW_NAND2 U26 ( .A(n160), .B(A[11]), .Z(n161) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n158), .C(n161), .D(n159), .Z(n162) );
    VMW_NAND2 U28 ( .A(n164), .B(B[14]), .Z(n163) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n166), .C(n162), .D(n157), .Z(n165) );
    VMW_NAND2 U30 ( .A(n166), .B(A[13]), .Z(n167) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n164), .C(n167), .D(n165), .Z(n168) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n169), .C(n168), .D(n163), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n158) );
    VMW_INV U34 ( .A(B[7]), .Z(n146) );
    VMW_INV U35 ( .A(A[7]), .Z(n149) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n151) );
    VMW_INV U39 ( .A(B[9]), .Z(n154) );
    VMW_INV U40 ( .A(A[4]), .Z(n127) );
    VMW_INV U41 ( .A(A[8]), .Z(n143) );
    VMW_INV U42 ( .A(A[14]), .Z(n164) );
    VMW_INV U43 ( .A(B[11]), .Z(n160) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n169) );
    VMW_INV U48 ( .A(B[13]), .Z(n166) );
    VMW_INV U49 ( .A(A[6]), .Z(n135) );
    VMW_INV U50 ( .A(A[2]), .Z(n119) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
        n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
        n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
        n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
        n217, n218;
    VMW_OAI21 U3 ( .A(B[15]), .B(n170), .C(n171), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n173), .B(B[2]), .Z(n172) );
    VMW_AO22 U5 ( .A(n175), .B(B[0]), .C(n176), .D(B[1]), .Z(n174) );
    VMW_OR2 U6 ( .A(B[2]), .B(n173), .Z(n177) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n176), .C(n177), .D(n174), .Z(n178) );
    VMW_NAND2 U8 ( .A(n180), .B(B[4]), .Z(n179) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n182), .C(n178), .D(n172), .Z(n181) );
    VMW_OR2 U10 ( .A(B[4]), .B(n180), .Z(n183) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n185), .C(n183), .D(n181), .Z(n184) );
    VMW_NAND2 U12 ( .A(n187), .B(B[6]), .Z(n186) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n189), .C(n184), .D(n179), .Z(n188) );
    VMW_OR2 U14 ( .A(B[6]), .B(n187), .Z(n190) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n192), .C(n190), .D(n188), .Z(n191) );
    VMW_NAND2 U16 ( .A(n194), .B(B[8]), .Z(n193) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n196), .C(n191), .D(n186), .Z(n195) );
    VMW_OR2 U18 ( .A(B[8]), .B(n194), .Z(n197) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n199), .C(n197), .D(n195), .Z(n198) );
    VMW_NAND2 U20 ( .A(n201), .B(B[10]), .Z(n200) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n203), .C(n198), .D(n193), .Z(n202) );
    VMW_NAND2 U22 ( .A(n203), .B(A[9]), .Z(n204) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n201), .C(n204), .D(n202), .Z(n205) );
    VMW_NAND2 U24 ( .A(n207), .B(B[12]), .Z(n206) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n209), .C(n205), .D(n200), .Z(n208) );
    VMW_NAND2 U26 ( .A(n209), .B(A[11]), .Z(n210) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n207), .C(n210), .D(n208), .Z(n211) );
    VMW_NAND2 U28 ( .A(n213), .B(B[14]), .Z(n212) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n215), .C(n211), .D(n206), .Z(n214) );
    VMW_NAND2 U30 ( .A(n215), .B(A[13]), .Z(n216) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n213), .C(n216), .D(n214), .Z(n217) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n218), .C(n217), .D(n212), .Z(n171) );
    VMW_INV U33 ( .A(A[12]), .Z(n207) );
    VMW_INV U34 ( .A(B[7]), .Z(n196) );
    VMW_INV U35 ( .A(A[7]), .Z(n199) );
    VMW_INV U36 ( .A(A[3]), .Z(n185) );
    VMW_INV U37 ( .A(B[3]), .Z(n182) );
    VMW_INV U38 ( .A(A[10]), .Z(n201) );
    VMW_INV U39 ( .A(B[9]), .Z(n203) );
    VMW_INV U40 ( .A(A[4]), .Z(n180) );
    VMW_INV U41 ( .A(A[8]), .Z(n194) );
    VMW_INV U42 ( .A(A[14]), .Z(n213) );
    VMW_INV U43 ( .A(B[11]), .Z(n209) );
    VMW_INV U44 ( .A(A[5]), .Z(n192) );
    VMW_INV U45 ( .A(B[5]), .Z(n189) );
    VMW_INV U46 ( .A(A[1]), .Z(n176) );
    VMW_INV U47 ( .A(B[15]), .Z(n218) );
    VMW_INV U48 ( .A(B[13]), .Z(n215) );
    VMW_INV U49 ( .A(A[6]), .Z(n187) );
    VMW_INV U50 ( .A(A[2]), .Z(n173) );
    VMW_INV U51 ( .A(A[0]), .Z(n175) );
    VMW_INV U52 ( .A(A[15]), .Z(n170) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267;
    VMW_OAI21 U3 ( .A(B[15]), .B(n219), .C(n220), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n222), .B(B[2]), .Z(n221) );
    VMW_AO22 U5 ( .A(n224), .B(B[0]), .C(n225), .D(B[1]), .Z(n223) );
    VMW_OR2 U6 ( .A(B[2]), .B(n222), .Z(n226) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n225), .C(n226), .D(n223), .Z(n227) );
    VMW_NAND2 U8 ( .A(n229), .B(B[4]), .Z(n228) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n231), .C(n227), .D(n221), .Z(n230) );
    VMW_OR2 U10 ( .A(B[4]), .B(n229), .Z(n232) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n234), .C(n232), .D(n230), .Z(n233) );
    VMW_NAND2 U12 ( .A(n236), .B(B[6]), .Z(n235) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n238), .C(n233), .D(n228), .Z(n237) );
    VMW_OR2 U14 ( .A(B[6]), .B(n236), .Z(n239) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n241), .C(n239), .D(n237), .Z(n240) );
    VMW_NAND2 U16 ( .A(n243), .B(B[8]), .Z(n242) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n245), .C(n240), .D(n235), .Z(n244) );
    VMW_OR2 U18 ( .A(B[8]), .B(n243), .Z(n246) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n248), .C(n246), .D(n244), .Z(n247) );
    VMW_NAND2 U20 ( .A(n250), .B(B[10]), .Z(n249) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n252), .C(n247), .D(n242), .Z(n251) );
    VMW_NAND2 U22 ( .A(n252), .B(A[9]), .Z(n253) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n250), .C(n253), .D(n251), .Z(n254) );
    VMW_NAND2 U24 ( .A(n256), .B(B[12]), .Z(n255) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n258), .C(n254), .D(n249), .Z(n257) );
    VMW_NAND2 U26 ( .A(n258), .B(A[11]), .Z(n259) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n256), .C(n259), .D(n257), .Z(n260) );
    VMW_NAND2 U28 ( .A(n262), .B(B[14]), .Z(n261) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n264), .C(n260), .D(n255), .Z(n263) );
    VMW_NAND2 U30 ( .A(n264), .B(A[13]), .Z(n265) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n262), .C(n265), .D(n263), .Z(n266) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n267), .C(n266), .D(n261), .Z(n220) );
    VMW_INV U33 ( .A(A[12]), .Z(n256) );
    VMW_INV U34 ( .A(B[7]), .Z(n245) );
    VMW_INV U35 ( .A(A[7]), .Z(n248) );
    VMW_INV U36 ( .A(A[3]), .Z(n234) );
    VMW_INV U37 ( .A(B[3]), .Z(n231) );
    VMW_INV U38 ( .A(A[10]), .Z(n250) );
    VMW_INV U39 ( .A(B[9]), .Z(n252) );
    VMW_INV U40 ( .A(A[4]), .Z(n229) );
    VMW_INV U41 ( .A(A[8]), .Z(n243) );
    VMW_INV U42 ( .A(A[14]), .Z(n262) );
    VMW_INV U43 ( .A(B[11]), .Z(n258) );
    VMW_INV U44 ( .A(A[5]), .Z(n241) );
    VMW_INV U45 ( .A(B[5]), .Z(n238) );
    VMW_INV U46 ( .A(A[1]), .Z(n225) );
    VMW_INV U47 ( .A(B[15]), .Z(n267) );
    VMW_INV U48 ( .A(B[13]), .Z(n264) );
    VMW_INV U49 ( .A(A[6]), .Z(n236) );
    VMW_INV U50 ( .A(A[2]), .Z(n222) );
    VMW_INV U51 ( .A(A[0]), .Z(n224) );
    VMW_INV U52 ( .A(A[15]), .Z(n219) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
        n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
        n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
        n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
        n315, n316;
    VMW_OAI21 U3 ( .A(B[15]), .B(n268), .C(n269), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n271), .B(B[2]), .Z(n270) );
    VMW_AO22 U5 ( .A(n273), .B(B[0]), .C(n274), .D(B[1]), .Z(n272) );
    VMW_OR2 U6 ( .A(B[2]), .B(n271), .Z(n275) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n274), .C(n275), .D(n272), .Z(n276) );
    VMW_NAND2 U8 ( .A(n278), .B(B[4]), .Z(n277) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n280), .C(n276), .D(n270), .Z(n279) );
    VMW_OR2 U10 ( .A(B[4]), .B(n278), .Z(n281) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n283), .C(n281), .D(n279), .Z(n282) );
    VMW_NAND2 U12 ( .A(n285), .B(B[6]), .Z(n284) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n287), .C(n282), .D(n277), .Z(n286) );
    VMW_OR2 U14 ( .A(B[6]), .B(n285), .Z(n288) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n290), .C(n288), .D(n286), .Z(n289) );
    VMW_NAND2 U16 ( .A(n292), .B(B[8]), .Z(n291) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n294), .C(n289), .D(n284), .Z(n293) );
    VMW_OR2 U18 ( .A(B[8]), .B(n292), .Z(n295) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n297), .C(n295), .D(n293), .Z(n296) );
    VMW_NAND2 U20 ( .A(n299), .B(B[10]), .Z(n298) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n301), .C(n296), .D(n291), .Z(n300) );
    VMW_NAND2 U22 ( .A(n301), .B(A[9]), .Z(n302) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n299), .C(n302), .D(n300), .Z(n303) );
    VMW_NAND2 U24 ( .A(n305), .B(B[12]), .Z(n304) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n307), .C(n303), .D(n298), .Z(n306) );
    VMW_NAND2 U26 ( .A(n307), .B(A[11]), .Z(n308) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n305), .C(n308), .D(n306), .Z(n309) );
    VMW_NAND2 U28 ( .A(n311), .B(B[14]), .Z(n310) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n313), .C(n309), .D(n304), .Z(n312) );
    VMW_NAND2 U30 ( .A(n313), .B(A[13]), .Z(n314) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n311), .C(n314), .D(n312), .Z(n315) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n316), .C(n315), .D(n310), .Z(n269) );
    VMW_INV U33 ( .A(A[12]), .Z(n305) );
    VMW_INV U34 ( .A(B[7]), .Z(n294) );
    VMW_INV U35 ( .A(A[7]), .Z(n297) );
    VMW_INV U36 ( .A(A[3]), .Z(n283) );
    VMW_INV U37 ( .A(B[3]), .Z(n280) );
    VMW_INV U38 ( .A(A[10]), .Z(n299) );
    VMW_INV U39 ( .A(B[9]), .Z(n301) );
    VMW_INV U40 ( .A(A[4]), .Z(n278) );
    VMW_INV U41 ( .A(A[8]), .Z(n292) );
    VMW_INV U42 ( .A(A[14]), .Z(n311) );
    VMW_INV U43 ( .A(B[11]), .Z(n307) );
    VMW_INV U44 ( .A(A[5]), .Z(n290) );
    VMW_INV U45 ( .A(B[5]), .Z(n287) );
    VMW_INV U46 ( .A(A[1]), .Z(n274) );
    VMW_INV U47 ( .A(B[15]), .Z(n316) );
    VMW_INV U48 ( .A(B[13]), .Z(n313) );
    VMW_INV U49 ( .A(A[6]), .Z(n285) );
    VMW_INV U50 ( .A(A[2]), .Z(n271) );
    VMW_INV U51 ( .A(A[0]), .Z(n273) );
    VMW_INV U52 ( .A(A[15]), .Z(n268) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
        n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
        n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
        n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
        n364, n365;
    VMW_OAI21 U3 ( .A(B[15]), .B(n317), .C(n318), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n320), .B(B[2]), .Z(n319) );
    VMW_AO22 U5 ( .A(n322), .B(B[0]), .C(n323), .D(B[1]), .Z(n321) );
    VMW_OR2 U6 ( .A(B[2]), .B(n320), .Z(n324) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n323), .C(n324), .D(n321), .Z(n325) );
    VMW_NAND2 U8 ( .A(n327), .B(B[4]), .Z(n326) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n329), .C(n325), .D(n319), .Z(n328) );
    VMW_OR2 U10 ( .A(B[4]), .B(n327), .Z(n330) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n332), .C(n330), .D(n328), .Z(n331) );
    VMW_NAND2 U12 ( .A(n334), .B(B[6]), .Z(n333) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n336), .C(n331), .D(n326), .Z(n335) );
    VMW_OR2 U14 ( .A(B[6]), .B(n334), .Z(n337) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n339), .C(n337), .D(n335), .Z(n338) );
    VMW_NAND2 U16 ( .A(n341), .B(B[8]), .Z(n340) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n343), .C(n338), .D(n333), .Z(n342) );
    VMW_OR2 U18 ( .A(B[8]), .B(n341), .Z(n344) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n346), .C(n344), .D(n342), .Z(n345) );
    VMW_NAND2 U20 ( .A(n348), .B(B[10]), .Z(n347) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n350), .C(n345), .D(n340), .Z(n349) );
    VMW_NAND2 U22 ( .A(n350), .B(A[9]), .Z(n351) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n348), .C(n351), .D(n349), .Z(n352) );
    VMW_NAND2 U24 ( .A(n354), .B(B[12]), .Z(n353) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n356), .C(n352), .D(n347), .Z(n355) );
    VMW_NAND2 U26 ( .A(n356), .B(A[11]), .Z(n357) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n354), .C(n357), .D(n355), .Z(n358) );
    VMW_NAND2 U28 ( .A(n360), .B(B[14]), .Z(n359) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n362), .C(n358), .D(n353), .Z(n361) );
    VMW_NAND2 U30 ( .A(n362), .B(A[13]), .Z(n363) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n360), .C(n363), .D(n361), .Z(n364) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n365), .C(n364), .D(n359), .Z(n318) );
    VMW_INV U33 ( .A(A[12]), .Z(n354) );
    VMW_INV U34 ( .A(B[7]), .Z(n343) );
    VMW_INV U35 ( .A(A[7]), .Z(n346) );
    VMW_INV U36 ( .A(A[3]), .Z(n332) );
    VMW_INV U37 ( .A(B[3]), .Z(n329) );
    VMW_INV U38 ( .A(A[10]), .Z(n348) );
    VMW_INV U39 ( .A(B[9]), .Z(n350) );
    VMW_INV U40 ( .A(A[4]), .Z(n327) );
    VMW_INV U41 ( .A(A[8]), .Z(n341) );
    VMW_INV U42 ( .A(A[14]), .Z(n360) );
    VMW_INV U43 ( .A(B[11]), .Z(n356) );
    VMW_INV U44 ( .A(A[5]), .Z(n339) );
    VMW_INV U45 ( .A(B[5]), .Z(n336) );
    VMW_INV U46 ( .A(A[1]), .Z(n323) );
    VMW_INV U47 ( .A(B[15]), .Z(n365) );
    VMW_INV U48 ( .A(B[13]), .Z(n362) );
    VMW_INV U49 ( .A(A[6]), .Z(n334) );
    VMW_INV U50 ( .A(A[2]), .Z(n320) );
    VMW_INV U51 ( .A(A[0]), .Z(n322) );
    VMW_INV U52 ( .A(A[15]), .Z(n317) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
        n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
        n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
        n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
        n413, n414;
    VMW_OAI21 U3 ( .A(B[15]), .B(n366), .C(n367), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n369), .B(B[2]), .Z(n368) );
    VMW_AO22 U5 ( .A(n371), .B(B[0]), .C(n372), .D(B[1]), .Z(n370) );
    VMW_OR2 U6 ( .A(B[2]), .B(n369), .Z(n373) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n372), .C(n373), .D(n370), .Z(n374) );
    VMW_NAND2 U8 ( .A(n376), .B(B[4]), .Z(n375) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n378), .C(n374), .D(n368), .Z(n377) );
    VMW_OR2 U10 ( .A(B[4]), .B(n376), .Z(n379) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n381), .C(n379), .D(n377), .Z(n380) );
    VMW_NAND2 U12 ( .A(n383), .B(B[6]), .Z(n382) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n385), .C(n380), .D(n375), .Z(n384) );
    VMW_OR2 U14 ( .A(B[6]), .B(n383), .Z(n386) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n388), .C(n386), .D(n384), .Z(n387) );
    VMW_NAND2 U16 ( .A(n390), .B(B[8]), .Z(n389) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n392), .C(n387), .D(n382), .Z(n391) );
    VMW_OR2 U18 ( .A(B[8]), .B(n390), .Z(n393) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n395), .C(n393), .D(n391), .Z(n394) );
    VMW_NAND2 U20 ( .A(n397), .B(B[10]), .Z(n396) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n399), .C(n394), .D(n389), .Z(n398) );
    VMW_NAND2 U22 ( .A(n399), .B(A[9]), .Z(n400) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n397), .C(n400), .D(n398), .Z(n401) );
    VMW_NAND2 U24 ( .A(n403), .B(B[12]), .Z(n402) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n405), .C(n401), .D(n396), .Z(n404) );
    VMW_NAND2 U26 ( .A(n405), .B(A[11]), .Z(n406) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n403), .C(n406), .D(n404), .Z(n407) );
    VMW_NAND2 U28 ( .A(n409), .B(B[14]), .Z(n408) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n411), .C(n407), .D(n402), .Z(n410) );
    VMW_NAND2 U30 ( .A(n411), .B(A[13]), .Z(n412) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n409), .C(n412), .D(n410), .Z(n413) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n414), .C(n413), .D(n408), .Z(n367) );
    VMW_INV U33 ( .A(A[12]), .Z(n403) );
    VMW_INV U34 ( .A(B[7]), .Z(n392) );
    VMW_INV U35 ( .A(A[7]), .Z(n395) );
    VMW_INV U36 ( .A(A[3]), .Z(n381) );
    VMW_INV U37 ( .A(B[3]), .Z(n378) );
    VMW_INV U38 ( .A(A[10]), .Z(n397) );
    VMW_INV U39 ( .A(B[9]), .Z(n399) );
    VMW_INV U40 ( .A(A[4]), .Z(n376) );
    VMW_INV U41 ( .A(A[8]), .Z(n390) );
    VMW_INV U42 ( .A(A[14]), .Z(n409) );
    VMW_INV U43 ( .A(B[11]), .Z(n405) );
    VMW_INV U44 ( .A(A[5]), .Z(n388) );
    VMW_INV U45 ( .A(B[5]), .Z(n385) );
    VMW_INV U46 ( .A(A[1]), .Z(n372) );
    VMW_INV U47 ( .A(B[15]), .Z(n414) );
    VMW_INV U48 ( .A(B[13]), .Z(n411) );
    VMW_INV U49 ( .A(A[6]), .Z(n383) );
    VMW_INV U50 ( .A(A[2]), .Z(n369) );
    VMW_INV U51 ( .A(A[0]), .Z(n371) );
    VMW_INV U52 ( .A(A[15]), .Z(n366) );
endmodule


module NodeAux_INDEGREE8_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [7:0] Nid;
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp240[2] , \temp334[3] , \temp424[2] , \temp604[10] , 
        \temp424[14] , n152, \temp694[10] , \temp604[3] , \temp784[12] , n112, 
        \temp424[10] , \temp604[14] , \temp424[6] , \temp240[6] , \temp334[7] , 
        \path[2] , \temp604[7] , \temp694[14] , \path[0] , \temp604[5] , 
        \temp784[14] , \temp424[4] , \temp240[4] , \temp334[5] , \temp424[12] , 
        \temp334[8] , n120, \temp784[10] , \temp240[9] , \temp424[9] , 
        \temp694[12] , \temp604[1] , \temp604[8] , \temp604[12] , \temp334[1] , 
        \temp424[0] , \temp240[0] , \temp240[14] , \temp514[3] , \temp334[10] , 
        \temp694[2] , \temp784[7] , \temp514[13] , \OutEdge166[13] , 
        \OutEdge166[3] , n128, \temp694[6] , \temp784[3] , \temp334[14] , 
        \temp514[7] , \OutEdge166[7] , \temp240[10] , \temp784[8] , 
        \temp514[15] , \OutEdge166[15] , \OutEdge166[5] , n96, \temp514[5] , 
        \temp240[12] , \temp784[1] , \temp694[4] , \temp514[8] , 
        \OutEdge166[11] , \OutEdge166[1] , \temp694[9] , \temp514[11] , 
        \temp334[12] , \temp694[0] , \temp784[5] , \temp514[1] , 
        \OutEdge166[8] , \temp514[9] , \OutEdge166[10] , \OutEdge166[0] , 
        \temp694[8] , \temp514[10] , \temp694[1] , \temp334[13] , \temp514[0] , 
        \temp784[4] , \OutEdge166[9] , \temp514[14] , \temp784[9] , n136, 
        \OutEdge166[14] , \OutEdge166[4] , \temp240[13] , \temp514[4] , 
        \temp784[0] , \temp694[5] , \temp784[2] , \temp334[15] , \temp694[7] , 
        \temp240[11] , \temp514[6] , n144, \OutEdge166[6] , \temp514[2] , n104, 
        \temp240[15] , \temp694[3] , \temp334[11] , \temp784[6] , 
        \temp514[12] , \OutEdge166[12] , \OutEdge166[2] , \temp334[9] , 
        \temp240[8] , \temp424[8] , \temp784[11] , \temp694[13] , \temp604[0] , 
        \temp604[13] , \temp604[9] , \temp334[0] , \temp240[1] , \temp424[1] , 
        \path[1] , \temp604[4] , \temp784[15] , \temp424[5] , \temp240[5] , 
        \temp334[4] , \temp424[13] , \temp424[11] , \temp604[15] , 
        \temp424[7] , \temp240[7] , \temp334[6] , \path[3] , \temp694[15] , 
        \temp604[6] , \temp334[2] , \temp424[3] , \temp240[3] , \temp604[11] , 
        \temp424[15] , \temp604[2] , \temp694[11] , \temp784[13] , n967, n968, 
        n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
        n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
        n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
        n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
        n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
        n1024, n1025, n1026;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U109 ( .Z(n1021) );
    VMW_PULLDOWN U110 ( .Z(n1020) );
    VMW_PULLDOWN U111 ( .Z(n1023) );
    VMW_PULLDOWN U112 ( .Z(n1024) );
    VMW_PULLDOWN U113 ( .Z(n1019) );
    VMW_PULLDOWN U114 ( .Z(n1026) );
    VMW_PULLDOWN U115 ( .Z(n1022) );
    VMW_PULLDOWN U116 ( .Z(n1025) );
    VMW_NOR2 U117 ( .A(Start), .B(n967), .Z(\OutEdge166[15] ) );
    VMW_NAND2 U118 ( .A(n968), .B(n969), .Z(\OutEdge166[14] ) );
    VMW_NAND2 U119 ( .A(n970), .B(n969), .Z(\OutEdge166[13] ) );
    VMW_NAND2 U120 ( .A(n971), .B(n969), .Z(\OutEdge166[12] ) );
    VMW_NAND2 U121 ( .A(n972), .B(n969), .Z(\OutEdge166[11] ) );
    VMW_NAND2 U122 ( .A(n973), .B(n969), .Z(\OutEdge166[10] ) );
    VMW_NAND2 U123 ( .A(n974), .B(n969), .Z(\OutEdge166[9] ) );
    VMW_NAND2 U124 ( .A(n975), .B(n969), .Z(\OutEdge166[8] ) );
    VMW_NAND2 U125 ( .A(n976), .B(n969), .Z(\OutEdge166[7] ) );
    VMW_NAND2 U126 ( .A(n977), .B(n969), .Z(\OutEdge166[6] ) );
    VMW_NAND2 U127 ( .A(n978), .B(n969), .Z(\OutEdge166[5] ) );
    VMW_NAND2 U128 ( .A(n979), .B(n969), .Z(\OutEdge166[4] ) );
    VMW_NAND2 U129 ( .A(n980), .B(n969), .Z(\OutEdge166[3] ) );
    VMW_NAND2 U130 ( .A(n981), .B(n969), .Z(\OutEdge166[2] ) );
    VMW_NAND2 U131 ( .A(n982), .B(n969), .Z(\OutEdge166[1] ) );
    VMW_NAND2 U132 ( .A(n983), .B(n969), .Z(\OutEdge166[0] ) );
    VMW_AO21 U133 ( .A(n984), .B(n985), .C(n986), .Z(n1018) );
    VMW_AO22 U134 ( .A(\path[3] ), .B(Start), .C(n987), .D(n988), .Z(n1017) );
    VMW_OR4 U135 ( .A(n136), .B(n128), .C(n987), .D(n990), .Z(n989) );
    VMW_OR2 U136 ( .A(n152), .B(n992), .Z(n991) );
    VMW_AO22 U137 ( .A(\temp694[15] ), .B(n993), .C(InEdges[111]), .D(n144), 
        .Z(\temp784[15] ) );
    VMW_OR2 U138 ( .A(n152), .B(n144), .Z(n990) );
    VMW_AND3 U139 ( .A(n969), .B(n994), .C(n995), .Z(n984) );
    VMW_AND4 U140 ( .A(n996), .B(n997), .C(n998), .D(n999), .Z(n987) );
    VMW_INV U141 ( .A(Start), .Z(n969) );
    VMW_OAI22 U142 ( .A(n989), .B(Start), .C(\path[2] ), .D(n969), .Z(n1000)
         );
    VMW_AO22 U143 ( .A(\path[1] ), .B(Start), .C(n990), .D(n969), .Z(n986) );
    VMW_OAI22 U144 ( .A(n991), .B(Start), .C(\path[0] ), .D(n969), .Z(n1001)
         );
    VMW_MUX2I U145 ( .A(\temp784[15] ), .B(InEdges[127]), .S(n152), .Z(n967)
         );
    VMW_NOR2 U146 ( .A(n990), .B(n1002), .Z(n988) );
    VMW_AND4 U147 ( .A(n1004), .B(n1005), .C(n1006), .D(n1007), .Z(n1003) );
    VMW_INV U148 ( .A(n120), .Z(n999) );
    VMW_INV U149 ( .A(n136), .Z(n994) );
    VMW_INV U150 ( .A(n112), .Z(n997) );
    VMW_OAI211 U151 ( .A(n96), .B(n104), .C(n997), .D(n999), .Z(n985) );
    VMW_AO21 U152 ( .A(n996), .B(n96), .C(n112), .Z(n1008) );
    VMW_AO21 U153 ( .A(n999), .B(n1008), .C(n128), .Z(n1009) );
    VMW_AOI21 U154 ( .A(n994), .B(n1009), .C(n144), .Z(n992) );
    VMW_AND5 U155 ( .A(n1010), .B(n1011), .C(n1012), .D(n1013), .E(n1003), .Z(
        n1014) );
    VMW_XNOR2 U156 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n1007) );
    VMW_XNOR2 U157 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n1006) );
    VMW_XNOR2 U158 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n1005) );
    VMW_XNOR2 U159 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n1004) );
    VMW_XNOR2 U160 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n1013) );
    VMW_XNOR2 U161 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n1012) );
    VMW_XNOR2 U162 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n1011) );
    VMW_XNOR2 U163 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n1010) );
    VMW_AO22 U164 ( .A(InEdges[9]), .B(n96), .C(OutEdge[9]), .D(n998), .Z(
        \temp240[9] ) );
    VMW_AO22 U165 ( .A(\temp240[9] ), .B(n996), .C(InEdges[25]), .D(n104), .Z(
        \temp334[9] ) );
    VMW_AO22 U166 ( .A(InEdges[41]), .B(n112), .C(\temp334[9] ), .D(n997), .Z(
        \temp424[9] ) );
    VMW_AO22 U167 ( .A(InEdges[57]), .B(n120), .C(\temp424[9] ), .D(n999), .Z(
        \temp514[9] ) );
    VMW_AO22 U168 ( .A(\temp514[9] ), .B(n995), .C(InEdges[73]), .D(n128), .Z(
        \temp604[9] ) );
    VMW_AO22 U169 ( .A(InEdges[89]), .B(n136), .C(\temp604[9] ), .D(n994), .Z(
        \temp694[9] ) );
    VMW_AO22 U170 ( .A(\temp694[9] ), .B(n993), .C(InEdges[105]), .D(n144), 
        .Z(\temp784[9] ) );
    VMW_AO22 U171 ( .A(InEdges[8]), .B(n96), .C(OutEdge[8]), .D(n998), .Z(
        \temp240[8] ) );
    VMW_AO22 U172 ( .A(\temp240[8] ), .B(n996), .C(InEdges[24]), .D(n104), .Z(
        \temp334[8] ) );
    VMW_AO22 U173 ( .A(InEdges[40]), .B(n112), .C(\temp334[8] ), .D(n997), .Z(
        \temp424[8] ) );
    VMW_AO22 U174 ( .A(InEdges[56]), .B(n120), .C(\temp424[8] ), .D(n999), .Z(
        \temp514[8] ) );
    VMW_AO22 U175 ( .A(\temp514[8] ), .B(n995), .C(InEdges[72]), .D(n128), .Z(
        \temp604[8] ) );
    VMW_AO22 U176 ( .A(InEdges[88]), .B(n136), .C(\temp604[8] ), .D(n994), .Z(
        \temp694[8] ) );
    VMW_AO22 U177 ( .A(\temp694[8] ), .B(n993), .C(InEdges[104]), .D(n144), 
        .Z(\temp784[8] ) );
    VMW_AO22 U178 ( .A(InEdges[7]), .B(n96), .C(OutEdge[7]), .D(n998), .Z(
        \temp240[7] ) );
    VMW_AO22 U179 ( .A(\temp240[7] ), .B(n996), .C(InEdges[23]), .D(n104), .Z(
        \temp334[7] ) );
    VMW_AO22 U180 ( .A(InEdges[39]), .B(n112), .C(\temp334[7] ), .D(n997), .Z(
        \temp424[7] ) );
    VMW_AO22 U181 ( .A(InEdges[55]), .B(n120), .C(\temp424[7] ), .D(n999), .Z(
        \temp514[7] ) );
    VMW_AO22 U182 ( .A(\temp514[7] ), .B(n995), .C(InEdges[71]), .D(n128), .Z(
        \temp604[7] ) );
    VMW_AO22 U183 ( .A(InEdges[87]), .B(n136), .C(\temp604[7] ), .D(n994), .Z(
        \temp694[7] ) );
    VMW_AO22 U184 ( .A(\temp694[7] ), .B(n993), .C(InEdges[103]), .D(n144), 
        .Z(\temp784[7] ) );
    VMW_AO22 U185 ( .A(InEdges[6]), .B(n96), .C(OutEdge[6]), .D(n998), .Z(
        \temp240[6] ) );
    VMW_AO22 U186 ( .A(\temp240[6] ), .B(n996), .C(InEdges[22]), .D(n104), .Z(
        \temp334[6] ) );
    VMW_AO22 U187 ( .A(InEdges[38]), .B(n112), .C(\temp334[6] ), .D(n997), .Z(
        \temp424[6] ) );
    VMW_AO22 U188 ( .A(InEdges[54]), .B(n120), .C(\temp424[6] ), .D(n999), .Z(
        \temp514[6] ) );
    VMW_AO22 U189 ( .A(\temp514[6] ), .B(n995), .C(InEdges[70]), .D(n128), .Z(
        \temp604[6] ) );
    VMW_AO22 U190 ( .A(InEdges[86]), .B(n136), .C(\temp604[6] ), .D(n994), .Z(
        \temp694[6] ) );
    VMW_AO22 U191 ( .A(\temp694[6] ), .B(n993), .C(InEdges[102]), .D(n144), 
        .Z(\temp784[6] ) );
    VMW_AO22 U192 ( .A(InEdges[5]), .B(n96), .C(OutEdge[5]), .D(n998), .Z(
        \temp240[5] ) );
    VMW_AO22 U193 ( .A(\temp240[5] ), .B(n996), .C(InEdges[21]), .D(n104), .Z(
        \temp334[5] ) );
    VMW_AO22 U194 ( .A(InEdges[37]), .B(n112), .C(\temp334[5] ), .D(n997), .Z(
        \temp424[5] ) );
    VMW_AO22 U195 ( .A(InEdges[53]), .B(n120), .C(\temp424[5] ), .D(n999), .Z(
        \temp514[5] ) );
    VMW_AO22 U196 ( .A(\temp514[5] ), .B(n995), .C(InEdges[69]), .D(n128), .Z(
        \temp604[5] ) );
    VMW_AO22 U197 ( .A(InEdges[85]), .B(n136), .C(\temp604[5] ), .D(n994), .Z(
        \temp694[5] ) );
    VMW_AO22 U198 ( .A(\temp694[5] ), .B(n993), .C(InEdges[101]), .D(n144), 
        .Z(\temp784[5] ) );
    VMW_AO22 U199 ( .A(InEdges[4]), .B(n96), .C(OutEdge[4]), .D(n998), .Z(
        \temp240[4] ) );
    VMW_AO22 U200 ( .A(\temp240[4] ), .B(n996), .C(InEdges[20]), .D(n104), .Z(
        \temp334[4] ) );
    VMW_AO22 U201 ( .A(InEdges[36]), .B(n112), .C(\temp334[4] ), .D(n997), .Z(
        \temp424[4] ) );
    VMW_AO22 U202 ( .A(InEdges[52]), .B(n120), .C(\temp424[4] ), .D(n999), .Z(
        \temp514[4] ) );
    VMW_AO22 U203 ( .A(\temp514[4] ), .B(n995), .C(InEdges[68]), .D(n128), .Z(
        \temp604[4] ) );
    VMW_AO22 U204 ( .A(InEdges[84]), .B(n136), .C(\temp604[4] ), .D(n994), .Z(
        \temp694[4] ) );
    VMW_AO22 U205 ( .A(\temp694[4] ), .B(n993), .C(InEdges[100]), .D(n144), 
        .Z(\temp784[4] ) );
    VMW_AO22 U206 ( .A(InEdges[3]), .B(n96), .C(OutEdge[3]), .D(n998), .Z(
        \temp240[3] ) );
    VMW_AO22 U207 ( .A(\temp240[3] ), .B(n996), .C(InEdges[19]), .D(n104), .Z(
        \temp334[3] ) );
    VMW_AO22 U208 ( .A(InEdges[35]), .B(n112), .C(\temp334[3] ), .D(n997), .Z(
        \temp424[3] ) );
    VMW_AO22 U209 ( .A(InEdges[51]), .B(n120), .C(\temp424[3] ), .D(n999), .Z(
        \temp514[3] ) );
    VMW_AO22 U210 ( .A(\temp514[3] ), .B(n995), .C(InEdges[67]), .D(n128), .Z(
        \temp604[3] ) );
    VMW_AO22 U211 ( .A(InEdges[83]), .B(n136), .C(\temp604[3] ), .D(n994), .Z(
        \temp694[3] ) );
    VMW_AO22 U212 ( .A(\temp694[3] ), .B(n993), .C(InEdges[99]), .D(n144), .Z(
        \temp784[3] ) );
    VMW_AO22 U213 ( .A(InEdges[2]), .B(n96), .C(OutEdge[2]), .D(n998), .Z(
        \temp240[2] ) );
    VMW_AO22 U214 ( .A(\temp240[2] ), .B(n996), .C(InEdges[18]), .D(n104), .Z(
        \temp334[2] ) );
    VMW_AO22 U215 ( .A(InEdges[34]), .B(n112), .C(\temp334[2] ), .D(n997), .Z(
        \temp424[2] ) );
    VMW_AO22 U216 ( .A(InEdges[50]), .B(n120), .C(\temp424[2] ), .D(n999), .Z(
        \temp514[2] ) );
    VMW_AO22 U217 ( .A(\temp514[2] ), .B(n995), .C(InEdges[66]), .D(n128), .Z(
        \temp604[2] ) );
    VMW_AO22 U218 ( .A(InEdges[82]), .B(n136), .C(\temp604[2] ), .D(n994), .Z(
        \temp694[2] ) );
    VMW_AO22 U219 ( .A(\temp694[2] ), .B(n993), .C(InEdges[98]), .D(n144), .Z(
        \temp784[2] ) );
    VMW_AO22 U220 ( .A(InEdges[1]), .B(n96), .C(OutEdge[1]), .D(n998), .Z(
        \temp240[1] ) );
    VMW_AO22 U221 ( .A(\temp240[1] ), .B(n996), .C(InEdges[17]), .D(n104), .Z(
        \temp334[1] ) );
    VMW_AO22 U222 ( .A(InEdges[33]), .B(n112), .C(\temp334[1] ), .D(n997), .Z(
        \temp424[1] ) );
    VMW_AO22 U223 ( .A(InEdges[49]), .B(n120), .C(\temp424[1] ), .D(n999), .Z(
        \temp514[1] ) );
    VMW_AO22 U224 ( .A(\temp514[1] ), .B(n995), .C(InEdges[65]), .D(n128), .Z(
        \temp604[1] ) );
    VMW_AO22 U225 ( .A(InEdges[81]), .B(n136), .C(\temp604[1] ), .D(n994), .Z(
        \temp694[1] ) );
    VMW_AO22 U226 ( .A(\temp694[1] ), .B(n993), .C(InEdges[97]), .D(n144), .Z(
        \temp784[1] ) );
    VMW_AO22 U227 ( .A(InEdges[15]), .B(n96), .C(OutEdge[15]), .D(n998), .Z(
        \temp240[15] ) );
    VMW_AO22 U228 ( .A(\temp240[15] ), .B(n996), .C(InEdges[31]), .D(n104), 
        .Z(\temp334[15] ) );
    VMW_AO22 U229 ( .A(InEdges[47]), .B(n112), .C(\temp334[15] ), .D(n997), 
        .Z(\temp424[15] ) );
    VMW_AO22 U230 ( .A(InEdges[63]), .B(n120), .C(\temp424[15] ), .D(n999), 
        .Z(\temp514[15] ) );
    VMW_AO22 U231 ( .A(\temp514[15] ), .B(n995), .C(InEdges[79]), .D(n128), 
        .Z(\temp604[15] ) );
    VMW_AO22 U232 ( .A(InEdges[95]), .B(n136), .C(\temp604[15] ), .D(n994), 
        .Z(\temp694[15] ) );
    VMW_AO22 U233 ( .A(InEdges[14]), .B(n96), .C(OutEdge[14]), .D(n998), .Z(
        \temp240[14] ) );
    VMW_AO22 U234 ( .A(\temp240[14] ), .B(n996), .C(InEdges[30]), .D(n104), 
        .Z(\temp334[14] ) );
    VMW_AO22 U235 ( .A(InEdges[46]), .B(n112), .C(\temp334[14] ), .D(n997), 
        .Z(\temp424[14] ) );
    VMW_AO22 U236 ( .A(InEdges[62]), .B(n120), .C(\temp424[14] ), .D(n999), 
        .Z(\temp514[14] ) );
    VMW_AO22 U237 ( .A(\temp514[14] ), .B(n995), .C(InEdges[78]), .D(n128), 
        .Z(\temp604[14] ) );
    VMW_AO22 U238 ( .A(InEdges[94]), .B(n136), .C(\temp604[14] ), .D(n994), 
        .Z(\temp694[14] ) );
    VMW_AO22 U239 ( .A(\temp694[14] ), .B(n993), .C(InEdges[110]), .D(n144), 
        .Z(\temp784[14] ) );
    VMW_AO22 U240 ( .A(InEdges[13]), .B(n96), .C(OutEdge[13]), .D(n998), .Z(
        \temp240[13] ) );
    VMW_AO22 U241 ( .A(\temp240[13] ), .B(n996), .C(InEdges[29]), .D(n104), 
        .Z(\temp334[13] ) );
    VMW_AO22 U242 ( .A(InEdges[45]), .B(n112), .C(\temp334[13] ), .D(n997), 
        .Z(\temp424[13] ) );
    VMW_AO22 U243 ( .A(InEdges[61]), .B(n120), .C(\temp424[13] ), .D(n999), 
        .Z(\temp514[13] ) );
    VMW_AO22 U244 ( .A(\temp514[13] ), .B(n995), .C(InEdges[77]), .D(n128), 
        .Z(\temp604[13] ) );
    VMW_AO22 U245 ( .A(InEdges[93]), .B(n136), .C(\temp604[13] ), .D(n994), 
        .Z(\temp694[13] ) );
    VMW_AO22 U246 ( .A(\temp694[13] ), .B(n993), .C(InEdges[109]), .D(n144), 
        .Z(\temp784[13] ) );
    VMW_AO22 U247 ( .A(InEdges[12]), .B(n96), .C(OutEdge[12]), .D(n998), .Z(
        \temp240[12] ) );
    VMW_AO22 U248 ( .A(\temp240[12] ), .B(n996), .C(InEdges[28]), .D(n104), 
        .Z(\temp334[12] ) );
    VMW_AO22 U249 ( .A(InEdges[44]), .B(n112), .C(\temp334[12] ), .D(n997), 
        .Z(\temp424[12] ) );
    VMW_AO22 U250 ( .A(InEdges[60]), .B(n120), .C(\temp424[12] ), .D(n999), 
        .Z(\temp514[12] ) );
    VMW_AO22 U251 ( .A(\temp514[12] ), .B(n995), .C(InEdges[76]), .D(n128), 
        .Z(\temp604[12] ) );
    VMW_AO22 U252 ( .A(InEdges[92]), .B(n136), .C(\temp604[12] ), .D(n994), 
        .Z(\temp694[12] ) );
    VMW_AO22 U253 ( .A(\temp694[12] ), .B(n993), .C(InEdges[108]), .D(n144), 
        .Z(\temp784[12] ) );
    VMW_AO22 U254 ( .A(InEdges[11]), .B(n96), .C(OutEdge[11]), .D(n998), .Z(
        \temp240[11] ) );
    VMW_AO22 U255 ( .A(\temp240[11] ), .B(n996), .C(InEdges[27]), .D(n104), 
        .Z(\temp334[11] ) );
    VMW_AO22 U256 ( .A(InEdges[43]), .B(n112), .C(\temp334[11] ), .D(n997), 
        .Z(\temp424[11] ) );
    VMW_AO22 U257 ( .A(InEdges[59]), .B(n120), .C(\temp424[11] ), .D(n999), 
        .Z(\temp514[11] ) );
    VMW_AO22 U258 ( .A(\temp514[11] ), .B(n995), .C(InEdges[75]), .D(n128), 
        .Z(\temp604[11] ) );
    VMW_AO22 U259 ( .A(InEdges[91]), .B(n136), .C(\temp604[11] ), .D(n994), 
        .Z(\temp694[11] ) );
    VMW_AO22 U260 ( .A(\temp694[11] ), .B(n993), .C(InEdges[107]), .D(n144), 
        .Z(\temp784[11] ) );
    VMW_AO22 U261 ( .A(InEdges[10]), .B(n96), .C(OutEdge[10]), .D(n998), .Z(
        \temp240[10] ) );
    VMW_AO22 U262 ( .A(\temp240[10] ), .B(n996), .C(InEdges[26]), .D(n104), 
        .Z(\temp334[10] ) );
    VMW_AO22 U263 ( .A(InEdges[42]), .B(n112), .C(\temp334[10] ), .D(n997), 
        .Z(\temp424[10] ) );
    VMW_AO22 U264 ( .A(InEdges[58]), .B(n120), .C(\temp424[10] ), .D(n999), 
        .Z(\temp514[10] ) );
    VMW_AO22 U265 ( .A(\temp514[10] ), .B(n995), .C(InEdges[74]), .D(n128), 
        .Z(\temp604[10] ) );
    VMW_AO22 U266 ( .A(InEdges[90]), .B(n136), .C(\temp604[10] ), .D(n994), 
        .Z(\temp694[10] ) );
    VMW_AO22 U267 ( .A(\temp694[10] ), .B(n993), .C(InEdges[106]), .D(n144), 
        .Z(\temp784[10] ) );
    VMW_AO22 U268 ( .A(InEdges[0]), .B(n96), .C(OutEdge[0]), .D(n998), .Z(
        \temp240[0] ) );
    VMW_AO22 U269 ( .A(\temp240[0] ), .B(n996), .C(InEdges[16]), .D(n104), .Z(
        \temp334[0] ) );
    VMW_AO22 U270 ( .A(InEdges[32]), .B(n112), .C(\temp334[0] ), .D(n997), .Z(
        \temp424[0] ) );
    VMW_AO22 U271 ( .A(InEdges[48]), .B(n120), .C(\temp424[0] ), .D(n999), .Z(
        \temp514[0] ) );
    VMW_AO22 U272 ( .A(\temp514[0] ), .B(n995), .C(InEdges[64]), .D(n128), .Z(
        \temp604[0] ) );
    VMW_AO22 U273 ( .A(InEdges[80]), .B(n136), .C(\temp604[0] ), .D(n994), .Z(
        \temp694[0] ) );
    VMW_AO22 U274 ( .A(\temp694[0] ), .B(n993), .C(InEdges[96]), .D(n144), .Z(
        \temp784[0] ) );
    VMW_MUX2I U275 ( .A(\temp784[9] ), .B(InEdges[121]), .S(n152), .Z(n974) );
    VMW_MUX2I U276 ( .A(\temp784[8] ), .B(InEdges[120]), .S(n152), .Z(n975) );
    VMW_MUX2I U277 ( .A(\temp784[7] ), .B(InEdges[119]), .S(n152), .Z(n976) );
    VMW_MUX2I U278 ( .A(\temp784[6] ), .B(InEdges[118]), .S(n152), .Z(n977) );
    VMW_MUX2I U279 ( .A(\temp784[5] ), .B(InEdges[117]), .S(n152), .Z(n978) );
    VMW_MUX2I U280 ( .A(\temp784[4] ), .B(InEdges[116]), .S(n152), .Z(n979) );
    VMW_MUX2I U281 ( .A(\temp784[3] ), .B(InEdges[115]), .S(n152), .Z(n980) );
    VMW_MUX2I U282 ( .A(\temp784[2] ), .B(InEdges[114]), .S(n152), .Z(n981) );
    VMW_MUX2I U283 ( .A(\temp784[1] ), .B(InEdges[113]), .S(n152), .Z(n982) );
    VMW_MUX2I U284 ( .A(\temp784[14] ), .B(InEdges[126]), .S(n152), .Z(n968)
         );
    VMW_MUX2I U285 ( .A(\temp784[13] ), .B(InEdges[125]), .S(n152), .Z(n970)
         );
    VMW_MUX2I U286 ( .A(\temp784[12] ), .B(InEdges[124]), .S(n152), .Z(n971)
         );
    VMW_MUX2I U287 ( .A(\temp784[11] ), .B(InEdges[123]), .S(n152), .Z(n972)
         );
    VMW_MUX2I U288 ( .A(\temp784[10] ), .B(InEdges[122]), .S(n152), .Z(n973)
         );
    VMW_MUX2I U289 ( .A(\temp784[0] ), .B(InEdges[112]), .S(n152), .Z(n983) );
    VMW_INV U290 ( .A(n96), .Z(n998) );
    VMW_INV U291 ( .A(n104), .Z(n996) );
    VMW_INV U292 ( .A(n128), .Z(n995) );
    VMW_INV U293 ( .A(n144), .Z(n993) );
    VMW_INV U294 ( .A(n984), .Z(n1002) );
    VMW_INV U295 ( .A(n1000), .Z(n1016) );
    VMW_INV U296 ( .A(n1001), .Z(n1015) );
    VMW_BUFIZ U297 ( .A(\path[3] ), .E(n1014), .Z(\PathData[3] ) );
    VMW_BUFIZ U298 ( .A(\path[1] ), .E(n1014), .Z(\PathData[1] ) );
    VMW_BUFIZ U299 ( .A(\path[0] ), .E(n1014), .Z(\PathData[0] ) );
    VMW_BUFIZ U300 ( .A(\path[2] ), .E(n1014), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n1015), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n1016), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n1017), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n1018), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge166[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge166[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge166[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge166[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge166[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge166[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge166[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge166[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge166[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge166[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge166[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge166[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge166[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge166[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge166[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge166[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_7 lte_55_2 ( .A({\temp334[15] , 
        \temp334[14] , \temp334[13] , \temp334[12] , \temp334[11] , 
        \temp334[10] , \temp334[9] , \temp334[8] , \temp334[7] , \temp334[6] , 
        \temp334[5] , \temp334[4] , \temp334[3] , \temp334[2] , \temp334[1] , 
        \temp334[0] }), .B(InEdges[47:32]), .LEQ(n1026), .TC(n1026), .GE_GT(
        n112) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_6 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n1025), .TC(n1025), .GE_GT(n96) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_5 lte_55_4 ( .A({\temp514[15] , 
        \temp514[14] , \temp514[13] , \temp514[12] , \temp514[11] , 
        \temp514[10] , \temp514[9] , \temp514[8] , \temp514[7] , \temp514[6] , 
        \temp514[5] , \temp514[4] , \temp514[3] , \temp514[2] , \temp514[1] , 
        \temp514[0] }), .B(InEdges[79:64]), .LEQ(n1024), .TC(n1024), .GE_GT(
        n128) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_4 lte_55_5 ( .A({\temp604[15] , 
        \temp604[14] , \temp604[13] , \temp604[12] , \temp604[11] , 
        \temp604[10] , \temp604[9] , \temp604[8] , \temp604[7] , \temp604[6] , 
        \temp604[5] , \temp604[4] , \temp604[3] , \temp604[2] , \temp604[1] , 
        \temp604[0] }), .B(InEdges[95:80]), .LEQ(n1023), .TC(n1023), .GE_GT(
        n136) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_3 lte_55_1 ( .A({\temp240[15] , 
        \temp240[14] , \temp240[13] , \temp240[12] , \temp240[11] , 
        \temp240[10] , \temp240[9] , \temp240[8] , \temp240[7] , \temp240[6] , 
        \temp240[5] , \temp240[4] , \temp240[3] , \temp240[2] , \temp240[1] , 
        \temp240[0] }), .B(InEdges[31:16]), .LEQ(n1022), .TC(n1022), .GE_GT(
        n104) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_2 lte_55_7 ( .A({\temp784[15] , 
        \temp784[14] , \temp784[13] , \temp784[12] , \temp784[11] , 
        \temp784[10] , \temp784[9] , \temp784[8] , \temp784[7] , \temp784[6] , 
        \temp784[5] , \temp784[4] , \temp784[3] , \temp784[2] , \temp784[1] , 
        \temp784[0] }), .B(InEdges[127:112]), .LEQ(n1021), .TC(n1021), .GE_GT(
        n152) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_1 lte_55_6 ( .A({\temp694[15] , 
        \temp694[14] , \temp694[13] , \temp694[12] , \temp694[11] , 
        \temp694[10] , \temp694[9] , \temp694[8] , \temp694[7] , \temp694[6] , 
        \temp694[5] , \temp694[4] , \temp694[3] , \temp694[2] , \temp694[1] , 
        \temp694[0] }), .B(InEdges[111:96]), .LEQ(n1020), .TC(n1020), .GE_GT(
        n144) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp424[15] , 
        \temp424[14] , \temp424[13] , \temp424[12] , \temp424[11] , 
        \temp424[10] , \temp424[9] , \temp424[8] , \temp424[7] , \temp424[6] , 
        \temp424[5] , \temp424[4] , \temp424[3] , \temp424[2] , \temp424[1] , 
        \temp424[0] }), .B(InEdges[63:48]), .LEQ(n1019), .TC(n1019), .GE_GT(
        n120) );
endmodule


module library ( InEdges, OutEdge, PathAddr, PathData, WeightAddr, WeightData, 
    Nid, Eid, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
input  [10:0] WeightAddr;
input  [10:0] Eid;
output [3:0] PathData;
input  [15:0] WeightData;
input  [7:0] Nid;
input  Start, Clk;
    EdgeAux edgeAux ( .Eid(Eid), .InEdge(InEdges[15:0]), .OutEdge(OutEdge), 
        .WeightAddr(WeightAddr), .WeightData(WeightData), .Clk(Clk) );
    NodeAux_INDEGREE8_SOURCE1 n_8_1 ( .Nid(Nid), .InEdges(InEdges), .OutEdge(
        OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(Start), 
        .Clk(Clk) );
    NodeAux_INDEGREE1_SOURCE0 n_1_0 ( .Nid(Nid), .InEdges(InEdges[15:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE2_SOURCE0 n_2_0 ( .Nid(Nid), .InEdges(InEdges[31:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE4_SOURCE0 n_4_0 ( .Nid(Nid), .InEdges(InEdges[63:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE5_SOURCE0 n_5_0 ( .Nid(Nid), .InEdges(InEdges[79:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE6_SOURCE0 n_6_0 ( .Nid(Nid), .InEdges(InEdges[95:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE7_SOURCE0 n_7_0 ( .Nid(Nid), .InEdges(InEdges[111:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE8_SOURCE0 n_8_0 ( .Nid(Nid), .InEdges(InEdges), .OutEdge(
        OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(Start), 
        .Clk(Clk) );
    NodeAux_INDEGREE3_SOURCE0 n_3_0 ( .Nid(Nid), .InEdges(InEdges[47:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
endmodule



module Node_NID0_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE1 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID0 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID3 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID4 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID5 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID6 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID7 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID1_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID8 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID9 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID2_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID10 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID11 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID12 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID13 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID14 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID15 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID3_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID16 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID17 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID4_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID18 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID19 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID20 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID21 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID22 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID23 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID24 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID25 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID5_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID26 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID27 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID28 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID29 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID30 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID6_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID31 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID32 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID33 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID34 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID35 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID7_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID36 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID37 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID38 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID39 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID40 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID41 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID8_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID42 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID43 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID9_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID44 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID45 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID10_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID46 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID47 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID48 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID49 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID50 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID51 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID52 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID53 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID11_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID54 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID55 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID56 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID57 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID58 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID12_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID59 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID60 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID61 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID62 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID63 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID64 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID13_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID65 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID14_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID66 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID67 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID68 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID69 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID70 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID71 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID72 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID73 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID15_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID74 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID75 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID76 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID77 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID78 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID79 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID80 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID16_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID81 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID82 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID17_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID83 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID84 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID18_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID85 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID19_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID86 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID87 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID88 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID89 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID20_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID90 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID91 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID92 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID21_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID93 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID94 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID95 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID96 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID97 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID98 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID22_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID99 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID100 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID101 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID102 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID23_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID103 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID24_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID104 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID105 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID106 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID107 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID25_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID108 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID109 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID110 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID26_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID111 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID112 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID113 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID114 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID115 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID27_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID116 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID117 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID118 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID119 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID120 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID121 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID122 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID123 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID28_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID124 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID125 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID126 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID127 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID128 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID129 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID130 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID29_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID131 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID132 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID133 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID134 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID30_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID135 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID136 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID137 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID138 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID139 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID140 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID141 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID31_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID142 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID143 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID144 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID145 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID146 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID147 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID148 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID149 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID32_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID150 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID33_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID151 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID152 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID153 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID154 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID34_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID155 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID156 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID157 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID158 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID159 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID160 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID161 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID35_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID162 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID163 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID164 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID165 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID166 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID167 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID36_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID168 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID169 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID170 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID171 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID172 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID173 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID174 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID37_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID175 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID176 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID177 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID38_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID178 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID39_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID179 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID180 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID181 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID182 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID183 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID184 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID185 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID40_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID186 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID187 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID188 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID189 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID190 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID191 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID192 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID41_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID193 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID194 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID42_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID195 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID196 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID43_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID197 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID198 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID199 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID200 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID201 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID202 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID203 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID204 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID44_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID205 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID206 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID207 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID208 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID45_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID209 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID210 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID211 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID212 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID46_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID213 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID214 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID215 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID216 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID217 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID218 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID47_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID219 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID220 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID221 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID222 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID223 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID48_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID224 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID225 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID226 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID227 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID49_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID228 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID50_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID229 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID230 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID231 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID232 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID51_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID233 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID234 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID235 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID236 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID52_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID237 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID238 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID239 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID240 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID241 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID242 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID243 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID244 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID53_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID245 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID54_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID246 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID247 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID248 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID249 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID250 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID251 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID252 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID253 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID55_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID254 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID255 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID56_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID256 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID257 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID57_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID258 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID259 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID260 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID261 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID262 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID263 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID264 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID265 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID58_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID266 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID267 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID268 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID269 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID270 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID271 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID272 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID273 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID59_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID274 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID275 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID60_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID276 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID277 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID278 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID279 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID280 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID281 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID282 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID61_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID283 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID284 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID285 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID286 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID287 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID62_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID288 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID289 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID290 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID291 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID63_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID292 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID293 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID294 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID295 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID296 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID297 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID64_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID298 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID299 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID300 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID301 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID302 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID303 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID304 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID65_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID305 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID306 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID307 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID308 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID309 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID66_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID310 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID311 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID312 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID313 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID67_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID314 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID68_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID315 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID316 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID317 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID318 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID319 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID320 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID321 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID322 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID69_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID323 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID324 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID325 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID326 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID327 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID328 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID329 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID330 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID70_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID331 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID332 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID71_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID333 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID334 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID335 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID72_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID336 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID337 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID338 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID339 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID340 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID341 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID73_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID342 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID343 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID344 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID345 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID346 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID347 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID348 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID74_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID349 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID350 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID351 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID352 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID353 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID75_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID354 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID355 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID356 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID357 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID358 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID359 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID76_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID360 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID361 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID362 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID363 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID77_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID364 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID365 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID366 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID78_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID367 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID368 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID369 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID370 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID371 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID79_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID372 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID373 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID374 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID375 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID80_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID376 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID377 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID81_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID378 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID379 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID380 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID381 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID382 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID82_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID383 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID384 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID83_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID385 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID386 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID387 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID388 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID84_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID389 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID390 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID391 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID392 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID393 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID85_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID394 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID395 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID396 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID86_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID397 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID398 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID399 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID400 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID87_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID401 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID402 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID403 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID404 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID405 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID406 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID407 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID408 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID88_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID409 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID410 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID89_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID411 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID412 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID90_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID413 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID414 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID415 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID91_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID416 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID417 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID418 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID419 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID92_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID420 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID421 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID422 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID423 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID424 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID425 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID426 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID427 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID93_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID428 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID429 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID430 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID431 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID432 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID433 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID434 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID435 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID94_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID436 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID437 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID438 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID95_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID439 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID440 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID441 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID442 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID443 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID444 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID445 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID446 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID96_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID447 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID97_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID448 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID449 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID450 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID451 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID452 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID453 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID454 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID98_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID455 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID99_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID456 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID457 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID100_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID458 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID459 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID460 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID101_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID461 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID462 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID102_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID463 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID464 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID465 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID466 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID467 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID468 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID469 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID470 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID103_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID471 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID472 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID473 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID474 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID475 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID476 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID477 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID104_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID478 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID479 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID480 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID481 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID482 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID483 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID105_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID484 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID485 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID106_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID486 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID487 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID488 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID489 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID490 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID491 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID107_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID492 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID493 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID494 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID108_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID495 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID496 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID497 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID498 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID109_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID499 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID110_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID500 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID501 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID502 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID503 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID111_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID504 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID505 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID112_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID506 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID507 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID113_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID508 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID509 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID510 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID114_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID511 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID512 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID513 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID514 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID515 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID115_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID516 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID517 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID518 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID116_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID519 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID520 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID521 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID522 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID523 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID117_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID524 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID525 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID526 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID527 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID118_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID528 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID529 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID530 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID531 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID119_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID532 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID533 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID534 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID535 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID536 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID537 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID538 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID539 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID120_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID540 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID541 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID542 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID543 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID544 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID545 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID546 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID547 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID121_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID548 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID549 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID122_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID550 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID551 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID552 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID553 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID554 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID555 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID123_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID556 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID557 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID558 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID559 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID560 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID124_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID561 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID562 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID563 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID564 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID125_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID565 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID566 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID567 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID568 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID569 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID126_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID570 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID571 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID572 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID573 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID127_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID574 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID575 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID576 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID577 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID578 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID128_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID579 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID580 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID581 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID129_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID582 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID130_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID583 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID584 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID585 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID586 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID587 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID588 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID131_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID589 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID590 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID591 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID132_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID592 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID593 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID594 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID595 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID596 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID597 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID598 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID599 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID133_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID600 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID601 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID602 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID603 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID604 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID605 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID606 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID607 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID134_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID608 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID609 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID610 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID611 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID612 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID613 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID614 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID135_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID615 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID616 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID617 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID618 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID619 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID620 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID136_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID621 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID622 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID623 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID624 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID625 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID626 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID627 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID137_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID628 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID138_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID629 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID630 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID631 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID632 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID139_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID633 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID634 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID635 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID636 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID637 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID638 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID140_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID639 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID640 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID641 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID642 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID141_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID643 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID644 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID645 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID646 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID647 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID648 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID649 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID650 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID142_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID651 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID652 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID653 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID654 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID143_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID655 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID656 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID657 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID658 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID659 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID660 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID661 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID662 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID144_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID663 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID664 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID665 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID666 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID667 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID668 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID669 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID145_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID670 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID671 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID672 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID673 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID674 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID675 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID676 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID677 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID146_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID678 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID679 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID147_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID680 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID681 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID148_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID682 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID149_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID683 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID684 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID685 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID686 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID687 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID688 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID689 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID150_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID690 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID691 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID692 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID151_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID693 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID694 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID695 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID696 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID697 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID698 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID699 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID700 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID152_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID701 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID702 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID703 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID704 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID705 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID706 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID707 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID708 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID153_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID709 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID710 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID711 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID712 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID713 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID714 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID715 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID716 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID154_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID717 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID718 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID719 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID720 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID155_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID721 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID722 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID723 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID724 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID725 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID726 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID727 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID156_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID728 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID729 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID730 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID731 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID732 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID733 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID734 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID157_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID735 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID736 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID737 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID738 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID739 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID740 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID741 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID742 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID158_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID743 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID744 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID745 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID159_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID746 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID747 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID748 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID160_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID749 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID750 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID751 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID752 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID753 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID754 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID161_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID755 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID756 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID757 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID758 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID162_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID759 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID760 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID761 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID762 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID763 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID764 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID163_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID765 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID766 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID767 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID768 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID769 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID770 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID771 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID772 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID164_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID773 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID774 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID775 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID776 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID777 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID778 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID165_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID779 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID780 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID781 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID166_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID782 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID783 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID784 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID785 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID167_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID786 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID168_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID787 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID788 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID789 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID790 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID169_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID791 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID792 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID793 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID794 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID170_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID795 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID796 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID171_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID797 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID798 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID799 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID800 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID172_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID801 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID802 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID803 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID804 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID805 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID173_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID806 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID174_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID807 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID808 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID809 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID175_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID810 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID811 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID812 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID176_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID813 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID177_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID814 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID815 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID178_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID816 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID817 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID179_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID818 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID819 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID820 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID821 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID180_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID822 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID823 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID824 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID825 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID826 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID827 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID828 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID829 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID181_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID830 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID831 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID832 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID833 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID834 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID835 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID836 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID182_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID837 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID838 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID183_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID839 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID184_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID840 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID841 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID842 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID843 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID844 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID845 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID185_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID846 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID847 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID848 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID849 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID850 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID851 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID852 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID186_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID853 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID854 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID855 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID856 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID857 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID187_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID858 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID859 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID860 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID861 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID862 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID863 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID864 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID865 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID188_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID866 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID867 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID189_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID868 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID869 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID870 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID871 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID872 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID190_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID873 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID874 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID875 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID876 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID191_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID877 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID878 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID879 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID880 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID192_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID881 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID882 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID883 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID884 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID885 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID193_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID886 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID887 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID888 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID889 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID890 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID891 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID194_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID892 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID893 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID894 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID895 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID195_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID896 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID897 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID196_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID898 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID899 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID197_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID900 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID901 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID902 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID903 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID904 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID905 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID906 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID198_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID907 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID908 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID909 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID199_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID910 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID911 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID912 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID913 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID914 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID915 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID200_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID916 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID917 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID201_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID918 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID202_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID919 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID920 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID203_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID921 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID922 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID923 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID924 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID925 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID926 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID204_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID927 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID928 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID929 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID930 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID205_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID931 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID206_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID932 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID933 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID934 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID935 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID936 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID937 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID207_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID938 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID939 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID940 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID941 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID942 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID943 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID944 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID208_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID945 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID946 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID209_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID947 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID948 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID949 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID950 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID951 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID952 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID953 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID954 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID210_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID955 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID956 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID957 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID211_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID958 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID959 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID960 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID961 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID962 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID963 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID964 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID212_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID965 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID966 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID213_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID967 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID214_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID968 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID969 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID970 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID971 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID972 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID215_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID973 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID974 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID975 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID976 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID216_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID977 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID217_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID978 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID979 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID980 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID981 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID982 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID983 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID218_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID984 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID985 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID219_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID986 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID220_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID987 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID988 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID989 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID990 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID991 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID992 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID221_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID993 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID994 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID995 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID222_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID996 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID997 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID998 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID223_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID999 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1000 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID224_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1001 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1002 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1003 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1004 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1005 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1006 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1007 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID225_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1008 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1009 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1010 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID226_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1011 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1012 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID227_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1013 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1014 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1015 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1016 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1017 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1018 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1019 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID228_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1020 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1021 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1022 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1023 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID229_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1024 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1025 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID230_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1026 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1027 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1028 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1029 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID231_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1030 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1031 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1032 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1033 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1034 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1035 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID232_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1036 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1037 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1038 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1039 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1040 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1041 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID233_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1042 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1043 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1044 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1045 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID234_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1046 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1047 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1048 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1049 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1050 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1051 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID235_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1052 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1053 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1054 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1055 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1056 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1057 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID236_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1058 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1059 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1060 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1061 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1062 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1063 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1064 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1065 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID237_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1066 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1067 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1068 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1069 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID238_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1070 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1071 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID239_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1072 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1073 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1074 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1075 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1076 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID240_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1077 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID241_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1078 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1079 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1080 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID242_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1081 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1082 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1083 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1084 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1085 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1086 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1087 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID243_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1088 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID244_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1089 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1090 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1091 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1092 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1093 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1094 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1095 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1096 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID245_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1097 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1098 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1099 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1100 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1101 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID246_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1102 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID247_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1103 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1104 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1105 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1106 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1107 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1108 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID248_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1109 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1110 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID249_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1111 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1112 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1113 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1114 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1115 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1116 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1117 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID250_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1118 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID251_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1119 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1120 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1121 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID252_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1122 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1123 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1124 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1125 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1126 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1127 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID253_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1128 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1129 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1130 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1131 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID254_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1132 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1133 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID255_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [7:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1134 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1135 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1136 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1137 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1138 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1139 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [10:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module graph ( WeightAddr, WeightData, PathAddr, PathData, Start, Clk );
input  [10:0] WeightAddr;
input  [15:0] WeightData;
input  [7:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire [127:0] In0;
    wire [15:0] Out0;
    wire [31:0] In1;
    wire [15:0] Out1;
    wire [95:0] In2;
    wire [15:0] Out2;
    wire [31:0] In3;
    wire [15:0] Out3;
    wire [127:0] In4;
    wire [15:0] Out4;
    wire [79:0] In5;
    wire [15:0] Out5;
    wire [79:0] In6;
    wire [15:0] Out6;
    wire [95:0] In7;
    wire [15:0] Out7;
    wire [31:0] In8;
    wire [15:0] Out8;
    wire [31:0] In9;
    wire [15:0] Out9;
    wire [127:0] In10;
    wire [15:0] Out10;
    wire [79:0] In11;
    wire [15:0] Out11;
    wire [95:0] In12;
    wire [15:0] Out12;
    wire [15:0] In13;
    wire [15:0] Out13;
    wire [127:0] In14;
    wire [15:0] Out14;
    wire [111:0] In15;
    wire [15:0] Out15;
    wire [31:0] In16;
    wire [15:0] Out16;
    wire [31:0] In17;
    wire [15:0] Out17;
    wire [15:0] In18;
    wire [15:0] Out18;
    wire [63:0] In19;
    wire [15:0] Out19;
    wire [47:0] In20;
    wire [15:0] Out20;
    wire [95:0] In21;
    wire [15:0] Out21;
    wire [63:0] In22;
    wire [15:0] Out22;
    wire [15:0] In23;
    wire [15:0] Out23;
    wire [63:0] In24;
    wire [15:0] Out24;
    wire [47:0] In25;
    wire [15:0] Out25;
    wire [79:0] In26;
    wire [15:0] Out26;
    wire [127:0] In27;
    wire [15:0] Out27;
    wire [111:0] In28;
    wire [15:0] Out28;
    wire [63:0] In29;
    wire [15:0] Out29;
    wire [111:0] In30;
    wire [15:0] Out30;
    wire [127:0] In31;
    wire [15:0] Out31;
    wire [15:0] In32;
    wire [15:0] Out32;
    wire [63:0] In33;
    wire [15:0] Out33;
    wire [111:0] In34;
    wire [15:0] Out34;
    wire [95:0] In35;
    wire [15:0] Out35;
    wire [111:0] In36;
    wire [15:0] Out36;
    wire [47:0] In37;
    wire [15:0] Out37;
    wire [15:0] In38;
    wire [15:0] Out38;
    wire [111:0] In39;
    wire [15:0] Out39;
    wire [111:0] In40;
    wire [15:0] Out40;
    wire [31:0] In41;
    wire [15:0] Out41;
    wire [31:0] In42;
    wire [15:0] Out42;
    wire [127:0] In43;
    wire [15:0] Out43;
    wire [63:0] In44;
    wire [15:0] Out44;
    wire [63:0] In45;
    wire [15:0] Out45;
    wire [95:0] In46;
    wire [15:0] Out46;
    wire [79:0] In47;
    wire [15:0] Out47;
    wire [63:0] In48;
    wire [15:0] Out48;
    wire [15:0] In49;
    wire [15:0] Out49;
    wire [63:0] In50;
    wire [15:0] Out50;
    wire [63:0] In51;
    wire [15:0] Out51;
    wire [127:0] In52;
    wire [15:0] Out52;
    wire [15:0] In53;
    wire [15:0] Out53;
    wire [127:0] In54;
    wire [15:0] Out54;
    wire [31:0] In55;
    wire [15:0] Out55;
    wire [31:0] In56;
    wire [15:0] Out56;
    wire [127:0] In57;
    wire [15:0] Out57;
    wire [127:0] In58;
    wire [15:0] Out58;
    wire [31:0] In59;
    wire [15:0] Out59;
    wire [111:0] In60;
    wire [15:0] Out60;
    wire [79:0] In61;
    wire [15:0] Out61;
    wire [63:0] In62;
    wire [15:0] Out62;
    wire [95:0] In63;
    wire [15:0] Out63;
    wire [111:0] In64;
    wire [15:0] Out64;
    wire [79:0] In65;
    wire [15:0] Out65;
    wire [63:0] In66;
    wire [15:0] Out66;
    wire [15:0] In67;
    wire [15:0] Out67;
    wire [127:0] In68;
    wire [15:0] Out68;
    wire [127:0] In69;
    wire [15:0] Out69;
    wire [31:0] In70;
    wire [15:0] Out70;
    wire [47:0] In71;
    wire [15:0] Out71;
    wire [95:0] In72;
    wire [15:0] Out72;
    wire [111:0] In73;
    wire [15:0] Out73;
    wire [79:0] In74;
    wire [15:0] Out74;
    wire [95:0] In75;
    wire [15:0] Out75;
    wire [63:0] In76;
    wire [15:0] Out76;
    wire [47:0] In77;
    wire [15:0] Out77;
    wire [79:0] In78;
    wire [15:0] Out78;
    wire [63:0] In79;
    wire [15:0] Out79;
    wire [31:0] In80;
    wire [15:0] Out80;
    wire [79:0] In81;
    wire [15:0] Out81;
    wire [31:0] In82;
    wire [15:0] Out82;
    wire [63:0] In83;
    wire [15:0] Out83;
    wire [79:0] In84;
    wire [15:0] Out84;
    wire [47:0] In85;
    wire [15:0] Out85;
    wire [63:0] In86;
    wire [15:0] Out86;
    wire [127:0] In87;
    wire [15:0] Out87;
    wire [31:0] In88;
    wire [15:0] Out88;
    wire [31:0] In89;
    wire [15:0] Out89;
    wire [47:0] In90;
    wire [15:0] Out90;
    wire [63:0] In91;
    wire [15:0] Out91;
    wire [127:0] In92;
    wire [15:0] Out92;
    wire [127:0] In93;
    wire [15:0] Out93;
    wire [47:0] In94;
    wire [15:0] Out94;
    wire [127:0] In95;
    wire [15:0] Out95;
    wire [15:0] In96;
    wire [15:0] Out96;
    wire [111:0] In97;
    wire [15:0] Out97;
    wire [15:0] In98;
    wire [15:0] Out98;
    wire [31:0] In99;
    wire [15:0] Out99;
    wire [47:0] In100;
    wire [15:0] Out100;
    wire [31:0] In101;
    wire [15:0] Out101;
    wire [127:0] In102;
    wire [15:0] Out102;
    wire [111:0] In103;
    wire [15:0] Out103;
    wire [95:0] In104;
    wire [15:0] Out104;
    wire [31:0] In105;
    wire [15:0] Out105;
    wire [95:0] In106;
    wire [15:0] Out106;
    wire [47:0] In107;
    wire [15:0] Out107;
    wire [63:0] In108;
    wire [15:0] Out108;
    wire [15:0] In109;
    wire [15:0] Out109;
    wire [63:0] In110;
    wire [15:0] Out110;
    wire [31:0] In111;
    wire [15:0] Out111;
    wire [31:0] In112;
    wire [15:0] Out112;
    wire [47:0] In113;
    wire [15:0] Out113;
    wire [79:0] In114;
    wire [15:0] Out114;
    wire [47:0] In115;
    wire [15:0] Out115;
    wire [79:0] In116;
    wire [15:0] Out116;
    wire [63:0] In117;
    wire [15:0] Out117;
    wire [63:0] In118;
    wire [15:0] Out118;
    wire [127:0] In119;
    wire [15:0] Out119;
    wire [127:0] In120;
    wire [15:0] Out120;
    wire [31:0] In121;
    wire [15:0] Out121;
    wire [95:0] In122;
    wire [15:0] Out122;
    wire [79:0] In123;
    wire [15:0] Out123;
    wire [63:0] In124;
    wire [15:0] Out124;
    wire [79:0] In125;
    wire [15:0] Out125;
    wire [63:0] In126;
    wire [15:0] Out126;
    wire [79:0] In127;
    wire [15:0] Out127;
    wire [47:0] In128;
    wire [15:0] Out128;
    wire [15:0] In129;
    wire [15:0] Out129;
    wire [95:0] In130;
    wire [15:0] Out130;
    wire [47:0] In131;
    wire [15:0] Out131;
    wire [127:0] In132;
    wire [15:0] Out132;
    wire [127:0] In133;
    wire [15:0] Out133;
    wire [111:0] In134;
    wire [15:0] Out134;
    wire [95:0] In135;
    wire [15:0] Out135;
    wire [111:0] In136;
    wire [15:0] Out136;
    wire [15:0] In137;
    wire [15:0] Out137;
    wire [63:0] In138;
    wire [15:0] Out138;
    wire [95:0] In139;
    wire [15:0] Out139;
    wire [63:0] In140;
    wire [15:0] Out140;
    wire [127:0] In141;
    wire [15:0] Out141;
    wire [63:0] In142;
    wire [15:0] Out142;
    wire [127:0] In143;
    wire [15:0] Out143;
    wire [111:0] In144;
    wire [15:0] Out144;
    wire [127:0] In145;
    wire [15:0] Out145;
    wire [31:0] In146;
    wire [15:0] Out146;
    wire [31:0] In147;
    wire [15:0] Out147;
    wire [15:0] In148;
    wire [15:0] Out148;
    wire [111:0] In149;
    wire [15:0] Out149;
    wire [47:0] In150;
    wire [15:0] Out150;
    wire [127:0] In151;
    wire [15:0] Out151;
    wire [127:0] In152;
    wire [15:0] Out152;
    wire [127:0] In153;
    wire [15:0] Out153;
    wire [63:0] In154;
    wire [15:0] Out154;
    wire [111:0] In155;
    wire [15:0] Out155;
    wire [111:0] In156;
    wire [15:0] Out156;
    wire [127:0] In157;
    wire [15:0] Out157;
    wire [47:0] In158;
    wire [15:0] Out158;
    wire [47:0] In159;
    wire [15:0] Out159;
    wire [95:0] In160;
    wire [15:0] Out160;
    wire [63:0] In161;
    wire [15:0] Out161;
    wire [95:0] In162;
    wire [15:0] Out162;
    wire [127:0] In163;
    wire [15:0] Out163;
    wire [95:0] In164;
    wire [15:0] Out164;
    wire [47:0] In165;
    wire [15:0] Out165;
    wire [63:0] In166;
    wire [15:0] Out166;
    wire [15:0] In167;
    wire [15:0] Out167;
    wire [63:0] In168;
    wire [15:0] Out168;
    wire [63:0] In169;
    wire [15:0] Out169;
    wire [31:0] In170;
    wire [15:0] Out170;
    wire [63:0] In171;
    wire [15:0] Out171;
    wire [79:0] In172;
    wire [15:0] Out172;
    wire [15:0] In173;
    wire [15:0] Out173;
    wire [47:0] In174;
    wire [15:0] Out174;
    wire [47:0] In175;
    wire [15:0] Out175;
    wire [15:0] In176;
    wire [15:0] Out176;
    wire [31:0] In177;
    wire [15:0] Out177;
    wire [31:0] In178;
    wire [15:0] Out178;
    wire [63:0] In179;
    wire [15:0] Out179;
    wire [127:0] In180;
    wire [15:0] Out180;
    wire [111:0] In181;
    wire [15:0] Out181;
    wire [31:0] In182;
    wire [15:0] Out182;
    wire [15:0] In183;
    wire [15:0] Out183;
    wire [95:0] In184;
    wire [15:0] Out184;
    wire [111:0] In185;
    wire [15:0] Out185;
    wire [79:0] In186;
    wire [15:0] Out186;
    wire [127:0] In187;
    wire [15:0] Out187;
    wire [31:0] In188;
    wire [15:0] Out188;
    wire [79:0] In189;
    wire [15:0] Out189;
    wire [63:0] In190;
    wire [15:0] Out190;
    wire [63:0] In191;
    wire [15:0] Out191;
    wire [79:0] In192;
    wire [15:0] Out192;
    wire [95:0] In193;
    wire [15:0] Out193;
    wire [63:0] In194;
    wire [15:0] Out194;
    wire [31:0] In195;
    wire [15:0] Out195;
    wire [31:0] In196;
    wire [15:0] Out196;
    wire [111:0] In197;
    wire [15:0] Out197;
    wire [47:0] In198;
    wire [15:0] Out198;
    wire [95:0] In199;
    wire [15:0] Out199;
    wire [31:0] In200;
    wire [15:0] Out200;
    wire [15:0] In201;
    wire [15:0] Out201;
    wire [31:0] In202;
    wire [15:0] Out202;
    wire [95:0] In203;
    wire [15:0] Out203;
    wire [63:0] In204;
    wire [15:0] Out204;
    wire [15:0] In205;
    wire [15:0] Out205;
    wire [95:0] In206;
    wire [15:0] Out206;
    wire [111:0] In207;
    wire [15:0] Out207;
    wire [31:0] In208;
    wire [15:0] Out208;
    wire [127:0] In209;
    wire [15:0] Out209;
    wire [47:0] In210;
    wire [15:0] Out210;
    wire [111:0] In211;
    wire [15:0] Out211;
    wire [31:0] In212;
    wire [15:0] Out212;
    wire [15:0] In213;
    wire [15:0] Out213;
    wire [79:0] In214;
    wire [15:0] Out214;
    wire [63:0] In215;
    wire [15:0] Out215;
    wire [15:0] In216;
    wire [15:0] Out216;
    wire [95:0] In217;
    wire [15:0] Out217;
    wire [31:0] In218;
    wire [15:0] Out218;
    wire [15:0] In219;
    wire [15:0] Out219;
    wire [95:0] In220;
    wire [15:0] Out220;
    wire [47:0] In221;
    wire [15:0] Out221;
    wire [47:0] In222;
    wire [15:0] Out222;
    wire [31:0] In223;
    wire [15:0] Out223;
    wire [111:0] In224;
    wire [15:0] Out224;
    wire [47:0] In225;
    wire [15:0] Out225;
    wire [31:0] In226;
    wire [15:0] Out226;
    wire [111:0] In227;
    wire [15:0] Out227;
    wire [63:0] In228;
    wire [15:0] Out228;
    wire [31:0] In229;
    wire [15:0] Out229;
    wire [63:0] In230;
    wire [15:0] Out230;
    wire [95:0] In231;
    wire [15:0] Out231;
    wire [95:0] In232;
    wire [15:0] Out232;
    wire [63:0] In233;
    wire [15:0] Out233;
    wire [95:0] In234;
    wire [15:0] Out234;
    wire [95:0] In235;
    wire [15:0] Out235;
    wire [127:0] In236;
    wire [15:0] Out236;
    wire [63:0] In237;
    wire [15:0] Out237;
    wire [31:0] In238;
    wire [15:0] Out238;
    wire [79:0] In239;
    wire [15:0] Out239;
    wire [15:0] In240;
    wire [15:0] Out240;
    wire [47:0] In241;
    wire [15:0] Out241;
    wire [111:0] In242;
    wire [15:0] Out242;
    wire [15:0] In243;
    wire [15:0] Out243;
    wire [127:0] In244;
    wire [15:0] Out244;
    wire [79:0] In245;
    wire [15:0] Out245;
    wire [15:0] In246;
    wire [15:0] Out246;
    wire [95:0] In247;
    wire [15:0] Out247;
    wire [31:0] In248;
    wire [15:0] Out248;
    wire [111:0] In249;
    wire [15:0] Out249;
    wire [15:0] In250;
    wire [15:0] Out250;
    wire [47:0] In251;
    wire [15:0] Out251;
    wire [95:0] In252;
    wire [15:0] Out252;
    wire [63:0] In253;
    wire [15:0] Out253;
    wire [31:0] In254;
    wire [15:0] Out254;
    wire [95:0] In255;
    wire [15:0] Out255;

    Node_NID0_INDEGREE8 n0 ( .InEdges(In0), .OutEdge(Out0),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID0 e0 ( .InEdge(Out23), .OutEdge(In0[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1 e1 ( .InEdge(Out179), .OutEdge(In0[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2 e2 ( .InEdge(Out140), .OutEdge(In0[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID3 e3 ( .InEdge(Out152), .OutEdge(In0[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID4 e4 ( .InEdge(Out67), .OutEdge(In0[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID5 e5 ( .InEdge(Out216), .OutEdge(In0[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID6 e6 ( .InEdge(Out130), .OutEdge(In0[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID7 e7 ( .InEdge(Out217), .OutEdge(In0[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID1_INDEGREE2 n1 ( .InEdges(In1), .OutEdge(Out1),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID8 e8 ( .InEdge(Out17), .OutEdge(In1[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID9 e9 ( .InEdge(Out84), .OutEdge(In1[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID2_INDEGREE6 n2 ( .InEdges(In2), .OutEdge(Out2),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID10 e10 ( .InEdge(Out98), .OutEdge(In2[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID11 e11 ( .InEdge(Out72), .OutEdge(In2[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID12 e12 ( .InEdge(Out153), .OutEdge(In2[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID13 e13 ( .InEdge(Out136), .OutEdge(In2[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID14 e14 ( .InEdge(Out107), .OutEdge(In2[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID15 e15 ( .InEdge(Out88), .OutEdge(In2[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID3_INDEGREE2 n3 ( .InEdges(In3), .OutEdge(Out3),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID16 e16 ( .InEdge(Out229), .OutEdge(In3[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID17 e17 ( .InEdge(Out13), .OutEdge(In3[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID4_INDEGREE8 n4 ( .InEdges(In4), .OutEdge(Out4),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID18 e18 ( .InEdge(Out156), .OutEdge(In4[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID19 e19 ( .InEdge(Out20), .OutEdge(In4[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID20 e20 ( .InEdge(Out132), .OutEdge(In4[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID21 e21 ( .InEdge(Out57), .OutEdge(In4[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID22 e22 ( .InEdge(Out2), .OutEdge(In4[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID23 e23 ( .InEdge(Out12), .OutEdge(In4[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID24 e24 ( .InEdge(Out237), .OutEdge(In4[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID25 e25 ( .InEdge(Out209), .OutEdge(In4[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID5_INDEGREE5 n5 ( .InEdges(In5), .OutEdge(Out5),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID26 e26 ( .InEdge(Out176), .OutEdge(In5[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID27 e27 ( .InEdge(Out197), .OutEdge(In5[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID28 e28 ( .InEdge(Out72), .OutEdge(In5[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID29 e29 ( .InEdge(Out202), .OutEdge(In5[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID30 e30 ( .InEdge(Out103), .OutEdge(In5[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID6_INDEGREE5 n6 ( .InEdges(In6), .OutEdge(Out6),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID31 e31 ( .InEdge(Out161), .OutEdge(In6[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID32 e32 ( .InEdge(Out247), .OutEdge(In6[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID33 e33 ( .InEdge(Out57), .OutEdge(In6[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID34 e34 ( .InEdge(Out155), .OutEdge(In6[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID35 e35 ( .InEdge(Out138), .OutEdge(In6[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID7_INDEGREE6 n7 ( .InEdges(In7), .OutEdge(Out7),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID36 e36 ( .InEdge(Out195), .OutEdge(In7[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID37 e37 ( .InEdge(Out250), .OutEdge(In7[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID38 e38 ( .InEdge(Out228), .OutEdge(In7[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID39 e39 ( .InEdge(Out243), .OutEdge(In7[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID40 e40 ( .InEdge(Out165), .OutEdge(In7[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID41 e41 ( .InEdge(Out254), .OutEdge(In7[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID8_INDEGREE2 n8 ( .InEdges(In8), .OutEdge(Out8),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID42 e42 ( .InEdge(Out12), .OutEdge(In8[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID43 e43 ( .InEdge(Out32), .OutEdge(In8[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID9_INDEGREE2 n9 ( .InEdges(In9), .OutEdge(Out9),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID44 e44 ( .InEdge(Out97), .OutEdge(In9[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID45 e45 ( .InEdge(Out152), .OutEdge(In9[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID10_INDEGREE8 n10 ( .InEdges(In10), .OutEdge(Out10),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID46 e46 ( .InEdge(Out192), .OutEdge(In10[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID47 e47 ( .InEdge(Out30), .OutEdge(In10[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID48 e48 ( .InEdge(Out195), .OutEdge(In10[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID49 e49 ( .InEdge(Out129), .OutEdge(In10[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID50 e50 ( .InEdge(Out233), .OutEdge(In10[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID51 e51 ( .InEdge(Out54), .OutEdge(In10[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID52 e52 ( .InEdge(Out25), .OutEdge(In10[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID53 e53 ( .InEdge(Out161), .OutEdge(In10[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID11_INDEGREE5 n11 ( .InEdges(In11), .OutEdge(Out11),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID54 e54 ( .InEdge(Out246), .OutEdge(In11[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID55 e55 ( .InEdge(Out178), .OutEdge(In11[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID56 e56 ( .InEdge(Out80), .OutEdge(In11[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID57 e57 ( .InEdge(Out200), .OutEdge(In11[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID58 e58 ( .InEdge(Out85), .OutEdge(In11[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID12_INDEGREE6 n12 ( .InEdges(In12), .OutEdge(Out12),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID59 e59 ( .InEdge(Out97), .OutEdge(In12[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID60 e60 ( .InEdge(Out31), .OutEdge(In12[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID61 e61 ( .InEdge(Out189), .OutEdge(In12[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID62 e62 ( .InEdge(Out136), .OutEdge(In12[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID63 e63 ( .InEdge(Out221), .OutEdge(In12[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID64 e64 ( .InEdge(Out76), .OutEdge(In12[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID13_INDEGREE1 n13 ( .InEdges(In13), .OutEdge(Out13),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID65 e65 ( .InEdge(Out120), .OutEdge(In13[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID14_INDEGREE8 n14 ( .InEdges(In14), .OutEdge(Out14),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID66 e66 ( .InEdge(Out70), .OutEdge(In14[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID67 e67 ( .InEdge(Out245), .OutEdge(In14[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID68 e68 ( .InEdge(Out91), .OutEdge(In14[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID69 e69 ( .InEdge(Out41), .OutEdge(In14[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID70 e70 ( .InEdge(Out161), .OutEdge(In14[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID71 e71 ( .InEdge(Out94), .OutEdge(In14[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID72 e72 ( .InEdge(Out7), .OutEdge(In14[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID73 e73 ( .InEdge(Out52), .OutEdge(In14[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID15_INDEGREE7 n15 ( .InEdges(In15), .OutEdge(Out15),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID74 e74 ( .InEdge(Out83), .OutEdge(In15[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID75 e75 ( .InEdge(Out135), .OutEdge(In15[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID76 e76 ( .InEdge(Out230), .OutEdge(In15[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID77 e77 ( .InEdge(Out18), .OutEdge(In15[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID78 e78 ( .InEdge(Out2), .OutEdge(In15[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID79 e79 ( .InEdge(Out54), .OutEdge(In15[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID80 e80 ( .InEdge(Out196), .OutEdge(In15[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID16_INDEGREE2 n16 ( .InEdges(In16), .OutEdge(Out16),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID81 e81 ( .InEdge(Out79), .OutEdge(In16[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID82 e82 ( .InEdge(Out8), .OutEdge(In16[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID17_INDEGREE2 n17 ( .InEdges(In17), .OutEdge(Out17),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID83 e83 ( .InEdge(Out180), .OutEdge(In17[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID84 e84 ( .InEdge(Out101), .OutEdge(In17[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID18_INDEGREE1 n18 ( .InEdges(In18), .OutEdge(Out18),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID85 e85 ( .InEdge(Out183), .OutEdge(In18[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID19_INDEGREE4 n19 ( .InEdges(In19), .OutEdge(Out19),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID86 e86 ( .InEdge(Out79), .OutEdge(In19[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID87 e87 ( .InEdge(Out24), .OutEdge(In19[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID88 e88 ( .InEdge(Out235), .OutEdge(In19[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID89 e89 ( .InEdge(Out238), .OutEdge(In19[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID20_INDEGREE3 n20 ( .InEdges(In20), .OutEdge(Out20),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID90 e90 ( .InEdge(Out173), .OutEdge(In20[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID91 e91 ( .InEdge(Out223), .OutEdge(In20[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID92 e92 ( .InEdge(Out140), .OutEdge(In20[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID21_INDEGREE6 n21 ( .InEdges(In21), .OutEdge(Out21),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID93 e93 ( .InEdge(Out140), .OutEdge(In21[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID94 e94 ( .InEdge(Out177), .OutEdge(In21[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID95 e95 ( .InEdge(Out33), .OutEdge(In21[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID96 e96 ( .InEdge(Out3), .OutEdge(In21[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID97 e97 ( .InEdge(Out58), .OutEdge(In21[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID98 e98 ( .InEdge(Out51), .OutEdge(In21[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID22_INDEGREE4 n22 ( .InEdges(In22), .OutEdge(Out22),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID99 e99 ( .InEdge(Out72), .OutEdge(In22[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID100 e100 ( .InEdge(Out140), .OutEdge(In22[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID101 e101 ( .InEdge(Out242), .OutEdge(In22[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID102 e102 ( .InEdge(Out47), .OutEdge(In22[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID23_INDEGREE1 n23 ( .InEdges(In23), .OutEdge(Out23),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID103 e103 ( .InEdge(Out72), .OutEdge(In23[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID24_INDEGREE4 n24 ( .InEdges(In24), .OutEdge(Out24),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID104 e104 ( .InEdge(Out215), .OutEdge(In24[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID105 e105 ( .InEdge(Out128), .OutEdge(In24[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID106 e106 ( .InEdge(Out113), .OutEdge(In24[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID107 e107 ( .InEdge(Out79), .OutEdge(In24[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID25_INDEGREE3 n25 ( .InEdges(In25), .OutEdge(Out25),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID108 e108 ( .InEdge(Out155), .OutEdge(In25[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID109 e109 ( .InEdge(Out196), .OutEdge(In25[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID110 e110 ( .InEdge(Out158), .OutEdge(In25[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID26_INDEGREE5 n26 ( .InEdges(In26), .OutEdge(Out26),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID111 e111 ( .InEdge(Out27), .OutEdge(In26[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID112 e112 ( .InEdge(Out115), .OutEdge(In26[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID113 e113 ( .InEdge(Out147), .OutEdge(In26[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID114 e114 ( .InEdge(Out171), .OutEdge(In26[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID115 e115 ( .InEdge(Out232), .OutEdge(In26[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID27_INDEGREE8 n27 ( .InEdges(In27), .OutEdge(Out27),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID116 e116 ( .InEdge(Out232), .OutEdge(In27[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID117 e117 ( .InEdge(Out149), .OutEdge(In27[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID118 e118 ( .InEdge(Out240), .OutEdge(In27[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID119 e119 ( .InEdge(Out21), .OutEdge(In27[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID120 e120 ( .InEdge(Out185), .OutEdge(In27[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID121 e121 ( .InEdge(Out100), .OutEdge(In27[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID122 e122 ( .InEdge(Out87), .OutEdge(In27[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID123 e123 ( .InEdge(Out196), .OutEdge(In27[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID28_INDEGREE7 n28 ( .InEdges(In28), .OutEdge(Out28),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID124 e124 ( .InEdge(Out57), .OutEdge(In28[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID125 e125 ( .InEdge(Out1), .OutEdge(In28[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID126 e126 ( .InEdge(Out50), .OutEdge(In28[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID127 e127 ( .InEdge(Out252), .OutEdge(In28[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID128 e128 ( .InEdge(Out104), .OutEdge(In28[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID129 e129 ( .InEdge(Out250), .OutEdge(In28[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID130 e130 ( .InEdge(Out24), .OutEdge(In28[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID29_INDEGREE4 n29 ( .InEdges(In29), .OutEdge(Out29),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID131 e131 ( .InEdge(Out248), .OutEdge(In29[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID132 e132 ( .InEdge(Out104), .OutEdge(In29[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID133 e133 ( .InEdge(Out202), .OutEdge(In29[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID134 e134 ( .InEdge(Out31), .OutEdge(In29[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID30_INDEGREE7 n30 ( .InEdges(In30), .OutEdge(Out30),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID135 e135 ( .InEdge(Out157), .OutEdge(In30[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID136 e136 ( .InEdge(Out26), .OutEdge(In30[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID137 e137 ( .InEdge(Out37), .OutEdge(In30[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID138 e138 ( .InEdge(Out219), .OutEdge(In30[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID139 e139 ( .InEdge(Out200), .OutEdge(In30[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID140 e140 ( .InEdge(Out202), .OutEdge(In30[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID141 e141 ( .InEdge(Out152), .OutEdge(In30[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID31_INDEGREE8 n31 ( .InEdges(In31), .OutEdge(Out31),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID142 e142 ( .InEdge(Out222), .OutEdge(In31[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID143 e143 ( .InEdge(Out157), .OutEdge(In31[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID144 e144 ( .InEdge(Out60), .OutEdge(In31[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID145 e145 ( .InEdge(Out197), .OutEdge(In31[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID146 e146 ( .InEdge(Out58), .OutEdge(In31[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID147 e147 ( .InEdge(Out175), .OutEdge(In31[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID148 e148 ( .InEdge(Out25), .OutEdge(In31[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID149 e149 ( .InEdge(Out38), .OutEdge(In31[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID32_INDEGREE1 n32 ( .InEdges(In32), .OutEdge(Out32),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID150 e150 ( .InEdge(Out96), .OutEdge(In32[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID33_INDEGREE4 n33 ( .InEdges(In33), .OutEdge(Out33),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID151 e151 ( .InEdge(Out96), .OutEdge(In33[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID152 e152 ( .InEdge(Out179), .OutEdge(In33[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID153 e153 ( .InEdge(Out195), .OutEdge(In33[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID154 e154 ( .InEdge(Out232), .OutEdge(In33[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID34_INDEGREE7 n34 ( .InEdges(In34), .OutEdge(Out34),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID155 e155 ( .InEdge(Out118), .OutEdge(In34[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID156 e156 ( .InEdge(Out247), .OutEdge(In34[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID157 e157 ( .InEdge(Out185), .OutEdge(In34[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID158 e158 ( .InEdge(Out98), .OutEdge(In34[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID159 e159 ( .InEdge(Out16), .OutEdge(In34[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID160 e160 ( .InEdge(Out2), .OutEdge(In34[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID161 e161 ( .InEdge(Out201), .OutEdge(In34[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID35_INDEGREE6 n35 ( .InEdges(In35), .OutEdge(Out35),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID162 e162 ( .InEdge(Out3), .OutEdge(In35[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID163 e163 ( .InEdge(Out129), .OutEdge(In35[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID164 e164 ( .InEdge(Out127), .OutEdge(In35[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID165 e165 ( .InEdge(Out135), .OutEdge(In35[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID166 e166 ( .InEdge(Out163), .OutEdge(In35[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID167 e167 ( .InEdge(Out219), .OutEdge(In35[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID36_INDEGREE7 n36 ( .InEdges(In36), .OutEdge(Out36),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID168 e168 ( .InEdge(Out5), .OutEdge(In36[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID169 e169 ( .InEdge(Out12), .OutEdge(In36[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID170 e170 ( .InEdge(Out32), .OutEdge(In36[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID171 e171 ( .InEdge(Out238), .OutEdge(In36[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID172 e172 ( .InEdge(Out113), .OutEdge(In36[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID173 e173 ( .InEdge(Out237), .OutEdge(In36[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID174 e174 ( .InEdge(Out112), .OutEdge(In36[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID37_INDEGREE3 n37 ( .InEdges(In37), .OutEdge(Out37),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID175 e175 ( .InEdge(Out71), .OutEdge(In37[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID176 e176 ( .InEdge(Out62), .OutEdge(In37[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID177 e177 ( .InEdge(Out244), .OutEdge(In37[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID38_INDEGREE1 n38 ( .InEdges(In38), .OutEdge(Out38),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID178 e178 ( .InEdge(Out141), .OutEdge(In38[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID39_INDEGREE7 n39 ( .InEdges(In39), .OutEdge(Out39),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID179 e179 ( .InEdge(Out27), .OutEdge(In39[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID180 e180 ( .InEdge(Out238), .OutEdge(In39[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID181 e181 ( .InEdge(Out187), .OutEdge(In39[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID182 e182 ( .InEdge(Out163), .OutEdge(In39[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID183 e183 ( .InEdge(Out146), .OutEdge(In39[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID184 e184 ( .InEdge(Out231), .OutEdge(In39[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID185 e185 ( .InEdge(Out35), .OutEdge(In39[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID40_INDEGREE7 n40 ( .InEdges(In40), .OutEdge(Out40),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID186 e186 ( .InEdge(Out175), .OutEdge(In40[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID187 e187 ( .InEdge(Out116), .OutEdge(In40[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID188 e188 ( .InEdge(Out150), .OutEdge(In40[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID189 e189 ( .InEdge(Out8), .OutEdge(In40[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID190 e190 ( .InEdge(Out240), .OutEdge(In40[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID191 e191 ( .InEdge(Out84), .OutEdge(In40[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID192 e192 ( .InEdge(Out56), .OutEdge(In40[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID41_INDEGREE2 n41 ( .InEdges(In41), .OutEdge(Out41),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID193 e193 ( .InEdge(Out106), .OutEdge(In41[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID194 e194 ( .InEdge(Out136), .OutEdge(In41[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID42_INDEGREE2 n42 ( .InEdges(In42), .OutEdge(Out42),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID195 e195 ( .InEdge(Out28), .OutEdge(In42[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID196 e196 ( .InEdge(Out88), .OutEdge(In42[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID43_INDEGREE8 n43 ( .InEdges(In43), .OutEdge(Out43),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID197 e197 ( .InEdge(Out134), .OutEdge(In43[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID198 e198 ( .InEdge(Out29), .OutEdge(In43[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID199 e199 ( .InEdge(Out17), .OutEdge(In43[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID200 e200 ( .InEdge(Out10), .OutEdge(In43[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID201 e201 ( .InEdge(Out63), .OutEdge(In43[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID202 e202 ( .InEdge(Out219), .OutEdge(In43[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID203 e203 ( .InEdge(Out78), .OutEdge(In43[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID204 e204 ( .InEdge(Out181), .OutEdge(In43[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID44_INDEGREE4 n44 ( .InEdges(In44), .OutEdge(Out44),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID205 e205 ( .InEdge(Out235), .OutEdge(In44[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID206 e206 ( .InEdge(Out31), .OutEdge(In44[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID207 e207 ( .InEdge(Out238), .OutEdge(In44[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID208 e208 ( .InEdge(Out11), .OutEdge(In44[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID45_INDEGREE4 n45 ( .InEdges(In45), .OutEdge(Out45),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID209 e209 ( .InEdge(Out70), .OutEdge(In45[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID210 e210 ( .InEdge(Out18), .OutEdge(In45[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID211 e211 ( .InEdge(Out125), .OutEdge(In45[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID212 e212 ( .InEdge(Out9), .OutEdge(In45[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID46_INDEGREE6 n46 ( .InEdges(In46), .OutEdge(Out46),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID213 e213 ( .InEdge(Out136), .OutEdge(In46[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID214 e214 ( .InEdge(Out126), .OutEdge(In46[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID215 e215 ( .InEdge(Out109), .OutEdge(In46[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID216 e216 ( .InEdge(Out217), .OutEdge(In46[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID217 e217 ( .InEdge(Out119), .OutEdge(In46[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID218 e218 ( .InEdge(Out252), .OutEdge(In46[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID47_INDEGREE5 n47 ( .InEdges(In47), .OutEdge(Out47),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID219 e219 ( .InEdge(Out117), .OutEdge(In47[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID220 e220 ( .InEdge(Out59), .OutEdge(In47[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID221 e221 ( .InEdge(Out179), .OutEdge(In47[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID222 e222 ( .InEdge(Out4), .OutEdge(In47[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID223 e223 ( .InEdge(Out24), .OutEdge(In47[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID48_INDEGREE4 n48 ( .InEdges(In48), .OutEdge(Out48),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID224 e224 ( .InEdge(Out144), .OutEdge(In48[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID225 e225 ( .InEdge(Out173), .OutEdge(In48[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID226 e226 ( .InEdge(Out80), .OutEdge(In48[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID227 e227 ( .InEdge(Out27), .OutEdge(In48[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID49_INDEGREE1 n49 ( .InEdges(In49), .OutEdge(Out49),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID228 e228 ( .InEdge(Out61), .OutEdge(In49[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID50_INDEGREE4 n50 ( .InEdges(In50), .OutEdge(Out50),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID229 e229 ( .InEdge(Out203), .OutEdge(In50[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID230 e230 ( .InEdge(Out191), .OutEdge(In50[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID231 e231 ( .InEdge(Out218), .OutEdge(In50[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID232 e232 ( .InEdge(Out79), .OutEdge(In50[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID51_INDEGREE4 n51 ( .InEdges(In51), .OutEdge(Out51),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID233 e233 ( .InEdge(Out213), .OutEdge(In51[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID234 e234 ( .InEdge(Out169), .OutEdge(In51[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID235 e235 ( .InEdge(Out179), .OutEdge(In51[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID236 e236 ( .InEdge(Out28), .OutEdge(In51[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID52_INDEGREE8 n52 ( .InEdges(In52), .OutEdge(Out52),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID237 e237 ( .InEdge(Out64), .OutEdge(In52[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID238 e238 ( .InEdge(Out9), .OutEdge(In52[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID239 e239 ( .InEdge(Out135), .OutEdge(In52[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID240 e240 ( .InEdge(Out229), .OutEdge(In52[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID241 e241 ( .InEdge(Out209), .OutEdge(In52[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID242 e242 ( .InEdge(Out126), .OutEdge(In52[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID243 e243 ( .InEdge(Out233), .OutEdge(In52[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID244 e244 ( .InEdge(Out76), .OutEdge(In52[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID53_INDEGREE1 n53 ( .InEdges(In53), .OutEdge(Out53),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID245 e245 ( .InEdge(Out128), .OutEdge(In53[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID54_INDEGREE8 n54 ( .InEdges(In54), .OutEdge(Out54),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID246 e246 ( .InEdge(Out14), .OutEdge(In54[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID247 e247 ( .InEdge(Out254), .OutEdge(In54[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID248 e248 ( .InEdge(Out51), .OutEdge(In54[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID249 e249 ( .InEdge(Out122), .OutEdge(In54[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID250 e250 ( .InEdge(Out56), .OutEdge(In54[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID251 e251 ( .InEdge(Out59), .OutEdge(In54[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID252 e252 ( .InEdge(Out104), .OutEdge(In54[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID253 e253 ( .InEdge(Out188), .OutEdge(In54[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID55_INDEGREE2 n55 ( .InEdges(In55), .OutEdge(Out55),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID254 e254 ( .InEdge(Out54), .OutEdge(In55[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID255 e255 ( .InEdge(Out129), .OutEdge(In55[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID56_INDEGREE2 n56 ( .InEdges(In56), .OutEdge(Out56),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID256 e256 ( .InEdge(Out210), .OutEdge(In56[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID257 e257 ( .InEdge(Out140), .OutEdge(In56[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID57_INDEGREE8 n57 ( .InEdges(In57), .OutEdge(Out57),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID258 e258 ( .InEdge(Out22), .OutEdge(In57[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID259 e259 ( .InEdge(Out99), .OutEdge(In57[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID260 e260 ( .InEdge(Out84), .OutEdge(In57[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID261 e261 ( .InEdge(Out20), .OutEdge(In57[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID262 e262 ( .InEdge(Out209), .OutEdge(In57[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID263 e263 ( .InEdge(Out139), .OutEdge(In57[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID264 e264 ( .InEdge(Out12), .OutEdge(In57[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID265 e265 ( .InEdge(Out250), .OutEdge(In57[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID58_INDEGREE8 n58 ( .InEdges(In58), .OutEdge(Out58),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID266 e266 ( .InEdge(Out110), .OutEdge(In58[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID267 e267 ( .InEdge(Out37), .OutEdge(In58[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID268 e268 ( .InEdge(Out91), .OutEdge(In58[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID269 e269 ( .InEdge(Out89), .OutEdge(In58[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID270 e270 ( .InEdge(Out93), .OutEdge(In58[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID271 e271 ( .InEdge(Out127), .OutEdge(In58[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID272 e272 ( .InEdge(Out61), .OutEdge(In58[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID273 e273 ( .InEdge(Out134), .OutEdge(In58[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID59_INDEGREE2 n59 ( .InEdges(In59), .OutEdge(Out59),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID274 e274 ( .InEdge(Out177), .OutEdge(In59[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID275 e275 ( .InEdge(Out97), .OutEdge(In59[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID60_INDEGREE7 n60 ( .InEdges(In60), .OutEdge(Out60),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID276 e276 ( .InEdge(Out40), .OutEdge(In60[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID277 e277 ( .InEdge(Out75), .OutEdge(In60[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID278 e278 ( .InEdge(Out135), .OutEdge(In60[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID279 e279 ( .InEdge(Out207), .OutEdge(In60[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID280 e280 ( .InEdge(Out87), .OutEdge(In60[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID281 e281 ( .InEdge(Out208), .OutEdge(In60[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID282 e282 ( .InEdge(Out103), .OutEdge(In60[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID61_INDEGREE5 n61 ( .InEdges(In61), .OutEdge(Out61),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID283 e283 ( .InEdge(Out65), .OutEdge(In61[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID284 e284 ( .InEdge(Out248), .OutEdge(In61[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID285 e285 ( .InEdge(Out199), .OutEdge(In61[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID286 e286 ( .InEdge(Out11), .OutEdge(In61[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID287 e287 ( .InEdge(Out136), .OutEdge(In61[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID62_INDEGREE4 n62 ( .InEdges(In62), .OutEdge(Out62),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID288 e288 ( .InEdge(Out103), .OutEdge(In62[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID289 e289 ( .InEdge(Out148), .OutEdge(In62[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID290 e290 ( .InEdge(Out222), .OutEdge(In62[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID291 e291 ( .InEdge(Out183), .OutEdge(In62[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID63_INDEGREE6 n63 ( .InEdges(In63), .OutEdge(Out63),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID292 e292 ( .InEdge(Out237), .OutEdge(In63[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID293 e293 ( .InEdge(Out144), .OutEdge(In63[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID294 e294 ( .InEdge(Out218), .OutEdge(In63[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID295 e295 ( .InEdge(Out22), .OutEdge(In63[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID296 e296 ( .InEdge(Out189), .OutEdge(In63[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID297 e297 ( .InEdge(Out235), .OutEdge(In63[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID64_INDEGREE7 n64 ( .InEdges(In64), .OutEdge(Out64),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID298 e298 ( .InEdge(Out79), .OutEdge(In64[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID299 e299 ( .InEdge(Out234), .OutEdge(In64[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID300 e300 ( .InEdge(Out140), .OutEdge(In64[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID301 e301 ( .InEdge(Out87), .OutEdge(In64[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID302 e302 ( .InEdge(Out139), .OutEdge(In64[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID303 e303 ( .InEdge(Out41), .OutEdge(In64[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID304 e304 ( .InEdge(Out137), .OutEdge(In64[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID65_INDEGREE5 n65 ( .InEdges(In65), .OutEdge(Out65),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID305 e305 ( .InEdge(Out118), .OutEdge(In65[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID306 e306 ( .InEdge(Out75), .OutEdge(In65[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID307 e307 ( .InEdge(Out141), .OutEdge(In65[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID308 e308 ( .InEdge(Out186), .OutEdge(In65[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID309 e309 ( .InEdge(Out41), .OutEdge(In65[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID66_INDEGREE4 n66 ( .InEdges(In66), .OutEdge(Out66),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID310 e310 ( .InEdge(Out150), .OutEdge(In66[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID311 e311 ( .InEdge(Out4), .OutEdge(In66[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID312 e312 ( .InEdge(Out67), .OutEdge(In66[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID313 e313 ( .InEdge(Out64), .OutEdge(In66[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID67_INDEGREE1 n67 ( .InEdges(In67), .OutEdge(Out67),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID314 e314 ( .InEdge(Out98), .OutEdge(In67[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID68_INDEGREE8 n68 ( .InEdges(In68), .OutEdge(Out68),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID315 e315 ( .InEdge(Out247), .OutEdge(In68[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID316 e316 ( .InEdge(Out189), .OutEdge(In68[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID317 e317 ( .InEdge(Out90), .OutEdge(In68[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID318 e318 ( .InEdge(Out119), .OutEdge(In68[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID319 e319 ( .InEdge(Out192), .OutEdge(In68[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID320 e320 ( .InEdge(Out97), .OutEdge(In68[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID321 e321 ( .InEdge(Out206), .OutEdge(In68[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID322 e322 ( .InEdge(Out146), .OutEdge(In68[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID69_INDEGREE8 n69 ( .InEdges(In69), .OutEdge(Out69),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID323 e323 ( .InEdge(Out56), .OutEdge(In69[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID324 e324 ( .InEdge(Out170), .OutEdge(In69[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID325 e325 ( .InEdge(Out96), .OutEdge(In69[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID326 e326 ( .InEdge(Out9), .OutEdge(In69[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID327 e327 ( .InEdge(Out76), .OutEdge(In69[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID328 e328 ( .InEdge(Out95), .OutEdge(In69[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID329 e329 ( .InEdge(Out203), .OutEdge(In69[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID330 e330 ( .InEdge(Out136), .OutEdge(In69[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID70_INDEGREE2 n70 ( .InEdges(In70), .OutEdge(Out70),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID331 e331 ( .InEdge(Out88), .OutEdge(In70[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID332 e332 ( .InEdge(Out226), .OutEdge(In70[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID71_INDEGREE3 n71 ( .InEdges(In71), .OutEdge(Out71),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID333 e333 ( .InEdge(Out148), .OutEdge(In71[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID334 e334 ( .InEdge(Out4), .OutEdge(In71[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID335 e335 ( .InEdge(Out230), .OutEdge(In71[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID72_INDEGREE6 n72 ( .InEdges(In72), .OutEdge(Out72),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID336 e336 ( .InEdge(Out164), .OutEdge(In72[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID337 e337 ( .InEdge(Out10), .OutEdge(In72[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID338 e338 ( .InEdge(Out69), .OutEdge(In72[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID339 e339 ( .InEdge(Out206), .OutEdge(In72[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID340 e340 ( .InEdge(Out184), .OutEdge(In72[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID341 e341 ( .InEdge(Out183), .OutEdge(In72[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID73_INDEGREE7 n73 ( .InEdges(In73), .OutEdge(Out73),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID342 e342 ( .InEdge(Out39), .OutEdge(In73[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID343 e343 ( .InEdge(Out107), .OutEdge(In73[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID344 e344 ( .InEdge(Out92), .OutEdge(In73[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID345 e345 ( .InEdge(Out129), .OutEdge(In73[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID346 e346 ( .InEdge(Out75), .OutEdge(In73[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID347 e347 ( .InEdge(Out238), .OutEdge(In73[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID348 e348 ( .InEdge(Out247), .OutEdge(In73[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID74_INDEGREE5 n74 ( .InEdges(In74), .OutEdge(Out74),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID349 e349 ( .InEdge(Out115), .OutEdge(In74[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID350 e350 ( .InEdge(Out239), .OutEdge(In74[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID351 e351 ( .InEdge(Out86), .OutEdge(In74[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID352 e352 ( .InEdge(Out102), .OutEdge(In74[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID353 e353 ( .InEdge(Out88), .OutEdge(In74[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID75_INDEGREE6 n75 ( .InEdges(In75), .OutEdge(Out75),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID354 e354 ( .InEdge(Out253), .OutEdge(In75[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID355 e355 ( .InEdge(Out248), .OutEdge(In75[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID356 e356 ( .InEdge(Out185), .OutEdge(In75[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID357 e357 ( .InEdge(Out21), .OutEdge(In75[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID358 e358 ( .InEdge(Out214), .OutEdge(In75[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID359 e359 ( .InEdge(Out145), .OutEdge(In75[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID76_INDEGREE4 n76 ( .InEdges(In76), .OutEdge(Out76),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID360 e360 ( .InEdge(Out185), .OutEdge(In76[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID361 e361 ( .InEdge(Out167), .OutEdge(In76[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID362 e362 ( .InEdge(Out102), .OutEdge(In76[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID363 e363 ( .InEdge(Out236), .OutEdge(In76[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID77_INDEGREE3 n77 ( .InEdges(In77), .OutEdge(Out77),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID364 e364 ( .InEdge(Out110), .OutEdge(In77[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID365 e365 ( .InEdge(Out206), .OutEdge(In77[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID366 e366 ( .InEdge(Out103), .OutEdge(In77[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID78_INDEGREE5 n78 ( .InEdges(In78), .OutEdge(Out78),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID367 e367 ( .InEdge(Out28), .OutEdge(In78[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID368 e368 ( .InEdge(Out85), .OutEdge(In78[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID369 e369 ( .InEdge(Out90), .OutEdge(In78[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID370 e370 ( .InEdge(Out12), .OutEdge(In78[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID371 e371 ( .InEdge(Out132), .OutEdge(In78[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID79_INDEGREE4 n79 ( .InEdges(In79), .OutEdge(Out79),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID372 e372 ( .InEdge(Out207), .OutEdge(In79[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID373 e373 ( .InEdge(Out3), .OutEdge(In79[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID374 e374 ( .InEdge(Out43), .OutEdge(In79[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID375 e375 ( .InEdge(Out74), .OutEdge(In79[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID80_INDEGREE2 n80 ( .InEdges(In80), .OutEdge(Out80),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID376 e376 ( .InEdge(Out196), .OutEdge(In80[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID377 e377 ( .InEdge(Out119), .OutEdge(In80[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID81_INDEGREE5 n81 ( .InEdges(In81), .OutEdge(Out81),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID378 e378 ( .InEdge(Out12), .OutEdge(In81[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID379 e379 ( .InEdge(Out190), .OutEdge(In81[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID380 e380 ( .InEdge(Out238), .OutEdge(In81[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID381 e381 ( .InEdge(Out144), .OutEdge(In81[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID382 e382 ( .InEdge(Out230), .OutEdge(In81[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID82_INDEGREE2 n82 ( .InEdges(In82), .OutEdge(Out82),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID383 e383 ( .InEdge(Out124), .OutEdge(In82[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID384 e384 ( .InEdge(Out84), .OutEdge(In82[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID83_INDEGREE4 n83 ( .InEdges(In83), .OutEdge(Out83),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID385 e385 ( .InEdge(Out160), .OutEdge(In83[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID386 e386 ( .InEdge(Out21), .OutEdge(In83[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID387 e387 ( .InEdge(Out221), .OutEdge(In83[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID388 e388 ( .InEdge(Out39), .OutEdge(In83[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID84_INDEGREE5 n84 ( .InEdges(In84), .OutEdge(Out84),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID389 e389 ( .InEdge(Out177), .OutEdge(In84[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID390 e390 ( .InEdge(Out93), .OutEdge(In84[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID391 e391 ( .InEdge(Out173), .OutEdge(In84[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID392 e392 ( .InEdge(Out234), .OutEdge(In84[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID393 e393 ( .InEdge(Out241), .OutEdge(In84[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID85_INDEGREE3 n85 ( .InEdges(In85), .OutEdge(Out85),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID394 e394 ( .InEdge(Out134), .OutEdge(In85[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID395 e395 ( .InEdge(Out91), .OutEdge(In85[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID396 e396 ( .InEdge(Out143), .OutEdge(In85[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID86_INDEGREE4 n86 ( .InEdges(In86), .OutEdge(Out86),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID397 e397 ( .InEdge(Out101), .OutEdge(In86[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID398 e398 ( .InEdge(Out207), .OutEdge(In86[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID399 e399 ( .InEdge(Out19), .OutEdge(In86[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID400 e400 ( .InEdge(Out79), .OutEdge(In86[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID87_INDEGREE8 n87 ( .InEdges(In87), .OutEdge(Out87),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID401 e401 ( .InEdge(Out251), .OutEdge(In87[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID402 e402 ( .InEdge(Out24), .OutEdge(In87[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID403 e403 ( .InEdge(Out147), .OutEdge(In87[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID404 e404 ( .InEdge(Out91), .OutEdge(In87[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID405 e405 ( .InEdge(Out243), .OutEdge(In87[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID406 e406 ( .InEdge(Out76), .OutEdge(In87[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID407 e407 ( .InEdge(Out77), .OutEdge(In87[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID408 e408 ( .InEdge(Out116), .OutEdge(In87[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID88_INDEGREE2 n88 ( .InEdges(In88), .OutEdge(Out88),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID409 e409 ( .InEdge(Out65), .OutEdge(In88[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID410 e410 ( .InEdge(Out111), .OutEdge(In88[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID89_INDEGREE2 n89 ( .InEdges(In89), .OutEdge(Out89),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID411 e411 ( .InEdge(Out48), .OutEdge(In89[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID412 e412 ( .InEdge(Out152), .OutEdge(In89[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID90_INDEGREE3 n90 ( .InEdges(In90), .OutEdge(Out90),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID413 e413 ( .InEdge(Out48), .OutEdge(In90[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID414 e414 ( .InEdge(Out186), .OutEdge(In90[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID415 e415 ( .InEdge(Out200), .OutEdge(In90[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID91_INDEGREE4 n91 ( .InEdges(In91), .OutEdge(Out91),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID416 e416 ( .InEdge(Out244), .OutEdge(In91[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID417 e417 ( .InEdge(Out30), .OutEdge(In91[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID418 e418 ( .InEdge(Out92), .OutEdge(In91[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID419 e419 ( .InEdge(Out192), .OutEdge(In91[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID92_INDEGREE8 n92 ( .InEdges(In92), .OutEdge(Out92),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID420 e420 ( .InEdge(Out69), .OutEdge(In92[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID421 e421 ( .InEdge(Out147), .OutEdge(In92[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID422 e422 ( .InEdge(Out199), .OutEdge(In92[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID423 e423 ( .InEdge(Out240), .OutEdge(In92[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID424 e424 ( .InEdge(Out101), .OutEdge(In92[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID425 e425 ( .InEdge(Out246), .OutEdge(In92[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID426 e426 ( .InEdge(Out56), .OutEdge(In92[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID427 e427 ( .InEdge(Out55), .OutEdge(In92[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID93_INDEGREE8 n93 ( .InEdges(In93), .OutEdge(Out93),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID428 e428 ( .InEdge(Out205), .OutEdge(In93[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID429 e429 ( .InEdge(Out180), .OutEdge(In93[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID430 e430 ( .InEdge(Out10), .OutEdge(In93[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID431 e431 ( .InEdge(Out61), .OutEdge(In93[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID432 e432 ( .InEdge(Out250), .OutEdge(In93[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID433 e433 ( .InEdge(Out66), .OutEdge(In93[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID434 e434 ( .InEdge(Out68), .OutEdge(In93[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID435 e435 ( .InEdge(Out155), .OutEdge(In93[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID94_INDEGREE3 n94 ( .InEdges(In94), .OutEdge(Out94),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID436 e436 ( .InEdge(Out173), .OutEdge(In94[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID437 e437 ( .InEdge(Out183), .OutEdge(In94[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID438 e438 ( .InEdge(Out110), .OutEdge(In94[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID95_INDEGREE8 n95 ( .InEdges(In95), .OutEdge(Out95),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID439 e439 ( .InEdge(Out151), .OutEdge(In95[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID440 e440 ( .InEdge(Out31), .OutEdge(In95[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID441 e441 ( .InEdge(Out246), .OutEdge(In95[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID442 e442 ( .InEdge(Out25), .OutEdge(In95[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID443 e443 ( .InEdge(Out190), .OutEdge(In95[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID444 e444 ( .InEdge(Out52), .OutEdge(In95[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID445 e445 ( .InEdge(Out23), .OutEdge(In95[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID446 e446 ( .InEdge(Out178), .OutEdge(In95[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID96_INDEGREE1 n96 ( .InEdges(In96), .OutEdge(Out96),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID447 e447 ( .InEdge(Out207), .OutEdge(In96[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID97_INDEGREE7 n97 ( .InEdges(In97), .OutEdge(Out97),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID448 e448 ( .InEdge(Out131), .OutEdge(In97[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID449 e449 ( .InEdge(Out151), .OutEdge(In97[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID450 e450 ( .InEdge(Out2), .OutEdge(In97[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID451 e451 ( .InEdge(Out136), .OutEdge(In97[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID452 e452 ( .InEdge(Out255), .OutEdge(In97[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID453 e453 ( .InEdge(Out110), .OutEdge(In97[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID454 e454 ( .InEdge(Out157), .OutEdge(In97[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID98_INDEGREE1 n98 ( .InEdges(In98), .OutEdge(Out98),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID455 e455 ( .InEdge(Out111), .OutEdge(In98[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID99_INDEGREE2 n99 ( .InEdges(In99), .OutEdge(Out99),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID456 e456 ( .InEdge(Out36), .OutEdge(In99[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID457 e457 ( .InEdge(Out14), .OutEdge(In99[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID100_INDEGREE3 n100 ( .InEdges(In100), .OutEdge(Out100),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID458 e458 ( .InEdge(Out31), .OutEdge(In100[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID459 e459 ( .InEdge(Out200), .OutEdge(In100[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID460 e460 ( .InEdge(Out52), .OutEdge(In100[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID101_INDEGREE2 n101 ( .InEdges(In101), .OutEdge(Out101),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID461 e461 ( .InEdge(Out112), .OutEdge(In101[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID462 e462 ( .InEdge(Out167), .OutEdge(In101[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID102_INDEGREE8 n102 ( .InEdges(In102), .OutEdge(Out102),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID463 e463 ( .InEdge(Out33), .OutEdge(In102[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID464 e464 ( .InEdge(Out126), .OutEdge(In102[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID465 e465 ( .InEdge(Out163), .OutEdge(In102[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID466 e466 ( .InEdge(Out113), .OutEdge(In102[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID467 e467 ( .InEdge(Out8), .OutEdge(In102[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID468 e468 ( .InEdge(Out32), .OutEdge(In102[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID469 e469 ( .InEdge(Out28), .OutEdge(In102[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID470 e470 ( .InEdge(Out250), .OutEdge(In102[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID103_INDEGREE7 n103 ( .InEdges(In103), .OutEdge(Out103),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID471 e471 ( .InEdge(Out227), .OutEdge(In103[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID472 e472 ( .InEdge(Out86), .OutEdge(In103[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID473 e473 ( .InEdge(Out155), .OutEdge(In103[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID474 e474 ( .InEdge(Out120), .OutEdge(In103[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID475 e475 ( .InEdge(Out140), .OutEdge(In103[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID476 e476 ( .InEdge(Out149), .OutEdge(In103[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID477 e477 ( .InEdge(Out214), .OutEdge(In103[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID104_INDEGREE6 n104 ( .InEdges(In104), .OutEdge(Out104),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID478 e478 ( .InEdge(Out212), .OutEdge(In104[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID479 e479 ( .InEdge(Out24), .OutEdge(In104[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID480 e480 ( .InEdge(Out242), .OutEdge(In104[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID481 e481 ( .InEdge(Out109), .OutEdge(In104[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID482 e482 ( .InEdge(Out139), .OutEdge(In104[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID483 e483 ( .InEdge(Out34), .OutEdge(In104[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID105_INDEGREE2 n105 ( .InEdges(In105), .OutEdge(Out105),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID484 e484 ( .InEdge(Out77), .OutEdge(In105[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID485 e485 ( .InEdge(Out244), .OutEdge(In105[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID106_INDEGREE6 n106 ( .InEdges(In106), .OutEdge(Out106),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID486 e486 ( .InEdge(Out15), .OutEdge(In106[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID487 e487 ( .InEdge(Out126), .OutEdge(In106[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID488 e488 ( .InEdge(Out98), .OutEdge(In106[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID489 e489 ( .InEdge(Out189), .OutEdge(In106[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID490 e490 ( .InEdge(Out234), .OutEdge(In106[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID491 e491 ( .InEdge(Out253), .OutEdge(In106[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID107_INDEGREE3 n107 ( .InEdges(In107), .OutEdge(Out107),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID492 e492 ( .InEdge(Out132), .OutEdge(In107[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID493 e493 ( .InEdge(Out84), .OutEdge(In107[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID494 e494 ( .InEdge(Out29), .OutEdge(In107[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID108_INDEGREE4 n108 ( .InEdges(In108), .OutEdge(Out108),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID495 e495 ( .InEdge(Out232), .OutEdge(In108[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID496 e496 ( .InEdge(Out48), .OutEdge(In108[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID497 e497 ( .InEdge(Out233), .OutEdge(In108[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID498 e498 ( .InEdge(Out59), .OutEdge(In108[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID109_INDEGREE1 n109 ( .InEdges(In109), .OutEdge(Out109),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID499 e499 ( .InEdge(Out122), .OutEdge(In109[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID110_INDEGREE4 n110 ( .InEdges(In110), .OutEdge(Out110),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID500 e500 ( .InEdge(Out218), .OutEdge(In110[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID501 e501 ( .InEdge(Out231), .OutEdge(In110[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID502 e502 ( .InEdge(Out184), .OutEdge(In110[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID503 e503 ( .InEdge(Out243), .OutEdge(In110[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID111_INDEGREE2 n111 ( .InEdges(In111), .OutEdge(Out111),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID504 e504 ( .InEdge(Out17), .OutEdge(In111[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID505 e505 ( .InEdge(Out101), .OutEdge(In111[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID112_INDEGREE2 n112 ( .InEdges(In112), .OutEdge(Out112),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID506 e506 ( .InEdge(Out75), .OutEdge(In112[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID507 e507 ( .InEdge(Out71), .OutEdge(In112[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID113_INDEGREE3 n113 ( .InEdges(In113), .OutEdge(Out113),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID508 e508 ( .InEdge(Out54), .OutEdge(In113[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID509 e509 ( .InEdge(Out233), .OutEdge(In113[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID510 e510 ( .InEdge(Out48), .OutEdge(In113[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID114_INDEGREE5 n114 ( .InEdges(In114), .OutEdge(Out114),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID511 e511 ( .InEdge(Out167), .OutEdge(In114[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID512 e512 ( .InEdge(Out220), .OutEdge(In114[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID513 e513 ( .InEdge(Out129), .OutEdge(In114[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID514 e514 ( .InEdge(Out84), .OutEdge(In114[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID515 e515 ( .InEdge(Out34), .OutEdge(In114[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID115_INDEGREE3 n115 ( .InEdges(In115), .OutEdge(Out115),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID516 e516 ( .InEdge(Out151), .OutEdge(In115[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID517 e517 ( .InEdge(Out113), .OutEdge(In115[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID518 e518 ( .InEdge(Out203), .OutEdge(In115[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID116_INDEGREE5 n116 ( .InEdges(In116), .OutEdge(Out116),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID519 e519 ( .InEdge(Out160), .OutEdge(In116[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID520 e520 ( .InEdge(Out204), .OutEdge(In116[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID521 e521 ( .InEdge(Out233), .OutEdge(In116[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID522 e522 ( .InEdge(Out22), .OutEdge(In116[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID523 e523 ( .InEdge(Out128), .OutEdge(In116[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID117_INDEGREE4 n117 ( .InEdges(In117), .OutEdge(Out117),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID524 e524 ( .InEdge(Out153), .OutEdge(In117[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID525 e525 ( .InEdge(Out22), .OutEdge(In117[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID526 e526 ( .InEdge(Out137), .OutEdge(In117[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID527 e527 ( .InEdge(Out144), .OutEdge(In117[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID118_INDEGREE4 n118 ( .InEdges(In118), .OutEdge(Out118),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID528 e528 ( .InEdge(Out182), .OutEdge(In118[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID529 e529 ( .InEdge(Out222), .OutEdge(In118[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID530 e530 ( .InEdge(Out232), .OutEdge(In118[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID531 e531 ( .InEdge(Out91), .OutEdge(In118[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID119_INDEGREE8 n119 ( .InEdges(In119), .OutEdge(Out119),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID532 e532 ( .InEdge(Out103), .OutEdge(In119[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID533 e533 ( .InEdge(Out217), .OutEdge(In119[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID534 e534 ( .InEdge(Out36), .OutEdge(In119[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID535 e535 ( .InEdge(Out111), .OutEdge(In119[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID536 e536 ( .InEdge(Out215), .OutEdge(In119[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID537 e537 ( .InEdge(Out228), .OutEdge(In119[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID538 e538 ( .InEdge(Out253), .OutEdge(In119[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID539 e539 ( .InEdge(Out86), .OutEdge(In119[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID120_INDEGREE8 n120 ( .InEdges(In120), .OutEdge(Out120),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID540 e540 ( .InEdge(Out121), .OutEdge(In120[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID541 e541 ( .InEdge(Out209), .OutEdge(In120[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID542 e542 ( .InEdge(Out51), .OutEdge(In120[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID543 e543 ( .InEdge(Out175), .OutEdge(In120[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID544 e544 ( .InEdge(Out102), .OutEdge(In120[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID545 e545 ( .InEdge(Out44), .OutEdge(In120[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID546 e546 ( .InEdge(Out228), .OutEdge(In120[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID547 e547 ( .InEdge(Out57), .OutEdge(In120[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID121_INDEGREE2 n121 ( .InEdges(In121), .OutEdge(Out121),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID548 e548 ( .InEdge(Out57), .OutEdge(In121[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID549 e549 ( .InEdge(Out233), .OutEdge(In121[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID122_INDEGREE6 n122 ( .InEdges(In122), .OutEdge(Out122),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID550 e550 ( .InEdge(Out167), .OutEdge(In122[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID551 e551 ( .InEdge(Out217), .OutEdge(In122[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID552 e552 ( .InEdge(Out48), .OutEdge(In122[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID553 e553 ( .InEdge(Out183), .OutEdge(In122[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID554 e554 ( .InEdge(Out200), .OutEdge(In122[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID555 e555 ( .InEdge(Out99), .OutEdge(In122[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID123_INDEGREE5 n123 ( .InEdges(In123), .OutEdge(Out123),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID556 e556 ( .InEdge(Out171), .OutEdge(In123[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID557 e557 ( .InEdge(Out141), .OutEdge(In123[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID558 e558 ( .InEdge(Out101), .OutEdge(In123[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID559 e559 ( .InEdge(Out10), .OutEdge(In123[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID560 e560 ( .InEdge(Out58), .OutEdge(In123[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID124_INDEGREE4 n124 ( .InEdges(In124), .OutEdge(Out124),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID561 e561 ( .InEdge(Out30), .OutEdge(In124[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID562 e562 ( .InEdge(Out145), .OutEdge(In124[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID563 e563 ( .InEdge(Out168), .OutEdge(In124[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID564 e564 ( .InEdge(Out97), .OutEdge(In124[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID125_INDEGREE5 n125 ( .InEdges(In125), .OutEdge(Out125),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID565 e565 ( .InEdge(Out216), .OutEdge(In125[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID566 e566 ( .InEdge(Out140), .OutEdge(In125[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID567 e567 ( .InEdge(Out95), .OutEdge(In125[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID568 e568 ( .InEdge(Out62), .OutEdge(In125[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID569 e569 ( .InEdge(Out238), .OutEdge(In125[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID126_INDEGREE4 n126 ( .InEdges(In126), .OutEdge(Out126),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID570 e570 ( .InEdge(Out144), .OutEdge(In126[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID571 e571 ( .InEdge(Out139), .OutEdge(In126[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID572 e572 ( .InEdge(Out222), .OutEdge(In126[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID573 e573 ( .InEdge(Out65), .OutEdge(In126[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID127_INDEGREE5 n127 ( .InEdges(In127), .OutEdge(Out127),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID574 e574 ( .InEdge(Out147), .OutEdge(In127[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID575 e575 ( .InEdge(Out36), .OutEdge(In127[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID576 e576 ( .InEdge(Out69), .OutEdge(In127[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID577 e577 ( .InEdge(Out137), .OutEdge(In127[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID578 e578 ( .InEdge(Out179), .OutEdge(In127[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID128_INDEGREE3 n128 ( .InEdges(In128), .OutEdge(Out128),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID579 e579 ( .InEdge(Out45), .OutEdge(In128[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID580 e580 ( .InEdge(Out55), .OutEdge(In128[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID581 e581 ( .InEdge(Out24), .OutEdge(In128[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID129_INDEGREE1 n129 ( .InEdges(In129), .OutEdge(Out129),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID582 e582 ( .InEdge(Out114), .OutEdge(In129[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID130_INDEGREE6 n130 ( .InEdges(In130), .OutEdge(Out130),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID583 e583 ( .InEdge(Out194), .OutEdge(In130[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID584 e584 ( .InEdge(Out188), .OutEdge(In130[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID585 e585 ( .InEdge(Out139), .OutEdge(In130[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID586 e586 ( .InEdge(Out32), .OutEdge(In130[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID587 e587 ( .InEdge(Out236), .OutEdge(In130[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID588 e588 ( .InEdge(Out239), .OutEdge(In130[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID131_INDEGREE3 n131 ( .InEdges(In131), .OutEdge(Out131),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID589 e589 ( .InEdge(Out243), .OutEdge(In131[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID590 e590 ( .InEdge(Out85), .OutEdge(In131[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID591 e591 ( .InEdge(Out26), .OutEdge(In131[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID132_INDEGREE8 n132 ( .InEdges(In132), .OutEdge(Out132),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID592 e592 ( .InEdge(Out188), .OutEdge(In132[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID593 e593 ( .InEdge(Out190), .OutEdge(In132[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID594 e594 ( .InEdge(Out80), .OutEdge(In132[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID595 e595 ( .InEdge(Out252), .OutEdge(In132[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID596 e596 ( .InEdge(Out232), .OutEdge(In132[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID597 e597 ( .InEdge(Out75), .OutEdge(In132[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID598 e598 ( .InEdge(Out150), .OutEdge(In132[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID599 e599 ( .InEdge(Out147), .OutEdge(In132[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID133_INDEGREE8 n133 ( .InEdges(In133), .OutEdge(Out133),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID600 e600 ( .InEdge(Out3), .OutEdge(In133[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID601 e601 ( .InEdge(Out8), .OutEdge(In133[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID602 e602 ( .InEdge(Out206), .OutEdge(In133[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID603 e603 ( .InEdge(Out17), .OutEdge(In133[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID604 e604 ( .InEdge(Out196), .OutEdge(In133[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID605 e605 ( .InEdge(Out101), .OutEdge(In133[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID606 e606 ( .InEdge(Out65), .OutEdge(In133[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID607 e607 ( .InEdge(Out66), .OutEdge(In133[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID134_INDEGREE7 n134 ( .InEdges(In134), .OutEdge(Out134),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID608 e608 ( .InEdge(Out143), .OutEdge(In134[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID609 e609 ( .InEdge(Out206), .OutEdge(In134[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID610 e610 ( .InEdge(Out23), .OutEdge(In134[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID611 e611 ( .InEdge(Out198), .OutEdge(In134[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID612 e612 ( .InEdge(Out20), .OutEdge(In134[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID613 e613 ( .InEdge(Out211), .OutEdge(In134[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID614 e614 ( .InEdge(Out248), .OutEdge(In134[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID135_INDEGREE6 n135 ( .InEdges(In135), .OutEdge(Out135),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID615 e615 ( .InEdge(Out177), .OutEdge(In135[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID616 e616 ( .InEdge(Out15), .OutEdge(In135[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID617 e617 ( .InEdge(Out115), .OutEdge(In135[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID618 e618 ( .InEdge(Out53), .OutEdge(In135[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID619 e619 ( .InEdge(Out130), .OutEdge(In135[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID620 e620 ( .InEdge(Out58), .OutEdge(In135[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID136_INDEGREE7 n136 ( .InEdges(In136), .OutEdge(Out136),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID621 e621 ( .InEdge(Out80), .OutEdge(In136[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID622 e622 ( .InEdge(Out86), .OutEdge(In136[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID623 e623 ( .InEdge(Out23), .OutEdge(In136[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID624 e624 ( .InEdge(Out154), .OutEdge(In136[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID625 e625 ( .InEdge(Out3), .OutEdge(In136[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID626 e626 ( .InEdge(Out179), .OutEdge(In136[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID627 e627 ( .InEdge(Out166), .OutEdge(In136[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID137_INDEGREE1 n137 ( .InEdges(In137), .OutEdge(Out137),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID628 e628 ( .InEdge(Out128), .OutEdge(In137[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID138_INDEGREE4 n138 ( .InEdges(In138), .OutEdge(Out138),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID629 e629 ( .InEdge(Out93), .OutEdge(In138[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID630 e630 ( .InEdge(Out40), .OutEdge(In138[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID631 e631 ( .InEdge(Out96), .OutEdge(In138[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID632 e632 ( .InEdge(Out59), .OutEdge(In138[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID139_INDEGREE6 n139 ( .InEdges(In139), .OutEdge(Out139),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID633 e633 ( .InEdge(Out204), .OutEdge(In139[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID634 e634 ( .InEdge(Out189), .OutEdge(In139[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID635 e635 ( .InEdge(Out134), .OutEdge(In139[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID636 e636 ( .InEdge(Out88), .OutEdge(In139[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID637 e637 ( .InEdge(Out37), .OutEdge(In139[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID638 e638 ( .InEdge(Out91), .OutEdge(In139[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID140_INDEGREE4 n140 ( .InEdges(In140), .OutEdge(Out140),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID639 e639 ( .InEdge(Out183), .OutEdge(In140[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID640 e640 ( .InEdge(Out37), .OutEdge(In140[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID641 e641 ( .InEdge(Out173), .OutEdge(In140[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID642 e642 ( .InEdge(Out85), .OutEdge(In140[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID141_INDEGREE8 n141 ( .InEdges(In141), .OutEdge(Out141),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID643 e643 ( .InEdge(Out249), .OutEdge(In141[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID644 e644 ( .InEdge(Out78), .OutEdge(In141[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID645 e645 ( .InEdge(Out175), .OutEdge(In141[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID646 e646 ( .InEdge(Out64), .OutEdge(In141[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID647 e647 ( .InEdge(Out176), .OutEdge(In141[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID648 e648 ( .InEdge(Out51), .OutEdge(In141[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID649 e649 ( .InEdge(Out60), .OutEdge(In141[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID650 e650 ( .InEdge(Out109), .OutEdge(In141[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID142_INDEGREE4 n142 ( .InEdges(In142), .OutEdge(Out142),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID651 e651 ( .InEdge(Out118), .OutEdge(In142[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID652 e652 ( .InEdge(Out143), .OutEdge(In142[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID653 e653 ( .InEdge(Out141), .OutEdge(In142[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID654 e654 ( .InEdge(Out23), .OutEdge(In142[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID143_INDEGREE8 n143 ( .InEdges(In143), .OutEdge(Out143),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID655 e655 ( .InEdge(Out223), .OutEdge(In143[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID656 e656 ( .InEdge(Out128), .OutEdge(In143[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID657 e657 ( .InEdge(Out96), .OutEdge(In143[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID658 e658 ( .InEdge(Out74), .OutEdge(In143[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID659 e659 ( .InEdge(Out212), .OutEdge(In143[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID660 e660 ( .InEdge(Out139), .OutEdge(In143[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID661 e661 ( .InEdge(Out124), .OutEdge(In143[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID662 e662 ( .InEdge(Out40), .OutEdge(In143[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID144_INDEGREE7 n144 ( .InEdges(In144), .OutEdge(Out144),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID663 e663 ( .InEdge(Out195), .OutEdge(In144[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID664 e664 ( .InEdge(Out89), .OutEdge(In144[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID665 e665 ( .InEdge(Out42), .OutEdge(In144[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID666 e666 ( .InEdge(Out167), .OutEdge(In144[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID667 e667 ( .InEdge(Out217), .OutEdge(In144[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID668 e668 ( .InEdge(Out232), .OutEdge(In144[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID669 e669 ( .InEdge(Out186), .OutEdge(In144[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID145_INDEGREE8 n145 ( .InEdges(In145), .OutEdge(Out145),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID670 e670 ( .InEdge(Out58), .OutEdge(In145[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID671 e671 ( .InEdge(Out242), .OutEdge(In145[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID672 e672 ( .InEdge(Out165), .OutEdge(In145[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID673 e673 ( .InEdge(Out197), .OutEdge(In145[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID674 e674 ( .InEdge(Out12), .OutEdge(In145[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID675 e675 ( .InEdge(Out210), .OutEdge(In145[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID676 e676 ( .InEdge(Out51), .OutEdge(In145[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID677 e677 ( .InEdge(Out247), .OutEdge(In145[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID146_INDEGREE2 n146 ( .InEdges(In146), .OutEdge(Out146),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID678 e678 ( .InEdge(Out37), .OutEdge(In146[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID679 e679 ( .InEdge(Out64), .OutEdge(In146[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID147_INDEGREE2 n147 ( .InEdges(In147), .OutEdge(Out147),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID680 e680 ( .InEdge(Out80), .OutEdge(In147[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID681 e681 ( .InEdge(Out242), .OutEdge(In147[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID148_INDEGREE1 n148 ( .InEdges(In148), .OutEdge(Out148),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID682 e682 ( .InEdge(Out9), .OutEdge(In148[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID149_INDEGREE7 n149 ( .InEdges(In149), .OutEdge(Out149),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID683 e683 ( .InEdge(Out59), .OutEdge(In149[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID684 e684 ( .InEdge(Out24), .OutEdge(In149[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID685 e685 ( .InEdge(Out83), .OutEdge(In149[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID686 e686 ( .InEdge(Out201), .OutEdge(In149[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID687 e687 ( .InEdge(Out186), .OutEdge(In149[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID688 e688 ( .InEdge(Out80), .OutEdge(In149[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID689 e689 ( .InEdge(Out99), .OutEdge(In149[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID150_INDEGREE3 n150 ( .InEdges(In150), .OutEdge(Out150),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID690 e690 ( .InEdge(Out40), .OutEdge(In150[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID691 e691 ( .InEdge(Out251), .OutEdge(In150[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID692 e692 ( .InEdge(Out120), .OutEdge(In150[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID151_INDEGREE8 n151 ( .InEdges(In151), .OutEdge(Out151),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID693 e693 ( .InEdge(Out124), .OutEdge(In151[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID694 e694 ( .InEdge(Out30), .OutEdge(In151[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID695 e695 ( .InEdge(Out79), .OutEdge(In151[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID696 e696 ( .InEdge(Out250), .OutEdge(In151[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID697 e697 ( .InEdge(Out192), .OutEdge(In151[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID698 e698 ( .InEdge(Out144), .OutEdge(In151[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID699 e699 ( .InEdge(Out128), .OutEdge(In151[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID700 e700 ( .InEdge(Out41), .OutEdge(In151[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID152_INDEGREE8 n152 ( .InEdges(In152), .OutEdge(Out152),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID701 e701 ( .InEdge(Out239), .OutEdge(In152[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID702 e702 ( .InEdge(Out211), .OutEdge(In152[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID703 e703 ( .InEdge(Out161), .OutEdge(In152[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID704 e704 ( .InEdge(Out113), .OutEdge(In152[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID705 e705 ( .InEdge(Out204), .OutEdge(In152[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID706 e706 ( .InEdge(Out20), .OutEdge(In152[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID707 e707 ( .InEdge(Out94), .OutEdge(In152[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID708 e708 ( .InEdge(Out134), .OutEdge(In152[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID153_INDEGREE8 n153 ( .InEdges(In153), .OutEdge(Out153),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID709 e709 ( .InEdge(Out41), .OutEdge(In153[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID710 e710 ( .InEdge(Out174), .OutEdge(In153[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID711 e711 ( .InEdge(Out71), .OutEdge(In153[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID712 e712 ( .InEdge(Out133), .OutEdge(In153[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID713 e713 ( .InEdge(Out91), .OutEdge(In153[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID714 e714 ( .InEdge(Out32), .OutEdge(In153[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID715 e715 ( .InEdge(Out14), .OutEdge(In153[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID716 e716 ( .InEdge(Out254), .OutEdge(In153[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID154_INDEGREE4 n154 ( .InEdges(In154), .OutEdge(Out154),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID717 e717 ( .InEdge(Out185), .OutEdge(In154[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID718 e718 ( .InEdge(Out43), .OutEdge(In154[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID719 e719 ( .InEdge(Out18), .OutEdge(In154[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID720 e720 ( .InEdge(Out192), .OutEdge(In154[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID155_INDEGREE7 n155 ( .InEdges(In155), .OutEdge(Out155),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID721 e721 ( .InEdge(Out119), .OutEdge(In155[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID722 e722 ( .InEdge(Out10), .OutEdge(In155[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID723 e723 ( .InEdge(Out222), .OutEdge(In155[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID724 e724 ( .InEdge(Out72), .OutEdge(In155[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID725 e725 ( .InEdge(Out131), .OutEdge(In155[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID726 e726 ( .InEdge(Out46), .OutEdge(In155[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID727 e727 ( .InEdge(Out232), .OutEdge(In155[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID156_INDEGREE7 n156 ( .InEdges(In156), .OutEdge(Out156),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID728 e728 ( .InEdge(Out134), .OutEdge(In156[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID729 e729 ( .InEdge(Out69), .OutEdge(In156[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID730 e730 ( .InEdge(Out143), .OutEdge(In156[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID731 e731 ( .InEdge(Out203), .OutEdge(In156[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID732 e732 ( .InEdge(Out17), .OutEdge(In156[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID733 e733 ( .InEdge(Out251), .OutEdge(In156[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID734 e734 ( .InEdge(Out107), .OutEdge(In156[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID157_INDEGREE8 n157 ( .InEdges(In157), .OutEdge(Out157),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID735 e735 ( .InEdge(Out38), .OutEdge(In157[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID736 e736 ( .InEdge(Out118), .OutEdge(In157[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID737 e737 ( .InEdge(Out147), .OutEdge(In157[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID738 e738 ( .InEdge(Out108), .OutEdge(In157[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID739 e739 ( .InEdge(Out129), .OutEdge(In157[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID740 e740 ( .InEdge(Out158), .OutEdge(In157[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID741 e741 ( .InEdge(Out119), .OutEdge(In157[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID742 e742 ( .InEdge(Out122), .OutEdge(In157[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID158_INDEGREE3 n158 ( .InEdges(In158), .OutEdge(Out158),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID743 e743 ( .InEdge(Out74), .OutEdge(In158[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID744 e744 ( .InEdge(Out144), .OutEdge(In158[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID745 e745 ( .InEdge(Out104), .OutEdge(In158[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID159_INDEGREE3 n159 ( .InEdges(In159), .OutEdge(Out159),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID746 e746 ( .InEdge(Out121), .OutEdge(In159[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID747 e747 ( .InEdge(Out203), .OutEdge(In159[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID748 e748 ( .InEdge(Out182), .OutEdge(In159[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID160_INDEGREE6 n160 ( .InEdges(In160), .OutEdge(Out160),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID749 e749 ( .InEdge(Out5), .OutEdge(In160[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID750 e750 ( .InEdge(Out132), .OutEdge(In160[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID751 e751 ( .InEdge(Out220), .OutEdge(In160[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID752 e752 ( .InEdge(Out131), .OutEdge(In160[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID753 e753 ( .InEdge(Out77), .OutEdge(In160[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID754 e754 ( .InEdge(Out206), .OutEdge(In160[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID161_INDEGREE4 n161 ( .InEdges(In161), .OutEdge(Out161),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID755 e755 ( .InEdge(Out81), .OutEdge(In161[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID756 e756 ( .InEdge(Out137), .OutEdge(In161[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID757 e757 ( .InEdge(Out63), .OutEdge(In161[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID758 e758 ( .InEdge(Out114), .OutEdge(In161[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID162_INDEGREE6 n162 ( .InEdges(In162), .OutEdge(Out162),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID759 e759 ( .InEdge(Out125), .OutEdge(In162[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID760 e760 ( .InEdge(Out70), .OutEdge(In162[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID761 e761 ( .InEdge(Out20), .OutEdge(In162[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID762 e762 ( .InEdge(Out171), .OutEdge(In162[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID763 e763 ( .InEdge(Out40), .OutEdge(In162[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID764 e764 ( .InEdge(Out252), .OutEdge(In162[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID163_INDEGREE8 n163 ( .InEdges(In163), .OutEdge(Out163),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID765 e765 ( .InEdge(Out51), .OutEdge(In163[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID766 e766 ( .InEdge(Out209), .OutEdge(In163[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID767 e767 ( .InEdge(Out95), .OutEdge(In163[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID768 e768 ( .InEdge(Out142), .OutEdge(In163[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID769 e769 ( .InEdge(Out148), .OutEdge(In163[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID770 e770 ( .InEdge(Out171), .OutEdge(In163[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID771 e771 ( .InEdge(Out111), .OutEdge(In163[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID772 e772 ( .InEdge(Out161), .OutEdge(In163[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID164_INDEGREE6 n164 ( .InEdges(In164), .OutEdge(Out164),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID773 e773 ( .InEdge(Out109), .OutEdge(In164[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID774 e774 ( .InEdge(Out105), .OutEdge(In164[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID775 e775 ( .InEdge(Out62), .OutEdge(In164[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID776 e776 ( .InEdge(Out223), .OutEdge(In164[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID777 e777 ( .InEdge(Out86), .OutEdge(In164[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID778 e778 ( .InEdge(Out144), .OutEdge(In164[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID165_INDEGREE3 n165 ( .InEdges(In165), .OutEdge(Out165),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID779 e779 ( .InEdge(Out230), .OutEdge(In165[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID780 e780 ( .InEdge(Out44), .OutEdge(In165[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID781 e781 ( .InEdge(Out10), .OutEdge(In165[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID166_INDEGREE4 n166 ( .InEdges(In166), .OutEdge(Out166),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID782 e782 ( .InEdge(Out247), .OutEdge(In166[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID783 e783 ( .InEdge(Out237), .OutEdge(In166[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID784 e784 ( .InEdge(Out229), .OutEdge(In166[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID785 e785 ( .InEdge(Out80), .OutEdge(In166[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID167_INDEGREE1 n167 ( .InEdges(In167), .OutEdge(Out167),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID786 e786 ( .InEdge(Out244), .OutEdge(In167[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID168_INDEGREE4 n168 ( .InEdges(In168), .OutEdge(Out168),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID787 e787 ( .InEdge(Out174), .OutEdge(In168[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID788 e788 ( .InEdge(Out153), .OutEdge(In168[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID789 e789 ( .InEdge(Out189), .OutEdge(In168[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID790 e790 ( .InEdge(Out62), .OutEdge(In168[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID169_INDEGREE4 n169 ( .InEdges(In169), .OutEdge(Out169),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID791 e791 ( .InEdge(Out206), .OutEdge(In169[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID792 e792 ( .InEdge(Out2), .OutEdge(In169[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID793 e793 ( .InEdge(Out55), .OutEdge(In169[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID794 e794 ( .InEdge(Out177), .OutEdge(In169[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID170_INDEGREE2 n170 ( .InEdges(In170), .OutEdge(Out170),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID795 e795 ( .InEdge(Out179), .OutEdge(In170[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID796 e796 ( .InEdge(Out142), .OutEdge(In170[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID171_INDEGREE4 n171 ( .InEdges(In171), .OutEdge(Out171),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID797 e797 ( .InEdge(Out254), .OutEdge(In171[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID798 e798 ( .InEdge(Out154), .OutEdge(In171[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID799 e799 ( .InEdge(Out101), .OutEdge(In171[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID800 e800 ( .InEdge(Out163), .OutEdge(In171[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID172_INDEGREE5 n172 ( .InEdges(In172), .OutEdge(Out172),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID801 e801 ( .InEdge(Out119), .OutEdge(In172[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID802 e802 ( .InEdge(Out115), .OutEdge(In172[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID803 e803 ( .InEdge(Out76), .OutEdge(In172[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID804 e804 ( .InEdge(Out21), .OutEdge(In172[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID805 e805 ( .InEdge(Out195), .OutEdge(In172[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID173_INDEGREE1 n173 ( .InEdges(In173), .OutEdge(Out173),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID806 e806 ( .InEdge(Out98), .OutEdge(In173[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID174_INDEGREE3 n174 ( .InEdges(In174), .OutEdge(Out174),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID807 e807 ( .InEdge(Out201), .OutEdge(In174[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID808 e808 ( .InEdge(Out150), .OutEdge(In174[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID809 e809 ( .InEdge(Out18), .OutEdge(In174[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID175_INDEGREE3 n175 ( .InEdges(In175), .OutEdge(Out175),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID810 e810 ( .InEdge(Out54), .OutEdge(In175[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID811 e811 ( .InEdge(Out197), .OutEdge(In175[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID812 e812 ( .InEdge(Out248), .OutEdge(In175[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID176_INDEGREE1 n176 ( .InEdges(In176), .OutEdge(Out176),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID813 e813 ( .InEdge(Out52), .OutEdge(In176[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID177_INDEGREE2 n177 ( .InEdges(In177), .OutEdge(Out177),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID814 e814 ( .InEdge(Out69), .OutEdge(In177[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID815 e815 ( .InEdge(Out116), .OutEdge(In177[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID178_INDEGREE2 n178 ( .InEdges(In178), .OutEdge(Out178),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID816 e816 ( .InEdge(Out237), .OutEdge(In178[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID817 e817 ( .InEdge(Out115), .OutEdge(In178[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID179_INDEGREE4 n179 ( .InEdges(In179), .OutEdge(Out179),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID818 e818 ( .InEdge(Out208), .OutEdge(In179[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID819 e819 ( .InEdge(Out58), .OutEdge(In179[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID820 e820 ( .InEdge(Out243), .OutEdge(In179[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID821 e821 ( .InEdge(Out201), .OutEdge(In179[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID180_INDEGREE8 n180 ( .InEdges(In180), .OutEdge(Out180),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID822 e822 ( .InEdge(Out177), .OutEdge(In180[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID823 e823 ( .InEdge(Out118), .OutEdge(In180[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID824 e824 ( .InEdge(Out242), .OutEdge(In180[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID825 e825 ( .InEdge(Out220), .OutEdge(In180[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID826 e826 ( .InEdge(Out37), .OutEdge(In180[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID827 e827 ( .InEdge(Out69), .OutEdge(In180[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID828 e828 ( .InEdge(Out114), .OutEdge(In180[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID829 e829 ( .InEdge(Out72), .OutEdge(In180[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID181_INDEGREE7 n181 ( .InEdges(In181), .OutEdge(Out181),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID830 e830 ( .InEdge(Out187), .OutEdge(In181[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID831 e831 ( .InEdge(Out10), .OutEdge(In181[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID832 e832 ( .InEdge(Out86), .OutEdge(In181[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID833 e833 ( .InEdge(Out173), .OutEdge(In181[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID834 e834 ( .InEdge(Out186), .OutEdge(In181[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID835 e835 ( .InEdge(Out114), .OutEdge(In181[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID836 e836 ( .InEdge(Out255), .OutEdge(In181[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID182_INDEGREE2 n182 ( .InEdges(In182), .OutEdge(Out182),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID837 e837 ( .InEdge(Out113), .OutEdge(In182[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID838 e838 ( .InEdge(Out5), .OutEdge(In182[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID183_INDEGREE1 n183 ( .InEdges(In183), .OutEdge(Out183),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID839 e839 ( .InEdge(Out71), .OutEdge(In183[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID184_INDEGREE6 n184 ( .InEdges(In184), .OutEdge(Out184),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID840 e840 ( .InEdge(Out134), .OutEdge(In184[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID841 e841 ( .InEdge(Out173), .OutEdge(In184[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID842 e842 ( .InEdge(Out27), .OutEdge(In184[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID843 e843 ( .InEdge(Out38), .OutEdge(In184[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID844 e844 ( .InEdge(Out74), .OutEdge(In184[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID845 e845 ( .InEdge(Out219), .OutEdge(In184[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID185_INDEGREE7 n185 ( .InEdges(In185), .OutEdge(Out185),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID846 e846 ( .InEdge(Out169), .OutEdge(In185[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID847 e847 ( .InEdge(Out130), .OutEdge(In185[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID848 e848 ( .InEdge(Out60), .OutEdge(In185[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID849 e849 ( .InEdge(Out238), .OutEdge(In185[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID850 e850 ( .InEdge(Out66), .OutEdge(In185[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID851 e851 ( .InEdge(Out183), .OutEdge(In185[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID852 e852 ( .InEdge(Out119), .OutEdge(In185[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID186_INDEGREE5 n186 ( .InEdges(In186), .OutEdge(Out186),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID853 e853 ( .InEdge(Out110), .OutEdge(In186[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID854 e854 ( .InEdge(Out254), .OutEdge(In186[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID855 e855 ( .InEdge(Out243), .OutEdge(In186[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID856 e856 ( .InEdge(Out212), .OutEdge(In186[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID857 e857 ( .InEdge(Out26), .OutEdge(In186[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID187_INDEGREE8 n187 ( .InEdges(In187), .OutEdge(Out187),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID858 e858 ( .InEdge(Out141), .OutEdge(In187[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID859 e859 ( .InEdge(Out160), .OutEdge(In187[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID860 e860 ( .InEdge(Out237), .OutEdge(In187[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID861 e861 ( .InEdge(Out122), .OutEdge(In187[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID862 e862 ( .InEdge(Out65), .OutEdge(In187[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID863 e863 ( .InEdge(Out194), .OutEdge(In187[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID864 e864 ( .InEdge(Out19), .OutEdge(In187[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID865 e865 ( .InEdge(Out235), .OutEdge(In187[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID188_INDEGREE2 n188 ( .InEdges(In188), .OutEdge(Out188),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID866 e866 ( .InEdge(Out96), .OutEdge(In188[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID867 e867 ( .InEdge(Out92), .OutEdge(In188[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID189_INDEGREE5 n189 ( .InEdges(In189), .OutEdge(Out189),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID868 e868 ( .InEdge(Out21), .OutEdge(In189[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID869 e869 ( .InEdge(Out138), .OutEdge(In189[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID870 e870 ( .InEdge(Out197), .OutEdge(In189[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID871 e871 ( .InEdge(Out95), .OutEdge(In189[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID872 e872 ( .InEdge(Out12), .OutEdge(In189[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID190_INDEGREE4 n190 ( .InEdges(In190), .OutEdge(Out190),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID873 e873 ( .InEdge(Out199), .OutEdge(In190[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID874 e874 ( .InEdge(Out65), .OutEdge(In190[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID875 e875 ( .InEdge(Out142), .OutEdge(In190[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID876 e876 ( .InEdge(Out111), .OutEdge(In190[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID191_INDEGREE4 n191 ( .InEdges(In191), .OutEdge(Out191),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID877 e877 ( .InEdge(Out239), .OutEdge(In191[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID878 e878 ( .InEdge(Out244), .OutEdge(In191[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID879 e879 ( .InEdge(Out221), .OutEdge(In191[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID880 e880 ( .InEdge(Out41), .OutEdge(In191[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID192_INDEGREE5 n192 ( .InEdges(In192), .OutEdge(Out192),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID881 e881 ( .InEdge(Out74), .OutEdge(In192[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID882 e882 ( .InEdge(Out113), .OutEdge(In192[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID883 e883 ( .InEdge(Out212), .OutEdge(In192[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID884 e884 ( .InEdge(Out5), .OutEdge(In192[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID885 e885 ( .InEdge(Out80), .OutEdge(In192[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID193_INDEGREE6 n193 ( .InEdges(In193), .OutEdge(Out193),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID886 e886 ( .InEdge(Out167), .OutEdge(In193[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID887 e887 ( .InEdge(Out124), .OutEdge(In193[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID888 e888 ( .InEdge(Out103), .OutEdge(In193[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID889 e889 ( .InEdge(Out153), .OutEdge(In193[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID890 e890 ( .InEdge(Out100), .OutEdge(In193[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID891 e891 ( .InEdge(Out158), .OutEdge(In193[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID194_INDEGREE4 n194 ( .InEdges(In194), .OutEdge(Out194),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID892 e892 ( .InEdge(Out187), .OutEdge(In194[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID893 e893 ( .InEdge(Out46), .OutEdge(In194[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID894 e894 ( .InEdge(Out32), .OutEdge(In194[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID895 e895 ( .InEdge(Out167), .OutEdge(In194[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID195_INDEGREE2 n195 ( .InEdges(In195), .OutEdge(Out195),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID896 e896 ( .InEdge(Out79), .OutEdge(In195[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID897 e897 ( .InEdge(Out176), .OutEdge(In195[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID196_INDEGREE2 n196 ( .InEdges(In196), .OutEdge(Out196),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID898 e898 ( .InEdge(Out102), .OutEdge(In196[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID899 e899 ( .InEdge(Out189), .OutEdge(In196[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID197_INDEGREE7 n197 ( .InEdges(In197), .OutEdge(Out197),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID900 e900 ( .InEdge(Out195), .OutEdge(In197[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID901 e901 ( .InEdge(Out8), .OutEdge(In197[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID902 e902 ( .InEdge(Out2), .OutEdge(In197[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID903 e903 ( .InEdge(Out111), .OutEdge(In197[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID904 e904 ( .InEdge(Out94), .OutEdge(In197[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID905 e905 ( .InEdge(Out57), .OutEdge(In197[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID906 e906 ( .InEdge(Out72), .OutEdge(In197[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID198_INDEGREE3 n198 ( .InEdges(In198), .OutEdge(Out198),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID907 e907 ( .InEdge(Out118), .OutEdge(In198[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID908 e908 ( .InEdge(Out71), .OutEdge(In198[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID909 e909 ( .InEdge(Out11), .OutEdge(In198[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID199_INDEGREE6 n199 ( .InEdges(In199), .OutEdge(Out199),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID910 e910 ( .InEdge(Out171), .OutEdge(In199[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID911 e911 ( .InEdge(Out17), .OutEdge(In199[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID912 e912 ( .InEdge(Out127), .OutEdge(In199[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID913 e913 ( .InEdge(Out115), .OutEdge(In199[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID914 e914 ( .InEdge(Out167), .OutEdge(In199[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID915 e915 ( .InEdge(Out26), .OutEdge(In199[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID200_INDEGREE2 n200 ( .InEdges(In200), .OutEdge(Out200),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID916 e916 ( .InEdge(Out51), .OutEdge(In200[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID917 e917 ( .InEdge(Out166), .OutEdge(In200[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID201_INDEGREE1 n201 ( .InEdges(In201), .OutEdge(Out201),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID918 e918 ( .InEdge(Out82), .OutEdge(In201[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID202_INDEGREE2 n202 ( .InEdges(In202), .OutEdge(Out202),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID919 e919 ( .InEdge(Out138), .OutEdge(In202[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID920 e920 ( .InEdge(Out136), .OutEdge(In202[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID203_INDEGREE6 n203 ( .InEdges(In203), .OutEdge(Out203),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID921 e921 ( .InEdge(Out173), .OutEdge(In203[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID922 e922 ( .InEdge(Out57), .OutEdge(In203[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID923 e923 ( .InEdge(Out60), .OutEdge(In203[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID924 e924 ( .InEdge(Out167), .OutEdge(In203[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID925 e925 ( .InEdge(Out208), .OutEdge(In203[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID926 e926 ( .InEdge(Out15), .OutEdge(In203[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID204_INDEGREE4 n204 ( .InEdges(In204), .OutEdge(Out204),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID927 e927 ( .InEdge(Out5), .OutEdge(In204[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID928 e928 ( .InEdge(Out224), .OutEdge(In204[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID929 e929 ( .InEdge(Out79), .OutEdge(In204[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID930 e930 ( .InEdge(Out125), .OutEdge(In204[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID205_INDEGREE1 n205 ( .InEdges(In205), .OutEdge(Out205),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID931 e931 ( .InEdge(Out161), .OutEdge(In205[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID206_INDEGREE6 n206 ( .InEdges(In206), .OutEdge(Out206),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID932 e932 ( .InEdge(Out41), .OutEdge(In206[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID933 e933 ( .InEdge(Out237), .OutEdge(In206[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID934 e934 ( .InEdge(Out93), .OutEdge(In206[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID935 e935 ( .InEdge(Out239), .OutEdge(In206[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID936 e936 ( .InEdge(Out118), .OutEdge(In206[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID937 e937 ( .InEdge(Out23), .OutEdge(In206[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID207_INDEGREE7 n207 ( .InEdges(In207), .OutEdge(Out207),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID938 e938 ( .InEdge(Out24), .OutEdge(In207[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID939 e939 ( .InEdge(Out19), .OutEdge(In207[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID940 e940 ( .InEdge(Out159), .OutEdge(In207[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID941 e941 ( .InEdge(Out69), .OutEdge(In207[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID942 e942 ( .InEdge(Out48), .OutEdge(In207[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID943 e943 ( .InEdge(Out106), .OutEdge(In207[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID944 e944 ( .InEdge(Out79), .OutEdge(In207[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID208_INDEGREE2 n208 ( .InEdges(In208), .OutEdge(Out208),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID945 e945 ( .InEdge(Out0), .OutEdge(In208[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID946 e946 ( .InEdge(Out54), .OutEdge(In208[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID209_INDEGREE8 n209 ( .InEdges(In209), .OutEdge(Out209),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID947 e947 ( .InEdge(Out221), .OutEdge(In209[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID948 e948 ( .InEdge(Out10), .OutEdge(In209[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID949 e949 ( .InEdge(Out146), .OutEdge(In209[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID950 e950 ( .InEdge(Out237), .OutEdge(In209[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID951 e951 ( .InEdge(Out212), .OutEdge(In209[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID952 e952 ( .InEdge(Out118), .OutEdge(In209[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID953 e953 ( .InEdge(Out169), .OutEdge(In209[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID954 e954 ( .InEdge(Out167), .OutEdge(In209[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID210_INDEGREE3 n210 ( .InEdges(In210), .OutEdge(Out210),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID955 e955 ( .InEdge(Out133), .OutEdge(In210[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID956 e956 ( .InEdge(Out47), .OutEdge(In210[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID957 e957 ( .InEdge(Out5), .OutEdge(In210[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID211_INDEGREE7 n211 ( .InEdges(In211), .OutEdge(Out211),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID958 e958 ( .InEdge(Out248), .OutEdge(In211[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID959 e959 ( .InEdge(Out5), .OutEdge(In211[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID960 e960 ( .InEdge(Out31), .OutEdge(In211[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID961 e961 ( .InEdge(Out46), .OutEdge(In211[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID962 e962 ( .InEdge(Out122), .OutEdge(In211[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID963 e963 ( .InEdge(Out22), .OutEdge(In211[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID964 e964 ( .InEdge(Out214), .OutEdge(In211[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID212_INDEGREE2 n212 ( .InEdges(In212), .OutEdge(Out212),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID965 e965 ( .InEdge(Out67), .OutEdge(In212[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID966 e966 ( .InEdge(Out202), .OutEdge(In212[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID213_INDEGREE1 n213 ( .InEdges(In213), .OutEdge(Out213),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID967 e967 ( .InEdge(Out189), .OutEdge(In213[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID214_INDEGREE5 n214 ( .InEdges(In214), .OutEdge(Out214),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID968 e968 ( .InEdge(Out145), .OutEdge(In214[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID969 e969 ( .InEdge(Out34), .OutEdge(In214[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID970 e970 ( .InEdge(Out155), .OutEdge(In214[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID971 e971 ( .InEdge(Out182), .OutEdge(In214[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID972 e972 ( .InEdge(Out250), .OutEdge(In214[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID215_INDEGREE4 n215 ( .InEdges(In215), .OutEdge(Out215),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID973 e973 ( .InEdge(Out157), .OutEdge(In215[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID974 e974 ( .InEdge(Out200), .OutEdge(In215[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID975 e975 ( .InEdge(Out80), .OutEdge(In215[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID976 e976 ( .InEdge(Out114), .OutEdge(In215[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID216_INDEGREE1 n216 ( .InEdges(In216), .OutEdge(Out216),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID977 e977 ( .InEdge(Out116), .OutEdge(In216[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID217_INDEGREE6 n217 ( .InEdges(In217), .OutEdge(Out217),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID978 e978 ( .InEdge(Out189), .OutEdge(In217[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID979 e979 ( .InEdge(Out212), .OutEdge(In217[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID980 e980 ( .InEdge(Out178), .OutEdge(In217[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID981 e981 ( .InEdge(Out238), .OutEdge(In217[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID982 e982 ( .InEdge(Out109), .OutEdge(In217[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID983 e983 ( .InEdge(Out148), .OutEdge(In217[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID218_INDEGREE2 n218 ( .InEdges(In218), .OutEdge(Out218),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID984 e984 ( .InEdge(Out50), .OutEdge(In218[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID985 e985 ( .InEdge(Out7), .OutEdge(In218[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID219_INDEGREE1 n219 ( .InEdges(In219), .OutEdge(Out219),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID986 e986 ( .InEdge(Out73), .OutEdge(In219[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID220_INDEGREE6 n220 ( .InEdges(In220), .OutEdge(Out220),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID987 e987 ( .InEdge(Out151), .OutEdge(In220[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID988 e988 ( .InEdge(Out76), .OutEdge(In220[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID989 e989 ( .InEdge(Out62), .OutEdge(In220[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID990 e990 ( .InEdge(Out247), .OutEdge(In220[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID991 e991 ( .InEdge(Out90), .OutEdge(In220[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID992 e992 ( .InEdge(Out224), .OutEdge(In220[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID221_INDEGREE3 n221 ( .InEdges(In221), .OutEdge(Out221),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID993 e993 ( .InEdge(Out41), .OutEdge(In221[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID994 e994 ( .InEdge(Out60), .OutEdge(In221[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID995 e995 ( .InEdge(Out217), .OutEdge(In221[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID222_INDEGREE3 n222 ( .InEdges(In222), .OutEdge(Out222),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID996 e996 ( .InEdge(Out108), .OutEdge(In222[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID997 e997 ( .InEdge(Out210), .OutEdge(In222[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID998 e998 ( .InEdge(Out137), .OutEdge(In222[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID223_INDEGREE2 n223 ( .InEdges(In223), .OutEdge(Out223),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID999 e999 ( .InEdge(Out55), .OutEdge(In223[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1000 e1000 ( .InEdge(Out70), .OutEdge(In223[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID224_INDEGREE7 n224 ( .InEdges(In224), .OutEdge(Out224),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1001 e1001 ( .InEdge(Out63), .OutEdge(In224[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1002 e1002 ( .InEdge(Out252), .OutEdge(In224[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1003 e1003 ( .InEdge(Out174), .OutEdge(In224[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1004 e1004 ( .InEdge(Out206), .OutEdge(In224[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1005 e1005 ( .InEdge(Out86), .OutEdge(In224[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1006 e1006 ( .InEdge(Out84), .OutEdge(In224[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1007 e1007 ( .InEdge(Out47), .OutEdge(In224[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID225_INDEGREE3 n225 ( .InEdges(In225), .OutEdge(Out225),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1008 e1008 ( .InEdge(Out223), .OutEdge(In225[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1009 e1009 ( .InEdge(Out54), .OutEdge(In225[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1010 e1010 ( .InEdge(Out254), .OutEdge(In225[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID226_INDEGREE2 n226 ( .InEdges(In226), .OutEdge(Out226),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1011 e1011 ( .InEdge(Out140), .OutEdge(In226[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1012 e1012 ( .InEdge(Out27), .OutEdge(In226[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID227_INDEGREE7 n227 ( .InEdges(In227), .OutEdge(Out227),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1013 e1013 ( .InEdge(Out89), .OutEdge(In227[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1014 e1014 ( .InEdge(Out117), .OutEdge(In227[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1015 e1015 ( .InEdge(Out15), .OutEdge(In227[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1016 e1016 ( .InEdge(Out87), .OutEdge(In227[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1017 e1017 ( .InEdge(Out11), .OutEdge(In227[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1018 e1018 ( .InEdge(Out203), .OutEdge(In227[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1019 e1019 ( .InEdge(Out126), .OutEdge(In227[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID228_INDEGREE4 n228 ( .InEdges(In228), .OutEdge(Out228),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1020 e1020 ( .InEdge(Out71), .OutEdge(In228[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1021 e1021 ( .InEdge(Out179), .OutEdge(In228[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1022 e1022 ( .InEdge(Out227), .OutEdge(In228[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1023 e1023 ( .InEdge(Out183), .OutEdge(In228[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID229_INDEGREE2 n229 ( .InEdges(In229), .OutEdge(Out229),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1024 e1024 ( .InEdge(Out110), .OutEdge(In229[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1025 e1025 ( .InEdge(Out25), .OutEdge(In229[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID230_INDEGREE4 n230 ( .InEdges(In230), .OutEdge(Out230),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1026 e1026 ( .InEdge(Out40), .OutEdge(In230[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1027 e1027 ( .InEdge(Out91), .OutEdge(In230[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1028 e1028 ( .InEdge(Out85), .OutEdge(In230[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1029 e1029 ( .InEdge(Out29), .OutEdge(In230[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID231_INDEGREE6 n231 ( .InEdges(In231), .OutEdge(Out231),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1030 e1030 ( .InEdge(Out93), .OutEdge(In231[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1031 e1031 ( .InEdge(Out11), .OutEdge(In231[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1032 e1032 ( .InEdge(Out150), .OutEdge(In231[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1033 e1033 ( .InEdge(Out139), .OutEdge(In231[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1034 e1034 ( .InEdge(Out80), .OutEdge(In231[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1035 e1035 ( .InEdge(Out85), .OutEdge(In231[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID232_INDEGREE6 n232 ( .InEdges(In232), .OutEdge(Out232),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1036 e1036 ( .InEdge(Out195), .OutEdge(In232[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1037 e1037 ( .InEdge(Out179), .OutEdge(In232[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1038 e1038 ( .InEdge(Out146), .OutEdge(In232[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1039 e1039 ( .InEdge(Out126), .OutEdge(In232[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1040 e1040 ( .InEdge(Out62), .OutEdge(In232[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1041 e1041 ( .InEdge(Out242), .OutEdge(In232[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID233_INDEGREE4 n233 ( .InEdges(In233), .OutEdge(Out233),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1042 e1042 ( .InEdge(Out185), .OutEdge(In233[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1043 e1043 ( .InEdge(Out227), .OutEdge(In233[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1044 e1044 ( .InEdge(Out112), .OutEdge(In233[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1045 e1045 ( .InEdge(Out172), .OutEdge(In233[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID234_INDEGREE6 n234 ( .InEdges(In234), .OutEdge(Out234),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1046 e1046 ( .InEdge(Out24), .OutEdge(In234[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1047 e1047 ( .InEdge(Out23), .OutEdge(In234[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1048 e1048 ( .InEdge(Out180), .OutEdge(In234[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1049 e1049 ( .InEdge(Out160), .OutEdge(In234[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1050 e1050 ( .InEdge(Out61), .OutEdge(In234[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1051 e1051 ( .InEdge(Out172), .OutEdge(In234[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID235_INDEGREE6 n235 ( .InEdges(In235), .OutEdge(Out235),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1052 e1052 ( .InEdge(Out238), .OutEdge(In235[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1053 e1053 ( .InEdge(Out248), .OutEdge(In235[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1054 e1054 ( .InEdge(Out156), .OutEdge(In235[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1055 e1055 ( .InEdge(Out135), .OutEdge(In235[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1056 e1056 ( .InEdge(Out116), .OutEdge(In235[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1057 e1057 ( .InEdge(Out132), .OutEdge(In235[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID236_INDEGREE8 n236 ( .InEdges(In236), .OutEdge(Out236),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1058 e1058 ( .InEdge(Out227), .OutEdge(In236[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1059 e1059 ( .InEdge(Out47), .OutEdge(In236[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1060 e1060 ( .InEdge(Out30), .OutEdge(In236[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1061 e1061 ( .InEdge(Out67), .OutEdge(In236[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1062 e1062 ( .InEdge(Out28), .OutEdge(In236[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1063 e1063 ( .InEdge(Out140), .OutEdge(In236[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1064 e1064 ( .InEdge(Out121), .OutEdge(In236[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1065 e1065 ( .InEdge(Out210), .OutEdge(In236[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID237_INDEGREE4 n237 ( .InEdges(In237), .OutEdge(Out237),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1066 e1066 ( .InEdge(Out41), .OutEdge(In237[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1067 e1067 ( .InEdge(Out84), .OutEdge(In237[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1068 e1068 ( .InEdge(Out201), .OutEdge(In237[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1069 e1069 ( .InEdge(Out71), .OutEdge(In237[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID238_INDEGREE2 n238 ( .InEdges(In238), .OutEdge(Out238),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1070 e1070 ( .InEdge(Out65), .OutEdge(In238[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1071 e1071 ( .InEdge(Out34), .OutEdge(In238[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID239_INDEGREE5 n239 ( .InEdges(In239), .OutEdge(Out239),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1072 e1072 ( .InEdge(Out201), .OutEdge(In239[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1073 e1073 ( .InEdge(Out142), .OutEdge(In239[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1074 e1074 ( .InEdge(Out140), .OutEdge(In239[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1075 e1075 ( .InEdge(Out93), .OutEdge(In239[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1076 e1076 ( .InEdge(Out52), .OutEdge(In239[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID240_INDEGREE1 n240 ( .InEdges(In240), .OutEdge(Out240),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1077 e1077 ( .InEdge(Out129), .OutEdge(In240[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID241_INDEGREE3 n241 ( .InEdges(In241), .OutEdge(Out241),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1078 e1078 ( .InEdge(Out232), .OutEdge(In241[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1079 e1079 ( .InEdge(Out15), .OutEdge(In241[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1080 e1080 ( .InEdge(Out148), .OutEdge(In241[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID242_INDEGREE7 n242 ( .InEdges(In242), .OutEdge(Out242),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1081 e1081 ( .InEdge(Out104), .OutEdge(In242[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1082 e1082 ( .InEdge(Out215), .OutEdge(In242[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1083 e1083 ( .InEdge(Out96), .OutEdge(In242[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1084 e1084 ( .InEdge(Out139), .OutEdge(In242[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1085 e1085 ( .InEdge(Out174), .OutEdge(In242[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1086 e1086 ( .InEdge(Out49), .OutEdge(In242[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1087 e1087 ( .InEdge(Out248), .OutEdge(In242[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID243_INDEGREE1 n243 ( .InEdges(In243), .OutEdge(Out243),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1088 e1088 ( .InEdge(Out147), .OutEdge(In243[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID244_INDEGREE8 n244 ( .InEdges(In244), .OutEdge(Out244),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1089 e1089 ( .InEdge(Out60), .OutEdge(In244[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1090 e1090 ( .InEdge(Out193), .OutEdge(In244[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1091 e1091 ( .InEdge(Out183), .OutEdge(In244[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1092 e1092 ( .InEdge(Out246), .OutEdge(In244[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1093 e1093 ( .InEdge(Out106), .OutEdge(In244[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1094 e1094 ( .InEdge(Out9), .OutEdge(In244[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1095 e1095 ( .InEdge(Out199), .OutEdge(In244[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1096 e1096 ( .InEdge(Out151), .OutEdge(In244[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID245_INDEGREE5 n245 ( .InEdges(In245), .OutEdge(Out245),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1097 e1097 ( .InEdge(Out238), .OutEdge(In245[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1098 e1098 ( .InEdge(Out114), .OutEdge(In245[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1099 e1099 ( .InEdge(Out29), .OutEdge(In245[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1100 e1100 ( .InEdge(Out105), .OutEdge(In245[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1101 e1101 ( .InEdge(Out223), .OutEdge(In245[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID246_INDEGREE1 n246 ( .InEdges(In246), .OutEdge(Out246),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1102 e1102 ( .InEdge(Out150), .OutEdge(In246[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID247_INDEGREE6 n247 ( .InEdges(In247), .OutEdge(Out247),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1103 e1103 ( .InEdge(Out111), .OutEdge(In247[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1104 e1104 ( .InEdge(Out67), .OutEdge(In247[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1105 e1105 ( .InEdge(Out189), .OutEdge(In247[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1106 e1106 ( .InEdge(Out198), .OutEdge(In247[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1107 e1107 ( .InEdge(Out53), .OutEdge(In247[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1108 e1108 ( .InEdge(Out230), .OutEdge(In247[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID248_INDEGREE2 n248 ( .InEdges(In248), .OutEdge(Out248),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1109 e1109 ( .InEdge(Out101), .OutEdge(In248[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1110 e1110 ( .InEdge(Out237), .OutEdge(In248[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID249_INDEGREE7 n249 ( .InEdges(In249), .OutEdge(Out249),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1111 e1111 ( .InEdge(Out24), .OutEdge(In249[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1112 e1112 ( .InEdge(Out95), .OutEdge(In249[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1113 e1113 ( .InEdge(Out200), .OutEdge(In249[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1114 e1114 ( .InEdge(Out165), .OutEdge(In249[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1115 e1115 ( .InEdge(Out56), .OutEdge(In249[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1116 e1116 ( .InEdge(Out69), .OutEdge(In249[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1117 e1117 ( .InEdge(Out184), .OutEdge(In249[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID250_INDEGREE1 n250 ( .InEdges(In250), .OutEdge(Out250),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1118 e1118 ( .InEdge(Out184), .OutEdge(In250[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID251_INDEGREE3 n251 ( .InEdges(In251), .OutEdge(Out251),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1119 e1119 ( .InEdge(Out226), .OutEdge(In251[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1120 e1120 ( .InEdge(Out150), .OutEdge(In251[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1121 e1121 ( .InEdge(Out110), .OutEdge(In251[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID252_INDEGREE6 n252 ( .InEdges(In252), .OutEdge(Out252),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1122 e1122 ( .InEdge(Out32), .OutEdge(In252[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1123 e1123 ( .InEdge(Out225), .OutEdge(In252[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1124 e1124 ( .InEdge(Out117), .OutEdge(In252[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1125 e1125 ( .InEdge(Out14), .OutEdge(In252[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1126 e1126 ( .InEdge(Out145), .OutEdge(In252[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1127 e1127 ( .InEdge(Out159), .OutEdge(In252[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID253_INDEGREE4 n253 ( .InEdges(In253), .OutEdge(Out253),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1128 e1128 ( .InEdge(Out50), .OutEdge(In253[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1129 e1129 ( .InEdge(Out144), .OutEdge(In253[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1130 e1130 ( .InEdge(Out83), .OutEdge(In253[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1131 e1131 ( .InEdge(Out99), .OutEdge(In253[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID254_INDEGREE2 n254 ( .InEdges(In254), .OutEdge(Out254),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1132 e1132 ( .InEdge(Out255), .OutEdge(In254[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1133 e1133 ( .InEdge(Out184), .OutEdge(In254[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID255_INDEGREE6 n255 ( .InEdges(In255), .OutEdge(Out255),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1134 e1134 ( .InEdge(Out55), .OutEdge(In255[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1135 e1135 ( .InEdge(Out33), .OutEdge(In255[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1136 e1136 ( .InEdge(Out200), .OutEdge(In255[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1137 e1137 ( .InEdge(Out57), .OutEdge(In255[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1138 e1138 ( .InEdge(Out199), .OutEdge(In255[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1139 e1139 ( .InEdge(Out16), .OutEdge(In255[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
endmodule
