
module Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Load, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
input  [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  Clk, Reset, RD, WR, ScanEnable, Load;
    wire \Out[31] , \Out[5] , n175, n190, n217, n182, n222, n167, n205, n199, 
        n185, n160, n219, n169, n210, n202, n224, n172, n203, n197, \Out[24] , 
        \Out[17] , n161, n184, \Out[30] , n196, n218, \Out[29] , \Out[22] , 
        \Out[20] , \Out[13] , \Out[8] , \Out[1] , n173, n168, n211, \Out[11] , 
        n216, \Out[2] , n183, \Out[18] , \Out[3] , n174, n191, \Out[26] , 
        \Out[15] , n166, n223, \Out[7] , n204, n198, n193, \Out[27] , 
        \Out[14] , n214, n176, \Out[23] , \Out[10] , \Out[6] , n188, n206, 
        n221, \Out[28] , \Out[19] , n164, n181, \Out[0] , n186, \Out[21] , 
        \Out[12] , \Out[9] , n163, n178, n213, n201, \Out[25] , \Out[16] , 
        \Out[4] , n171, n208, n194, n179, n200, n162, n187, n209, n195, n170, 
        n212, n215, n192, n189, n177, n180, n165, n220, n207;
    assign ScanOut[31] = \Out[31] ;
    assign ScanOut[30] = \Out[30] ;
    assign ScanOut[29] = \Out[29] ;
    assign ScanOut[28] = \Out[28] ;
    assign ScanOut[27] = \Out[27] ;
    assign ScanOut[26] = \Out[26] ;
    assign ScanOut[25] = \Out[25] ;
    assign ScanOut[24] = \Out[24] ;
    assign ScanOut[23] = \Out[23] ;
    assign ScanOut[22] = \Out[22] ;
    assign ScanOut[21] = \Out[21] ;
    assign ScanOut[20] = \Out[20] ;
    assign ScanOut[19] = \Out[19] ;
    assign ScanOut[18] = \Out[18] ;
    assign ScanOut[17] = \Out[17] ;
    assign ScanOut[16] = \Out[16] ;
    assign ScanOut[15] = \Out[15] ;
    assign ScanOut[14] = \Out[14] ;
    assign ScanOut[13] = \Out[13] ;
    assign ScanOut[12] = \Out[12] ;
    assign ScanOut[11] = \Out[11] ;
    assign ScanOut[10] = \Out[10] ;
    assign ScanOut[9] = \Out[9] ;
    assign ScanOut[8] = \Out[8] ;
    assign ScanOut[7] = \Out[7] ;
    assign ScanOut[6] = \Out[6] ;
    assign ScanOut[5] = \Out[5] ;
    assign ScanOut[4] = \Out[4] ;
    assign ScanOut[3] = \Out[3] ;
    assign ScanOut[2] = \Out[2] ;
    assign ScanOut[1] = \Out[1] ;
    assign ScanOut[0] = \Out[0] ;
    assign Out[31] = \Out[31] ;
    assign Out[30] = \Out[30] ;
    assign Out[29] = \Out[29] ;
    assign Out[28] = \Out[28] ;
    assign Out[27] = \Out[27] ;
    assign Out[26] = \Out[26] ;
    assign Out[25] = \Out[25] ;
    assign Out[24] = \Out[24] ;
    assign Out[23] = \Out[23] ;
    assign Out[22] = \Out[22] ;
    assign Out[21] = \Out[21] ;
    assign Out[20] = \Out[20] ;
    assign Out[19] = \Out[19] ;
    assign Out[18] = \Out[18] ;
    assign Out[17] = \Out[17] ;
    assign Out[16] = \Out[16] ;
    assign Out[15] = \Out[15] ;
    assign Out[14] = \Out[14] ;
    assign Out[13] = \Out[13] ;
    assign Out[12] = \Out[12] ;
    assign Out[11] = \Out[11] ;
    assign Out[10] = \Out[10] ;
    assign Out[9] = \Out[9] ;
    assign Out[8] = \Out[8] ;
    assign Out[7] = \Out[7] ;
    assign Out[6] = \Out[6] ;
    assign Out[5] = \Out[5] ;
    assign Out[4] = \Out[4] ;
    assign Out[3] = \Out[3] ;
    assign Out[2] = \Out[2] ;
    assign Out[1] = \Out[1] ;
    assign Out[0] = \Out[0] ;
    VMW_AO21 U54 ( .A(\Out[27] ), .B(n160), .C(n188), .Z(n197) );
    VMW_AO21 U73 ( .A(ScanIn[26]), .B(ScanEnable), .C(Reset), .Z(n187) );
    VMW_AO21 U68 ( .A(ScanIn[30]), .B(ScanEnable), .C(Reset), .Z(n191) );
    VMW_AO21 U28 ( .A(\Out[1] ), .B(n160), .C(n162), .Z(n223) );
    VMW_AO21 U33 ( .A(\Out[6] ), .B(n160), .C(n167), .Z(n218) );
    VMW_AO21 U34 ( .A(\Out[7] ), .B(n160), .C(n168), .Z(n217) );
    VMW_AO21 U41 ( .A(\Out[14] ), .B(n160), .C(n175), .Z(n210) );
    VMW_AO21 U46 ( .A(\Out[19] ), .B(n160), .C(n180), .Z(n205) );
    VMW_AO21 U61 ( .A(ScanIn[8]), .B(ScanEnable), .C(Reset), .Z(n169) );
    VMW_AO21 U84 ( .A(ScanIn[16]), .B(ScanEnable), .C(Reset), .Z(n177) );
    VMW_AO21 U66 ( .A(ScanIn[3]), .B(ScanEnable), .C(Reset), .Z(n164) );
    VMW_AO21 U83 ( .A(ScanIn[17]), .B(ScanEnable), .C(Reset), .Z(n178) );
    VMW_AO21 U35 ( .A(\Out[8] ), .B(n160), .C(n169), .Z(n216) );
    VMW_AO21 U48 ( .A(\Out[21] ), .B(n160), .C(n182), .Z(n203) );
    VMW_AO21 U53 ( .A(\Out[26] ), .B(n160), .C(n187), .Z(n198) );
    VMW_AO21 U91 ( .A(ScanIn[0]), .B(ScanEnable), .C(Reset), .Z(n161) );
    VMW_AO21 U74 ( .A(ScanIn[25]), .B(ScanEnable), .C(Reset), .Z(n186) );
    VMW_FD \Out_reg[25]  ( .D(n199), .CP(Clk), .Q(\Out[25] ) );
    VMW_FD \Out_reg[16]  ( .D(n208), .CP(Clk), .Q(\Out[16] ) );
    VMW_AO21 U27 ( .A(\Out[0] ), .B(n160), .C(n161), .Z(n224) );
    VMW_AO21 U40 ( .A(\Out[13] ), .B(n160), .C(n174), .Z(n211) );
    VMW_AO21 U82 ( .A(ScanIn[18]), .B(ScanEnable), .C(Reset), .Z(n179) );
    VMW_FD \Out_reg[5]  ( .D(n219), .CP(Clk), .Q(\Out[5] ) );
    VMW_AO21 U52 ( .A(\Out[25] ), .B(n160), .C(n186), .Z(n199) );
    VMW_AO21 U67 ( .A(ScanIn[31]), .B(ScanEnable), .C(Reset), .Z(n192) );
    VMW_AO21 U75 ( .A(ScanIn[24]), .B(ScanEnable), .C(Reset), .Z(n185) );
    VMW_FD \Out_reg[12]  ( .D(n212), .CP(Clk), .Q(\Out[12] ) );
    VMW_AO21 U90 ( .A(ScanIn[10]), .B(ScanEnable), .C(Reset), .Z(n171) );
    VMW_FD \Out_reg[21]  ( .D(n203), .CP(Clk), .Q(\Out[21] ) );
    VMW_FD \Out_reg[8]  ( .D(n216), .CP(Clk), .Q(\Out[8] ) );
    VMW_AO21 U29 ( .A(\Out[2] ), .B(n160), .C(n163), .Z(n222) );
    VMW_AO21 U47 ( .A(\Out[20] ), .B(n160), .C(n181), .Z(n204) );
    VMW_AO21 U49 ( .A(\Out[22] ), .B(n160), .C(n183), .Z(n202) );
    VMW_FD \Out_reg[31]  ( .D(n193), .CP(Clk), .Q(\Out[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n196), .CP(Clk), .Q(\Out[28] ) );
    VMW_FD \Out_reg[1]  ( .D(n223), .CP(Clk), .Q(\Out[1] ) );
    VMW_AO21 U55 ( .A(\Out[28] ), .B(n160), .C(n189), .Z(n196) );
    VMW_AO21 U69 ( .A(ScanIn[2]), .B(ScanEnable), .C(Reset), .Z(n163) );
    VMW_FD \Out_reg[19]  ( .D(n205), .CP(Clk), .Q(\Out[19] ) );
    VMW_AO21 U72 ( .A(ScanIn[27]), .B(ScanEnable), .C(Reset), .Z(n188) );
    VMW_FD \Out_reg[3]  ( .D(n221), .CP(Clk), .Q(\Out[3] ) );
    VMW_FD \Out_reg[23]  ( .D(n201), .CP(Clk), .Q(\Out[23] ) );
    VMW_FD \Out_reg[10]  ( .D(n214), .CP(Clk), .Q(\Out[10] ) );
    VMW_AO21 U60 ( .A(ScanIn[9]), .B(ScanEnable), .C(Reset), .Z(n170) );
    VMW_FD \Out_reg[7]  ( .D(n217), .CP(Clk), .Q(\Out[7] ) );
    VMW_AO21 U32 ( .A(\Out[5] ), .B(n160), .C(n166), .Z(n219) );
    VMW_AO21 U85 ( .A(ScanIn[15]), .B(ScanEnable), .C(Reset), .Z(n176) );
    VMW_FD \Out_reg[27]  ( .D(n197), .CP(Clk), .Q(\Out[27] ) );
    VMW_FD \Out_reg[14]  ( .D(n210), .CP(Clk), .Q(\Out[14] ) );
    VMW_AO21 U30 ( .A(\Out[3] ), .B(n160), .C(n164), .Z(n221) );
    VMW_AO21 U39 ( .A(\Out[12] ), .B(n160), .C(n173), .Z(n212) );
    VMW_AO21 U57 ( .A(\Out[30] ), .B(n160), .C(n191), .Z(n194) );
    VMW_FD \Out_reg[6]  ( .D(n218), .CP(Clk), .Q(\Out[6] ) );
    VMW_AO21 U70 ( .A(ScanIn[29]), .B(ScanEnable), .C(Reset), .Z(n190) );
    VMW_AO21 U79 ( .A(ScanIn[20]), .B(ScanEnable), .C(Reset), .Z(n181) );
    VMW_FD \Out_reg[26]  ( .D(n198), .CP(Clk), .Q(\Out[26] ) );
    VMW_FD \Out_reg[15]  ( .D(n209), .CP(Clk), .Q(\Out[15] ) );
    VMW_FD \Out_reg[18]  ( .D(n206), .CP(Clk), .Q(\Out[18] ) );
    VMW_AO21 U31 ( .A(\Out[4] ), .B(n160), .C(n165), .Z(n220) );
    VMW_AO21 U36 ( .A(\Out[9] ), .B(n160), .C(n170), .Z(n215) );
    VMW_AO21 U37 ( .A(\Out[10] ), .B(n160), .C(n171), .Z(n214) );
    VMW_AO21 U42 ( .A(\Out[15] ), .B(n160), .C(n176), .Z(n209) );
    VMW_AO21 U45 ( .A(\Out[18] ), .B(n160), .C(n179), .Z(n206) );
    VMW_AO21 U87 ( .A(ScanIn[13]), .B(ScanEnable), .C(Reset), .Z(n174) );
    VMW_FD \Out_reg[2]  ( .D(n222), .CP(Clk), .Q(\Out[2] ) );
    VMW_FD \Out_reg[11]  ( .D(n213), .CP(Clk), .Q(\Out[11] ) );
    VMW_AO21 U62 ( .A(ScanIn[7]), .B(ScanEnable), .C(Reset), .Z(n168) );
    VMW_FD \Out_reg[22]  ( .D(n202), .CP(Clk), .Q(\Out[22] ) );
    VMW_AO21 U65 ( .A(ScanIn[4]), .B(ScanEnable), .C(Reset), .Z(n165) );
    VMW_FD \Out_reg[20]  ( .D(n204), .CP(Clk), .Q(\Out[20] ) );
    VMW_FD \Out_reg[13]  ( .D(n211), .CP(Clk), .Q(\Out[13] ) );
    VMW_AO21 U80 ( .A(ScanIn[1]), .B(ScanEnable), .C(Reset), .Z(n162) );
    VMW_FD \Out_reg[9]  ( .D(n215), .CP(Clk), .Q(\Out[9] ) );
    VMW_AO21 U50 ( .A(\Out[23] ), .B(n160), .C(n184), .Z(n201) );
    VMW_NOR2 U59 ( .A(ScanEnable), .B(Load), .Z(n160) );
    VMW_FD \Out_reg[30]  ( .D(n194), .CP(Clk), .Q(\Out[30] ) );
    VMW_FD \Out_reg[0]  ( .D(n224), .CP(Clk), .Q(\Out[0] ) );
    VMW_FD \Out_reg[29]  ( .D(n195), .CP(Clk), .Q(\Out[29] ) );
    VMW_AO21 U77 ( .A(ScanIn[22]), .B(ScanEnable), .C(Reset), .Z(n183) );
    VMW_AO21 U89 ( .A(ScanIn[11]), .B(ScanEnable), .C(Reset), .Z(n172) );
    VMW_FD \Out_reg[24]  ( .D(n200), .CP(Clk), .Q(\Out[24] ) );
    VMW_FD \Out_reg[17]  ( .D(n207), .CP(Clk), .Q(\Out[17] ) );
    VMW_FD \Out_reg[4]  ( .D(n220), .CP(Clk), .Q(\Out[4] ) );
    VMW_AO21 U58 ( .A(\Out[31] ), .B(n160), .C(n192), .Z(n193) );
    VMW_AO21 U38 ( .A(\Out[11] ), .B(n160), .C(n172), .Z(n213) );
    VMW_AO21 U43 ( .A(\Out[16] ), .B(n160), .C(n177), .Z(n208) );
    VMW_AO21 U64 ( .A(ScanIn[5]), .B(ScanEnable), .C(Reset), .Z(n166) );
    VMW_AO21 U81 ( .A(ScanIn[19]), .B(ScanEnable), .C(Reset), .Z(n180) );
    VMW_AO21 U51 ( .A(\Out[24] ), .B(n160), .C(n185), .Z(n200) );
    VMW_AO21 U76 ( .A(ScanIn[23]), .B(ScanEnable), .C(Reset), .Z(n184) );
    VMW_AO21 U88 ( .A(ScanIn[12]), .B(ScanEnable), .C(Reset), .Z(n173) );
    VMW_AO21 U44 ( .A(\Out[17] ), .B(n160), .C(n178), .Z(n207) );
    VMW_AO21 U56 ( .A(\Out[29] ), .B(n160), .C(n190), .Z(n195) );
    VMW_AO21 U71 ( .A(ScanIn[28]), .B(ScanEnable), .C(Reset), .Z(n189) );
    VMW_AO21 U63 ( .A(ScanIn[6]), .B(ScanEnable), .C(Reset), .Z(n167) );
    VMW_AO21 U86 ( .A(ScanIn[14]), .B(ScanEnable), .C(Reset), .Z(n175) );
    VMW_AO21 U78 ( .A(ScanIn[21]), .B(ScanEnable), .C(Reset), .Z(n182) );
endmodule


module Merge_Node_DWIDTH32_DW01_cmp2_32_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n55, n72, n97, n20, n69, n100, n112, n32, n29, n85, n47, n60, 
        n109, n40, n67, n82, n99, n27, n35, n49, n115, n107, n90, n52, n75, 
        n98, n114, n34, n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, 
        n101, n21, n46, n54, n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, 
        n113, n94, n23, n103, n16, n111, n31, n36, n44, n63, n86, n43, n64, 
        n81, n58, n104, n18, n24, n88, n37, n51, n93, n59, n76, n80, n42, n65, 
        n19, n50, n77, n89, n92, n25, n102, n105, n22, n39, n95, n45, n57, n62, 
        n87, n17, n30, n79, n110;
    VMW_AO21 U3 ( .A(n15), .B(A[31]), .C(n16), .Z(GE_GT) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n18), .C(B[0]), .Z(n19) );
    VMW_AO22 U6 ( .A(A[2]), .B(n21), .C(n19), .D(A[0]), .Z(n20) );
    VMW_OR2 U14 ( .A(B[6]), .B(n30), .Z(n33) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n46), .C(n41), .D(n36), .Z(n45) );
    VMW_OR2 U54 ( .A(B[26]), .B(n96), .Z(n99) );
    VMW_INV U73 ( .A(B[27]), .Z(n105) );
    VMW_INV U96 ( .A(n115), .Z(n16) );
    VMW_INV U68 ( .A(A[30]), .Z(n110) );
    VMW_NAND2 U28 ( .A(n56), .B(B[14]), .Z(n55) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n64), .C(n60), .D(n55), .Z(n63) );
    VMW_OAI22 U7 ( .A(n17), .B(n20), .C(A[2]), .D(n21), .Z(n22) );
    VMW_NAND2 U8 ( .A(n24), .B(B[4]), .Z(n23) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n32), .C(n28), .D(n23), .Z(n31) );
    VMW_OR2 U34 ( .A(B[16]), .B(n62), .Z(n65) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n74), .D(n68), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_OAI211 U61 ( .A(A[29]), .B(n112), .C(n107), .D(n102), .Z(n111) );
    VMW_INV U84 ( .A(A[4]), .Z(n24) );
    VMW_INV U101 ( .A(A[6]), .Z(n30) );
    VMW_INV U66 ( .A(B[7]), .Z(n39) );
    VMW_INV U83 ( .A(B[15]), .Z(n64) );
    VMW_INV U98 ( .A(B[13]), .Z(n58) );
    VMW_NAND2 U26 ( .A(n52), .B(A[11]), .Z(n53) );
    VMW_NAND2 U48 ( .A(n90), .B(B[24]), .Z(n89) );
    VMW_AO21 U9 ( .A(B[3]), .B(n26), .C(n22), .Z(n25) );
    VMW_NAND2 U12 ( .A(n30), .B(B[6]), .Z(n29) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n67), .C(n65), .D(n63), .Z(n66) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n98), .C(n94), .D(n89), .Z(n97) );
    VMW_INV U91 ( .A(A[28]), .Z(n103) );
    VMW_INV U74 ( .A(A[3]), .Z(n26) );
    VMW_INV U99 ( .A(A[26]), .Z(n96) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n50), .C(n53), .D(n51), .Z(n54) );
    VMW_NAND2 U40 ( .A(n77), .B(B[20]), .Z(n76) );
    VMW_INV U82 ( .A(A[15]), .Z(n67) );
    VMW_NAND2 U52 ( .A(n96), .B(B[26]), .Z(n95) );
    VMW_INV U67 ( .A(A[7]), .Z(n42) );
    VMW_INV U75 ( .A(B[25]), .Z(n98) );
    VMW_INV U90 ( .A(B[11]), .Z(n52) );
    VMW_NAND2 U20 ( .A(n44), .B(B[10]), .Z(n43) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n92), .C(n88), .D(n83), .Z(n91) );
    VMW_INV U69 ( .A(B[17]), .Z(n72) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n58), .C(n54), .D(n49), .Z(n57) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n101), .C(n99), .D(n97), .Z(n100) );
    VMW_INV U72 ( .A(A[27]), .Z(n108) );
    VMW_INV U97 ( .A(A[16]), .Z(n62) );
    VMW_NAND2 U60 ( .A(n110), .B(B[30]), .Z(n109) );
    VMW_INV U100 ( .A(B[23]), .Z(n92) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n35), .C(n33), .D(n31), .Z(n34) );
    VMW_INV U85 ( .A(A[24]), .Z(n90) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n39), .C(n34), .D(n29), .Z(n38) );
    VMW_NAND2 U22 ( .A(n46), .B(A[9]), .Z(n47) );
    VMW_NAND2 U32 ( .A(n62), .B(B[16]), .Z(n61) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n75), .C(n73), .D(n71), .Z(n74) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_INV U70 ( .A(A[17]), .Z(n75) );
    VMW_INV U95 ( .A(B[31]), .Z(n15) );
    VMW_NAND2 U30 ( .A(n58), .B(A[13]), .Z(n59) );
    VMW_INV U79 ( .A(A[10]), .Z(n44) );
    VMW_INV U87 ( .A(B[21]), .Z(n86) );
    VMW_OR2 U10 ( .A(B[4]), .B(n24), .Z(n27) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n76), .Z(n85) );
    VMW_NAND2 U62 ( .A(n112), .B(A[29]), .Z(n113) );
    VMW_INV U65 ( .A(A[12]), .Z(n50) );
    VMW_INV U102 ( .A(B[2]), .Z(n21) );
    VMW_INV U80 ( .A(B[9]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n26), .C(n27), .D(n25), .Z(n28) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n42), .C(n40), .D(n38), .Z(n41) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n52), .C(n48), .D(n43), .Z(n51) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n72), .C(n66), .D(n61), .Z(n71) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n108), .C(n106), .D(n104), .Z(n107) );
    VMW_INV U89 ( .A(A[14]), .Z(n56) );
    VMW_NAND2 U50 ( .A(n92), .B(A[23]), .Z(n93) );
    VMW_INV U77 ( .A(A[20]), .Z(n77) );
    VMW_INV U92 ( .A(A[5]), .Z(n35) );
    VMW_OR2 U58 ( .A(B[28]), .B(n103), .Z(n106) );
    VMW_NAND2 U36 ( .A(n69), .B(B[18]), .Z(n68) );
    VMW_INV U81 ( .A(B[29]), .Z(n112) );
    VMW_NOR2 U4 ( .A(n18), .B(B[1]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n37), .Z(n40) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n77), .C(n81), .D(n79), .Z(n82) );
    VMW_OAI211 U64 ( .A(A[31]), .B(n15), .C(n114), .D(n109), .Z(n115) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n90), .C(n93), .D(n91), .Z(n94) );
    VMW_INV U76 ( .A(A[25]), .Z(n101) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n44), .C(n47), .D(n45), .Z(n48) );
    VMW_NAND2 U24 ( .A(n50), .B(B[12]), .Z(n49) );
    VMW_INV U88 ( .A(A[18]), .Z(n69) );
    VMW_INV U93 ( .A(B[5]), .Z(n32) );
    VMW_OR2 U38 ( .A(B[18]), .B(n69), .Z(n73) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n103), .B(B[28]), .Z(n102) );
    VMW_INV U94 ( .A(A[1]), .Z(n18) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_OAI211 U63 ( .A(B[30]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_INV U86 ( .A(A[8]), .Z(n37) );
    VMW_NAND2 U16 ( .A(n37), .B(B[8]), .Z(n36) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n56), .C(n59), .D(n57), .Z(n60) );
    VMW_INV U78 ( .A(B[19]), .Z(n80) );
endmodule


module Merge_Node_DWIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n190, n149, n152, n175, n127, n135, n205, n199, n140, n167, n182, 
        n129, n185, n147, n160, n120, n132, n202, n169, n210, n155, n172, n197, 
        n133, n203, n146, n161, n121, n128, n184, n154, n196, n168, n173, n211, 
        n126, n148, n153, n174, n183, n191, n166, n141, n118, n134, n204, n193, 
        n198, n151, n176, n124, n188, n206, n136, n143, n158, n144, n163, n164, 
        n181, n186, n178, n116, n123, n131, n201, n213, n171, n156, n117, n138, 
        n194, n208, n130, n179, n200, n145, n162, n187, n195, n139, n209, n170, 
        n157, n122, n125, n212, n189, n150, n177, n192, n119, n142, n180, n165, 
        n159, n137, n207;
    VMW_OAI21 U3 ( .A(A[31]), .B(n116), .C(n117), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n119), .C(B[0]), .Z(n120) );
    VMW_AO22 U6 ( .A(A[2]), .B(n122), .C(n120), .D(A[0]), .Z(n121) );
    VMW_OR2 U14 ( .A(B[6]), .B(n131), .Z(n134) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n147), .C(n142), .D(n137), .Z(n146) );
    VMW_OR2 U54 ( .A(B[26]), .B(n195), .Z(n198) );
    VMW_INV U73 ( .A(B[27]), .Z(n204) );
    VMW_INV U96 ( .A(A[16]), .Z(n163) );
    VMW_INV U68 ( .A(A[30]), .Z(n212) );
    VMW_NAND2 U28 ( .A(n157), .B(B[14]), .Z(n156) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n165), .C(n161), .D(n156), .Z(n164) );
    VMW_OAI22 U7 ( .A(n118), .B(n121), .C(A[2]), .D(n122), .Z(n123) );
    VMW_NAND2 U8 ( .A(n125), .B(B[4]), .Z(n124) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n133), .C(n129), .D(n124), .Z(n132) );
    VMW_OR2 U34 ( .A(B[16]), .B(n163), .Z(n166) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n179), .C(n174), .D(n169), .Z(n178) );
    VMW_NAND2 U46 ( .A(n185), .B(A[21]), .Z(n186) );
    VMW_NAND2 U61 ( .A(n209), .B(A[29]), .Z(n210) );
    VMW_INV U84 ( .A(A[4]), .Z(n125) );
    VMW_INV U101 ( .A(B[2]), .Z(n122) );
    VMW_INV U66 ( .A(B[7]), .Z(n140) );
    VMW_INV U83 ( .A(B[15]), .Z(n165) );
    VMW_INV U98 ( .A(A[26]), .Z(n195) );
    VMW_NAND2 U26 ( .A(n153), .B(A[11]), .Z(n154) );
    VMW_NAND2 U48 ( .A(n189), .B(B[24]), .Z(n188) );
    VMW_AO21 U9 ( .A(B[3]), .B(n127), .C(n123), .Z(n126) );
    VMW_NAND2 U12 ( .A(n131), .B(B[6]), .Z(n130) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n168), .C(n166), .D(n164), .Z(n167) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n197), .C(n193), .D(n188), .Z(n196) );
    VMW_INV U91 ( .A(A[28]), .Z(n202) );
    VMW_INV U74 ( .A(A[3]), .Z(n127) );
    VMW_INV U99 ( .A(B[23]), .Z(n191) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n151), .C(n154), .D(n152), .Z(n155) );
    VMW_NAND2 U40 ( .A(n177), .B(B[20]), .Z(n176) );
    VMW_INV U82 ( .A(A[15]), .Z(n168) );
    VMW_NAND2 U52 ( .A(n195), .B(B[26]), .Z(n194) );
    VMW_INV U67 ( .A(A[7]), .Z(n143) );
    VMW_INV U75 ( .A(B[25]), .Z(n197) );
    VMW_INV U90 ( .A(B[11]), .Z(n153) );
    VMW_NAND2 U20 ( .A(n145), .B(B[10]), .Z(n144) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n191), .C(n187), .D(n182), .Z(n190) );
    VMW_INV U69 ( .A(B[17]), .Z(n172) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n159), .C(n155), .D(n150), .Z(n158) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n183), .C(n186), .D(n184), .Z(n187) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n200), .C(n198), .D(n196), .Z(n199) );
    VMW_INV U72 ( .A(A[27]), .Z(n207) );
    VMW_INV U97 ( .A(B[13]), .Z(n159) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n209), .C(n206), .D(n201), .Z(n208) );
    VMW_INV U100 ( .A(A[6]), .Z(n131) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n136), .C(n134), .D(n132), .Z(n135) );
    VMW_INV U85 ( .A(A[24]), .Z(n189) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n140), .C(n135), .D(n130), .Z(n139) );
    VMW_NAND2 U22 ( .A(n147), .B(A[9]), .Z(n148) );
    VMW_NAND2 U32 ( .A(n163), .B(B[16]), .Z(n162) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n175), .C(n173), .D(n171), .Z(n174) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n204), .C(n199), .D(n194), .Z(n203) );
    VMW_INV U70 ( .A(A[17]), .Z(n175) );
    VMW_INV U95 ( .A(B[31]), .Z(n116) );
    VMW_NAND2 U30 ( .A(n159), .B(A[13]), .Z(n160) );
    VMW_INV U79 ( .A(A[10]), .Z(n145) );
    VMW_INV U87 ( .A(B[21]), .Z(n185) );
    VMW_OR2 U10 ( .A(B[4]), .B(n125), .Z(n128) );
    VMW_NAND2 U42 ( .A(n179), .B(A[19]), .Z(n180) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n185), .C(n181), .D(n176), .Z(n184) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n212), .C(n210), .D(n208), .Z(n211) );
    VMW_INV U65 ( .A(A[12]), .Z(n151) );
    VMW_INV U80 ( .A(B[9]), .Z(n147) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n127), .C(n128), .D(n126), .Z(n129) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n143), .C(n141), .D(n139), .Z(n142) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n153), .C(n149), .D(n144), .Z(n152) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n172), .C(n167), .D(n162), .Z(n171) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n207), .C(n205), .D(n203), .Z(n206) );
    VMW_INV U89 ( .A(A[14]), .Z(n157) );
    VMW_NAND2 U50 ( .A(n191), .B(A[23]), .Z(n192) );
    VMW_INV U77 ( .A(A[20]), .Z(n177) );
    VMW_INV U92 ( .A(A[5]), .Z(n136) );
    VMW_OR2 U58 ( .A(B[28]), .B(n202), .Z(n205) );
    VMW_NAND2 U36 ( .A(n170), .B(B[18]), .Z(n169) );
    VMW_INV U81 ( .A(B[29]), .Z(n209) );
    VMW_NOR2 U4 ( .A(n119), .B(B[1]), .Z(n118) );
    VMW_OR2 U18 ( .A(B[8]), .B(n138), .Z(n141) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n177), .C(n180), .D(n178), .Z(n181) );
    VMW_AO22 U64 ( .A(n211), .B(n213), .C(A[31]), .D(n116), .Z(n117) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n189), .C(n192), .D(n190), .Z(n193) );
    VMW_INV U76 ( .A(A[25]), .Z(n200) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n145), .C(n148), .D(n146), .Z(n149) );
    VMW_NAND2 U24 ( .A(n151), .B(B[12]), .Z(n150) );
    VMW_INV U88 ( .A(A[18]), .Z(n170) );
    VMW_INV U93 ( .A(B[5]), .Z(n133) );
    VMW_OR2 U38 ( .A(B[18]), .B(n170), .Z(n173) );
    VMW_NAND2 U44 ( .A(n183), .B(B[22]), .Z(n182) );
    VMW_NAND2 U56 ( .A(n202), .B(B[28]), .Z(n201) );
    VMW_INV U94 ( .A(A[1]), .Z(n119) );
    VMW_INV U71 ( .A(A[22]), .Z(n183) );
    VMW_NAND2 U63 ( .A(n212), .B(B[30]), .Z(n213) );
    VMW_INV U86 ( .A(A[8]), .Z(n138) );
    VMW_NAND2 U16 ( .A(n138), .B(B[8]), .Z(n137) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n157), .C(n160), .D(n158), .Z(n161) );
    VMW_INV U78 ( .A(B[19]), .Z(n179) );
endmodule


module Merge_Node_DWIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, Load, 
    Out, In1, In2, Read1, Read2 );
input  [14:0] Addr;
input  [31:0] DataIn;
input  [31:0] DataOut;
input  [31:0] In1;
output [31:0] Out;
input  [31:0] In2;
input  Clk, Reset, RD, WR, Load;
output Read1, Read2;
    wire n337, n339, n217, n287, n330, n317, n245, n262, n279, n230, n222, 
        n219, n257, n270, n239, n295, n305, n322, n292, n325, n302, n250, n277, 
        n225, n289, n319, n237, n259, n265, n242, n336, n218, n224, n280, n310, 
        n251, n276, n288, n318, n293, n303, n324, n338, n216, n231, n236, n243, 
        n264, n281, n311, n258, n278, n223, n238, n244, n263, n286, n316, n294, 
        n331, n304, n323, n256, n271, n70, n215, n214, n228, n284, n333, n314, 
        n246, n261, n221, n233, n328, n226, n248, n254, n268, n78, n273, n253, 
        n291, n296, n321, n301, n306, n326, n274, n227, n234, n241, n298, n308, 
        n266, n283, n313, n334, n249, n252, n275, n282, n290, n300, n327, n312, 
        n335, n235, n240, n267, n299, n309, n232, n329, n247, n260, n332, n229, 
        n285, n315, n297, n307, n320, n255, n272, n220, n269;
    VMW_PULLDOWN U36 ( .Z(n337) );
    VMW_PULLUP U37 ( .Z(n336) );
    VMW_PULLUP U39 ( .Z(n338) );
    VMW_OAI21 U40 ( .A(n70), .B(n215), .C(Load), .Z(n214) );
    VMW_AO21 U41 ( .A(n215), .B(n217), .C(Reset), .Z(n216) );
    VMW_AOI211 U46 ( .A(n219), .B(In2[5]), .C(n228), .D(n216), .Z(n227) );
    VMW_AOI211 U54 ( .A(n219), .B(In2[27]), .C(n244), .D(n216), .Z(n243) );
    VMW_AOI211 U73 ( .A(n219), .B(In2[0]), .C(n282), .D(n216), .Z(n281) );
    VMW_AO22 U113 ( .A(Out[22]), .B(n293), .C(n294), .D(In1[22]), .Z(n254) );
    VMW_INV U134 ( .A(n225), .Z(n329) );
    VMW_AOI211 U61 ( .A(n219), .B(In2[20]), .C(n258), .D(n216), .Z(n257) );
    VMW_AOI211 U68 ( .A(n219), .B(In2[14]), .C(n272), .D(n216), .Z(n271) );
    VMW_AO22 U96 ( .A(Out[9]), .B(n293), .C(n294), .D(In1[9]), .Z(n220) );
    VMW_AO22 U108 ( .A(Out[27]), .B(n293), .C(n294), .D(In1[27]), .Z(n244) );
    VMW_INV U141 ( .A(n239), .Z(n306) );
    Merge_Node_DWIDTH32_DW01_cmp2_32_1 r140 ( .A(In1), .B(In2), .LEQ(n338), 
        .TC(n339), .GE_GT(n70) );
    VMW_AND4 U84 ( .A(In2[23]), .B(In2[22]), .C(In2[21]), .D(In2[20]), .Z(n285
        ) );
    VMW_INV U148 ( .A(n253), .Z(n313) );
    VMW_INV U153 ( .A(n263), .Z(n317) );
    VMW_AO22 U101 ( .A(Out[4]), .B(n293), .C(n294), .D(In1[4]), .Z(n230) );
    VMW_AO22 U126 ( .A(Out[10]), .B(n293), .C(n294), .D(In1[10]), .Z(n280) );
    VMW_AOI211 U48 ( .A(n219), .B(In2[3]), .C(n232), .D(n216), .Z(n231) );
    VMW_AOI211 U66 ( .A(n219), .B(In2[16]), .C(n268), .D(n216), .Z(n267) );
    VMW_AO22 U106 ( .A(Out[29]), .B(n293), .C(n294), .D(In1[29]), .Z(n240) );
    VMW_AO22 U121 ( .A(Out[15]), .B(n293), .C(n294), .D(In1[15]), .Z(n270) );
    VMW_AND4 U83 ( .A(In2[19]), .B(In2[18]), .C(In2[17]), .D(In2[16]), .Z(n286
        ) );
    VMW_AO22 U98 ( .A(Out[7]), .B(n293), .C(n294), .D(In1[7]), .Z(n224) );
    VMW_OAI21 U128 ( .A(n78), .B(n217), .C(Load), .Z(n303) );
    VMW_INV U154 ( .A(n265), .Z(n318) );
    VMW_AOI211 U53 ( .A(n219), .B(In2[28]), .C(n242), .D(n216), .Z(n241) );
    VMW_AND4 U91 ( .A(n302), .B(n301), .C(n300), .D(n299), .Z(n292) );
    VMW_INV U146 ( .A(n249), .Z(n311) );
    VMW_INV U161 ( .A(n279), .Z(n325) );
    VMW_AND5 U74 ( .A(n283), .B(n284), .C(n285), .D(n286), .E(n287), .Z(n217)
         );
    VMW_AO22 U114 ( .A(Out[21]), .B(n293), .C(n294), .D(In1[21]), .Z(n256) );
    VMW_INV U133 ( .A(n223), .Z(n328) );
    VMW_AND4 U82 ( .A(n298), .B(n297), .C(n296), .D(n295), .Z(n287) );
    VMW_AO22 U99 ( .A(Out[6]), .B(n293), .C(n294), .D(In1[6]), .Z(n226) );
    VMW_INV U155 ( .A(n267), .Z(n319) );
    VMW_FD \Out_reg[16]  ( .D(n319), .CP(Clk), .Q(Out[16]) );
    VMW_FD \Out_reg[25]  ( .D(n310), .CP(Clk), .Q(Out[25]) );
    VMW_FD \Out_reg[5]  ( .D(n330), .CP(Clk), .Q(Out[5]) );
    VMW_AOI211 U47 ( .A(n219), .B(In2[4]), .C(n230), .D(n216), .Z(n229) );
    VMW_AOI211 U49 ( .A(n219), .B(In2[31]), .C(n234), .D(n216), .Z(n233) );
    VMW_AOI211 U52 ( .A(n219), .B(In2[29]), .C(n240), .D(n216), .Z(n239) );
    VMW_AOI211 U67 ( .A(n219), .B(In2[15]), .C(n270), .D(n216), .Z(n269) );
    VMW_AO22 U107 ( .A(Out[28]), .B(n293), .C(n294), .D(In1[28]), .Z(n242) );
    VMW_AO22 U120 ( .A(Out[16]), .B(n293), .C(n294), .D(In1[16]), .Z(n268) );
    VMW_AND5 U75 ( .A(n288), .B(n289), .C(n290), .D(n291), .E(n292), .Z(n215)
         );
    VMW_AO22 U115 ( .A(Out[20]), .B(n293), .C(n294), .D(In1[20]), .Z(n258) );
    VMW_INV U132 ( .A(n221), .Z(n327) );
    VMW_FD \Out_reg[12]  ( .D(n323), .CP(Clk), .Q(Out[12]) );
    VMW_AND4 U90 ( .A(In1[15]), .B(In1[14]), .C(In1[13]), .D(In1[12]), .Z(n302
        ) );
    VMW_FD \Out_reg[21]  ( .D(n314), .CP(Clk), .Q(Out[21]) );
    VMW_INV U129 ( .A(n214), .Z(Read1) );
    VMW_INV U147 ( .A(n251), .Z(n312) );
    VMW_FD \Out_reg[8]  ( .D(n327), .CP(Clk), .Q(Out[8]) );
    VMW_INV U160 ( .A(n277), .Z(n324) );
    VMW_FD \Out_reg[31]  ( .D(n304), .CP(Clk), .Q(Out[31]) );
    VMW_FD \Out_reg[28]  ( .D(n307), .CP(Clk), .Q(Out[28]) );
    VMW_FD \Out_reg[1]  ( .D(n334), .CP(Clk), .Q(Out[1]) );
    VMW_AOI211 U55 ( .A(n219), .B(In2[26]), .C(n246), .D(n216), .Z(n245) );
    VMW_AOI211 U69 ( .A(n219), .B(In2[13]), .C(n274), .D(n216), .Z(n273) );
    VMW_AO22 U109 ( .A(Out[26]), .B(n293), .C(n294), .D(In1[26]), .Z(n246) );
    VMW_FD \Out_reg[19]  ( .D(n316), .CP(Clk), .Q(Out[19]) );
    VMW_AOI211 U72 ( .A(n219), .B(In2[10]), .C(n280), .D(n216), .Z(n279) );
    VMW_AO22 U97 ( .A(Out[8]), .B(n293), .C(n294), .D(In1[8]), .Z(n222) );
    VMW_INV U140 ( .A(n237), .Z(n333) );
    VMW_FD \Out_reg[3]  ( .D(n332), .CP(Clk), .Q(Out[3]) );
    VMW_AO22 U112 ( .A(Out[23]), .B(n293), .C(n294), .D(In1[23]), .Z(n252) );
    VMW_INV U135 ( .A(n227), .Z(n330) );
    VMW_FD \Out_reg[10]  ( .D(n325), .CP(Clk), .Q(Out[10]) );
    VMW_FD \Out_reg[23]  ( .D(n312), .CP(Clk), .Q(Out[23]) );
    VMW_AOI211 U60 ( .A(n219), .B(In2[21]), .C(n256), .D(n216), .Z(n255) );
    VMW_FD \Out_reg[7]  ( .D(n328), .CP(Clk), .Q(Out[7]) );
    VMW_AO22 U100 ( .A(Out[5]), .B(n293), .C(n294), .D(In1[5]), .Z(n228) );
    VMW_AO22 U127 ( .A(Out[0]), .B(n293), .C(n294), .D(In1[0]), .Z(n282) );
    VMW_AOI211 U57 ( .A(n219), .B(In2[24]), .C(n250), .D(n216), .Z(n249) );
    VMW_AND4 U85 ( .A(In2[27]), .B(In2[26]), .C(In2[25]), .D(In2[24]), .Z(n284
        ) );
    VMW_INV U149 ( .A(n255), .Z(n314) );
    VMW_INV U137 ( .A(n231), .Z(n332) );
    VMW_INV U152 ( .A(n261), .Z(n316) );
    VMW_FD \Out_reg[27]  ( .D(n308), .CP(Clk), .Q(Out[27]) );
    VMW_FD \Out_reg[14]  ( .D(n321), .CP(Clk), .Q(Out[14]) );
    VMW_FD \Out_reg[6]  ( .D(n329), .CP(Clk), .Q(Out[6]) );
    VMW_AOI211 U70 ( .A(n219), .B(In2[12]), .C(n276), .D(n216), .Z(n275) );
    VMW_AO22 U110 ( .A(Out[25]), .B(n293), .C(n294), .D(In1[25]), .Z(n248) );
    VMW_INV U159 ( .A(n275), .Z(n323) );
    VMW_AOI211 U42 ( .A(n219), .B(In2[9]), .C(n220), .D(n216), .Z(n218) );
    VMW_AOI211 U45 ( .A(n219), .B(In2[6]), .C(n226), .D(n216), .Z(n225) );
    VMW_AND4 U79 ( .A(In2[7]), .B(In2[6]), .C(In2[5]), .D(In2[4]), .Z(n296) );
    VMW_AND4 U95 ( .A(In1[31]), .B(In1[30]), .C(In1[29]), .D(In1[28]), .Z(n288
        ) );
    VMW_AO22 U119 ( .A(Out[17]), .B(n293), .C(n294), .D(In1[17]), .Z(n266) );
    VMW_INV U142 ( .A(n241), .Z(n307) );
    VMW_FD \Out_reg[26]  ( .D(n309), .CP(Clk), .Q(Out[26]) );
    VMW_FD \Out_reg[15]  ( .D(n320), .CP(Clk), .Q(Out[15]) );
    VMW_FD \Out_reg[18]  ( .D(n317), .CP(Clk), .Q(Out[18]) );
    VMW_AND4 U87 ( .A(In1[3]), .B(In1[2]), .C(In1[1]), .D(In1[0]), .Z(n299) );
    VMW_INV U150 ( .A(n257), .Z(n315) );
    VMW_FD \Out_reg[2]  ( .D(n333), .CP(Clk), .Q(Out[2]) );
    VMW_AO22 U125 ( .A(Out[11]), .B(n293), .C(n294), .D(In1[11]), .Z(n278) );
    VMW_FD \Out_reg[11]  ( .D(n324), .CP(Clk), .Q(Out[11]) );
    VMW_AOI211 U62 ( .A(n219), .B(In2[1]), .C(n260), .D(n216), .Z(n259) );
    VMW_FD \Out_reg[22]  ( .D(n313), .CP(Clk), .Q(Out[22]) );
    VMW_AOI211 U65 ( .A(n219), .B(In2[17]), .C(n266), .D(n216), .Z(n265) );
    VMW_AO22 U102 ( .A(Out[3]), .B(n293), .C(n294), .D(In1[3]), .Z(n232) );
    VMW_AO22 U105 ( .A(Out[2]), .B(n293), .C(n294), .D(In1[2]), .Z(n238) );
    VMW_FD \Out_reg[20]  ( .D(n315), .CP(Clk), .Q(Out[20]) );
    VMW_FD \Out_reg[13]  ( .D(n322), .CP(Clk), .Q(Out[13]) );
    VMW_AND4 U80 ( .A(In2[11]), .B(In2[10]), .C(In2[9]), .D(In2[8]), .Z(n297)
         );
    VMW_AO22 U122 ( .A(Out[14]), .B(n293), .C(n294), .D(In1[14]), .Z(n272) );
    VMW_INV U157 ( .A(n271), .Z(n321) );
    VMW_FD \Out_reg[9]  ( .D(n326), .CP(Clk), .Q(Out[9]) );
    VMW_AOI211 U50 ( .A(n219), .B(In2[30]), .C(n236), .D(n216), .Z(n235) );
    VMW_AOI211 U59 ( .A(n219), .B(In2[22]), .C(n254), .D(n216), .Z(n253) );
    VMW_INV U139 ( .A(n235), .Z(n305) );
    VMW_FD \Out_reg[30]  ( .D(n305), .CP(Clk), .Q(Out[30]) );
    VMW_FD \Out_reg[0]  ( .D(n335), .CP(Clk), .Q(Out[0]) );
    VMW_FD \Out_reg[29]  ( .D(n306), .CP(Clk), .Q(Out[29]) );
    VMW_AND2 U77 ( .A(n70), .B(Load), .Z(n294) );
    VMW_AND4 U89 ( .A(In1[11]), .B(In1[10]), .C(In1[9]), .D(In1[8]), .Z(n301)
         );
    VMW_AND4 U92 ( .A(In1[19]), .B(In1[18]), .C(In1[17]), .D(In1[16]), .Z(n291
        ) );
    VMW_INV U145 ( .A(n247), .Z(n310) );
    VMW_INV U162 ( .A(n281), .Z(n335) );
    VMW_FD \Out_reg[24]  ( .D(n311), .CP(Clk), .Q(Out[24]) );
    VMW_FD \Out_reg[17]  ( .D(n318), .CP(Clk), .Q(Out[17]) );
    VMW_AO22 U117 ( .A(Out[19]), .B(n293), .C(n294), .D(In1[19]), .Z(n262) );
    VMW_FD \Out_reg[4]  ( .D(n331), .CP(Clk), .Q(Out[4]) );
    VMW_AOI211 U58 ( .A(n219), .B(In2[23]), .C(n252), .D(n216), .Z(n251) );
    VMW_INV U130 ( .A(Load), .Z(n293) );
    VMW_INV U138 ( .A(n233), .Z(n304) );
    VMW_INV U156 ( .A(n269), .Z(n320) );
    VMW_PULLDOWN U38 ( .Z(n339) );
    VMW_AOI211 U43 ( .A(n219), .B(In2[8]), .C(n222), .D(n216), .Z(n221) );
    VMW_AOI211 U64 ( .A(n219), .B(In2[18]), .C(n264), .D(n216), .Z(n263) );
    VMW_AND4 U81 ( .A(In2[15]), .B(In2[14]), .C(In2[13]), .D(In2[12]), .Z(n298
        ) );
    VMW_AO22 U104 ( .A(Out[30]), .B(n293), .C(n294), .D(In1[30]), .Z(n236) );
    VMW_AOI211 U51 ( .A(n219), .B(In2[2]), .C(n238), .D(n216), .Z(n237) );
    VMW_NOR2 U76 ( .A(n293), .B(n70), .Z(n219) );
    VMW_AO22 U116 ( .A(Out[1]), .B(n293), .C(n294), .D(In1[1]), .Z(n260) );
    VMW_AO22 U123 ( .A(Out[13]), .B(n293), .C(n294), .D(In1[13]), .Z(n274) );
    VMW_AND4 U88 ( .A(In1[7]), .B(In1[6]), .C(In1[5]), .D(In1[4]), .Z(n300) );
    VMW_AND4 U93 ( .A(In1[23]), .B(In1[22]), .C(In1[21]), .D(In1[20]), .Z(n290
        ) );
    VMW_INV U131 ( .A(n218), .Z(n326) );
    VMW_INV U143 ( .A(n243), .Z(n308) );
    VMW_INV U144 ( .A(n245), .Z(n309) );
    VMW_INV U163 ( .A(n303), .Z(Read2) );
    VMW_INV U158 ( .A(n273), .Z(n322) );
    VMW_AOI211 U44 ( .A(n219), .B(In2[7]), .C(n224), .D(n216), .Z(n223) );
    VMW_AOI211 U56 ( .A(n219), .B(In2[25]), .C(n248), .D(n216), .Z(n247) );
    VMW_AND4 U94 ( .A(In1[27]), .B(In1[26]), .C(In1[25]), .D(In1[24]), .Z(n289
        ) );
    VMW_INV U136 ( .A(n229), .Z(n331) );
    VMW_AOI211 U71 ( .A(n219), .B(In2[11]), .C(n278), .D(n216), .Z(n277) );
    VMW_AO22 U111 ( .A(Out[24]), .B(n293), .C(n294), .D(In1[24]), .Z(n250) );
    VMW_AO22 U124 ( .A(Out[12]), .B(n293), .C(n294), .D(In1[12]), .Z(n276) );
    Merge_Node_DWIDTH32_DW01_cmp2_32_0 lte_86 ( .A(In1), .B(In2), .LEQ(n336), 
        .TC(n337), .LT_LE(n78) );
    VMW_AOI211 U63 ( .A(n219), .B(In2[19]), .C(n262), .D(n216), .Z(n261) );
    VMW_AND4 U78 ( .A(In2[3]), .B(In2[2]), .C(In2[1]), .D(In2[0]), .Z(n295) );
    VMW_AND4 U86 ( .A(In2[31]), .B(In2[30]), .C(In2[29]), .D(In2[28]), .Z(n283
        ) );
    VMW_AO22 U103 ( .A(Out[31]), .B(n293), .C(n294), .D(In1[31]), .Z(n234) );
    VMW_AO22 U118 ( .A(Out[18]), .B(n293), .C(n294), .D(In1[18]), .Z(n264) );
    VMW_INV U151 ( .A(n259), .Z(n334) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_1 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n112, n32, n29, n85, n47, n60, n109, 
        n40, n67, n82, n99, n27, n35, n49, n107, n90, n52, n75, n98, n114, n34, 
        n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, n21, n46, n54, 
        n96, n73, n61, n28, n84, n33, n38, n56, n71, n113, n94, n23, n103, n16, 
        n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, n58, n104, n18, n24, 
        n88, n37, n51, n93, n59, n76, n80, n42, n65, n19, n50, n77, n89, n92, 
        n25, n102, n105, n22, n39, n95, n45, n57, n70, n62, n87, n17, n30, n79, 
        n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n18), .C(B[0]), .Z(n19) );
    VMW_AO22 U6 ( .A(A[2]), .B(n21), .C(n19), .D(A[0]), .Z(n20) );
    VMW_OR2 U14 ( .A(B[6]), .B(n30), .Z(n33) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n46), .C(n41), .D(n36), .Z(n45) );
    VMW_OR2 U54 ( .A(B[26]), .B(n94), .Z(n97) );
    VMW_INV U73 ( .A(B[27]), .Z(n104) );
    VMW_INV U96 ( .A(A[16]), .Z(n62) );
    VMW_INV U68 ( .A(A[30]), .Z(n113) );
    VMW_NAND2 U28 ( .A(n56), .B(B[14]), .Z(n55) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n64), .C(n60), .D(n55), .Z(n63) );
    VMW_OAI22 U7 ( .A(n17), .B(n20), .C(A[2]), .D(n21), .Z(n22) );
    VMW_NAND2 U8 ( .A(n24), .B(B[4]), .Z(n23) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n32), .C(n28), .D(n23), .Z(n31) );
    VMW_OR2 U34 ( .A(B[16]), .B(n62), .Z(n65) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n78), .C(n73), .D(n68), .Z(n77) );
    VMW_NAND2 U46 ( .A(n84), .B(A[21]), .Z(n85) );
    VMW_NAND2 U61 ( .A(n110), .B(A[29]), .Z(n111) );
    VMW_INV U84 ( .A(A[4]), .Z(n24) );
    VMW_INV U101 ( .A(B[2]), .Z(n21) );
    VMW_INV U66 ( .A(B[7]), .Z(n39) );
    VMW_INV U83 ( .A(B[15]), .Z(n64) );
    VMW_INV U98 ( .A(A[26]), .Z(n94) );
    VMW_NAND2 U26 ( .A(n52), .B(A[11]), .Z(n53) );
    VMW_NAND2 U48 ( .A(n88), .B(B[24]), .Z(n87) );
    VMW_AO21 U9 ( .A(B[3]), .B(n26), .C(n22), .Z(n25) );
    VMW_NAND2 U12 ( .A(n30), .B(B[6]), .Z(n29) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n67), .C(n65), .D(n63), .Z(n66) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n96), .C(n92), .D(n87), .Z(n95) );
    VMW_INV U91 ( .A(A[28]), .Z(n102) );
    VMW_INV U74 ( .A(A[3]), .Z(n26) );
    VMW_INV U99 ( .A(B[23]), .Z(n90) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n50), .C(n53), .D(n51), .Z(n54) );
    VMW_NAND2 U40 ( .A(n76), .B(B[20]), .Z(n75) );
    VMW_INV U82 ( .A(A[15]), .Z(n67) );
    VMW_NAND2 U52 ( .A(n94), .B(B[26]), .Z(n93) );
    VMW_INV U67 ( .A(A[7]), .Z(n42) );
    VMW_INV U75 ( .A(B[25]), .Z(n96) );
    VMW_INV U90 ( .A(B[11]), .Z(n52) );
    VMW_NAND2 U20 ( .A(n44), .B(B[10]), .Z(n43) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n90), .C(n86), .D(n81), .Z(n89) );
    VMW_INV U69 ( .A(B[17]), .Z(n71) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n58), .C(n54), .D(n49), .Z(n57) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n82), .C(n85), .D(n83), .Z(n86) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n99), .C(n97), .D(n95), .Z(n98) );
    VMW_INV U72 ( .A(A[27]), .Z(n107) );
    VMW_INV U97 ( .A(B[13]), .Z(n58) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n110), .C(n106), .D(n101), .Z(n109) );
    VMW_INV U100 ( .A(A[6]), .Z(n30) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n35), .C(n33), .D(n31), .Z(n34) );
    VMW_INV U85 ( .A(A[24]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n39), .C(n34), .D(n29), .Z(n38) );
    VMW_NAND2 U22 ( .A(n46), .B(A[9]), .Z(n47) );
    VMW_NAND2 U32 ( .A(n62), .B(B[16]), .Z(n61) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n74), .C(n72), .D(n70), .Z(n73) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n104), .C(n98), .D(n93), .Z(n103) );
    VMW_INV U70 ( .A(A[17]), .Z(n74) );
    VMW_INV U95 ( .A(B[31]), .Z(n15) );
    VMW_NAND2 U30 ( .A(n58), .B(A[13]), .Z(n59) );
    VMW_INV U79 ( .A(A[10]), .Z(n44) );
    VMW_INV U87 ( .A(B[21]), .Z(n84) );
    VMW_OR2 U10 ( .A(B[4]), .B(n24), .Z(n27) );
    VMW_NAND2 U42 ( .A(n78), .B(A[19]), .Z(n79) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n84), .C(n80), .D(n75), .Z(n83) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n113), .C(n111), .D(n109), .Z(n112) );
    VMW_INV U65 ( .A(A[12]), .Z(n50) );
    VMW_INV U80 ( .A(B[9]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n26), .C(n27), .D(n25), .Z(n28) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n42), .C(n40), .D(n38), .Z(n41) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n52), .C(n48), .D(n43), .Z(n51) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n71), .C(n66), .D(n61), .Z(n70) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n107), .C(n105), .D(n103), .Z(n106) );
    VMW_INV U89 ( .A(A[14]), .Z(n56) );
    VMW_NAND2 U50 ( .A(n90), .B(A[23]), .Z(n91) );
    VMW_INV U77 ( .A(A[20]), .Z(n76) );
    VMW_INV U92 ( .A(A[5]), .Z(n35) );
    VMW_OR2 U58 ( .A(B[28]), .B(n102), .Z(n105) );
    VMW_NAND2 U36 ( .A(n69), .B(B[18]), .Z(n68) );
    VMW_INV U81 ( .A(B[29]), .Z(n110) );
    VMW_NOR2 U4 ( .A(n18), .B(B[1]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n37), .Z(n40) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n76), .C(n79), .D(n77), .Z(n80) );
    VMW_AO22 U64 ( .A(n112), .B(n114), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n88), .C(n91), .D(n89), .Z(n92) );
    VMW_INV U76 ( .A(A[25]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n44), .C(n47), .D(n45), .Z(n48) );
    VMW_NAND2 U24 ( .A(n50), .B(B[12]), .Z(n49) );
    VMW_INV U88 ( .A(A[18]), .Z(n69) );
    VMW_INV U93 ( .A(B[5]), .Z(n32) );
    VMW_OR2 U38 ( .A(B[18]), .B(n69), .Z(n72) );
    VMW_NAND2 U44 ( .A(n82), .B(B[22]), .Z(n81) );
    VMW_NAND2 U56 ( .A(n102), .B(B[28]), .Z(n101) );
    VMW_INV U94 ( .A(A[1]), .Z(n18) );
    VMW_INV U71 ( .A(A[22]), .Z(n82) );
    VMW_NAND2 U63 ( .A(n113), .B(B[30]), .Z(n114) );
    VMW_INV U86 ( .A(A[8]), .Z(n37) );
    VMW_NAND2 U16 ( .A(n37), .B(B[8]), .Z(n36) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n56), .C(n59), .D(n57), .Z(n60) );
    VMW_INV U78 ( .A(B[19]), .Z(n78) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_0 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n115, n190, n149, n152, n175, n127, n135, n205, n199, n140, n167, 
        n182, n129, n185, n147, n160, n132, n202, n120, n169, n210, n155, n172, 
        n197, n133, n203, n146, n161, n121, n128, n184, n154, n196, n168, n173, 
        n211, n126, n148, n153, n174, n183, n191, n166, n141, n118, n134, n204, 
        n193, n198, n151, n176, n124, n188, n206, n136, n144, n143, n158, n164, 
        n163, n181, n186, n178, n116, n123, n131, n201, n213, n171, n156, n117, 
        n138, n194, n208, n130, n179, n200, n145, n162, n187, n195, n139, n209, 
        n170, n157, n122, n125, n212, n189, n150, n177, n192, n119, n142, n180, 
        n165, n159, n137, n207;
    VMW_AO21 U3 ( .A(n115), .B(A[31]), .C(n116), .Z(GE_GT) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n118), .C(B[0]), .Z(n119) );
    VMW_AO22 U6 ( .A(A[2]), .B(n121), .C(n119), .D(A[0]), .Z(n120) );
    VMW_OR2 U14 ( .A(B[6]), .B(n130), .Z(n133) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n146), .C(n141), .D(n136), .Z(n145) );
    VMW_OR2 U54 ( .A(B[26]), .B(n194), .Z(n197) );
    VMW_INV U73 ( .A(B[27]), .Z(n203) );
    VMW_INV U96 ( .A(n213), .Z(n116) );
    VMW_INV U68 ( .A(A[30]), .Z(n208) );
    VMW_NAND2 U28 ( .A(n156), .B(B[14]), .Z(n155) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_OAI22 U7 ( .A(n117), .B(n120), .C(A[2]), .D(n121), .Z(n122) );
    VMW_NAND2 U8 ( .A(n124), .B(B[4]), .Z(n123) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n132), .C(n128), .D(n123), .Z(n131) );
    VMW_OR2 U34 ( .A(B[16]), .B(n162), .Z(n165) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n178), .C(n173), .D(n168), .Z(n177) );
    VMW_NAND2 U46 ( .A(n184), .B(A[21]), .Z(n185) );
    VMW_OAI211 U61 ( .A(A[29]), .B(n210), .C(n205), .D(n200), .Z(n209) );
    VMW_INV U84 ( .A(A[4]), .Z(n124) );
    VMW_INV U101 ( .A(A[6]), .Z(n130) );
    VMW_INV U66 ( .A(B[7]), .Z(n139) );
    VMW_INV U83 ( .A(B[15]), .Z(n164) );
    VMW_INV U98 ( .A(B[13]), .Z(n158) );
    VMW_NAND2 U26 ( .A(n152), .B(A[11]), .Z(n153) );
    VMW_NAND2 U48 ( .A(n188), .B(B[24]), .Z(n187) );
    VMW_AO21 U9 ( .A(B[3]), .B(n126), .C(n122), .Z(n125) );
    VMW_NAND2 U12 ( .A(n130), .B(B[6]), .Z(n129) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n167), .C(n165), .D(n163), .Z(n166) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n196), .C(n192), .D(n187), .Z(n195) );
    VMW_INV U91 ( .A(A[28]), .Z(n201) );
    VMW_INV U74 ( .A(A[3]), .Z(n126) );
    VMW_INV U99 ( .A(A[26]), .Z(n194) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U40 ( .A(n176), .B(B[20]), .Z(n175) );
    VMW_INV U82 ( .A(A[15]), .Z(n167) );
    VMW_NAND2 U52 ( .A(n194), .B(B[26]), .Z(n193) );
    VMW_INV U67 ( .A(A[7]), .Z(n142) );
    VMW_INV U75 ( .A(B[25]), .Z(n196) );
    VMW_INV U90 ( .A(B[11]), .Z(n152) );
    VMW_NAND2 U20 ( .A(n144), .B(B[10]), .Z(n143) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n190), .C(n186), .D(n181), .Z(n189) );
    VMW_INV U69 ( .A(B[17]), .Z(n171) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n182), .C(n185), .D(n183), .Z(n186) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n199), .C(n197), .D(n195), .Z(n198) );
    VMW_INV U72 ( .A(A[27]), .Z(n206) );
    VMW_INV U97 ( .A(A[16]), .Z(n162) );
    VMW_NAND2 U60 ( .A(n208), .B(B[30]), .Z(n207) );
    VMW_INV U100 ( .A(B[23]), .Z(n190) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n135), .C(n133), .D(n131), .Z(n134) );
    VMW_INV U85 ( .A(A[24]), .Z(n188) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n139), .C(n134), .D(n129), .Z(n138) );
    VMW_NAND2 U22 ( .A(n146), .B(A[9]), .Z(n147) );
    VMW_NAND2 U32 ( .A(n162), .B(B[16]), .Z(n161) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n174), .C(n172), .D(n170), .Z(n173) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n203), .C(n198), .D(n193), .Z(n202) );
    VMW_INV U70 ( .A(A[17]), .Z(n174) );
    VMW_INV U95 ( .A(B[31]), .Z(n115) );
    VMW_NAND2 U30 ( .A(n158), .B(A[13]), .Z(n159) );
    VMW_INV U79 ( .A(A[10]), .Z(n144) );
    VMW_INV U87 ( .A(B[21]), .Z(n184) );
    VMW_OR2 U10 ( .A(B[4]), .B(n124), .Z(n127) );
    VMW_NAND2 U42 ( .A(n178), .B(A[19]), .Z(n179) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n184), .C(n180), .D(n175), .Z(n183) );
    VMW_NAND2 U62 ( .A(n210), .B(A[29]), .Z(n211) );
    VMW_INV U65 ( .A(A[12]), .Z(n150) );
    VMW_INV U102 ( .A(B[2]), .Z(n121) );
    VMW_INV U80 ( .A(B[9]), .Z(n146) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n126), .C(n127), .D(n125), .Z(n128) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n142), .C(n140), .D(n138), .Z(n141) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n152), .C(n148), .D(n143), .Z(n151) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n171), .C(n166), .D(n161), .Z(n170) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n206), .C(n204), .D(n202), .Z(n205) );
    VMW_INV U89 ( .A(A[14]), .Z(n156) );
    VMW_NAND2 U50 ( .A(n190), .B(A[23]), .Z(n191) );
    VMW_INV U77 ( .A(A[20]), .Z(n176) );
    VMW_INV U92 ( .A(A[5]), .Z(n135) );
    VMW_OR2 U58 ( .A(B[28]), .B(n201), .Z(n204) );
    VMW_NAND2 U36 ( .A(n169), .B(B[18]), .Z(n168) );
    VMW_INV U81 ( .A(B[29]), .Z(n210) );
    VMW_NOR2 U4 ( .A(n118), .B(B[1]), .Z(n117) );
    VMW_OR2 U18 ( .A(B[8]), .B(n137), .Z(n140) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n176), .C(n179), .D(n177), .Z(n180) );
    VMW_OAI211 U64 ( .A(A[31]), .B(n115), .C(n212), .D(n207), .Z(n213) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n188), .C(n191), .D(n189), .Z(n192) );
    VMW_INV U76 ( .A(A[25]), .Z(n199) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n144), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U24 ( .A(n150), .B(B[12]), .Z(n149) );
    VMW_INV U88 ( .A(A[18]), .Z(n169) );
    VMW_INV U93 ( .A(B[5]), .Z(n132) );
    VMW_OR2 U38 ( .A(B[18]), .B(n169), .Z(n172) );
    VMW_NAND2 U44 ( .A(n182), .B(B[22]), .Z(n181) );
    VMW_NAND2 U56 ( .A(n201), .B(B[28]), .Z(n200) );
    VMW_INV U94 ( .A(A[1]), .Z(n118) );
    VMW_INV U71 ( .A(A[22]), .Z(n182) );
    VMW_OAI211 U63 ( .A(B[30]), .B(n208), .C(n211), .D(n209), .Z(n212) );
    VMW_INV U86 ( .A(A[8]), .Z(n137) );
    VMW_NAND2 U16 ( .A(n137), .B(B[8]), .Z(n136) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_INV U78 ( .A(B[19]), .Z(n178) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, In1, In2, Read1, 
    Read2, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] In1;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In2;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Read1, Read2;
    wire \Out[31] , n100, n245, n287, n317, n330, n262, n279, n362, n345, n357, 
        n339, n270, n257, n295, n305, n322, n292, n325, n302, n250, n277, n350, 
        n289, n319, n259, n342, n365, n265, n359, n356, \Out[5] , n280, n310, 
        n337, n288, n318, n351, \Out[24] , \Out[17] , n276, n251, \Out[30] , 
        n293, n303, n324, n281, n336, n311, \Out[29] , \Out[8] , \Out[1] , 
        n358, n243, n264, n258, n343, n364, \Out[20] , \Out[13] , \Out[26] , 
        \Out[22] , \Out[11] , \Out[18] , \Out[3] , n344, n278, n363, n244, 
        n263, n286, n316, n331, \Out[15] , n294, n304, n323, n256, n108, n271, 
        \Out[27] , \Out[14] , \Out[7] , n338, n284, n314, n333, n246, n261, 
        n361, n346, \Out[6] , n328, \Out[28] , \Out[23] , \Out[10] , \Out[19] , 
        \Out[2] , n268, n354, n368, n254, n273, n321, n306, n296, \Out[9] , 
        \Out[0] , n291, n301, n326, n348, n274, n253, n248, n353, \Out[25] , 
        \Out[21] , \Out[12] , \Out[16] , \Out[4] , n366, n298, n308, n341, 
        n266, n283, n313, n334, n249, n352, n349, n252, n275, n282, n290, n300, 
        n312, n327, n335, n267, n315, n367, n340, n299, n309, n329, n360, n347, 
        n247, n260, n332, n285, n269, n255, n297, n307, n320, n272, n355;
    assign ScanEnable = WR;
    assign DataOut[31] = \Out[31] ;
    assign DataOut[30] = \Out[30] ;
    assign DataOut[29] = \Out[29] ;
    assign DataOut[28] = \Out[28] ;
    assign DataOut[27] = \Out[27] ;
    assign DataOut[26] = \Out[26] ;
    assign DataOut[25] = \Out[25] ;
    assign DataOut[24] = \Out[24] ;
    assign DataOut[23] = \Out[23] ;
    assign DataOut[22] = \Out[22] ;
    assign DataOut[21] = \Out[21] ;
    assign DataOut[20] = \Out[20] ;
    assign DataOut[19] = \Out[19] ;
    assign DataOut[18] = \Out[18] ;
    assign DataOut[17] = \Out[17] ;
    assign DataOut[16] = \Out[16] ;
    assign DataOut[15] = \Out[15] ;
    assign DataOut[14] = \Out[14] ;
    assign DataOut[13] = \Out[13] ;
    assign DataOut[12] = \Out[12] ;
    assign DataOut[11] = \Out[11] ;
    assign DataOut[10] = \Out[10] ;
    assign DataOut[9] = \Out[9] ;
    assign DataOut[8] = \Out[8] ;
    assign DataOut[7] = \Out[7] ;
    assign DataOut[6] = \Out[6] ;
    assign DataOut[5] = \Out[5] ;
    assign DataOut[4] = \Out[4] ;
    assign DataOut[3] = \Out[3] ;
    assign DataOut[2] = \Out[2] ;
    assign DataOut[1] = \Out[1] ;
    assign DataOut[0] = \Out[0] ;
    assign Out[31] = \Out[31] ;
    assign Out[30] = \Out[30] ;
    assign Out[29] = \Out[29] ;
    assign Out[28] = \Out[28] ;
    assign Out[27] = \Out[27] ;
    assign Out[26] = \Out[26] ;
    assign Out[25] = \Out[25] ;
    assign Out[24] = \Out[24] ;
    assign Out[23] = \Out[23] ;
    assign Out[22] = \Out[22] ;
    assign Out[21] = \Out[21] ;
    assign Out[20] = \Out[20] ;
    assign Out[19] = \Out[19] ;
    assign Out[18] = \Out[18] ;
    assign Out[17] = \Out[17] ;
    assign Out[16] = \Out[16] ;
    assign Out[15] = \Out[15] ;
    assign Out[14] = \Out[14] ;
    assign Out[13] = \Out[13] ;
    assign Out[12] = \Out[12] ;
    assign Out[11] = \Out[11] ;
    assign Out[10] = \Out[10] ;
    assign Out[9] = \Out[9] ;
    assign Out[8] = \Out[8] ;
    assign Out[7] = \Out[7] ;
    assign Out[6] = \Out[6] ;
    assign Out[5] = \Out[5] ;
    assign Out[4] = \Out[4] ;
    assign Out[3] = \Out[3] ;
    assign Out[2] = \Out[2] ;
    assign Out[1] = \Out[1] ;
    assign Out[0] = \Out[0] ;
    VMW_AND2 U54 ( .A(DataIn[24]), .B(ScanEnable), .Z(ScanOut[24]) );
    VMW_AND2 U73 ( .A(DataIn[5]), .B(ScanEnable), .Z(ScanOut[5]) );
    VMW_AND5 U113 ( .A(n317), .B(n318), .C(n319), .D(n320), .E(n321), .Z(n246)
         );
    VMW_AO22 U134 ( .A(\Out[9] ), .B(n322), .C(n323), .D(In1[9]), .Z(n249) );
    VMW_AND2 U68 ( .A(DataIn[10]), .B(ScanEnable), .Z(ScanOut[10]) );
    VMW_AOI211 U96 ( .A(n248), .B(In2[23]), .C(n281), .D(n245), .Z(n280) );
    VMW_INV U198 ( .A(n306), .Z(n353) );
    VMW_AOI211 U108 ( .A(n248), .B(In2[12]), .C(n305), .D(n245), .Z(n304) );
    VMW_AO22 U141 ( .A(\Out[31] ), .B(n322), .C(n323), .D(In1[31]), .Z(n263)
         );
    VMW_OAI21 U166 ( .A(n108), .B(n246), .C(RD), .Z(n332) );
    VMW_INV U183 ( .A(n276), .Z(n339) );
    VMW_OAI21 U46 ( .A(n100), .B(n244), .C(RD), .Z(n243) );
    VMW_AND2 U61 ( .A(DataIn[17]), .B(ScanEnable), .Z(ScanOut[17]) );
    VMW_AOI211 U84 ( .A(n248), .B(In2[5]), .C(n257), .D(n245), .Z(n256) );
    VMW_AO22 U148 ( .A(\Out[25] ), .B(n322), .C(n323), .D(In1[25]), .Z(n277)
         );
    VMW_AO22 U153 ( .A(\Out[20] ), .B(n322), .C(n323), .D(In1[20]), .Z(n287)
         );
    VMW_INV U174 ( .A(n258), .Z(n360) );
    VMW_INV U191 ( .A(n292), .Z(n346) );
    VMW_AOI211 U101 ( .A(n248), .B(In2[19]), .C(n291), .D(n245), .Z(n290) );
    VMW_AND4 U126 ( .A(In1[7]), .B(In1[6]), .C(In1[5]), .D(In1[4]), .Z(n329)
         );
    VMW_AND2 U48 ( .A(DataIn[30]), .B(ScanEnable), .Z(ScanOut[30]) );
    VMW_AND2 U66 ( .A(DataIn[12]), .B(ScanEnable), .Z(ScanOut[12]) );
    VMW_AOI211 U106 ( .A(n248), .B(In2[14]), .C(n301), .D(n245), .Z(n300) );
    VMW_AND4 U121 ( .A(In2[19]), .B(In2[18]), .C(In2[17]), .D(In2[16]), .Z(
        n320) );
    VMW_AOI211 U83 ( .A(n248), .B(In2[6]), .C(n255), .D(n245), .Z(n254) );
    VMW_INV U168 ( .A(RD), .Z(n322) );
    VMW_AOI211 U98 ( .A(n248), .B(In2[21]), .C(n285), .D(n245), .Z(n284) );
    VMW_AND4 U128 ( .A(In1[15]), .B(In1[14]), .C(In1[13]), .D(In1[12]), .Z(
        n331) );
    VMW_AO22 U154 ( .A(\Out[1] ), .B(n322), .C(n323), .D(In1[1]), .Z(n289) );
    VMW_INV U173 ( .A(n256), .Z(n359) );
    VMW_INV U184 ( .A(n278), .Z(n340) );
    VMW_INV U196 ( .A(n302), .Z(n351) );
    VMW_AND2 U53 ( .A(DataIn[25]), .B(ScanEnable), .Z(ScanOut[25]) );
    VMW_AOI211 U91 ( .A(n248), .B(In2[28]), .C(n271), .D(n245), .Z(n270) );
    VMW_AO22 U146 ( .A(\Out[27] ), .B(n322), .C(n323), .D(In1[27]), .Z(n273)
         );
    VMW_AO22 U161 ( .A(\Out[13] ), .B(n322), .C(n323), .D(In1[13]), .Z(n303)
         );
    VMW_AND2 U74 ( .A(DataIn[4]), .B(ScanEnable), .Z(ScanOut[4]) );
    VMW_NOR2 U114 ( .A(n322), .B(n100), .Z(n248) );
    VMW_AND4 U133 ( .A(In1[31]), .B(In1[30]), .C(In1[29]), .D(In1[28]), .Z(
        n312) );
    VMW_AOI211 U99 ( .A(n248), .B(In2[20]), .C(n287), .D(n245), .Z(n286) );
    VMW_INV U197 ( .A(n304), .Z(n352) );
    VMW_AO22 U155 ( .A(\Out[19] ), .B(n322), .C(n323), .D(In1[19]), .Z(n291)
         );
    VMW_FD \Out_reg[16]  ( .D(n348), .CP(Clk), .Q(\Out[16] ) );
    VMW_INV U172 ( .A(n254), .Z(n358) );
    VMW_FD \Out_reg[25]  ( .D(n339), .CP(Clk), .Q(\Out[25] ) );
    VMW_AND2 U47 ( .A(DataIn[31]), .B(ScanEnable), .Z(ScanOut[31]) );
    VMW_AND2 U49 ( .A(DataIn[29]), .B(ScanEnable), .Z(ScanOut[29]) );
    VMW_AND2 U52 ( .A(DataIn[26]), .B(ScanEnable), .Z(ScanOut[26]) );
    VMW_AND2 U67 ( .A(DataIn[11]), .B(ScanEnable), .Z(ScanOut[11]) );
    VMW_AOI211 U82 ( .A(n248), .B(In2[7]), .C(n253), .D(n245), .Z(n252) );
    VMW_INV U169 ( .A(n247), .Z(n355) );
    VMW_AOI211 U107 ( .A(n248), .B(In2[13]), .C(n303), .D(n245), .Z(n302) );
    VMW_AND4 U120 ( .A(n327), .B(n326), .C(n325), .D(n324), .Z(n321) );
    VMW_FD \Out_reg[5]  ( .D(n359), .CP(Clk), .Q(\Out[5] ) );
    VMW_AND2 U75 ( .A(DataIn[3]), .B(ScanEnable), .Z(ScanOut[3]) );
    VMW_AND2 U115 ( .A(n100), .B(RD), .Z(n323) );
    VMW_AND4 U132 ( .A(In1[27]), .B(In1[26]), .C(In1[25]), .D(In1[24]), .Z(
        n313) );
    VMW_FD \Out_reg[12]  ( .D(n352), .CP(Clk), .Q(\Out[12] ) );
    VMW_AOI211 U90 ( .A(n248), .B(In2[29]), .C(n269), .D(n245), .Z(n268) );
    VMW_FD \Out_reg[21]  ( .D(n343), .CP(Clk), .Q(\Out[21] ) );
    VMW_AND4 U129 ( .A(n331), .B(n330), .C(n329), .D(n328), .Z(n316) );
    VMW_AO22 U147 ( .A(\Out[26] ), .B(n322), .C(n323), .D(In1[26]), .Z(n275)
         );
    VMW_FD \Out_reg[8]  ( .D(n356), .CP(Clk), .Q(\Out[8] ) );
    VMW_AO22 U160 ( .A(\Out[14] ), .B(n322), .C(n323), .D(In1[14]), .Z(n301)
         );
    VMW_INV U185 ( .A(n280), .Z(n341) );
    VMW_FD \Out_reg[31]  ( .D(n333), .CP(Clk), .Q(\Out[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n336), .CP(Clk), .Q(\Out[28] ) );
    VMW_FD \Out_reg[1]  ( .D(n363), .CP(Clk), .Q(\Out[1] ) );
    VMW_AND2 U55 ( .A(DataIn[23]), .B(ScanEnable), .Z(ScanOut[23]) );
    VMW_AND2 U69 ( .A(ScanEnable), .B(DataIn[9]), .Z(ScanOut[9]) );
    VMW_AOI211 U109 ( .A(n248), .B(In2[11]), .C(n307), .D(n245), .Z(n306) );
    VMW_INV U182 ( .A(n274), .Z(n338) );
    VMW_FD \Out_reg[19]  ( .D(n345), .CP(Clk), .Q(\Out[19] ) );
    VMW_AND2 U72 ( .A(DataIn[6]), .B(ScanEnable), .Z(ScanOut[6]) );
    VMW_AOI211 U97 ( .A(n248), .B(In2[22]), .C(n283), .D(n245), .Z(n282) );
    VMW_AO22 U140 ( .A(\Out[3] ), .B(n322), .C(n323), .D(In1[3]), .Z(n261) );
    VMW_INV U167 ( .A(n243), .Z(Read1) );
    VMW_FD \Out_reg[3]  ( .D(n361), .CP(Clk), .Q(\Out[3] ) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_0 r141 ( .A(In1), .B(
        In2), .LEQ(n365), .TC(n366), .GE_GT(n100) );
    VMW_AND5 U112 ( .A(n312), .B(n313), .C(n314), .D(n315), .E(n316), .Z(n244)
         );
    VMW_AO22 U135 ( .A(\Out[8] ), .B(n322), .C(n323), .D(In1[8]), .Z(n251) );
    VMW_FD \Out_reg[10]  ( .D(n354), .CP(Clk), .Q(\Out[10] ) );
    VMW_FD \Out_reg[23]  ( .D(n341), .CP(Clk), .Q(\Out[23] ) );
    VMW_AND2 U60 ( .A(DataIn[18]), .B(ScanEnable), .Z(ScanOut[18]) );
    VMW_INV U199 ( .A(n308), .Z(n354) );
    VMW_FD \Out_reg[7]  ( .D(n357), .CP(Clk), .Q(\Out[7] ) );
    VMW_AOI211 U100 ( .A(n248), .B(In2[1]), .C(n289), .D(n245), .Z(n288) );
    VMW_AND4 U127 ( .A(In1[11]), .B(In1[10]), .C(In1[9]), .D(In1[8]), .Z(n330)
         );
    VMW_AOI211 U85 ( .A(n248), .B(In2[4]), .C(n259), .D(n245), .Z(n258) );
    VMW_AO22 U149 ( .A(\Out[24] ), .B(n322), .C(n323), .D(In1[24]), .Z(n279)
         );
    VMW_AO22 U152 ( .A(\Out[21] ), .B(n322), .C(n323), .D(In1[21]), .Z(n285)
         );
    VMW_INV U175 ( .A(n260), .Z(n361) );
    VMW_FD \Out_reg[14]  ( .D(n350), .CP(Clk), .Q(\Out[14] ) );
    VMW_FD \Out_reg[27]  ( .D(n337), .CP(Clk), .Q(\Out[27] ) );
    VMW_PULLDOWN U42 ( .Z(n366) );
    VMW_PULLUP U45 ( .Z(n367) );
    VMW_AND2 U57 ( .A(DataIn[21]), .B(ScanEnable), .Z(ScanOut[21]) );
    VMW_AO22 U137 ( .A(\Out[6] ), .B(n322), .C(n323), .D(In1[6]), .Z(n255) );
    VMW_INV U190 ( .A(n290), .Z(n345) );
    VMW_FD \Out_reg[6]  ( .D(n358), .CP(Clk), .Q(\Out[6] ) );
    VMW_AND2 U70 ( .A(DataIn[8]), .B(ScanEnable), .Z(ScanOut[8]) );
    VMW_AO21 U79 ( .A(n246), .B(n244), .C(Reset), .Z(n245) );
    VMW_AOI211 U95 ( .A(n248), .B(In2[24]), .C(n279), .D(n245), .Z(n278) );
    VMW_AOI211 U110 ( .A(n248), .B(In2[10]), .C(n309), .D(n245), .Z(n308) );
    VMW_AO22 U159 ( .A(\Out[15] ), .B(n322), .C(n323), .D(In1[15]), .Z(n299)
         );
    VMW_AND4 U119 ( .A(In2[15]), .B(In2[14]), .C(In2[13]), .D(In2[12]), .Z(
        n327) );
    VMW_AO22 U142 ( .A(\Out[30] ), .B(n322), .C(n323), .D(In1[30]), .Z(n265)
         );
    VMW_AO22 U165 ( .A(\Out[0] ), .B(n322), .C(n323), .D(In1[0]), .Z(n311) );
    VMW_INV U180 ( .A(n270), .Z(n336) );
    VMW_FD \Out_reg[26]  ( .D(n338), .CP(Clk), .Q(\Out[26] ) );
    VMW_FD \Out_reg[15]  ( .D(n349), .CP(Clk), .Q(\Out[15] ) );
    VMW_INV U192 ( .A(n294), .Z(n347) );
    VMW_FD \Out_reg[18]  ( .D(n346), .CP(Clk), .Q(\Out[18] ) );
    VMW_AOI211 U87 ( .A(n248), .B(In2[31]), .C(n263), .D(n245), .Z(n262) );
    VMW_AO22 U150 ( .A(\Out[23] ), .B(n322), .C(n323), .D(In1[23]), .Z(n281)
         );
    VMW_INV U177 ( .A(n264), .Z(n334) );
    VMW_FD \Out_reg[2]  ( .D(n362), .CP(Clk), .Q(\Out[2] ) );
    VMW_AND4 U125 ( .A(In1[3]), .B(In1[2]), .C(In1[1]), .D(In1[0]), .Z(n328)
         );
    VMW_FD \Out_reg[11]  ( .D(n353), .CP(Clk), .Q(\Out[11] ) );
    VMW_AND2 U62 ( .A(DataIn[16]), .B(ScanEnable), .Z(ScanOut[16]) );
    VMW_FD \Out_reg[22]  ( .D(n342), .CP(Clk), .Q(\Out[22] ) );
    VMW_AND2 U65 ( .A(DataIn[13]), .B(ScanEnable), .Z(ScanOut[13]) );
    VMW_AOI211 U102 ( .A(n248), .B(In2[18]), .C(n293), .D(n245), .Z(n292) );
    VMW_AOI211 U105 ( .A(n248), .B(In2[15]), .C(n299), .D(n245), .Z(n298) );
    VMW_INV U189 ( .A(n288), .Z(n363) );
    VMW_FD \Out_reg[20]  ( .D(n344), .CP(Clk), .Q(\Out[20] ) );
    VMW_FD \Out_reg[13]  ( .D(n351), .CP(Clk), .Q(\Out[13] ) );
    VMW_PULLUP U43 ( .Z(n365) );
    VMW_AND2 U50 ( .A(DataIn[28]), .B(ScanEnable), .Z(ScanOut[28]) );
    VMW_AND2 U59 ( .A(DataIn[19]), .B(ScanEnable), .Z(ScanOut[19]) );
    VMW_AOI211 U80 ( .A(n248), .B(In2[9]), .C(n249), .D(n245), .Z(n247) );
    VMW_AND4 U122 ( .A(In2[23]), .B(In2[22]), .C(In2[21]), .D(In2[20]), .Z(
        n319) );
    VMW_AO22 U139 ( .A(\Out[4] ), .B(n322), .C(n323), .D(In1[4]), .Z(n259) );
    VMW_AO22 U157 ( .A(\Out[17] ), .B(n322), .C(n323), .D(In1[17]), .Z(n295)
         );
    VMW_INV U170 ( .A(n250), .Z(n356) );
    VMW_FD \Out_reg[9]  ( .D(n355), .CP(Clk), .Q(\Out[9] ) );
    VMW_INV U195 ( .A(n300), .Z(n350) );
    VMW_FD \Out_reg[30]  ( .D(n334), .CP(Clk), .Q(\Out[30] ) );
    VMW_FD \Out_reg[0]  ( .D(n364), .CP(Clk), .Q(\Out[0] ) );
    VMW_FD \Out_reg[29]  ( .D(n335), .CP(Clk), .Q(\Out[29] ) );
    VMW_AND2 U77 ( .A(DataIn[1]), .B(ScanEnable), .Z(ScanOut[1]) );
    VMW_AOI211 U89 ( .A(n248), .B(In2[2]), .C(n267), .D(n245), .Z(n266) );
    VMW_INV U187 ( .A(n284), .Z(n343) );
    VMW_AOI211 U92 ( .A(n248), .B(In2[27]), .C(n273), .D(n245), .Z(n272) );
    VMW_AO22 U145 ( .A(\Out[28] ), .B(n322), .C(n323), .D(In1[28]), .Z(n271)
         );
    VMW_AO22 U162 ( .A(\Out[12] ), .B(n322), .C(n323), .D(In1[12]), .Z(n305)
         );
    VMW_INV U179 ( .A(n268), .Z(n335) );
    VMW_FD \Out_reg[24]  ( .D(n340), .CP(Clk), .Q(\Out[24] ) );
    VMW_FD \Out_reg[17]  ( .D(n347), .CP(Clk), .Q(\Out[17] ) );
    VMW_AND4 U117 ( .A(In2[7]), .B(In2[6]), .C(In2[5]), .D(In2[4]), .Z(n325)
         );
    VMW_FD \Out_reg[4]  ( .D(n360), .CP(Clk), .Q(\Out[4] ) );
    VMW_INV U200 ( .A(n310), .Z(n364) );
    VMW_AND2 U58 ( .A(DataIn[20]), .B(ScanEnable), .Z(ScanOut[20]) );
    VMW_AND4 U130 ( .A(In1[19]), .B(In1[18]), .C(In1[17]), .D(In1[16]), .Z(
        n315) );
    VMW_AO22 U138 ( .A(\Out[5] ), .B(n322), .C(n323), .D(In1[5]), .Z(n257) );
    VMW_INV U194 ( .A(n298), .Z(n349) );
    VMW_AND2 U64 ( .A(DataIn[14]), .B(ScanEnable), .Z(ScanOut[14]) );
    VMW_AOI211 U81 ( .A(n248), .B(In2[8]), .C(n251), .D(n245), .Z(n250) );
    VMW_AO22 U156 ( .A(\Out[18] ), .B(n322), .C(n323), .D(In1[18]), .Z(n293)
         );
    VMW_INV U171 ( .A(n252), .Z(n357) );
    VMW_AOI211 U104 ( .A(n248), .B(In2[16]), .C(n297), .D(n245), .Z(n296) );
    VMW_PULLDOWN U44 ( .Z(n368) );
    VMW_AND2 U51 ( .A(DataIn[27]), .B(ScanEnable), .Z(ScanOut[27]) );
    VMW_AND2 U76 ( .A(DataIn[2]), .B(ScanEnable), .Z(ScanOut[2]) );
    VMW_AND4 U116 ( .A(In2[3]), .B(In2[2]), .C(In2[1]), .D(In2[0]), .Z(n324)
         );
    VMW_AND4 U123 ( .A(In2[27]), .B(In2[26]), .C(In2[25]), .D(In2[24]), .Z(
        n318) );
    VMW_AND2 U56 ( .A(DataIn[22]), .B(ScanEnable), .Z(ScanOut[22]) );
    VMW_AOI211 U88 ( .A(n248), .B(In2[30]), .C(n265), .D(n245), .Z(n264) );
    VMW_AOI211 U93 ( .A(n248), .B(In2[26]), .C(n275), .D(n245), .Z(n274) );
    VMW_AND4 U131 ( .A(In1[23]), .B(In1[22]), .C(In1[21]), .D(In1[20]), .Z(
        n314) );
    VMW_INV U201 ( .A(n332), .Z(Read2) );
    VMW_INV U178 ( .A(n266), .Z(n362) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_1 lte_43 ( .A(In1), 
        .B(In2), .LEQ(n367), .TC(n368), .LT_LE(n108) );
    VMW_AOI211 U94 ( .A(n248), .B(In2[25]), .C(n277), .D(n245), .Z(n276) );
    VMW_AO22 U143 ( .A(\Out[2] ), .B(n322), .C(n323), .D(In1[2]), .Z(n267) );
    VMW_AO22 U144 ( .A(\Out[29] ), .B(n322), .C(n323), .D(In1[29]), .Z(n269)
         );
    VMW_AO22 U163 ( .A(\Out[11] ), .B(n322), .C(n323), .D(In1[11]), .Z(n307)
         );
    VMW_INV U181 ( .A(n272), .Z(n337) );
    VMW_INV U186 ( .A(n282), .Z(n342) );
    VMW_AO22 U158 ( .A(\Out[16] ), .B(n322), .C(n323), .D(In1[16]), .Z(n297)
         );
    VMW_AO22 U164 ( .A(\Out[10] ), .B(n322), .C(n323), .D(In1[10]), .Z(n309)
         );
    VMW_AO22 U136 ( .A(\Out[7] ), .B(n322), .C(n323), .D(In1[7]), .Z(n253) );
    VMW_AND2 U71 ( .A(DataIn[7]), .B(ScanEnable), .Z(ScanOut[7]) );
    VMW_AOI211 U111 ( .A(n248), .B(In2[0]), .C(n311), .D(n245), .Z(n310) );
    VMW_AND4 U124 ( .A(In2[31]), .B(In2[30]), .C(In2[29]), .D(In2[28]), .Z(
        n317) );
    VMW_AND2 U63 ( .A(DataIn[15]), .B(ScanEnable), .Z(ScanOut[15]) );
    VMW_AND2 U78 ( .A(DataIn[0]), .B(ScanEnable), .Z(ScanOut[0]) );
    VMW_AOI211 U86 ( .A(n248), .B(In2[3]), .C(n261), .D(n245), .Z(n260) );
    VMW_AOI211 U103 ( .A(n248), .B(In2[17]), .C(n295), .D(n245), .Z(n294) );
    VMW_INV U188 ( .A(n286), .Z(n344) );
    VMW_AND4 U118 ( .A(In2[11]), .B(In2[10]), .C(In2[9]), .D(In2[8]), .Z(n326)
         );
    VMW_AO22 U151 ( .A(\Out[22] ), .B(n322), .C(n323), .D(In1[22]), .Z(n283)
         );
    VMW_INV U176 ( .A(n262), .Z(n333) );
    VMW_INV U193 ( .A(n296), .Z(n348) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \ScanLink0[13] , \Level4Out0[18] , \ScanLink0[20] , \ScanLink1[19] , 
        \Level1Out1[7] , \Level1Out2[23] , \Level1Out2[10] , \Level1Out6[21] , 
        \Level2Out0[0] , \Level1Out2[4] , \ScanLink4[22] , \ScanLink4[11] , 
        \Level1Out6[12] , \Level1Load7[0] , \Level1Out7[9] , \Level4Out4[30] , 
        \Level4Out4[29] , \Level4Out4[6] , \ScanLink5[31] , \ScanLink5[28] , 
        \Level1Out7[18] , \Level2Out6[20] , \Level2Out6[13] , \Level2Out2[22] , 
        \ScanLink0[30] , \ScanLink1[23] , \ScanLink1[10] , \Level1Out3[30] , 
        \ScanLink4[3] , \ScanLink7[0] , \Level1Out3[29] , \Level1Out3[20] , 
        \ScanLink5[21] , \ScanLink5[12] , \Level2Out2[11] , \ScanLink7[9] , 
        \Level1Out7[22] , \Level1Out7[11] , \Level2Out6[30] , \Level2Out6[29] , 
        \Level2Out2[18] , \Level1Out3[13] , \ScanLink1[7] , \ScanLink2[4] , 
        \Level1Out2[19] , \ScanLink0[29] , \ScanLink4[18] , \Level1Out4[3] , 
        \Level1Out7[0] , \Level4Out0[22] , \Level4Out0[11] , \Level4Out4[20] , 
        \Level4Out4[13] , \Level1Out6[31] , \Level1Out6[28] , \Level2Out0[9] , 
        \Level2Out6[7] , \ScanLink7[4] , \Level2Out2[26] , \Level2Out2[15] , 
        \ScanLink4[7] , \ScanLink0[17] , \ScanEnable[0] , \ScanLink2[9] , 
        \ScanLink4[26] , \ScanLink4[15] , \Level2Out6[24] , \Level2Out6[17] , 
        \Level4Out4[2] , \Level1Out6[25] , \Level1Out1[3] , \Level1Out2[0] , 
        \Level1Out6[16] , \Level2Out0[4] , \Level1Out2[27] , \Level1Out2[14] , 
        \ScanLink0[24] , \Level1Load2[0] , \Level1Out2[9] , \Level1Out4[7] , 
        \Level1Out7[4] , \Level2Out6[3] , \Level4Out4[24] , \Level4Out0[26] , 
        \Level4Out4[17] , \ScanLink1[27] , \ScanLink1[14] , \ScanLink1[3] , 
        \Level4Load0[0] , \Level4Out0[15] , \ScanLink2[0] , \Level1Out3[24] , 
        \ScanLink1[25] , \ScanLink1[16] , \Level1Out3[17] , \ScanLink5[25] , 
        \ScanLink5[16] , \Level1Out7[26] , \Level1Out7[15] , \ScanLink1[1] , 
        \ScanLink2[2] , \Level1Out1[8] , \Level1Out3[26] , \Level1Out3[15] , 
        \ScanLink5[27] , \ScanLink5[14] , \Level1Out7[24] , \Level1Out7[17] , 
        \Level1Out4[5] , \Level1Out7[6] , \Level4Out4[26] , \Level2Out6[1] , 
        \Level4Out4[15] , \Level4Out0[24] , \Level4Out4[9] , \Level1Out1[1] , 
        \ScanLink4[24] , \ScanLink4[17] , \Level4Out0[17] , \Level2Out6[8] , 
        \Level4Out4[0] , \Level1Out6[27] , \Level2Out0[6] , \Level1Out2[25] , 
        \Level1Out2[2] , \Level1Out6[14] , \Level1Out2[16] , \ScanLink0[15] , 
        \ScanLink0[26] , \Level2Out2[24] , \ScanLink0[18] , \ScanLink1[8] , 
        \ScanLink4[5] , \ScanLink7[6] , \Level2Out2[17] , \Level1Out2[31] , 
        \Level1Out2[28] , \Level2Out6[26] , \Level2Out6[15] , \Level4Out0[20] , 
        \ScanLink4[30] , \Level1Out4[1] , \Level4Out0[13] , \Level1Out7[2] , 
        \ScanLink4[29] , \Level2Out6[5] , \Level4Out4[22] , \ScanLink1[31] , 
        \ScanLink1[28] , \ScanLink1[21] , \ScanLink1[12] , \ScanLink1[5] , 
        \Level1Out3[22] , \ScanLink5[23] , \ScanLink5[10] , \Level1Out6[19] , 
        \Level4Out4[11] , \Level1Out7[20] , \Level2Out6[18] , \Level1Out7[13] , 
        \Level1Out3[11] , \ScanLink4[8] , \Level2Out2[30] , \Level2Out2[29] , 
        \ScanLink2[6] , \ScanLink5[19] , \Level1Out7[30] , \Level2Out6[22] , 
        \Level1Out7[29] , \Level2Load4[0] , \Level2Out6[11] , \Level1Out3[18] , 
        \ScanLink7[2] , \Level2Out2[20] , \Level2Out2[13] , \ScanLink0[11] , 
        \ScanLink4[1] , \ScanLink0[22] , \Level4Out0[30] , \Level4Out0[29] , 
        \Level1Out0[27] , \Level1Out0[14] , \Level1Out0[8] , \Level1Out1[5] , 
        \Level1Out2[21] , \Level1Out2[12] , \Level1Out2[6] , \Level1Out6[23] , 
        \Level1Out6[10] , \Level2Out0[2] , \ScanLink2[24] , \ScanLink4[20] , 
        \ScanLink4[13] , \Level4Out4[18] , \Level4Out4[4] , \Level1Out4[8] , 
        \ScanLink2[17] , \Level4Out0[4] , \Level2Out4[2] , \Level1Out5[5] , 
        \Level1Out4[25] , \Level1Out4[16] , \Level1Out6[6] , \ScanLink6[26] , 
        \ScanLink8[9] , \ScanLink0[1] , \ScanLink6[15] , \Level2Out4[17] , 
        \ScanLink3[2] , \Level2Out4[24] , \Level2Load0[0] , \ScanLink0[8] , 
        \ScanLink5[5] , \ScanLink6[6] , \ScanLink8[22] , \Level2Out0[15] , 
        \ScanLink8[11] , \Level2Out0[26] , \ScanLink7[25] , \ScanLink7[16] , 
        \Level1Out1[24] , \Level1Out1[17] , \Level1Out5[26] , \Level1Out5[15] , 
        \ScanLink8[18] , \ScanLink3[27] , \Level1Out0[1] , \ScanLink3[14] , 
        \Level1Out3[2] , \Level1Out1[30] , \Level1Out1[29] , \ScanLink8[26] , 
        \ScanLink8[0] , \Level2Out2[5] , \Level2Out0[11] , \ScanLink3[19] , 
        \ScanLink8[15] , \Level2Out0[22] , \ScanLink0[5] , \ScanLink3[6] , 
        \ScanLink5[8] , \ScanLink7[31] , \ScanLink7[28] , \Level2Out4[13] , 
        \Level1Out5[18] , \Level2Out4[20] , \ScanLink6[22] , \ScanLink6[11] , 
        \Level1Out0[23] , \Level1Out0[10] , \Level1Out4[21] , \Level1Out4[12] , 
        \Level1Out6[2] , \Level2Out4[6] , \Level1Out0[19] , \Level1Out0[5] , 
        \ScanLink2[20] , \Level1Out5[1] , \Level4Out0[0] , \ScanLink2[13] , 
        \Level2Out2[8] , \Level1Out4[31] , \Level1Out4[28] , \ScanLink6[18] , 
        \ScanLink8[4] , \ScanLink2[30] , \ScanLink2[29] , \Level1Out3[6] , 
        \Level4Out0[9] , \Level1Out5[8] , \Level2Out2[1] , \ScanLink3[23] , 
        \ScanLink3[10] , \Level1Out1[20] , \Level1Out1[13] , \Level1Out5[11] , 
        \Level2Out0[18] , \Level2Out4[30] , \Level2Out4[29] , \ScanLink3[21] , 
        \ScanLink5[1] , \Level1Out5[22] , \ScanLink6[2] , \ScanLink7[21] , 
        \ScanLink7[12] , \Level1Out1[22] , \Level1Out1[11] , \ScanLink3[12] , 
        \Level2Out0[30] , \Level2Out0[29] , \Level1Out4[19] , \ScanLink5[3] , 
        \Level1Out5[20] , \Level1Out5[13] , \ScanLink6[0] , \Level2Out4[18] , 
        \ScanLink7[23] , \ScanLink7[10] , \Level4Load4[0] , \Level1Out0[31] , 
        \Level1Out0[7] , \ScanLink2[18] , \Level1Out3[4] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink8[6] , \Level2Out2[3] , \Level1Out0[28] , 
        \ScanLink6[20] , \Level1Load6[0] , \Level1Out6[9] , \Level1Out4[10] , 
        \ScanLink6[13] , \Level1Out0[21] , \Level1Out0[12] , \Level1Out4[23] , 
        \Level2Out4[4] , \Level1Out5[3] , \Level1Out1[18] , \ScanLink2[22] , 
        \Level1Out6[0] , \ScanLink2[11] , \Level4Out0[2] , \ScanLink8[24] , 
        \Level2Out0[13] , \Level2Out0[20] , \ScanLink8[17] , \Level1Out0[3] , 
        \ScanLink0[7] , \ScanLink3[31] , \ScanLink3[28] , \Level1Out5[30] , 
        \Level1Out5[29] , \ScanLink6[9] , \ScanLink7[19] , \Level2Out4[11] , 
        \ScanLink3[4] , \Level2Out4[22] , \Level2Out4[9] , \Level1Out1[26] , 
        \Level1Out1[15] , \ScanLink3[9] , \Level1Out3[0] , \ScanLink5[7] , 
        \ScanLink8[2] , \Level2Out2[7] , \Level1Out5[17] , \ScanLink6[4] , 
        \ScanLink7[27] , \ScanLink7[14] , \Level1Out5[24] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink3[25] , \ScanLink3[16] , \ScanLink0[3] , 
        \ScanLink3[0] , \Level2Out4[26] , \Level2Out4[15] , \Level1Out0[25] , 
        \Level1Out0[16] , \ScanLink2[26] , \ScanLink8[20] , \ScanLink8[13] , 
        \Level2Out0[17] , \Level2Out0[24] , \Level4Out0[6] , \ScanLink2[15] , 
        \Level1Load3[0] , \Level1Out3[9] , \Level1Out6[4] , \Level2Out4[0] , 
        \Level1Out4[27] , \Level1Out4[14] , \Level1Out5[7] , \ScanLink6[24] , 
        \ScanLink6[17] , \Level1Out0[2] , \Level1Out3[1] , \ScanLink3[24] , 
        \ScanLink3[8] , \ScanLink8[3] , \Level2Out2[6] , \Level2Out4[8] , 
        \ScanLink5[6] , \Level1Out5[25] , \Level1Out5[16] , \ScanLink6[5] , 
        \ScanLink7[26] , \ScanLink7[15] , \ScanLink3[17] , \ScanLink0[2] , 
        \Level1Out1[27] , \Level1Out1[14] , \ScanLink8[31] , \ScanLink8[28] , 
        \Level2Out4[14] , \ScanLink3[1] , \ScanLink8[21] , \Level2Out0[16] , 
        \Level2Out4[27] , \ScanLink8[12] , \Level2Out0[25] , \Level1Out0[24] , 
        \Level1Out0[17] , \Level2Out4[1] , \Level1Out5[6] , \Level1Out6[5] , 
        \ScanLink2[27] , \ScanLink2[14] , \Level4Out0[7] , \Level1Out3[8] , 
        \ScanLink6[25] , \Level1Out1[23] , \Level1Out1[10] , \Level1Out4[26] , 
        \Level1Out4[15] , \ScanLink6[16] , \Level2Out0[31] , \Level2Out0[28] , 
        \Level2Load6[0] , \ScanLink3[20] , \ScanLink3[13] , \ScanLink5[2] , 
        \Level1Out5[21] , \Level1Out5[12] , \ScanLink6[1] , \ScanLink7[22] , 
        \ScanLink7[11] , \Level2Out4[19] , \Level1Out0[30] , \Level1Out0[29] , 
        \Level1Out4[18] , \ScanLink6[31] , \ScanLink6[28] , \ScanLink8[7] , 
        \Level1Out0[6] , \Level1Out6[8] , \ScanLink2[19] , \Level1Out3[5] , 
        \Level1Out4[22] , \Level1Out4[11] , \Level2Out2[2] , \ScanLink6[21] , 
        \ScanLink6[12] , \Level1Out0[20] , \Level1Out0[13] , \ScanLink2[23] , 
        \Level4Out0[3] , \ScanLink2[10] , \Level2Out4[5] , \Level1Out5[2] , 
        \Level1Out6[1] , \ScanLink3[30] , \ScanLink3[29] , \ScanLink0[6] , 
        \Level1Out1[19] , \ScanLink8[25] , \ScanLink8[16] , \Level2Out0[12] , 
        \ScanLink3[5] , \Level1Out5[31] , \Level2Out0[21] , \Level1Out5[28] , 
        \Level2Out4[23] , \Level2Out4[10] , \ScanLink6[8] , \ScanLink7[18] , 
        \ScanLink3[18] , \ScanLink0[4] , \Level1Out1[31] , \Level1Out1[28] , 
        \ScanLink8[27] , \Level2Out0[10] , \ScanLink8[14] , \Level2Out0[23] , 
        \Level2Out4[12] , \ScanLink3[7] , \Level1Out5[19] , \Level2Out4[21] , 
        \Level1Out4[20] , \Level1Out4[13] , \ScanLink5[9] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink6[23] , \Level1Out0[22] , \Level1Out0[11] , 
        \ScanLink2[21] , \ScanLink6[10] , \ScanLink2[12] , \Level2Out2[9] , 
        \Level4Out0[1] , \Level2Out4[7] , \Level1Out5[0] , \Level1Out6[3] , 
        \Level1Out0[18] , \Level1Out4[30] , \Level1Out4[29] , \ScanLink6[19] , 
        \ScanLink8[5] , \Level1Load5[0] , \Level1Out5[9] , \Level1Out0[4] , 
        \Level1Out3[7] , \Level1Out1[12] , \ScanLink2[31] , \ScanLink2[28] , 
        \Level2Out2[0] , \Level4Out0[8] , \Level1Out1[21] , \Level2Out0[19] , 
        \ScanLink3[22] , \ScanLink3[11] , \Level1Load0[0] , \Level1Out0[26] , 
        \Level1Out0[15] , \ScanLink5[0] , \ScanLink6[3] , \ScanLink7[20] , 
        \Level1Out5[23] , \Level1Out5[10] , \ScanLink7[13] , \Level2Out4[31] , 
        \Level2Out4[28] , \Level2Out4[3] , \Level1Out5[4] , \Level1Out6[7] , 
        \Level4Out0[5] , \Level1Out0[9] , \ScanLink2[25] , \ScanLink2[16] , 
        \ScanLink6[27] , \ScanLink6[14] , \ScanLink8[8] , \ScanLink0[0] , 
        \ScanLink3[3] , \Level1Out4[24] , \Level1Out4[17] , \Level2Out4[16] , 
        \Level2Out4[25] , \ScanLink8[23] , \ScanLink8[10] , \Level2Out0[14] , 
        \Level2Out0[27] , \ScanLink0[9] , \Level1Out5[14] , \ScanLink3[26] , 
        \ScanLink5[4] , \Level1Out5[27] , \ScanLink6[7] , \ScanLink7[24] , 
        \ScanLink7[17] , \Level1Out0[0] , \Level1Out1[25] , \Level1Out1[16] , 
        \ScanLink3[15] , \ScanLink8[19] , \ScanLink0[19] , \Level1Out3[3] , 
        \ScanLink8[1] , \Level2Out2[4] , \Level4Out0[21] , \Level1Out2[30] , 
        \Level4Out0[12] , \Level1Out2[29] , \ScanLink4[31] , \ScanLink4[28] , 
        \Level1Out6[18] , \Level1Out7[3] , \Level1Out4[0] , \Level4Out4[23] , 
        \ScanLink1[20] , \ScanLink1[13] , \ScanLink2[7] , \ScanLink5[22] , 
        \ScanLink5[11] , \Level1Out7[21] , \Level2Out6[4] , \Level4Out4[10] , 
        \Level1Out7[12] , \Level2Out6[19] , \ScanLink1[4] , \Level1Out3[23] , 
        \ScanLink4[9] , \Level1Out3[19] , \Level1Out3[10] , \ScanLink5[18] , 
        \Level2Out2[31] , \Level2Out2[28] , \Level1Out7[31] , \Level1Out7[28] , 
        \Level2Out6[23] , \Level2Out6[10] , \Level2Out2[21] , \ScanLink4[0] , 
        \ScanLink1[30] , \ScanLink7[3] , \Level2Out2[12] , \ScanLink1[29] , 
        \Level1Out2[20] , \Level1Out2[13] , \ScanLink0[10] , \ScanLink0[23] , 
        \Level4Out0[31] , \Level4Out0[28] , \ScanLink1[24] , \ScanLink1[17] , 
        \ScanLink1[0] , \Level1Out1[4] , \ScanLink4[21] , \ScanLink4[12] , 
        \Level4Out4[19] , \Level1Load4[0] , \Level4Out4[5] , \Level1Out4[9] , 
        \Level1Out6[22] , \Level2Out0[3] , \Level1Out2[7] , \Level1Out6[11] , 
        \Level1Out3[27] , \Level1Out3[14] , \ScanLink2[3] , \Level1Out4[4] , 
        \ScanLink5[26] , \ScanLink5[15] , \Level1Out7[25] , \Level1Out7[16] , 
        \Level1Out7[7] , \Level4Out4[27] , \Level2Out6[0] , \Level4Out4[8] , 
        \Level1Load1[0] , \Level1Out1[9] , \Level4Out4[14] , \Level4Out0[25] , 
        \Level4Out0[16] , \ScanLink0[14] , \Level1Out1[0] , \Level1Out2[3] , 
        \Level1Out6[26] , \Level2Out0[7] , \Level1Out6[15] , \ScanLink4[25] , 
        \ScanLink4[16] , \Level4Out4[1] , \Level2Out6[9] , \ScanLink0[27] , 
        \ScanLink1[9] , \Level1Out2[24] , \Level1Out2[17] , \ScanLink4[4] , 
        \ScanLink7[7] , \Level2Out2[25] , \Level2Out2[16] , \ScanLink2[8] , 
        \Level2Out6[27] , \Level2Out6[14] , \ScanLink4[6] , \Level2Out2[27] , 
        \Level1Out1[2] , \Level1Out6[24] , \ScanLink7[5] , \Level2Out0[5] , 
        \Level2Out2[14] , \Level2Out6[25] , \Level2Out6[16] , \Level1Out2[1] , 
        \Level1Out6[17] , \ScanLink4[27] , \ScanLink4[14] , \Level4Out4[3] , 
        \ScanLink0[16] , \ScanLink0[25] , \Level1Out2[26] , \Level1Out2[15] , 
        \Level1Out2[8] , \Level1Out4[6] , \Level1Out7[5] , \Level4Out4[25] , 
        \Level2Out6[2] , \Level4Out4[16] , \Level4Out0[27] , \Level4Out0[14] , 
        \ScanLink0[12] , \ScanLink1[26] , \ScanLink1[15] , \ScanLink2[1] , 
        \Level1Out3[25] , \Level1Out3[16] , \ScanLink1[2] , \Level1Out2[22] , 
        \ScanLink5[24] , \ScanLink5[17] , \Level1Out7[27] , \Level1Out7[14] , 
        \Level2Load2[0] , \Level1Out2[11] , \Level4Out0[19] , \ScanLink0[21] , 
        \Level1Out1[6] , \Level1Out2[5] , \ScanLink4[23] , \ScanLink4[10] , 
        \Level4Out4[7] , \Level4Out4[31] , \Level4Out4[28] , \Level1Out6[20] , 
        \Level1Out7[8] , \Level2Out0[1] , \Level1Out6[13] , \Level1Out3[31] , 
        \Level1Out3[28] , \ScanLink5[30] , \ScanLink5[29] , \Level1Out7[19] , 
        \Level2Out6[21] , \Level2Out2[23] , \Level2Out6[12] , \Level2Out2[10] , 
        \ScanLink4[2] , \ScanLink7[1] , \ScanLink0[31] , \ScanLink0[28] , 
        \ScanLink1[22] , \ScanLink1[18] , \ScanLink1[11] , \ScanLink1[6] , 
        \ScanLink5[20] , \ScanLink5[13] , \Level1Out7[23] , \Level1Out7[10] , 
        \Level2Out6[31] , \Level2Out6[28] , \ScanLink2[5] , \Level1Out3[21] , 
        \Level1Out3[12] , \ScanLink7[8] , \Level2Out2[19] , \Level1Out2[18] , 
        \Level4Out0[23] , \Level4Out0[10] , \ScanLink4[19] , \Level1Out4[2] , 
        \Level1Out6[30] , \Level1Out6[29] , \Level2Out0[8] , \Level1Out7[1] , 
        \Level4Out4[21] , \Level2Out6[6] , \Level4Out4[12] ;
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanOut({\ScanLink2[31] , 
        \ScanLink2[30] , \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , 
        \ScanLink2[26] , \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , 
        \ScanLink2[22] , \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , 
        \ScanLink2[18] , \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , 
        \ScanLink2[14] , \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , 
        \ScanLink2[10] , \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , 
        \ScanLink2[6] , \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , 
        \ScanLink2[2] , \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load1[0] ), .Out({
        \Level1Out1[31] , \Level1Out1[30] , \Level1Out1[29] , \Level1Out1[28] , 
        \Level1Out1[27] , \Level1Out1[26] , \Level1Out1[25] , \Level1Out1[24] , 
        \Level1Out1[23] , \Level1Out1[22] , \Level1Out1[21] , \Level1Out1[20] , 
        \Level1Out1[19] , \Level1Out1[18] , \Level1Out1[17] , \Level1Out1[16] , 
        \Level1Out1[15] , \Level1Out1[14] , \Level1Out1[13] , \Level1Out1[12] , 
        \Level1Out1[11] , \Level1Out1[10] , \Level1Out1[9] , \Level1Out1[8] , 
        \Level1Out1[7] , \Level1Out1[6] , \Level1Out1[5] , \Level1Out1[4] , 
        \Level1Out1[3] , \Level1Out1[2] , \Level1Out1[1] , \Level1Out1[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanOut({\ScanLink1[31] , 
        \ScanLink1[30] , \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , 
        \ScanLink1[26] , \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , 
        \ScanLink1[22] , \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , 
        \ScanLink1[18] , \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , 
        \ScanLink1[14] , \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , 
        \ScanLink1[10] , \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , 
        \ScanLink1[6] , \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , 
        \ScanLink1[2] , \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load0[0] ), .Out({
        \Level1Out0[31] , \Level1Out0[30] , \Level1Out0[29] , \Level1Out0[28] , 
        \Level1Out0[27] , \Level1Out0[26] , \Level1Out0[25] , \Level1Out0[24] , 
        \Level1Out0[23] , \Level1Out0[22] , \Level1Out0[21] , \Level1Out0[20] , 
        \Level1Out0[19] , \Level1Out0[18] , \Level1Out0[17] , \Level1Out0[16] , 
        \Level1Out0[15] , \Level1Out0[14] , \Level1Out0[13] , \Level1Out0[12] , 
        \Level1Out0[11] , \Level1Out0[10] , \Level1Out0[9] , \Level1Out0[8] , 
        \Level1Out0[7] , \Level1Out0[6] , \Level1Out0[5] , \Level1Out0[4] , 
        \Level1Out0[3] , \Level1Out0[2] , \Level1Out0[1] , \Level1Out0[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_6 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink6[31] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , 
        \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , 
        \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , 
        \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , 
        \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , 
        \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanOut({\ScanLink7[31] , 
        \ScanLink7[30] , \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , 
        \ScanLink7[26] , \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , 
        \ScanLink7[22] , \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , 
        \ScanLink7[18] , \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , 
        \ScanLink7[14] , \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , 
        \ScanLink7[10] , \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , 
        \ScanLink7[6] , \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , 
        \ScanLink7[2] , \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load6[0] ), .Out({
        \Level1Out6[31] , \Level1Out6[30] , \Level1Out6[29] , \Level1Out6[28] , 
        \Level1Out6[27] , \Level1Out6[26] , \Level1Out6[25] , \Level1Out6[24] , 
        \Level1Out6[23] , \Level1Out6[22] , \Level1Out6[21] , \Level1Out6[20] , 
        \Level1Out6[19] , \Level1Out6[18] , \Level1Out6[17] , \Level1Out6[16] , 
        \Level1Out6[15] , \Level1Out6[14] , \Level1Out6[13] , \Level1Out6[12] , 
        \Level1Out6[11] , \Level1Out6[10] , \Level1Out6[9] , \Level1Out6[8] , 
        \Level1Out6[7] , \Level1Out6[6] , \Level1Out6[5] , \Level1Out6[4] , 
        \Level1Out6[3] , \Level1Out6[2] , \Level1Out6[1] , \Level1Out6[0] })
         );
    Merge_Node_DWIDTH32 U_Merge_Node_0_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load0[0] ), .Out({\Level2Out0[31] , \Level2Out0[30] , 
        \Level2Out0[29] , \Level2Out0[28] , \Level2Out0[27] , \Level2Out0[26] , 
        \Level2Out0[25] , \Level2Out0[24] , \Level2Out0[23] , \Level2Out0[22] , 
        \Level2Out0[21] , \Level2Out0[20] , \Level2Out0[19] , \Level2Out0[18] , 
        \Level2Out0[17] , \Level2Out0[16] , \Level2Out0[15] , \Level2Out0[14] , 
        \Level2Out0[13] , \Level2Out0[12] , \Level2Out0[11] , \Level2Out0[10] , 
        \Level2Out0[9] , \Level2Out0[8] , \Level2Out0[7] , \Level2Out0[6] , 
        \Level2Out0[5] , \Level2Out0[4] , \Level2Out0[3] , \Level2Out0[2] , 
        \Level2Out0[1] , \Level2Out0[0] }), .In1({\Level1Out0[31] , 
        \Level1Out0[30] , \Level1Out0[29] , \Level1Out0[28] , \Level1Out0[27] , 
        \Level1Out0[26] , \Level1Out0[25] , \Level1Out0[24] , \Level1Out0[23] , 
        \Level1Out0[22] , \Level1Out0[21] , \Level1Out0[20] , \Level1Out0[19] , 
        \Level1Out0[18] , \Level1Out0[17] , \Level1Out0[16] , \Level1Out0[15] , 
        \Level1Out0[14] , \Level1Out0[13] , \Level1Out0[12] , \Level1Out0[11] , 
        \Level1Out0[10] , \Level1Out0[9] , \Level1Out0[8] , \Level1Out0[7] , 
        \Level1Out0[6] , \Level1Out0[5] , \Level1Out0[4] , \Level1Out0[3] , 
        \Level1Out0[2] , \Level1Out0[1] , \Level1Out0[0] }), .In2({
        \Level1Out1[31] , \Level1Out1[30] , \Level1Out1[29] , \Level1Out1[28] , 
        \Level1Out1[27] , \Level1Out1[26] , \Level1Out1[25] , \Level1Out1[24] , 
        \Level1Out1[23] , \Level1Out1[22] , \Level1Out1[21] , \Level1Out1[20] , 
        \Level1Out1[19] , \Level1Out1[18] , \Level1Out1[17] , \Level1Out1[16] , 
        \Level1Out1[15] , \Level1Out1[14] , \Level1Out1[13] , \Level1Out1[12] , 
        \Level1Out1[11] , \Level1Out1[10] , \Level1Out1[9] , \Level1Out1[8] , 
        \Level1Out1[7] , \Level1Out1[6] , \Level1Out1[5] , \Level1Out1[4] , 
        \Level1Out1[3] , \Level1Out1[2] , \Level1Out1[1] , \Level1Out1[0] }), 
        .Read1(\Level1Load0[0] ), .Read2(\Level1Load1[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_4_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load4[0] ), .Out({\Level4Out4[31] , \Level4Out4[30] , 
        \Level4Out4[29] , \Level4Out4[28] , \Level4Out4[27] , \Level4Out4[26] , 
        \Level4Out4[25] , \Level4Out4[24] , \Level4Out4[23] , \Level4Out4[22] , 
        \Level4Out4[21] , \Level4Out4[20] , \Level4Out4[19] , \Level4Out4[18] , 
        \Level4Out4[17] , \Level4Out4[16] , \Level4Out4[15] , \Level4Out4[14] , 
        \Level4Out4[13] , \Level4Out4[12] , \Level4Out4[11] , \Level4Out4[10] , 
        \Level4Out4[9] , \Level4Out4[8] , \Level4Out4[7] , \Level4Out4[6] , 
        \Level4Out4[5] , \Level4Out4[4] , \Level4Out4[3] , \Level4Out4[2] , 
        \Level4Out4[1] , \Level4Out4[0] }), .In1({\Level2Out4[31] , 
        \Level2Out4[30] , \Level2Out4[29] , \Level2Out4[28] , \Level2Out4[27] , 
        \Level2Out4[26] , \Level2Out4[25] , \Level2Out4[24] , \Level2Out4[23] , 
        \Level2Out4[22] , \Level2Out4[21] , \Level2Out4[20] , \Level2Out4[19] , 
        \Level2Out4[18] , \Level2Out4[17] , \Level2Out4[16] , \Level2Out4[15] , 
        \Level2Out4[14] , \Level2Out4[13] , \Level2Out4[12] , \Level2Out4[11] , 
        \Level2Out4[10] , \Level2Out4[9] , \Level2Out4[8] , \Level2Out4[7] , 
        \Level2Out4[6] , \Level2Out4[5] , \Level2Out4[4] , \Level2Out4[3] , 
        \Level2Out4[2] , \Level2Out4[1] , \Level2Out4[0] }), .In2({
        \Level2Out6[31] , \Level2Out6[30] , \Level2Out6[29] , \Level2Out6[28] , 
        \Level2Out6[27] , \Level2Out6[26] , \Level2Out6[25] , \Level2Out6[24] , 
        \Level2Out6[23] , \Level2Out6[22] , \Level2Out6[21] , \Level2Out6[20] , 
        \Level2Out6[19] , \Level2Out6[18] , \Level2Out6[17] , \Level2Out6[16] , 
        \Level2Out6[15] , \Level2Out6[14] , \Level2Out6[13] , \Level2Out6[12] , 
        \Level2Out6[11] , \Level2Out6[10] , \Level2Out6[9] , \Level2Out6[8] , 
        \Level2Out6[7] , \Level2Out6[6] , \Level2Out6[5] , \Level2Out6[4] , 
        \Level2Out6[3] , \Level2Out6[2] , \Level2Out6[1] , \Level2Out6[0] }), 
        .Read1(\Level2Load4[0] ), .Read2(\Level2Load6[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_7 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink7[31] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , 
        \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , 
        \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , 
        \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , 
        \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , 
        \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanOut({\ScanLink8[31] , 
        \ScanLink8[30] , \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , 
        \ScanLink8[26] , \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , 
        \ScanLink8[22] , \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , 
        \ScanLink8[18] , \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , 
        \ScanLink8[14] , \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , 
        \ScanLink8[10] , \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , 
        \ScanLink8[6] , \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , 
        \ScanLink8[2] , \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load7[0] ), .Out({
        \Level1Out7[31] , \Level1Out7[30] , \Level1Out7[29] , \Level1Out7[28] , 
        \Level1Out7[27] , \Level1Out7[26] , \Level1Out7[25] , \Level1Out7[24] , 
        \Level1Out7[23] , \Level1Out7[22] , \Level1Out7[21] , \Level1Out7[20] , 
        \Level1Out7[19] , \Level1Out7[18] , \Level1Out7[17] , \Level1Out7[16] , 
        \Level1Out7[15] , \Level1Out7[14] , \Level1Out7[13] , \Level1Out7[12] , 
        \Level1Out7[11] , \Level1Out7[10] , \Level1Out7[9] , \Level1Out7[8] , 
        \Level1Out7[7] , \Level1Out7[6] , \Level1Out7[5] , \Level1Out7[4] , 
        \Level1Out7[3] , \Level1Out7[2] , \Level1Out7[1] , \Level1Out7[0] })
         );
    Merge_Node_DWIDTH32 U_Merge_Node_0_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load0[0] ), .Out({\Level4Out0[31] , \Level4Out0[30] , 
        \Level4Out0[29] , \Level4Out0[28] , \Level4Out0[27] , \Level4Out0[26] , 
        \Level4Out0[25] , \Level4Out0[24] , \Level4Out0[23] , \Level4Out0[22] , 
        \Level4Out0[21] , \Level4Out0[20] , \Level4Out0[19] , \Level4Out0[18] , 
        \Level4Out0[17] , \Level4Out0[16] , \Level4Out0[15] , \Level4Out0[14] , 
        \Level4Out0[13] , \Level4Out0[12] , \Level4Out0[11] , \Level4Out0[10] , 
        \Level4Out0[9] , \Level4Out0[8] , \Level4Out0[7] , \Level4Out0[6] , 
        \Level4Out0[5] , \Level4Out0[4] , \Level4Out0[3] , \Level4Out0[2] , 
        \Level4Out0[1] , \Level4Out0[0] }), .In1({\Level2Out0[31] , 
        \Level2Out0[30] , \Level2Out0[29] , \Level2Out0[28] , \Level2Out0[27] , 
        \Level2Out0[26] , \Level2Out0[25] , \Level2Out0[24] , \Level2Out0[23] , 
        \Level2Out0[22] , \Level2Out0[21] , \Level2Out0[20] , \Level2Out0[19] , 
        \Level2Out0[18] , \Level2Out0[17] , \Level2Out0[16] , \Level2Out0[15] , 
        \Level2Out0[14] , \Level2Out0[13] , \Level2Out0[12] , \Level2Out0[11] , 
        \Level2Out0[10] , \Level2Out0[9] , \Level2Out0[8] , \Level2Out0[7] , 
        \Level2Out0[6] , \Level2Out0[5] , \Level2Out0[4] , \Level2Out0[3] , 
        \Level2Out0[2] , \Level2Out0[1] , \Level2Out0[0] }), .In2({
        \Level2Out2[31] , \Level2Out2[30] , \Level2Out2[29] , \Level2Out2[28] , 
        \Level2Out2[27] , \Level2Out2[26] , \Level2Out2[25] , \Level2Out2[24] , 
        \Level2Out2[23] , \Level2Out2[22] , \Level2Out2[21] , \Level2Out2[20] , 
        \Level2Out2[19] , \Level2Out2[18] , \Level2Out2[17] , \Level2Out2[16] , 
        \Level2Out2[15] , \Level2Out2[14] , \Level2Out2[13] , \Level2Out2[12] , 
        \Level2Out2[11] , \Level2Out2[10] , \Level2Out2[9] , \Level2Out2[8] , 
        \Level2Out2[7] , \Level2Out2[6] , \Level2Out2[5] , \Level2Out2[4] , 
        \Level2Out2[3] , \Level2Out2[2] , \Level2Out2[1] , \Level2Out2[0] }), 
        .Read1(\Level2Load0[0] ), .Read2(\Level2Load2[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_2 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanOut({\ScanLink3[31] , 
        \ScanLink3[30] , \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , 
        \ScanLink3[26] , \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , 
        \ScanLink3[22] , \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , 
        \ScanLink3[18] , \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , 
        \ScanLink3[14] , \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , 
        \ScanLink3[10] , \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , 
        \ScanLink3[6] , \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , 
        \ScanLink3[2] , \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load2[0] ), .Out({
        \Level1Out2[31] , \Level1Out2[30] , \Level1Out2[29] , \Level1Out2[28] , 
        \Level1Out2[27] , \Level1Out2[26] , \Level1Out2[25] , \Level1Out2[24] , 
        \Level1Out2[23] , \Level1Out2[22] , \Level1Out2[21] , \Level1Out2[20] , 
        \Level1Out2[19] , \Level1Out2[18] , \Level1Out2[17] , \Level1Out2[16] , 
        \Level1Out2[15] , \Level1Out2[14] , \Level1Out2[13] , \Level1Out2[12] , 
        \Level1Out2[11] , \Level1Out2[10] , \Level1Out2[9] , \Level1Out2[8] , 
        \Level1Out2[7] , \Level1Out2[6] , \Level1Out2[5] , \Level1Out2[4] , 
        \Level1Out2[3] , \Level1Out2[2] , \Level1Out2[1] , \Level1Out2[0] })
         );
    Merge_Node_DWIDTH32 U_Merge_Node_4_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load4[0] ), .Out({\Level2Out4[31] , \Level2Out4[30] , 
        \Level2Out4[29] , \Level2Out4[28] , \Level2Out4[27] , \Level2Out4[26] , 
        \Level2Out4[25] , \Level2Out4[24] , \Level2Out4[23] , \Level2Out4[22] , 
        \Level2Out4[21] , \Level2Out4[20] , \Level2Out4[19] , \Level2Out4[18] , 
        \Level2Out4[17] , \Level2Out4[16] , \Level2Out4[15] , \Level2Out4[14] , 
        \Level2Out4[13] , \Level2Out4[12] , \Level2Out4[11] , \Level2Out4[10] , 
        \Level2Out4[9] , \Level2Out4[8] , \Level2Out4[7] , \Level2Out4[6] , 
        \Level2Out4[5] , \Level2Out4[4] , \Level2Out4[3] , \Level2Out4[2] , 
        \Level2Out4[1] , \Level2Out4[0] }), .In1({\Level1Out4[31] , 
        \Level1Out4[30] , \Level1Out4[29] , \Level1Out4[28] , \Level1Out4[27] , 
        \Level1Out4[26] , \Level1Out4[25] , \Level1Out4[24] , \Level1Out4[23] , 
        \Level1Out4[22] , \Level1Out4[21] , \Level1Out4[20] , \Level1Out4[19] , 
        \Level1Out4[18] , \Level1Out4[17] , \Level1Out4[16] , \Level1Out4[15] , 
        \Level1Out4[14] , \Level1Out4[13] , \Level1Out4[12] , \Level1Out4[11] , 
        \Level1Out4[10] , \Level1Out4[9] , \Level1Out4[8] , \Level1Out4[7] , 
        \Level1Out4[6] , \Level1Out4[5] , \Level1Out4[4] , \Level1Out4[3] , 
        \Level1Out4[2] , \Level1Out4[1] , \Level1Out4[0] }), .In2({
        \Level1Out5[31] , \Level1Out5[30] , \Level1Out5[29] , \Level1Out5[28] , 
        \Level1Out5[27] , \Level1Out5[26] , \Level1Out5[25] , \Level1Out5[24] , 
        \Level1Out5[23] , \Level1Out5[22] , \Level1Out5[21] , \Level1Out5[20] , 
        \Level1Out5[19] , \Level1Out5[18] , \Level1Out5[17] , \Level1Out5[16] , 
        \Level1Out5[15] , \Level1Out5[14] , \Level1Out5[13] , \Level1Out5[12] , 
        \Level1Out5[11] , \Level1Out5[10] , \Level1Out5[9] , \Level1Out5[8] , 
        \Level1Out5[7] , \Level1Out5[6] , \Level1Out5[5] , \Level1Out5[4] , 
        \Level1Out5[3] , \Level1Out5[2] , \Level1Out5[1] , \Level1Out5[0] }), 
        .Read1(\Level1Load4[0] ), .Read2(\Level1Load5[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_3 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanOut({\ScanLink4[31] , 
        \ScanLink4[30] , \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , 
        \ScanLink4[26] , \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , 
        \ScanLink4[22] , \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , 
        \ScanLink4[18] , \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , 
        \ScanLink4[14] , \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , 
        \ScanLink4[10] , \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , 
        \ScanLink4[6] , \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , 
        \ScanLink4[2] , \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load3[0] ), .Out({
        \Level1Out3[31] , \Level1Out3[30] , \Level1Out3[29] , \Level1Out3[28] , 
        \Level1Out3[27] , \Level1Out3[26] , \Level1Out3[25] , \Level1Out3[24] , 
        \Level1Out3[23] , \Level1Out3[22] , \Level1Out3[21] , \Level1Out3[20] , 
        \Level1Out3[19] , \Level1Out3[18] , \Level1Out3[17] , \Level1Out3[16] , 
        \Level1Out3[15] , \Level1Out3[14] , \Level1Out3[13] , \Level1Out3[12] , 
        \Level1Out3[11] , \Level1Out3[10] , \Level1Out3[9] , \Level1Out3[8] , 
        \Level1Out3[7] , \Level1Out3[6] , \Level1Out3[5] , \Level1Out3[4] , 
        \Level1Out3[3] , \Level1Out3[2] , \Level1Out3[1] , \Level1Out3[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_4 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink4[31] , \ScanLink4[30] , 
        \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , 
        \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , 
        \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , 
        \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , 
        \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , 
        \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanOut({\ScanLink5[31] , 
        \ScanLink5[30] , \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , 
        \ScanLink5[26] , \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , 
        \ScanLink5[22] , \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , 
        \ScanLink5[18] , \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , 
        \ScanLink5[14] , \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , 
        \ScanLink5[10] , \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , 
        \ScanLink5[6] , \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , 
        \ScanLink5[2] , \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load4[0] ), .Out({
        \Level1Out4[31] , \Level1Out4[30] , \Level1Out4[29] , \Level1Out4[28] , 
        \Level1Out4[27] , \Level1Out4[26] , \Level1Out4[25] , \Level1Out4[24] , 
        \Level1Out4[23] , \Level1Out4[22] , \Level1Out4[21] , \Level1Out4[20] , 
        \Level1Out4[19] , \Level1Out4[18] , \Level1Out4[17] , \Level1Out4[16] , 
        \Level1Out4[15] , \Level1Out4[14] , \Level1Out4[13] , \Level1Out4[12] , 
        \Level1Out4[11] , \Level1Out4[10] , \Level1Out4[9] , \Level1Out4[8] , 
        \Level1Out4[7] , \Level1Out4[6] , \Level1Out4[5] , \Level1Out4[4] , 
        \Level1Out4[3] , \Level1Out4[2] , \Level1Out4[1] , \Level1Out4[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_5 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink5[31] , \ScanLink5[30] , 
        \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , 
        \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , 
        \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , 
        \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , 
        \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , 
        \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanOut({\ScanLink6[31] , 
        \ScanLink6[30] , \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , 
        \ScanLink6[26] , \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , 
        \ScanLink6[22] , \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , 
        \ScanLink6[18] , \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , 
        \ScanLink6[14] , \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , 
        \ScanLink6[10] , \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , 
        \ScanLink6[6] , \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , 
        \ScanLink6[2] , \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load5[0] ), .Out({
        \Level1Out5[31] , \Level1Out5[30] , \Level1Out5[29] , \Level1Out5[28] , 
        \Level1Out5[27] , \Level1Out5[26] , \Level1Out5[25] , \Level1Out5[24] , 
        \Level1Out5[23] , \Level1Out5[22] , \Level1Out5[21] , \Level1Out5[20] , 
        \Level1Out5[19] , \Level1Out5[18] , \Level1Out5[17] , \Level1Out5[16] , 
        \Level1Out5[15] , \Level1Out5[14] , \Level1Out5[13] , \Level1Out5[12] , 
        \Level1Out5[11] , \Level1Out5[10] , \Level1Out5[9] , \Level1Out5[8] , 
        \Level1Out5[7] , \Level1Out5[6] , \Level1Out5[5] , \Level1Out5[4] , 
        \Level1Out5[3] , \Level1Out5[2] , \Level1Out5[1] , \Level1Out5[0] })
         );
    Merge_Node_DWIDTH32 U_Merge_Node_6_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load6[0] ), .Out({\Level2Out6[31] , \Level2Out6[30] , 
        \Level2Out6[29] , \Level2Out6[28] , \Level2Out6[27] , \Level2Out6[26] , 
        \Level2Out6[25] , \Level2Out6[24] , \Level2Out6[23] , \Level2Out6[22] , 
        \Level2Out6[21] , \Level2Out6[20] , \Level2Out6[19] , \Level2Out6[18] , 
        \Level2Out6[17] , \Level2Out6[16] , \Level2Out6[15] , \Level2Out6[14] , 
        \Level2Out6[13] , \Level2Out6[12] , \Level2Out6[11] , \Level2Out6[10] , 
        \Level2Out6[9] , \Level2Out6[8] , \Level2Out6[7] , \Level2Out6[6] , 
        \Level2Out6[5] , \Level2Out6[4] , \Level2Out6[3] , \Level2Out6[2] , 
        \Level2Out6[1] , \Level2Out6[0] }), .In1({\Level1Out6[31] , 
        \Level1Out6[30] , \Level1Out6[29] , \Level1Out6[28] , \Level1Out6[27] , 
        \Level1Out6[26] , \Level1Out6[25] , \Level1Out6[24] , \Level1Out6[23] , 
        \Level1Out6[22] , \Level1Out6[21] , \Level1Out6[20] , \Level1Out6[19] , 
        \Level1Out6[18] , \Level1Out6[17] , \Level1Out6[16] , \Level1Out6[15] , 
        \Level1Out6[14] , \Level1Out6[13] , \Level1Out6[12] , \Level1Out6[11] , 
        \Level1Out6[10] , \Level1Out6[9] , \Level1Out6[8] , \Level1Out6[7] , 
        \Level1Out6[6] , \Level1Out6[5] , \Level1Out6[4] , \Level1Out6[3] , 
        \Level1Out6[2] , \Level1Out6[1] , \Level1Out6[0] }), .In2({
        \Level1Out7[31] , \Level1Out7[30] , \Level1Out7[29] , \Level1Out7[28] , 
        \Level1Out7[27] , \Level1Out7[26] , \Level1Out7[25] , \Level1Out7[24] , 
        \Level1Out7[23] , \Level1Out7[22] , \Level1Out7[21] , \Level1Out7[20] , 
        \Level1Out7[19] , \Level1Out7[18] , \Level1Out7[17] , \Level1Out7[16] , 
        \Level1Out7[15] , \Level1Out7[14] , \Level1Out7[13] , \Level1Out7[12] , 
        \Level1Out7[11] , \Level1Out7[10] , \Level1Out7[9] , \Level1Out7[8] , 
        \Level1Out7[7] , \Level1Out7[6] , \Level1Out7[5] , \Level1Out7[4] , 
        \Level1Out7[3] , \Level1Out7[2] , \Level1Out7[1] , \Level1Out7[0] }), 
        .Read1(\Level1Load6[0] ), .Read2(\Level1Load7[0] ) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Top_Node ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink8[31] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , 
        \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , 
        \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , 
        \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , 
        \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , 
        \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanOut({\ScanLink0[31] , 
        \ScanLink0[30] , \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , 
        \ScanLink0[26] , \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , 
        \ScanLink0[22] , \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , 
        \ScanLink0[18] , \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , 
        \ScanLink0[14] , \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , 
        \ScanLink0[10] , \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , 
        \ScanLink0[6] , \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , 
        \ScanLink0[2] , \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(
        \ScanEnable[0] ), .ScanId(1'b0), .Id(1'b1), .In1({\Level4Out0[31] , 
        \Level4Out0[30] , \Level4Out0[29] , \Level4Out0[28] , \Level4Out0[27] , 
        \Level4Out0[26] , \Level4Out0[25] , \Level4Out0[24] , \Level4Out0[23] , 
        \Level4Out0[22] , \Level4Out0[21] , \Level4Out0[20] , \Level4Out0[19] , 
        \Level4Out0[18] , \Level4Out0[17] , \Level4Out0[16] , \Level4Out0[15] , 
        \Level4Out0[14] , \Level4Out0[13] , \Level4Out0[12] , \Level4Out0[11] , 
        \Level4Out0[10] , \Level4Out0[9] , \Level4Out0[8] , \Level4Out0[7] , 
        \Level4Out0[6] , \Level4Out0[5] , \Level4Out0[4] , \Level4Out0[3] , 
        \Level4Out0[2] , \Level4Out0[1] , \Level4Out0[0] }), .In2({
        \Level4Out4[31] , \Level4Out4[30] , \Level4Out4[29] , \Level4Out4[28] , 
        \Level4Out4[27] , \Level4Out4[26] , \Level4Out4[25] , \Level4Out4[24] , 
        \Level4Out4[23] , \Level4Out4[22] , \Level4Out4[21] , \Level4Out4[20] , 
        \Level4Out4[19] , \Level4Out4[18] , \Level4Out4[17] , \Level4Out4[16] , 
        \Level4Out4[15] , \Level4Out4[14] , \Level4Out4[13] , \Level4Out4[12] , 
        \Level4Out4[11] , \Level4Out4[10] , \Level4Out4[9] , \Level4Out4[8] , 
        \Level4Out4[7] , \Level4Out4[6] , \Level4Out4[5] , \Level4Out4[4] , 
        \Level4Out4[3] , \Level4Out4[2] , \Level4Out4[1] , \Level4Out4[0] }), 
        .Read1(\Level4Load0[0] ), .Read2(\Level4Load4[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load2[0] ), .Out({\Level2Out2[31] , \Level2Out2[30] , 
        \Level2Out2[29] , \Level2Out2[28] , \Level2Out2[27] , \Level2Out2[26] , 
        \Level2Out2[25] , \Level2Out2[24] , \Level2Out2[23] , \Level2Out2[22] , 
        \Level2Out2[21] , \Level2Out2[20] , \Level2Out2[19] , \Level2Out2[18] , 
        \Level2Out2[17] , \Level2Out2[16] , \Level2Out2[15] , \Level2Out2[14] , 
        \Level2Out2[13] , \Level2Out2[12] , \Level2Out2[11] , \Level2Out2[10] , 
        \Level2Out2[9] , \Level2Out2[8] , \Level2Out2[7] , \Level2Out2[6] , 
        \Level2Out2[5] , \Level2Out2[4] , \Level2Out2[3] , \Level2Out2[2] , 
        \Level2Out2[1] , \Level2Out2[0] }), .In1({\Level1Out2[31] , 
        \Level1Out2[30] , \Level1Out2[29] , \Level1Out2[28] , \Level1Out2[27] , 
        \Level1Out2[26] , \Level1Out2[25] , \Level1Out2[24] , \Level1Out2[23] , 
        \Level1Out2[22] , \Level1Out2[21] , \Level1Out2[20] , \Level1Out2[19] , 
        \Level1Out2[18] , \Level1Out2[17] , \Level1Out2[16] , \Level1Out2[15] , 
        \Level1Out2[14] , \Level1Out2[13] , \Level1Out2[12] , \Level1Out2[11] , 
        \Level1Out2[10] , \Level1Out2[9] , \Level1Out2[8] , \Level1Out2[7] , 
        \Level1Out2[6] , \Level1Out2[5] , \Level1Out2[4] , \Level1Out2[3] , 
        \Level1Out2[2] , \Level1Out2[1] , \Level1Out2[0] }), .In2({
        \Level1Out3[31] , \Level1Out3[30] , \Level1Out3[29] , \Level1Out3[28] , 
        \Level1Out3[27] , \Level1Out3[26] , \Level1Out3[25] , \Level1Out3[24] , 
        \Level1Out3[23] , \Level1Out3[22] , \Level1Out3[21] , \Level1Out3[20] , 
        \Level1Out3[19] , \Level1Out3[18] , \Level1Out3[17] , \Level1Out3[16] , 
        \Level1Out3[15] , \Level1Out3[14] , \Level1Out3[13] , \Level1Out3[12] , 
        \Level1Out3[11] , \Level1Out3[10] , \Level1Out3[9] , \Level1Out3[8] , 
        \Level1Out3[7] , \Level1Out3[6] , \Level1Out3[5] , \Level1Out3[4] , 
        \Level1Out3[3] , \Level1Out3[2] , \Level1Out3[1] , \Level1Out3[0] }), 
        .Read1(\Level1Load2[0] ), .Read2(\Level1Load3[0] ) );
endmodule

