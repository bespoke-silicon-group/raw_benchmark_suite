
module EdgeAux_DW01_add_16_0 ( A, B, CI, SUM, CO );
input  [15:0] A;
input  [15:0] B;
output [15:0] SUM;
input  CI;
output CO;
    wire \carry[15] , \carry[13] , \carry[9] , \carry[4] , \carry[6] , 
        \carry[2] , \carry[14] , \carry[11] , \carry[10] , \carry[12] , 
        \carry[8] , \carry[7] , \carry[3] , \carry[5] , \carry[1] , n1;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_8 ( .CI(\carry[8] ), .A(A[8]), .B(B[8]), .S(SUM[8]), .CO(
        \carry[9] ) );
    VMW_FADD U1_11 ( .CI(\carry[11] ), .A(A[11]), .B(B[11]), .S(SUM[11]), .CO(
        \carry[12] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]), .CO(
        \carry[8] ) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_9 ( .CI(\carry[9] ), .A(A[9]), .B(B[9]), .S(SUM[9]), .CO(
        \carry[10] ) );
    VMW_FADD U1_10 ( .CI(\carry[10] ), .A(A[10]), .B(B[10]), .S(SUM[10]), .CO(
        \carry[11] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
    VMW_FADD U1_12 ( .CI(\carry[12] ), .A(A[12]), .B(B[12]), .S(SUM[12]), .CO(
        \carry[13] ) );
    VMW_FADD U1_15 ( .CI(\carry[15] ), .A(A[15]), .B(B[15]), .S(SUM[15]) );
    VMW_FADD U1_14 ( .CI(\carry[14] ), .A(A[14]), .B(B[14]), .S(SUM[14]), .CO(
        \carry[15] ) );
    VMW_FADD U1_13 ( .CI(\carry[13] ), .A(A[13]), .B(B[13]), .S(SUM[13]), .CO(
        \carry[14] ) );
endmodule


module EdgeAux ( Eid, InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [7:0] Eid;
input  [7:0] WeightAddr;
input  [15:0] InEdge;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire \Weight[11] , \Weight[6] , \Weight[15] , \Weight[2] , \Weight[0] , 
        \Weight[9] , \Weight[13] , \Weight[4] , \Weight[12] , \Weight[5] , 
        \Weight[1] , \Weight[8] , \Weight[14] , \Weight[3] , \Weight[10] , 
        \Weight[7] , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
        n101, n102, n103;
    VMW_PULLDOWN U15 ( .Z(n103) );
    VMW_AO22 U16 ( .A(\Weight[9] ), .B(n76), .C(WeightData[9]), .D(n77), .Z(
        n93) );
    VMW_AO22 U17 ( .A(\Weight[8] ), .B(n76), .C(WeightData[8]), .D(n77), .Z(
        n94) );
    VMW_AO22 U18 ( .A(\Weight[7] ), .B(n76), .C(WeightData[7]), .D(n77), .Z(
        n95) );
    VMW_AO22 U19 ( .A(\Weight[6] ), .B(n76), .C(WeightData[6]), .D(n77), .Z(
        n96) );
    VMW_AO22 U20 ( .A(\Weight[5] ), .B(n76), .C(WeightData[5]), .D(n77), .Z(
        n97) );
    VMW_AO22 U21 ( .A(\Weight[4] ), .B(n76), .C(WeightData[4]), .D(n77), .Z(
        n98) );
    VMW_AO22 U22 ( .A(\Weight[3] ), .B(n76), .C(WeightData[3]), .D(n77), .Z(
        n99) );
    VMW_AO22 U23 ( .A(\Weight[2] ), .B(n76), .C(WeightData[2]), .D(n77), .Z(
        n100) );
    VMW_AO22 U24 ( .A(\Weight[1] ), .B(n76), .C(WeightData[1]), .D(n77), .Z(
        n101) );
    VMW_AO22 U25 ( .A(\Weight[15] ), .B(n76), .C(WeightData[15]), .D(n77), .Z(
        n87) );
    VMW_AO22 U26 ( .A(\Weight[14] ), .B(n76), .C(WeightData[14]), .D(n77), .Z(
        n88) );
    VMW_AO22 U27 ( .A(\Weight[13] ), .B(n76), .C(WeightData[13]), .D(n77), .Z(
        n89) );
    VMW_AO22 U28 ( .A(\Weight[12] ), .B(n76), .C(WeightData[12]), .D(n77), .Z(
        n90) );
    VMW_AO22 U29 ( .A(\Weight[11] ), .B(n76), .C(WeightData[11]), .D(n77), .Z(
        n91) );
    VMW_AO22 U30 ( .A(\Weight[10] ), .B(n76), .C(WeightData[10]), .D(n77), .Z(
        n92) );
    VMW_AO22 U31 ( .A(\Weight[0] ), .B(n76), .C(WeightData[0]), .D(n77), .Z(
        n102) );
    VMW_AND4 U32 ( .A(n79), .B(n80), .C(n81), .D(n82), .Z(n78) );
    VMW_AND5 U33 ( .A(n83), .B(n84), .C(n85), .D(n86), .E(n78), .Z(n77) );
    VMW_XNOR2 U34 ( .A(WeightAddr[0]), .B(Eid[0]), .Z(n82) );
    VMW_XNOR2 U35 ( .A(WeightAddr[1]), .B(Eid[1]), .Z(n81) );
    VMW_XNOR2 U36 ( .A(WeightAddr[4]), .B(Eid[4]), .Z(n80) );
    VMW_XNOR2 U37 ( .A(WeightAddr[5]), .B(Eid[5]), .Z(n79) );
    VMW_XNOR2 U38 ( .A(WeightAddr[6]), .B(Eid[6]), .Z(n86) );
    VMW_XNOR2 U39 ( .A(WeightAddr[7]), .B(Eid[7]), .Z(n85) );
    VMW_XNOR2 U40 ( .A(WeightAddr[3]), .B(Eid[3]), .Z(n84) );
    VMW_XNOR2 U41 ( .A(WeightAddr[2]), .B(Eid[2]), .Z(n83) );
    VMW_INV U42 ( .A(n77), .Z(n76) );
    VMW_FD \Weight_reg[15]  ( .D(n87), .CP(Clk), .Q(\Weight[15] ) );
    VMW_FD \Weight_reg[14]  ( .D(n88), .CP(Clk), .Q(\Weight[14] ) );
    VMW_FD \Weight_reg[13]  ( .D(n89), .CP(Clk), .Q(\Weight[13] ) );
    VMW_FD \Weight_reg[12]  ( .D(n90), .CP(Clk), .Q(\Weight[12] ) );
    VMW_FD \Weight_reg[11]  ( .D(n91), .CP(Clk), .Q(\Weight[11] ) );
    VMW_FD \Weight_reg[10]  ( .D(n92), .CP(Clk), .Q(\Weight[10] ) );
    VMW_FD \Weight_reg[9]  ( .D(n93), .CP(Clk), .Q(\Weight[9] ) );
    VMW_FD \Weight_reg[8]  ( .D(n94), .CP(Clk), .Q(\Weight[8] ) );
    VMW_FD \Weight_reg[7]  ( .D(n95), .CP(Clk), .Q(\Weight[7] ) );
    VMW_FD \Weight_reg[6]  ( .D(n96), .CP(Clk), .Q(\Weight[6] ) );
    VMW_FD \Weight_reg[5]  ( .D(n97), .CP(Clk), .Q(\Weight[5] ) );
    VMW_FD \Weight_reg[4]  ( .D(n98), .CP(Clk), .Q(\Weight[4] ) );
    VMW_FD \Weight_reg[3]  ( .D(n99), .CP(Clk), .Q(\Weight[3] ) );
    VMW_FD \Weight_reg[2]  ( .D(n100), .CP(Clk), .Q(\Weight[2] ) );
    VMW_FD \Weight_reg[1]  ( .D(n101), .CP(Clk), .Q(\Weight[1] ) );
    VMW_FD \Weight_reg[0]  ( .D(n102), .CP(Clk), .Q(\Weight[0] ) );
    EdgeAux_DW01_add_16_0 add_92 ( .A({\Weight[15] , \Weight[14] , 
        \Weight[13] , \Weight[12] , \Weight[11] , \Weight[10] , \Weight[9] , 
        \Weight[8] , \Weight[7] , \Weight[6] , \Weight[5] , \Weight[4] , 
        \Weight[3] , \Weight[2] , \Weight[1] , \Weight[0] }), .B(InEdge), .CI(
        n103), .SUM(OutEdge) );
endmodule


module NodeAux_INDEGREE2_SOURCE1_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE2_SOURCE1_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n85) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n85), .D(n82), .Z(n86) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n86), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n93) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n93), .D(n90), .Z(n94) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n94), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n96), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n102), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n112) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n112), .D(n110), .Z(n113) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n114), .C(n113), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n114) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE2_SOURCE1 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp180[1] , \temp180[8] , \OutEdge106[5] , \temp180[5] , 
        \OutEdge106[8] , \OutEdge106[1] , \path[2] , \path[0] , 
        \OutEdge106[3] , \temp180[7] , \OutEdge106[7] , \temp180[3] , 
        \OutEdge106[13] , \temp180[12] , \temp180[10] , \OutEdge106[11] , 
        \OutEdge106[15] , \temp180[14] , n84, \OutEdge106[14] , \temp180[15] , 
        \temp180[11] , \OutEdge106[10] , \OutEdge106[12] , \temp180[13] , 
        \OutEdge106[6] , \temp180[2] , \path[1] , n92, \OutEdge106[2] , 
        \temp180[6] , \temp180[4] , \OutEdge106[9] , \OutEdge106[0] , 
        \temp180[0] , \temp180[9] , \OutEdge106[4] , n367, n368, n369, n370, 
        n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
        n383, n384;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U55 ( .Z(n383) );
    VMW_PULLDOWN U56 ( .Z(n384) );
    VMW_AO22 U57 ( .A(n367), .B(\temp180[15] ), .C(InEdges[31]), .D(n368), .Z(
        \OutEdge106[15] ) );
    VMW_AO22 U58 ( .A(n367), .B(\temp180[14] ), .C(InEdges[30]), .D(n368), .Z(
        \OutEdge106[14] ) );
    VMW_AO22 U59 ( .A(n367), .B(\temp180[13] ), .C(InEdges[29]), .D(n368), .Z(
        \OutEdge106[13] ) );
    VMW_AO22 U60 ( .A(n367), .B(\temp180[12] ), .C(InEdges[28]), .D(n368), .Z(
        \OutEdge106[12] ) );
    VMW_AO22 U61 ( .A(n367), .B(\temp180[11] ), .C(InEdges[27]), .D(n368), .Z(
        \OutEdge106[11] ) );
    VMW_AO22 U62 ( .A(n367), .B(\temp180[10] ), .C(InEdges[26]), .D(n368), .Z(
        \OutEdge106[10] ) );
    VMW_AO22 U63 ( .A(n367), .B(\temp180[9] ), .C(InEdges[25]), .D(n368), .Z(
        \OutEdge106[9] ) );
    VMW_AO22 U64 ( .A(n367), .B(\temp180[8] ), .C(InEdges[24]), .D(n368), .Z(
        \OutEdge106[8] ) );
    VMW_AO22 U65 ( .A(n367), .B(\temp180[7] ), .C(InEdges[23]), .D(n368), .Z(
        \OutEdge106[7] ) );
    VMW_AO22 U66 ( .A(n367), .B(\temp180[6] ), .C(InEdges[22]), .D(n368), .Z(
        \OutEdge106[6] ) );
    VMW_AO22 U67 ( .A(n367), .B(\temp180[5] ), .C(InEdges[21]), .D(n368), .Z(
        \OutEdge106[5] ) );
    VMW_AO22 U68 ( .A(n367), .B(\temp180[4] ), .C(InEdges[20]), .D(n368), .Z(
        \OutEdge106[4] ) );
    VMW_AO22 U69 ( .A(n367), .B(\temp180[3] ), .C(InEdges[19]), .D(n368), .Z(
        \OutEdge106[3] ) );
    VMW_AO22 U70 ( .A(n367), .B(\temp180[2] ), .C(InEdges[18]), .D(n368), .Z(
        \OutEdge106[2] ) );
    VMW_AO22 U71 ( .A(n367), .B(\temp180[1] ), .C(InEdges[17]), .D(n368), .Z(
        \OutEdge106[1] ) );
    VMW_AO22 U72 ( .A(n367), .B(\temp180[0] ), .C(InEdges[16]), .D(n368), .Z(
        \OutEdge106[0] ) );
    VMW_AO22 U73 ( .A(Start), .B(\path[1] ), .C(n369), .D(n367), .Z(n382) );
    VMW_AO22 U74 ( .A(\path[2] ), .B(Start), .C(n369), .D(n367), .Z(n381) );
    VMW_OR2 U75 ( .A(n368), .B(n370), .Z(n380) );
    VMW_AO22 U76 ( .A(InEdges[9]), .B(n84), .C(OutEdge[9]), .D(n369), .Z(
        \temp180[9] ) );
    VMW_AO22 U77 ( .A(InEdges[8]), .B(n84), .C(OutEdge[8]), .D(n369), .Z(
        \temp180[8] ) );
    VMW_AO22 U78 ( .A(InEdges[7]), .B(n84), .C(OutEdge[7]), .D(n369), .Z(
        \temp180[7] ) );
    VMW_AO22 U79 ( .A(InEdges[6]), .B(n84), .C(OutEdge[6]), .D(n369), .Z(
        \temp180[6] ) );
    VMW_AO22 U80 ( .A(InEdges[5]), .B(n84), .C(OutEdge[5]), .D(n369), .Z(
        \temp180[5] ) );
    VMW_AO22 U81 ( .A(InEdges[4]), .B(n84), .C(OutEdge[4]), .D(n369), .Z(
        \temp180[4] ) );
    VMW_AO22 U82 ( .A(InEdges[3]), .B(n84), .C(OutEdge[3]), .D(n369), .Z(
        \temp180[3] ) );
    VMW_AO22 U83 ( .A(InEdges[2]), .B(n84), .C(OutEdge[2]), .D(n369), .Z(
        \temp180[2] ) );
    VMW_AO22 U84 ( .A(InEdges[1]), .B(n84), .C(OutEdge[1]), .D(n369), .Z(
        \temp180[1] ) );
    VMW_AO22 U85 ( .A(InEdges[15]), .B(n84), .C(OutEdge[15]), .D(n369), .Z(
        \temp180[15] ) );
    VMW_AO22 U86 ( .A(InEdges[14]), .B(n84), .C(OutEdge[14]), .D(n369), .Z(
        \temp180[14] ) );
    VMW_AO22 U87 ( .A(InEdges[13]), .B(n84), .C(OutEdge[13]), .D(n369), .Z(
        \temp180[13] ) );
    VMW_AO22 U88 ( .A(InEdges[12]), .B(n84), .C(OutEdge[12]), .D(n369), .Z(
        \temp180[12] ) );
    VMW_AO22 U89 ( .A(InEdges[11]), .B(n84), .C(OutEdge[11]), .D(n369), .Z(
        \temp180[11] ) );
    VMW_AO22 U90 ( .A(InEdges[10]), .B(n84), .C(OutEdge[10]), .D(n369), .Z(
        \temp180[10] ) );
    VMW_AO22 U91 ( .A(InEdges[0]), .B(n84), .C(OutEdge[0]), .D(n369), .Z(
        \temp180[0] ) );
    VMW_NOR2 U92 ( .A(Start), .B(n92), .Z(n367) );
    VMW_AND2 U93 ( .A(n92), .B(n371), .Z(n368) );
    VMW_AO22 U94 ( .A(n369), .B(n371), .C(\path[0] ), .D(Start), .Z(n370) );
    VMW_AND3 U95 ( .A(n373), .B(n374), .C(n375), .Z(n372) );
    VMW_AND4 U96 ( .A(n376), .B(n377), .C(n378), .D(n372), .Z(n379) );
    VMW_XNOR2 U97 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n374) );
    VMW_XNOR2 U98 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n373) );
    VMW_XNOR2 U99 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n375) );
    VMW_XNOR2 U100 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n377) );
    VMW_XNOR2 U101 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n376) );
    VMW_XNOR2 U102 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n378) );
    VMW_INV U103 ( .A(n84), .Z(n369) );
    VMW_INV U104 ( .A(Start), .Z(n371) );
    VMW_BUFIZ U105 ( .A(\path[1] ), .E(n379), .Z(\PathData[1] ) );
    VMW_BUFIZ U106 ( .A(\path[0] ), .E(n379), .Z(\PathData[0] ) );
    VMW_BUFIZ U107 ( .A(\path[2] ), .E(n379), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n380), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n381), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n382), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge106[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge106[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge106[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge106[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge106[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge106[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge106[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge106[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge106[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge106[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge106[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge106[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge106[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge106[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge106[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge106[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE2_SOURCE1_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n384), .TC(n384), .GE_GT(n84) );
    NodeAux_INDEGREE2_SOURCE1_DW01_cmp2_16_0 lte_55_1 ( .A({\temp180[15] , 
        \temp180[14] , \temp180[13] , \temp180[12] , \temp180[11] , 
        \temp180[10] , \temp180[9] , \temp180[8] , \temp180[7] , \temp180[6] , 
        \temp180[5] , \temp180[4] , \temp180[3] , \temp180[2] , \temp180[1] , 
        \temp180[0] }), .B(InEdges[31:16]), .LEQ(n383), .TC(n383), .GE_GT(n92)
         );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n85) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n85), .D(n82), .Z(n86) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n86), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n93) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n93), .D(n90), .Z(n94) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n94), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n96), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n102), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n112) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n112), .D(n110), .Z(n113) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n114), .C(n113), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n114) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE2_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp180[1] , \temp180[8] , \OutEdge106[5] , \temp180[5] , 
        \OutEdge106[8] , \OutEdge106[1] , \path[2] , \path[0] , 
        \OutEdge106[3] , \temp180[7] , \OutEdge106[7] , \temp180[3] , 
        \OutEdge106[13] , \temp180[12] , \temp180[10] , \OutEdge106[11] , 
        \OutEdge106[15] , \temp180[14] , n84, \OutEdge106[14] , \temp180[15] , 
        \temp180[11] , \OutEdge106[10] , \OutEdge106[12] , \temp180[13] , 
        \OutEdge106[6] , \temp180[2] , \path[1] , n92, \OutEdge106[2] , 
        \temp180[6] , \temp180[4] , \OutEdge106[9] , \OutEdge106[0] , 
        \temp180[0] , \temp180[9] , \OutEdge106[4] , n367, n368, n369, n370, 
        n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
        n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
        n395, n396, n397, n398, n399, n400;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U55 ( .Z(n399) );
    VMW_PULLDOWN U56 ( .Z(n400) );
    VMW_NOR2 U57 ( .A(Start), .B(n367), .Z(\OutEdge106[15] ) );
    VMW_NAND2 U58 ( .A(n368), .B(n369), .Z(\OutEdge106[14] ) );
    VMW_NAND2 U59 ( .A(n370), .B(n369), .Z(\OutEdge106[13] ) );
    VMW_NAND2 U60 ( .A(n371), .B(n369), .Z(\OutEdge106[12] ) );
    VMW_NAND2 U61 ( .A(n372), .B(n369), .Z(\OutEdge106[11] ) );
    VMW_NAND2 U62 ( .A(n373), .B(n369), .Z(\OutEdge106[10] ) );
    VMW_NAND2 U63 ( .A(n374), .B(n369), .Z(\OutEdge106[9] ) );
    VMW_NAND2 U64 ( .A(n375), .B(n369), .Z(\OutEdge106[8] ) );
    VMW_NAND2 U65 ( .A(n376), .B(n369), .Z(\OutEdge106[7] ) );
    VMW_NAND2 U66 ( .A(n377), .B(n369), .Z(\OutEdge106[6] ) );
    VMW_NAND2 U67 ( .A(n378), .B(n369), .Z(\OutEdge106[5] ) );
    VMW_NAND2 U68 ( .A(n379), .B(n369), .Z(\OutEdge106[4] ) );
    VMW_NAND2 U69 ( .A(n380), .B(n369), .Z(\OutEdge106[3] ) );
    VMW_NAND2 U70 ( .A(n381), .B(n369), .Z(\OutEdge106[2] ) );
    VMW_NAND2 U71 ( .A(n382), .B(n369), .Z(\OutEdge106[1] ) );
    VMW_NAND2 U72 ( .A(n383), .B(n369), .Z(\OutEdge106[0] ) );
    VMW_AO21 U73 ( .A(Start), .B(\path[1] ), .C(n384), .Z(n398) );
    VMW_AO21 U74 ( .A(\path[2] ), .B(Start), .C(n384), .Z(n397) );
    VMW_OR2 U75 ( .A(n386), .B(n92), .Z(n385) );
    VMW_AO22 U76 ( .A(OutEdge[15]), .B(n386), .C(InEdges[15]), .D(n84), .Z(
        \temp180[15] ) );
    VMW_OAI22 U77 ( .A(\path[0] ), .B(n369), .C(n385), .D(Start), .Z(n387) );
    VMW_MUX2I U78 ( .A(\temp180[15] ), .B(InEdges[31]), .S(n92), .Z(n367) );
    VMW_AND3 U79 ( .A(n389), .B(n390), .C(n391), .Z(n388) );
    VMW_NOR3 U80 ( .A(Start), .B(n84), .C(n92), .Z(n384) );
    VMW_AND4 U81 ( .A(n392), .B(n393), .C(n394), .D(n388), .Z(n395) );
    VMW_XNOR2 U82 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n390) );
    VMW_XNOR2 U83 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n389) );
    VMW_XNOR2 U84 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n391) );
    VMW_XNOR2 U85 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n393) );
    VMW_XNOR2 U86 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n392) );
    VMW_XNOR2 U87 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n394) );
    VMW_AO22 U88 ( .A(OutEdge[9]), .B(n386), .C(InEdges[9]), .D(n84), .Z(
        \temp180[9] ) );
    VMW_AO22 U89 ( .A(OutEdge[8]), .B(n386), .C(InEdges[8]), .D(n84), .Z(
        \temp180[8] ) );
    VMW_AO22 U90 ( .A(OutEdge[7]), .B(n386), .C(InEdges[7]), .D(n84), .Z(
        \temp180[7] ) );
    VMW_AO22 U91 ( .A(OutEdge[6]), .B(n386), .C(InEdges[6]), .D(n84), .Z(
        \temp180[6] ) );
    VMW_AO22 U92 ( .A(OutEdge[5]), .B(n386), .C(InEdges[5]), .D(n84), .Z(
        \temp180[5] ) );
    VMW_AO22 U93 ( .A(OutEdge[4]), .B(n386), .C(InEdges[4]), .D(n84), .Z(
        \temp180[4] ) );
    VMW_AO22 U94 ( .A(OutEdge[3]), .B(n386), .C(InEdges[3]), .D(n84), .Z(
        \temp180[3] ) );
    VMW_AO22 U95 ( .A(OutEdge[2]), .B(n386), .C(InEdges[2]), .D(n84), .Z(
        \temp180[2] ) );
    VMW_AO22 U96 ( .A(OutEdge[1]), .B(n386), .C(InEdges[1]), .D(n84), .Z(
        \temp180[1] ) );
    VMW_AO22 U97 ( .A(OutEdge[14]), .B(n386), .C(InEdges[14]), .D(n84), .Z(
        \temp180[14] ) );
    VMW_AO22 U98 ( .A(OutEdge[13]), .B(n386), .C(InEdges[13]), .D(n84), .Z(
        \temp180[13] ) );
    VMW_AO22 U99 ( .A(OutEdge[12]), .B(n386), .C(InEdges[12]), .D(n84), .Z(
        \temp180[12] ) );
    VMW_AO22 U100 ( .A(OutEdge[11]), .B(n386), .C(InEdges[11]), .D(n84), .Z(
        \temp180[11] ) );
    VMW_AO22 U101 ( .A(OutEdge[10]), .B(n386), .C(InEdges[10]), .D(n84), .Z(
        \temp180[10] ) );
    VMW_AO22 U102 ( .A(OutEdge[0]), .B(n386), .C(InEdges[0]), .D(n84), .Z(
        \temp180[0] ) );
    VMW_MUX2I U103 ( .A(\temp180[9] ), .B(InEdges[25]), .S(n92), .Z(n374) );
    VMW_MUX2I U104 ( .A(\temp180[8] ), .B(InEdges[24]), .S(n92), .Z(n375) );
    VMW_MUX2I U105 ( .A(\temp180[7] ), .B(InEdges[23]), .S(n92), .Z(n376) );
    VMW_MUX2I U106 ( .A(\temp180[6] ), .B(InEdges[22]), .S(n92), .Z(n377) );
    VMW_MUX2I U107 ( .A(\temp180[5] ), .B(InEdges[21]), .S(n92), .Z(n378) );
    VMW_MUX2I U108 ( .A(\temp180[4] ), .B(InEdges[20]), .S(n92), .Z(n379) );
    VMW_MUX2I U109 ( .A(\temp180[3] ), .B(InEdges[19]), .S(n92), .Z(n380) );
    VMW_MUX2I U110 ( .A(\temp180[2] ), .B(InEdges[18]), .S(n92), .Z(n381) );
    VMW_MUX2I U111 ( .A(\temp180[1] ), .B(InEdges[17]), .S(n92), .Z(n382) );
    VMW_MUX2I U112 ( .A(\temp180[14] ), .B(InEdges[30]), .S(n92), .Z(n368) );
    VMW_MUX2I U113 ( .A(\temp180[13] ), .B(InEdges[29]), .S(n92), .Z(n370) );
    VMW_MUX2I U114 ( .A(\temp180[12] ), .B(InEdges[28]), .S(n92), .Z(n371) );
    VMW_MUX2I U115 ( .A(\temp180[11] ), .B(InEdges[27]), .S(n92), .Z(n372) );
    VMW_MUX2I U116 ( .A(\temp180[10] ), .B(InEdges[26]), .S(n92), .Z(n373) );
    VMW_MUX2I U117 ( .A(\temp180[0] ), .B(InEdges[16]), .S(n92), .Z(n383) );
    VMW_INV U118 ( .A(n84), .Z(n386) );
    VMW_INV U119 ( .A(Start), .Z(n369) );
    VMW_INV U120 ( .A(n387), .Z(n396) );
    VMW_BUFIZ U121 ( .A(\path[1] ), .E(n395), .Z(\PathData[1] ) );
    VMW_BUFIZ U122 ( .A(\path[0] ), .E(n395), .Z(\PathData[0] ) );
    VMW_BUFIZ U123 ( .A(\path[2] ), .E(n395), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n396), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n397), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n398), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge106[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge106[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge106[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge106[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge106[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge106[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge106[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge106[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge106[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge106[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge106[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge106[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge106[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge106[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge106[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge106[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n400), .TC(n400), .GE_GT(n84) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 lte_55_1 ( .A({\temp180[15] , 
        \temp180[14] , \temp180[13] , \temp180[12] , \temp180[11] , 
        \temp180[10] , \temp180[9] , \temp180[8] , \temp180[7] , \temp180[6] , 
        \temp180[5] , \temp180[4] , \temp180[3] , \temp180[2] , \temp180[1] , 
        \temp180[0] }), .B(InEdges[31:16]), .LEQ(n399), .TC(n399), .GE_GT(n92)
         );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, 
        n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, n107, 
        n108, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n104), .B(B[12]), .Z(n103) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n96), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n104), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n103), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n104) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
        n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
        n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
        n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
        n163, n164;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n119), .B(B[2]), .Z(n118) );
    VMW_AO22 U5 ( .A(n121), .B(B[0]), .C(n122), .D(B[1]), .Z(n120) );
    VMW_OR2 U6 ( .A(B[2]), .B(n119), .Z(n123) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n122), .C(n123), .D(n120), .Z(n124) );
    VMW_NAND2 U8 ( .A(n126), .B(B[4]), .Z(n125) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n128), .C(n124), .D(n118), .Z(n127) );
    VMW_OR2 U10 ( .A(B[4]), .B(n126), .Z(n129) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n131), .C(n129), .D(n127), .Z(n130) );
    VMW_NAND2 U12 ( .A(n133), .B(B[6]), .Z(n132) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n135), .C(n130), .D(n125), .Z(n134) );
    VMW_OR2 U14 ( .A(B[6]), .B(n133), .Z(n136) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n138), .C(n136), .D(n134), .Z(n137) );
    VMW_NAND2 U16 ( .A(n140), .B(B[8]), .Z(n139) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n142), .C(n137), .D(n132), .Z(n141) );
    VMW_OR2 U18 ( .A(B[8]), .B(n140), .Z(n143) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n145), .C(n143), .D(n141), .Z(n144) );
    VMW_NAND2 U20 ( .A(n147), .B(B[10]), .Z(n146) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n149), .C(n144), .D(n139), .Z(n148) );
    VMW_NAND2 U22 ( .A(n149), .B(A[9]), .Z(n150) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n147), .C(n150), .D(n148), .Z(n151) );
    VMW_NAND2 U24 ( .A(n153), .B(B[12]), .Z(n152) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n155), .C(n151), .D(n146), .Z(n154) );
    VMW_NAND2 U26 ( .A(n155), .B(A[11]), .Z(n156) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n153), .C(n156), .D(n154), .Z(n157) );
    VMW_NAND2 U28 ( .A(n159), .B(B[14]), .Z(n158) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n161), .C(n157), .D(n152), .Z(n160) );
    VMW_NAND2 U30 ( .A(n161), .B(A[13]), .Z(n162) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n159), .C(n162), .D(n160), .Z(n163) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n164), .C(n163), .D(n158), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n153) );
    VMW_INV U34 ( .A(B[7]), .Z(n142) );
    VMW_INV U35 ( .A(A[7]), .Z(n145) );
    VMW_INV U36 ( .A(A[3]), .Z(n131) );
    VMW_INV U37 ( .A(B[3]), .Z(n128) );
    VMW_INV U38 ( .A(A[10]), .Z(n147) );
    VMW_INV U39 ( .A(B[9]), .Z(n149) );
    VMW_INV U40 ( .A(A[4]), .Z(n126) );
    VMW_INV U41 ( .A(A[8]), .Z(n140) );
    VMW_INV U42 ( .A(A[14]), .Z(n159) );
    VMW_INV U43 ( .A(B[11]), .Z(n155) );
    VMW_INV U44 ( .A(A[5]), .Z(n138) );
    VMW_INV U45 ( .A(B[5]), .Z(n135) );
    VMW_INV U46 ( .A(A[1]), .Z(n122) );
    VMW_INV U47 ( .A(B[15]), .Z(n164) );
    VMW_INV U48 ( .A(B[13]), .Z(n161) );
    VMW_INV U49 ( .A(A[6]), .Z(n133) );
    VMW_INV U50 ( .A(A[2]), .Z(n119) );
    VMW_INV U51 ( .A(A[0]), .Z(n121) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE3_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp284[0] , \OutEdge116[6] , \temp284[9] , \temp284[11] , 
        \temp190[2] , \OutEdge116[2] , \temp284[4] , \temp190[6] , 
        \temp284[15] , \path[2] , \OutEdge116[9] , \path[0] , \temp190[4] , 
        \OutEdge116[0] , \temp284[6] , \temp284[13] , \temp190[0] , 
        \temp284[2] , \OutEdge116[4] , \temp190[9] , \temp190[10] , 
        \OutEdge116[11] , \OutEdge116[15] , \temp190[14] , \OutEdge116[13] , 
        \temp190[12] , n94, \OutEdge116[12] , \temp190[13] , n86, 
        \OutEdge116[14] , \temp190[15] , \temp190[11] , \OutEdge116[10] , 
        \temp284[12] , \temp190[1] , \temp284[3] , \OutEdge116[5] , 
        \temp190[8] , \path[1] , \OutEdge116[8] , \temp190[5] , 
        \OutEdge116[1] , \temp284[7] , n102, \OutEdge116[3] , \temp284[5] , 
        \temp190[7] , \temp284[14] , \temp284[1] , \OutEdge116[7] , 
        \temp284[8] , \temp284[10] , \temp190[3] , n467, n468, n469, n470, 
        n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
        n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U64 ( .Z(n503) );
    VMW_PULLDOWN U65 ( .Z(n505) );
    VMW_PULLDOWN U66 ( .Z(n504) );
    VMW_AND2 U67 ( .A(n467), .B(n468), .Z(\OutEdge116[15] ) );
    VMW_OR2 U68 ( .A(n469), .B(Start), .Z(\OutEdge116[14] ) );
    VMW_OR2 U69 ( .A(n470), .B(Start), .Z(\OutEdge116[13] ) );
    VMW_OR2 U70 ( .A(n471), .B(Start), .Z(\OutEdge116[12] ) );
    VMW_OR2 U71 ( .A(n472), .B(Start), .Z(\OutEdge116[11] ) );
    VMW_OR2 U72 ( .A(n473), .B(Start), .Z(\OutEdge116[10] ) );
    VMW_OR2 U73 ( .A(n474), .B(Start), .Z(\OutEdge116[9] ) );
    VMW_OR2 U74 ( .A(n475), .B(Start), .Z(\OutEdge116[8] ) );
    VMW_OR2 U75 ( .A(n476), .B(Start), .Z(\OutEdge116[7] ) );
    VMW_OR2 U76 ( .A(n477), .B(Start), .Z(\OutEdge116[6] ) );
    VMW_OR2 U77 ( .A(n478), .B(Start), .Z(\OutEdge116[5] ) );
    VMW_OR2 U78 ( .A(n479), .B(Start), .Z(\OutEdge116[4] ) );
    VMW_OR2 U79 ( .A(n480), .B(Start), .Z(\OutEdge116[3] ) );
    VMW_OR2 U80 ( .A(n481), .B(Start), .Z(\OutEdge116[2] ) );
    VMW_OR2 U81 ( .A(n482), .B(Start), .Z(\OutEdge116[1] ) );
    VMW_OR2 U82 ( .A(n483), .B(Start), .Z(\OutEdge116[0] ) );
    VMW_OR2 U83 ( .A(n484), .B(n485), .Z(n502) );
    VMW_AO22 U84 ( .A(\path[2] ), .B(Start), .C(n486), .D(n485), .Z(n501) );
    VMW_AO22 U85 ( .A(\temp190[15] ), .B(n487), .C(InEdges[31]), .D(n94), .Z(
        \temp284[15] ) );
    VMW_AND3 U86 ( .A(n467), .B(n488), .C(n487), .Z(n485) );
    VMW_INV U87 ( .A(Start), .Z(n467) );
    VMW_AO22 U88 ( .A(n490), .B(n467), .C(n491), .D(Start), .Z(n489) );
    VMW_AO22 U89 ( .A(\temp284[15] ), .B(n486), .C(InEdges[47]), .D(n102), .Z(
        n468) );
    VMW_AND3 U90 ( .A(n493), .B(n494), .C(n495), .Z(n492) );
    VMW_INV U91 ( .A(n102), .Z(n486) );
    VMW_AND4 U92 ( .A(n496), .B(n497), .C(n498), .D(n492), .Z(n499) );
    VMW_XNOR2 U93 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n494) );
    VMW_XNOR2 U94 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n493) );
    VMW_XNOR2 U95 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n495) );
    VMW_XNOR2 U96 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n497) );
    VMW_XNOR2 U97 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n496) );
    VMW_XNOR2 U98 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n498) );
    VMW_AO22 U99 ( .A(InEdges[9]), .B(n86), .C(OutEdge[9]), .D(n488), .Z(
        \temp190[9] ) );
    VMW_AO22 U100 ( .A(\temp190[9] ), .B(n487), .C(InEdges[25]), .D(n94), .Z(
        \temp284[9] ) );
    VMW_AO22 U101 ( .A(InEdges[8]), .B(n86), .C(OutEdge[8]), .D(n488), .Z(
        \temp190[8] ) );
    VMW_AO22 U102 ( .A(\temp190[8] ), .B(n487), .C(InEdges[24]), .D(n94), .Z(
        \temp284[8] ) );
    VMW_AO22 U103 ( .A(InEdges[7]), .B(n86), .C(OutEdge[7]), .D(n488), .Z(
        \temp190[7] ) );
    VMW_AO22 U104 ( .A(\temp190[7] ), .B(n487), .C(InEdges[23]), .D(n94), .Z(
        \temp284[7] ) );
    VMW_AO22 U105 ( .A(InEdges[6]), .B(n86), .C(OutEdge[6]), .D(n488), .Z(
        \temp190[6] ) );
    VMW_AO22 U106 ( .A(\temp190[6] ), .B(n487), .C(InEdges[22]), .D(n94), .Z(
        \temp284[6] ) );
    VMW_AO22 U107 ( .A(InEdges[5]), .B(n86), .C(OutEdge[5]), .D(n488), .Z(
        \temp190[5] ) );
    VMW_AO22 U108 ( .A(\temp190[5] ), .B(n487), .C(InEdges[21]), .D(n94), .Z(
        \temp284[5] ) );
    VMW_AO22 U109 ( .A(InEdges[4]), .B(n86), .C(OutEdge[4]), .D(n488), .Z(
        \temp190[4] ) );
    VMW_AO22 U110 ( .A(\temp190[4] ), .B(n487), .C(InEdges[20]), .D(n94), .Z(
        \temp284[4] ) );
    VMW_AO22 U111 ( .A(InEdges[3]), .B(n86), .C(OutEdge[3]), .D(n488), .Z(
        \temp190[3] ) );
    VMW_AO22 U112 ( .A(\temp190[3] ), .B(n487), .C(InEdges[19]), .D(n94), .Z(
        \temp284[3] ) );
    VMW_AO22 U113 ( .A(InEdges[2]), .B(n86), .C(OutEdge[2]), .D(n488), .Z(
        \temp190[2] ) );
    VMW_AO22 U114 ( .A(\temp190[2] ), .B(n487), .C(InEdges[18]), .D(n94), .Z(
        \temp284[2] ) );
    VMW_AO22 U115 ( .A(InEdges[1]), .B(n86), .C(OutEdge[1]), .D(n488), .Z(
        \temp190[1] ) );
    VMW_AO22 U116 ( .A(\temp190[1] ), .B(n487), .C(InEdges[17]), .D(n94), .Z(
        \temp284[1] ) );
    VMW_AO22 U117 ( .A(InEdges[15]), .B(n86), .C(OutEdge[15]), .D(n488), .Z(
        \temp190[15] ) );
    VMW_AO22 U118 ( .A(InEdges[14]), .B(n86), .C(OutEdge[14]), .D(n488), .Z(
        \temp190[14] ) );
    VMW_AO22 U119 ( .A(\temp190[14] ), .B(n487), .C(InEdges[30]), .D(n94), .Z(
        \temp284[14] ) );
    VMW_AO22 U120 ( .A(InEdges[13]), .B(n86), .C(OutEdge[13]), .D(n488), .Z(
        \temp190[13] ) );
    VMW_AO22 U121 ( .A(\temp190[13] ), .B(n487), .C(InEdges[29]), .D(n94), .Z(
        \temp284[13] ) );
    VMW_AO22 U122 ( .A(InEdges[12]), .B(n86), .C(OutEdge[12]), .D(n488), .Z(
        \temp190[12] ) );
    VMW_AO22 U123 ( .A(\temp190[12] ), .B(n487), .C(InEdges[28]), .D(n94), .Z(
        \temp284[12] ) );
    VMW_AO22 U124 ( .A(InEdges[11]), .B(n86), .C(OutEdge[11]), .D(n488), .Z(
        \temp190[11] ) );
    VMW_AO22 U125 ( .A(\temp190[11] ), .B(n487), .C(InEdges[27]), .D(n94), .Z(
        \temp284[11] ) );
    VMW_AO22 U126 ( .A(InEdges[10]), .B(n86), .C(OutEdge[10]), .D(n488), .Z(
        \temp190[10] ) );
    VMW_AO22 U127 ( .A(\temp190[10] ), .B(n487), .C(InEdges[26]), .D(n94), .Z(
        \temp284[10] ) );
    VMW_AO22 U128 ( .A(InEdges[0]), .B(n86), .C(OutEdge[0]), .D(n488), .Z(
        \temp190[0] ) );
    VMW_AO22 U129 ( .A(\temp190[0] ), .B(n487), .C(InEdges[16]), .D(n94), .Z(
        \temp284[0] ) );
    VMW_AO22 U130 ( .A(\path[1] ), .B(Start), .C(n102), .D(n467), .Z(n484) );
    VMW_AO21 U131 ( .A(n487), .B(n86), .C(n102), .Z(n490) );
    VMW_AO22 U132 ( .A(\temp284[9] ), .B(n486), .C(InEdges[41]), .D(n102), .Z(
        n474) );
    VMW_AO22 U133 ( .A(\temp284[8] ), .B(n486), .C(InEdges[40]), .D(n102), .Z(
        n475) );
    VMW_AO22 U134 ( .A(\temp284[7] ), .B(n486), .C(InEdges[39]), .D(n102), .Z(
        n476) );
    VMW_AO22 U135 ( .A(\temp284[6] ), .B(n486), .C(InEdges[38]), .D(n102), .Z(
        n477) );
    VMW_AO22 U136 ( .A(\temp284[5] ), .B(n486), .C(InEdges[37]), .D(n102), .Z(
        n478) );
    VMW_AO22 U137 ( .A(\temp284[4] ), .B(n486), .C(InEdges[36]), .D(n102), .Z(
        n479) );
    VMW_AO22 U138 ( .A(\temp284[3] ), .B(n486), .C(InEdges[35]), .D(n102), .Z(
        n480) );
    VMW_AO22 U139 ( .A(\temp284[2] ), .B(n486), .C(InEdges[34]), .D(n102), .Z(
        n481) );
    VMW_AO22 U140 ( .A(\temp284[1] ), .B(n486), .C(InEdges[33]), .D(n102), .Z(
        n482) );
    VMW_AO22 U141 ( .A(\temp284[14] ), .B(n486), .C(InEdges[46]), .D(n102), 
        .Z(n469) );
    VMW_AO22 U142 ( .A(\temp284[13] ), .B(n486), .C(InEdges[45]), .D(n102), 
        .Z(n470) );
    VMW_AO22 U143 ( .A(\temp284[12] ), .B(n486), .C(InEdges[44]), .D(n102), 
        .Z(n471) );
    VMW_AO22 U144 ( .A(\temp284[11] ), .B(n486), .C(InEdges[43]), .D(n102), 
        .Z(n472) );
    VMW_AO22 U145 ( .A(\temp284[10] ), .B(n486), .C(InEdges[42]), .D(n102), 
        .Z(n473) );
    VMW_AO22 U146 ( .A(\temp284[0] ), .B(n486), .C(InEdges[32]), .D(n102), .Z(
        n483) );
    VMW_INV U147 ( .A(n86), .Z(n488) );
    VMW_INV U148 ( .A(n94), .Z(n487) );
    VMW_INV U149 ( .A(n489), .Z(n500) );
    VMW_INV U150 ( .A(\path[0] ), .Z(n491) );
    VMW_BUFIZ U151 ( .A(\path[1] ), .E(n499), .Z(\PathData[1] ) );
    VMW_BUFIZ U152 ( .A(\path[0] ), .E(n499), .Z(\PathData[0] ) );
    VMW_BUFIZ U153 ( .A(\path[2] ), .E(n499), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n500), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n501), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n502), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge116[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge116[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge116[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge116[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge116[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge116[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge116[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge116[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge116[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge116[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge116[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge116[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge116[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge116[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge116[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge116[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp190[15] , 
        \temp190[14] , \temp190[13] , \temp190[12] , \temp190[11] , 
        \temp190[10] , \temp190[9] , \temp190[8] , \temp190[7] , \temp190[6] , 
        \temp190[5] , \temp190[4] , \temp190[3] , \temp190[2] , \temp190[1] , 
        \temp190[0] }), .B(InEdges[31:16]), .LEQ(n505), .TC(n505), .GE_GT(n94)
         );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n504), .TC(n504), .GE_GT(n86) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 lte_55_2 ( .A({\temp284[15] , 
        \temp284[14] , \temp284[13] , \temp284[12] , \temp284[11] , 
        \temp284[10] , \temp284[9] , \temp284[8] , \temp284[7] , \temp284[6] , 
        \temp284[5] , \temp284[4] , \temp284[3] , \temp284[2] , \temp284[1] , 
        \temp284[0] }), .B(InEdges[47:32]), .LEQ(n503), .TC(n503), .GE_GT(n102
        ) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, 
        n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, 
        n108, n109, n110, n111, n113, n114, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n95), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n113), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n113), .B(A[13]), .Z(n114) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n114), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n113) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
        n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
        n164, n165;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n127), .B(B[4]), .Z(n126) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n129), .C(n125), .D(n119), .Z(n128) );
    VMW_OR2 U10 ( .A(B[4]), .B(n127), .Z(n130) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n132), .C(n130), .D(n128), .Z(n131) );
    VMW_NAND2 U12 ( .A(n134), .B(B[6]), .Z(n133) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n136), .C(n131), .D(n126), .Z(n135) );
    VMW_OR2 U14 ( .A(B[6]), .B(n134), .Z(n137) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n139), .C(n137), .D(n135), .Z(n138) );
    VMW_NAND2 U16 ( .A(n141), .B(B[8]), .Z(n140) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n143), .C(n138), .D(n133), .Z(n142) );
    VMW_OR2 U18 ( .A(B[8]), .B(n141), .Z(n144) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n146), .C(n144), .D(n142), .Z(n145) );
    VMW_NAND2 U20 ( .A(n148), .B(B[10]), .Z(n147) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n150), .C(n145), .D(n140), .Z(n149) );
    VMW_NAND2 U22 ( .A(n150), .B(A[9]), .Z(n151) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n148), .C(n151), .D(n149), .Z(n152) );
    VMW_NAND2 U24 ( .A(n154), .B(B[12]), .Z(n153) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n156), .C(n152), .D(n147), .Z(n155) );
    VMW_NAND2 U26 ( .A(n156), .B(A[11]), .Z(n157) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n154), .C(n157), .D(n155), .Z(n158) );
    VMW_NAND2 U28 ( .A(n160), .B(B[14]), .Z(n159) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n162), .C(n158), .D(n153), .Z(n161) );
    VMW_NAND2 U30 ( .A(n162), .B(A[13]), .Z(n163) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n160), .C(n163), .D(n161), .Z(n164) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n165), .C(n164), .D(n159), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n154) );
    VMW_INV U34 ( .A(B[7]), .Z(n143) );
    VMW_INV U35 ( .A(A[7]), .Z(n146) );
    VMW_INV U36 ( .A(A[3]), .Z(n132) );
    VMW_INV U37 ( .A(B[3]), .Z(n129) );
    VMW_INV U38 ( .A(A[10]), .Z(n148) );
    VMW_INV U39 ( .A(B[9]), .Z(n150) );
    VMW_INV U40 ( .A(A[4]), .Z(n127) );
    VMW_INV U41 ( .A(A[8]), .Z(n141) );
    VMW_INV U42 ( .A(A[14]), .Z(n160) );
    VMW_INV U43 ( .A(B[11]), .Z(n156) );
    VMW_INV U44 ( .A(A[5]), .Z(n139) );
    VMW_INV U45 ( .A(B[5]), .Z(n136) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n165) );
    VMW_INV U48 ( .A(B[13]), .Z(n162) );
    VMW_INV U49 ( .A(A[6]), .Z(n134) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
        n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
        n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
        n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
        n213, n214;
    VMW_OAI21 U3 ( .A(B[15]), .B(n166), .C(n167), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n169), .B(B[2]), .Z(n168) );
    VMW_AO22 U5 ( .A(n171), .B(B[0]), .C(n172), .D(B[1]), .Z(n170) );
    VMW_OR2 U6 ( .A(B[2]), .B(n169), .Z(n173) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n172), .C(n173), .D(n170), .Z(n174) );
    VMW_NAND2 U8 ( .A(n176), .B(B[4]), .Z(n175) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n178), .C(n174), .D(n168), .Z(n177) );
    VMW_OR2 U10 ( .A(B[4]), .B(n176), .Z(n179) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n181), .C(n179), .D(n177), .Z(n180) );
    VMW_NAND2 U12 ( .A(n183), .B(B[6]), .Z(n182) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n185), .C(n180), .D(n175), .Z(n184) );
    VMW_OR2 U14 ( .A(B[6]), .B(n183), .Z(n186) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n188), .C(n186), .D(n184), .Z(n187) );
    VMW_NAND2 U16 ( .A(n190), .B(B[8]), .Z(n189) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n192), .C(n187), .D(n182), .Z(n191) );
    VMW_OR2 U18 ( .A(B[8]), .B(n190), .Z(n193) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n195), .C(n193), .D(n191), .Z(n194) );
    VMW_NAND2 U20 ( .A(n197), .B(B[10]), .Z(n196) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n199), .C(n194), .D(n189), .Z(n198) );
    VMW_NAND2 U22 ( .A(n199), .B(A[9]), .Z(n200) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n197), .C(n200), .D(n198), .Z(n201) );
    VMW_NAND2 U24 ( .A(n203), .B(B[12]), .Z(n202) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n205), .C(n201), .D(n196), .Z(n204) );
    VMW_NAND2 U26 ( .A(n205), .B(A[11]), .Z(n206) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n203), .C(n206), .D(n204), .Z(n207) );
    VMW_NAND2 U28 ( .A(n209), .B(B[14]), .Z(n208) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n211), .C(n207), .D(n202), .Z(n210) );
    VMW_NAND2 U30 ( .A(n211), .B(A[13]), .Z(n212) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n209), .C(n212), .D(n210), .Z(n213) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n214), .C(n213), .D(n208), .Z(n167) );
    VMW_INV U33 ( .A(A[12]), .Z(n203) );
    VMW_INV U34 ( .A(B[7]), .Z(n192) );
    VMW_INV U35 ( .A(A[7]), .Z(n195) );
    VMW_INV U36 ( .A(A[3]), .Z(n181) );
    VMW_INV U37 ( .A(B[3]), .Z(n178) );
    VMW_INV U38 ( .A(A[10]), .Z(n197) );
    VMW_INV U39 ( .A(B[9]), .Z(n199) );
    VMW_INV U40 ( .A(A[4]), .Z(n176) );
    VMW_INV U41 ( .A(A[8]), .Z(n190) );
    VMW_INV U42 ( .A(A[14]), .Z(n209) );
    VMW_INV U43 ( .A(B[11]), .Z(n205) );
    VMW_INV U44 ( .A(A[5]), .Z(n188) );
    VMW_INV U45 ( .A(B[5]), .Z(n185) );
    VMW_INV U46 ( .A(A[1]), .Z(n172) );
    VMW_INV U47 ( .A(B[15]), .Z(n214) );
    VMW_INV U48 ( .A(B[13]), .Z(n211) );
    VMW_INV U49 ( .A(A[6]), .Z(n183) );
    VMW_INV U50 ( .A(A[2]), .Z(n169) );
    VMW_INV U51 ( .A(A[0]), .Z(n171) );
    VMW_INV U52 ( .A(A[15]), .Z(n166) );
endmodule


module NodeAux_INDEGREE4_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp200[0] , \temp384[15] , \OutEdge126[12] , \temp200[15] , 
        \temp200[9] , \temp384[6] , \temp294[3] , n112, \temp294[13] , 
        \temp384[11] , \temp200[4] , \temp294[7] , \temp384[2] , \path[2] , 
        \temp200[11] , \temp200[13] , \path[0] , \temp294[5] , \temp384[0] , 
        \temp384[13] , \temp200[6] , \temp384[9] , \OutEdge126[14] , 
        \temp294[11] , \temp384[4] , \temp294[1] , \OutEdge126[10] , 
        \temp294[15] , \temp200[2] , \temp294[8] , \OutEdge126[8] , 
        \OutEdge126[1] , \OutEdge126[5] , n96, \OutEdge126[7] , 
        \OutEdge126[3] , \OutEdge126[2] , \OutEdge126[6] , \OutEdge126[4] , 
        n104, \OutEdge126[9] , n88, \OutEdge126[0] , \temp384[5] , 
        \temp294[0] , \OutEdge126[11] , \temp294[14] , \temp200[3] , 
        \temp294[9] , \path[1] , \temp200[12] , \temp294[4] , \temp384[1] , 
        \temp384[12] , \temp384[8] , \temp200[7] , \OutEdge126[15] , 
        \temp294[10] , \temp294[12] , \temp384[10] , \temp200[5] , 
        \temp294[6] , \temp384[3] , \temp200[10] , \temp200[1] , \temp384[14] , 
        \OutEdge126[13] , \temp200[14] , \temp384[7] , \temp200[8] , 
        \temp294[2] , n567, n568, n569, n570, n571, n572, n573, n574, n575, 
        n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
        n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
        n600, n601, n602, n603, n604, n605, n606, n607, n608, n609;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U73 ( .Z(n606) );
    VMW_PULLDOWN U74 ( .Z(n607) );
    VMW_PULLDOWN U75 ( .Z(n608) );
    VMW_PULLDOWN U76 ( .Z(n609) );
    VMW_NOR2 U77 ( .A(Start), .B(n567), .Z(\OutEdge126[15] ) );
    VMW_NAND2 U78 ( .A(n568), .B(n569), .Z(\OutEdge126[14] ) );
    VMW_NAND2 U79 ( .A(n570), .B(n569), .Z(\OutEdge126[13] ) );
    VMW_NAND2 U80 ( .A(n571), .B(n569), .Z(\OutEdge126[12] ) );
    VMW_NAND2 U81 ( .A(n572), .B(n569), .Z(\OutEdge126[11] ) );
    VMW_NAND2 U82 ( .A(n573), .B(n569), .Z(\OutEdge126[10] ) );
    VMW_NAND2 U83 ( .A(n574), .B(n569), .Z(\OutEdge126[9] ) );
    VMW_NAND2 U84 ( .A(n575), .B(n569), .Z(\OutEdge126[8] ) );
    VMW_NAND2 U85 ( .A(n576), .B(n569), .Z(\OutEdge126[7] ) );
    VMW_NAND2 U86 ( .A(n577), .B(n569), .Z(\OutEdge126[6] ) );
    VMW_NAND2 U87 ( .A(n578), .B(n569), .Z(\OutEdge126[5] ) );
    VMW_NAND2 U88 ( .A(n579), .B(n569), .Z(\OutEdge126[4] ) );
    VMW_NAND2 U89 ( .A(n580), .B(n569), .Z(\OutEdge126[3] ) );
    VMW_NAND2 U90 ( .A(n581), .B(n569), .Z(\OutEdge126[2] ) );
    VMW_NAND2 U91 ( .A(n582), .B(n569), .Z(\OutEdge126[1] ) );
    VMW_NAND2 U92 ( .A(n583), .B(n569), .Z(\OutEdge126[0] ) );
    VMW_OAI211 U93 ( .A(n96), .B(n88), .C(n585), .D(n586), .Z(n584) );
    VMW_NAND2 U94 ( .A(n585), .B(n588), .Z(n587) );
    VMW_AO22 U95 ( .A(\temp294[15] ), .B(n586), .C(InEdges[47]), .D(n104), .Z(
        \temp384[15] ) );
    VMW_INV U96 ( .A(n88), .Z(n589) );
    VMW_OAI22 U97 ( .A(n591), .B(Start), .C(\path[2] ), .D(n569), .Z(n590) );
    VMW_OAI22 U98 ( .A(n584), .B(Start), .C(\path[1] ), .D(n569), .Z(n592) );
    VMW_OAI22 U99 ( .A(n587), .B(Start), .C(\path[0] ), .D(n569), .Z(n593) );
    VMW_MUX2I U100 ( .A(\temp384[15] ), .B(InEdges[63]), .S(n112), .Z(n567) );
    VMW_AND3 U101 ( .A(n595), .B(n596), .C(n597), .Z(n594) );
    VMW_INV U102 ( .A(Start), .Z(n569) );
    VMW_INV U103 ( .A(n96), .Z(n598) );
    VMW_OAI21 U104 ( .A(n96), .B(n589), .C(n586), .Z(n588) );
    VMW_AND4 U105 ( .A(n599), .B(n600), .C(n601), .D(n594), .Z(n602) );
    VMW_XNOR2 U106 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n596) );
    VMW_XNOR2 U107 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n595) );
    VMW_XNOR2 U108 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n597) );
    VMW_XNOR2 U109 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n600) );
    VMW_XNOR2 U110 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n599) );
    VMW_XNOR2 U111 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n601) );
    VMW_AO22 U112 ( .A(InEdges[9]), .B(n88), .C(OutEdge[9]), .D(n589), .Z(
        \temp200[9] ) );
    VMW_AO22 U113 ( .A(InEdges[25]), .B(n96), .C(\temp200[9] ), .D(n598), .Z(
        \temp294[9] ) );
    VMW_AO22 U114 ( .A(\temp294[9] ), .B(n586), .C(InEdges[41]), .D(n104), .Z(
        \temp384[9] ) );
    VMW_AO22 U115 ( .A(InEdges[8]), .B(n88), .C(OutEdge[8]), .D(n589), .Z(
        \temp200[8] ) );
    VMW_AO22 U116 ( .A(InEdges[24]), .B(n96), .C(\temp200[8] ), .D(n598), .Z(
        \temp294[8] ) );
    VMW_AO22 U117 ( .A(\temp294[8] ), .B(n586), .C(InEdges[40]), .D(n104), .Z(
        \temp384[8] ) );
    VMW_AO22 U118 ( .A(InEdges[7]), .B(n88), .C(OutEdge[7]), .D(n589), .Z(
        \temp200[7] ) );
    VMW_AO22 U119 ( .A(InEdges[23]), .B(n96), .C(\temp200[7] ), .D(n598), .Z(
        \temp294[7] ) );
    VMW_AO22 U120 ( .A(\temp294[7] ), .B(n586), .C(InEdges[39]), .D(n104), .Z(
        \temp384[7] ) );
    VMW_AO22 U121 ( .A(InEdges[6]), .B(n88), .C(OutEdge[6]), .D(n589), .Z(
        \temp200[6] ) );
    VMW_AO22 U122 ( .A(InEdges[22]), .B(n96), .C(\temp200[6] ), .D(n598), .Z(
        \temp294[6] ) );
    VMW_AO22 U123 ( .A(\temp294[6] ), .B(n586), .C(InEdges[38]), .D(n104), .Z(
        \temp384[6] ) );
    VMW_AO22 U124 ( .A(InEdges[5]), .B(n88), .C(OutEdge[5]), .D(n589), .Z(
        \temp200[5] ) );
    VMW_AO22 U125 ( .A(InEdges[21]), .B(n96), .C(\temp200[5] ), .D(n598), .Z(
        \temp294[5] ) );
    VMW_AO22 U126 ( .A(\temp294[5] ), .B(n586), .C(InEdges[37]), .D(n104), .Z(
        \temp384[5] ) );
    VMW_AO22 U127 ( .A(InEdges[4]), .B(n88), .C(OutEdge[4]), .D(n589), .Z(
        \temp200[4] ) );
    VMW_AO22 U128 ( .A(InEdges[20]), .B(n96), .C(\temp200[4] ), .D(n598), .Z(
        \temp294[4] ) );
    VMW_AO22 U129 ( .A(\temp294[4] ), .B(n586), .C(InEdges[36]), .D(n104), .Z(
        \temp384[4] ) );
    VMW_AO22 U130 ( .A(InEdges[3]), .B(n88), .C(OutEdge[3]), .D(n589), .Z(
        \temp200[3] ) );
    VMW_AO22 U131 ( .A(InEdges[19]), .B(n96), .C(\temp200[3] ), .D(n598), .Z(
        \temp294[3] ) );
    VMW_AO22 U132 ( .A(\temp294[3] ), .B(n586), .C(InEdges[35]), .D(n104), .Z(
        \temp384[3] ) );
    VMW_AO22 U133 ( .A(InEdges[2]), .B(n88), .C(OutEdge[2]), .D(n589), .Z(
        \temp200[2] ) );
    VMW_AO22 U134 ( .A(InEdges[18]), .B(n96), .C(\temp200[2] ), .D(n598), .Z(
        \temp294[2] ) );
    VMW_AO22 U135 ( .A(\temp294[2] ), .B(n586), .C(InEdges[34]), .D(n104), .Z(
        \temp384[2] ) );
    VMW_AO22 U136 ( .A(InEdges[1]), .B(n88), .C(OutEdge[1]), .D(n589), .Z(
        \temp200[1] ) );
    VMW_AO22 U137 ( .A(InEdges[17]), .B(n96), .C(\temp200[1] ), .D(n598), .Z(
        \temp294[1] ) );
    VMW_AO22 U138 ( .A(\temp294[1] ), .B(n586), .C(InEdges[33]), .D(n104), .Z(
        \temp384[1] ) );
    VMW_AO22 U139 ( .A(InEdges[15]), .B(n88), .C(OutEdge[15]), .D(n589), .Z(
        \temp200[15] ) );
    VMW_AO22 U140 ( .A(InEdges[31]), .B(n96), .C(\temp200[15] ), .D(n598), .Z(
        \temp294[15] ) );
    VMW_AO22 U141 ( .A(InEdges[14]), .B(n88), .C(OutEdge[14]), .D(n589), .Z(
        \temp200[14] ) );
    VMW_AO22 U142 ( .A(InEdges[30]), .B(n96), .C(\temp200[14] ), .D(n598), .Z(
        \temp294[14] ) );
    VMW_AO22 U143 ( .A(\temp294[14] ), .B(n586), .C(InEdges[46]), .D(n104), 
        .Z(\temp384[14] ) );
    VMW_AO22 U144 ( .A(InEdges[13]), .B(n88), .C(OutEdge[13]), .D(n589), .Z(
        \temp200[13] ) );
    VMW_AO22 U145 ( .A(InEdges[29]), .B(n96), .C(\temp200[13] ), .D(n598), .Z(
        \temp294[13] ) );
    VMW_AO22 U146 ( .A(\temp294[13] ), .B(n586), .C(InEdges[45]), .D(n104), 
        .Z(\temp384[13] ) );
    VMW_AO22 U147 ( .A(InEdges[12]), .B(n88), .C(OutEdge[12]), .D(n589), .Z(
        \temp200[12] ) );
    VMW_AO22 U148 ( .A(InEdges[28]), .B(n96), .C(\temp200[12] ), .D(n598), .Z(
        \temp294[12] ) );
    VMW_AO22 U149 ( .A(\temp294[12] ), .B(n586), .C(InEdges[44]), .D(n104), 
        .Z(\temp384[12] ) );
    VMW_AO22 U150 ( .A(InEdges[11]), .B(n88), .C(OutEdge[11]), .D(n589), .Z(
        \temp200[11] ) );
    VMW_AO22 U151 ( .A(InEdges[27]), .B(n96), .C(\temp200[11] ), .D(n598), .Z(
        \temp294[11] ) );
    VMW_AO22 U152 ( .A(\temp294[11] ), .B(n586), .C(InEdges[43]), .D(n104), 
        .Z(\temp384[11] ) );
    VMW_AO22 U153 ( .A(InEdges[10]), .B(n88), .C(OutEdge[10]), .D(n589), .Z(
        \temp200[10] ) );
    VMW_AO22 U154 ( .A(InEdges[26]), .B(n96), .C(\temp200[10] ), .D(n598), .Z(
        \temp294[10] ) );
    VMW_AO22 U155 ( .A(\temp294[10] ), .B(n586), .C(InEdges[42]), .D(n104), 
        .Z(\temp384[10] ) );
    VMW_AO22 U156 ( .A(InEdges[0]), .B(n88), .C(OutEdge[0]), .D(n589), .Z(
        \temp200[0] ) );
    VMW_AO22 U157 ( .A(InEdges[16]), .B(n96), .C(\temp200[0] ), .D(n598), .Z(
        \temp294[0] ) );
    VMW_AO22 U158 ( .A(\temp294[0] ), .B(n586), .C(InEdges[32]), .D(n104), .Z(
        \temp384[0] ) );
    VMW_AND4 U159 ( .A(n598), .B(n586), .C(n589), .D(n585), .Z(n591) );
    VMW_MUX2I U160 ( .A(\temp384[9] ), .B(InEdges[57]), .S(n112), .Z(n574) );
    VMW_MUX2I U161 ( .A(\temp384[8] ), .B(InEdges[56]), .S(n112), .Z(n575) );
    VMW_MUX2I U162 ( .A(\temp384[7] ), .B(InEdges[55]), .S(n112), .Z(n576) );
    VMW_MUX2I U163 ( .A(\temp384[6] ), .B(InEdges[54]), .S(n112), .Z(n577) );
    VMW_MUX2I U164 ( .A(\temp384[5] ), .B(InEdges[53]), .S(n112), .Z(n578) );
    VMW_MUX2I U165 ( .A(\temp384[4] ), .B(InEdges[52]), .S(n112), .Z(n579) );
    VMW_MUX2I U166 ( .A(\temp384[3] ), .B(InEdges[51]), .S(n112), .Z(n580) );
    VMW_MUX2I U167 ( .A(\temp384[2] ), .B(InEdges[50]), .S(n112), .Z(n581) );
    VMW_MUX2I U168 ( .A(\temp384[1] ), .B(InEdges[49]), .S(n112), .Z(n582) );
    VMW_MUX2I U169 ( .A(\temp384[14] ), .B(InEdges[62]), .S(n112), .Z(n568) );
    VMW_MUX2I U170 ( .A(\temp384[13] ), .B(InEdges[61]), .S(n112), .Z(n570) );
    VMW_MUX2I U171 ( .A(\temp384[12] ), .B(InEdges[60]), .S(n112), .Z(n571) );
    VMW_MUX2I U172 ( .A(\temp384[11] ), .B(InEdges[59]), .S(n112), .Z(n572) );
    VMW_MUX2I U173 ( .A(\temp384[10] ), .B(InEdges[58]), .S(n112), .Z(n573) );
    VMW_MUX2I U174 ( .A(\temp384[0] ), .B(InEdges[48]), .S(n112), .Z(n583) );
    VMW_INV U175 ( .A(n104), .Z(n586) );
    VMW_INV U176 ( .A(n112), .Z(n585) );
    VMW_INV U177 ( .A(n590), .Z(n604) );
    VMW_INV U178 ( .A(n592), .Z(n605) );
    VMW_INV U179 ( .A(n593), .Z(n603) );
    VMW_BUFIZ U180 ( .A(\path[1] ), .E(n602), .Z(\PathData[1] ) );
    VMW_BUFIZ U181 ( .A(\path[0] ), .E(n602), .Z(\PathData[0] ) );
    VMW_BUFIZ U182 ( .A(\path[2] ), .E(n602), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n603), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n604), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n605), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge126[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge126[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge126[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge126[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge126[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge126[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge126[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge126[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge126[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge126[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge126[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge126[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge126[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge126[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge126[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge126[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n609), .TC(n609), .GE_GT(n88) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp200[15] , 
        \temp200[14] , \temp200[13] , \temp200[12] , \temp200[11] , 
        \temp200[10] , \temp200[9] , \temp200[8] , \temp200[7] , \temp200[6] , 
        \temp200[5] , \temp200[4] , \temp200[3] , \temp200[2] , \temp200[1] , 
        \temp200[0] }), .B(InEdges[31:16]), .LEQ(n608), .TC(n608), .GE_GT(n96)
         );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp294[15] , 
        \temp294[14] , \temp294[13] , \temp294[12] , \temp294[11] , 
        \temp294[10] , \temp294[9] , \temp294[8] , \temp294[7] , \temp294[6] , 
        \temp294[5] , \temp294[4] , \temp294[3] , \temp294[2] , \temp294[1] , 
        \temp294[0] }), .B(InEdges[47:32]), .LEQ(n607), .TC(n607), .GE_GT(n104
        ) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp384[15] , 
        \temp384[14] , \temp384[13] , \temp384[12] , \temp384[11] , 
        \temp384[10] , \temp384[9] , \temp384[8] , \temp384[7] , \temp384[6] , 
        \temp384[5] , \temp384[4] , \temp384[3] , \temp384[2] , \temp384[1] , 
        \temp384[0] }), .B(InEdges[63:48]), .LEQ(n606), .TC(n606), .GE_GT(n112
        ) );
endmodule


module library ( InEdges, OutEdge, PathAddr, PathData, WeightAddr, WeightData, 
    Nid, Eid, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
input  [7:0] WeightAddr;
input  [7:0] Eid;
output [2:0] PathData;
input  [15:0] WeightData;
input  [5:0] Nid;
input  Start, Clk;
    EdgeAux edgeAux ( .Eid(Eid), .InEdge(InEdges[15:0]), .OutEdge(OutEdge), 
        .WeightAddr(WeightAddr), .WeightData(WeightData), .Clk(Clk) );
    NodeAux_INDEGREE2_SOURCE1 n_2_1 ( .Nid(Nid), .InEdges(InEdges[31:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE4_SOURCE0 n_4_0 ( .Nid(Nid), .InEdges(InEdges), .OutEdge(
        OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(Start), 
        .Clk(Clk) );
    NodeAux_INDEGREE2_SOURCE0 n_2_0 ( .Nid(Nid), .InEdges(InEdges[31:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE3_SOURCE0 n_3_0 ( .Nid(Nid), .InEdges(InEdges[47:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
endmodule



module Node_NID0_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE1 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID0 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID1_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID3 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID4 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID2_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID5 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID6 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID7 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID3_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID8 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID9 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID10 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID4_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID11 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID12 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID13 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID5_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID14 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID15 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID16 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID6_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID17 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID18 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID19 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID7_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID20 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID21 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID8_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID22 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID23 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID24 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID9_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID25 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID26 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID27 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID28 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID10_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID29 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID30 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID31 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID32 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID11_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID33 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID34 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID35 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID36 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID12_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID37 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID38 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID39 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID40 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID13_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID41 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID42 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID43 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID44 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID14_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID45 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID46 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID47 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID48 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID15_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID49 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID50 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID51 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID16_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID52 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID53 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID54 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID17_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID55 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID56 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID57 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID58 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID18_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID59 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID60 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID61 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID62 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID19_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID63 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID64 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID65 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID66 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID20_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID67 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID68 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID69 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID70 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID21_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID71 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID72 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID73 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID74 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID22_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID75 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID76 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID77 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID78 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID23_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID79 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID80 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID81 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID24_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID82 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID83 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID84 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID25_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID85 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID86 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID87 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID88 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID26_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID89 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID90 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID91 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID92 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID27_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID93 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID94 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID95 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID96 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID28_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID97 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID98 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID99 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID100 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID29_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID101 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID102 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID103 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID104 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID30_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID105 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID106 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID107 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID108 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID31_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID109 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID110 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID111 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID32_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID112 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID113 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID114 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID33_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID115 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID116 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID117 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID118 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID34_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID119 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID120 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID121 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID122 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID35_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID123 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID124 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID125 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID126 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID36_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID127 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID128 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID129 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID130 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID37_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID131 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID132 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID133 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID134 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID38_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID135 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID136 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID137 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID138 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID39_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID139 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID140 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID141 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID40_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID142 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID143 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID144 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID41_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID145 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID146 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID147 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID148 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID42_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID149 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID150 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID151 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID152 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID43_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID153 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID154 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID155 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID156 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID44_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID157 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID158 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID159 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID160 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID45_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID161 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID162 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID163 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID164 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID46_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID165 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID166 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID167 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID168 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID47_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID169 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID170 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID171 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID48_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID172 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID173 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID174 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID49_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID175 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID176 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID177 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID178 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID50_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID179 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID180 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID181 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID182 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID51_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID183 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID184 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID185 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID186 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID52_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID187 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID188 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID189 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID190 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID53_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID191 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID192 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID193 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID194 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID54_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID195 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID196 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID197 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID198 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID55_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID199 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID200 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID201 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID56_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID202 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID203 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID57_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID204 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID205 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID206 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID58_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID207 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID208 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID209 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID59_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID210 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID211 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID212 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID60_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID213 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID214 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID215 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID61_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID216 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID217 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID218 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID62_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID219 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID220 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID221 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID63_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID222 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID223 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module graph ( WeightAddr, WeightData, PathAddr, PathData, Start, Clk );
input  [7:0] WeightAddr;
input  [15:0] WeightData;
input  [5:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire [31:0] In0;
    wire [15:0] Out0;
    wire [47:0] In1;
    wire [15:0] Out1;
    wire [47:0] In2;
    wire [15:0] Out2;
    wire [47:0] In3;
    wire [15:0] Out3;
    wire [47:0] In4;
    wire [15:0] Out4;
    wire [47:0] In5;
    wire [15:0] Out5;
    wire [47:0] In6;
    wire [15:0] Out6;
    wire [31:0] In7;
    wire [15:0] Out7;
    wire [47:0] In8;
    wire [15:0] Out8;
    wire [63:0] In9;
    wire [15:0] Out9;
    wire [63:0] In10;
    wire [15:0] Out10;
    wire [63:0] In11;
    wire [15:0] Out11;
    wire [63:0] In12;
    wire [15:0] Out12;
    wire [63:0] In13;
    wire [15:0] Out13;
    wire [63:0] In14;
    wire [15:0] Out14;
    wire [47:0] In15;
    wire [15:0] Out15;
    wire [47:0] In16;
    wire [15:0] Out16;
    wire [63:0] In17;
    wire [15:0] Out17;
    wire [63:0] In18;
    wire [15:0] Out18;
    wire [63:0] In19;
    wire [15:0] Out19;
    wire [63:0] In20;
    wire [15:0] Out20;
    wire [63:0] In21;
    wire [15:0] Out21;
    wire [63:0] In22;
    wire [15:0] Out22;
    wire [47:0] In23;
    wire [15:0] Out23;
    wire [47:0] In24;
    wire [15:0] Out24;
    wire [63:0] In25;
    wire [15:0] Out25;
    wire [63:0] In26;
    wire [15:0] Out26;
    wire [63:0] In27;
    wire [15:0] Out27;
    wire [63:0] In28;
    wire [15:0] Out28;
    wire [63:0] In29;
    wire [15:0] Out29;
    wire [63:0] In30;
    wire [15:0] Out30;
    wire [47:0] In31;
    wire [15:0] Out31;
    wire [47:0] In32;
    wire [15:0] Out32;
    wire [63:0] In33;
    wire [15:0] Out33;
    wire [63:0] In34;
    wire [15:0] Out34;
    wire [63:0] In35;
    wire [15:0] Out35;
    wire [63:0] In36;
    wire [15:0] Out36;
    wire [63:0] In37;
    wire [15:0] Out37;
    wire [63:0] In38;
    wire [15:0] Out38;
    wire [47:0] In39;
    wire [15:0] Out39;
    wire [47:0] In40;
    wire [15:0] Out40;
    wire [63:0] In41;
    wire [15:0] Out41;
    wire [63:0] In42;
    wire [15:0] Out42;
    wire [63:0] In43;
    wire [15:0] Out43;
    wire [63:0] In44;
    wire [15:0] Out44;
    wire [63:0] In45;
    wire [15:0] Out45;
    wire [63:0] In46;
    wire [15:0] Out46;
    wire [47:0] In47;
    wire [15:0] Out47;
    wire [47:0] In48;
    wire [15:0] Out48;
    wire [63:0] In49;
    wire [15:0] Out49;
    wire [63:0] In50;
    wire [15:0] Out50;
    wire [63:0] In51;
    wire [15:0] Out51;
    wire [63:0] In52;
    wire [15:0] Out52;
    wire [63:0] In53;
    wire [15:0] Out53;
    wire [63:0] In54;
    wire [15:0] Out54;
    wire [47:0] In55;
    wire [15:0] Out55;
    wire [31:0] In56;
    wire [15:0] Out56;
    wire [47:0] In57;
    wire [15:0] Out57;
    wire [47:0] In58;
    wire [15:0] Out58;
    wire [47:0] In59;
    wire [15:0] Out59;
    wire [47:0] In60;
    wire [15:0] Out60;
    wire [47:0] In61;
    wire [15:0] Out61;
    wire [47:0] In62;
    wire [15:0] Out62;
    wire [31:0] In63;
    wire [15:0] Out63;

    Node_NID0_INDEGREE2 n0 ( .InEdges(In0), .OutEdge(Out0),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID0 e0 ( .InEdge(Out8), .OutEdge(In0[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1 e1 ( .InEdge(Out1), .OutEdge(In0[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID1_INDEGREE3 n1 ( .InEdges(In1), .OutEdge(Out1),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2 e2 ( .InEdge(Out9), .OutEdge(In1[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID3 e3 ( .InEdge(Out2), .OutEdge(In1[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID4 e4 ( .InEdge(Out0), .OutEdge(In1[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID2_INDEGREE3 n2 ( .InEdges(In2), .OutEdge(Out2),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID5 e5 ( .InEdge(Out10), .OutEdge(In2[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID6 e6 ( .InEdge(Out3), .OutEdge(In2[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID7 e7 ( .InEdge(Out1), .OutEdge(In2[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID3_INDEGREE3 n3 ( .InEdges(In3), .OutEdge(Out3),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID8 e8 ( .InEdge(Out11), .OutEdge(In3[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID9 e9 ( .InEdge(Out4), .OutEdge(In3[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID10 e10 ( .InEdge(Out2), .OutEdge(In3[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID4_INDEGREE3 n4 ( .InEdges(In4), .OutEdge(Out4),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID11 e11 ( .InEdge(Out12), .OutEdge(In4[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID12 e12 ( .InEdge(Out5), .OutEdge(In4[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID13 e13 ( .InEdge(Out3), .OutEdge(In4[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID5_INDEGREE3 n5 ( .InEdges(In5), .OutEdge(Out5),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID14 e14 ( .InEdge(Out13), .OutEdge(In5[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID15 e15 ( .InEdge(Out6), .OutEdge(In5[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID16 e16 ( .InEdge(Out4), .OutEdge(In5[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID6_INDEGREE3 n6 ( .InEdges(In6), .OutEdge(Out6),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID17 e17 ( .InEdge(Out14), .OutEdge(In6[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID18 e18 ( .InEdge(Out7), .OutEdge(In6[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID19 e19 ( .InEdge(Out5), .OutEdge(In6[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID7_INDEGREE2 n7 ( .InEdges(In7), .OutEdge(Out7),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID20 e20 ( .InEdge(Out15), .OutEdge(In7[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID21 e21 ( .InEdge(Out6), .OutEdge(In7[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID8_INDEGREE3 n8 ( .InEdges(In8), .OutEdge(Out8),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID22 e22 ( .InEdge(Out16), .OutEdge(In8[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID23 e23 ( .InEdge(Out9), .OutEdge(In8[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID24 e24 ( .InEdge(Out0), .OutEdge(In8[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID9_INDEGREE4 n9 ( .InEdges(In9), .OutEdge(Out9),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID25 e25 ( .InEdge(Out17), .OutEdge(In9[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID26 e26 ( .InEdge(Out10), .OutEdge(In9[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID27 e27 ( .InEdge(Out8), .OutEdge(In9[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID28 e28 ( .InEdge(Out1), .OutEdge(In9[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID10_INDEGREE4 n10 ( .InEdges(In10), .OutEdge(Out10),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID29 e29 ( .InEdge(Out18), .OutEdge(In10[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID30 e30 ( .InEdge(Out11), .OutEdge(In10[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID31 e31 ( .InEdge(Out9), .OutEdge(In10[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID32 e32 ( .InEdge(Out2), .OutEdge(In10[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID11_INDEGREE4 n11 ( .InEdges(In11), .OutEdge(Out11),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID33 e33 ( .InEdge(Out19), .OutEdge(In11[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID34 e34 ( .InEdge(Out12), .OutEdge(In11[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID35 e35 ( .InEdge(Out10), .OutEdge(In11[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID36 e36 ( .InEdge(Out3), .OutEdge(In11[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID12_INDEGREE4 n12 ( .InEdges(In12), .OutEdge(Out12),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID37 e37 ( .InEdge(Out20), .OutEdge(In12[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID38 e38 ( .InEdge(Out13), .OutEdge(In12[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID39 e39 ( .InEdge(Out11), .OutEdge(In12[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID40 e40 ( .InEdge(Out4), .OutEdge(In12[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID13_INDEGREE4 n13 ( .InEdges(In13), .OutEdge(Out13),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID41 e41 ( .InEdge(Out21), .OutEdge(In13[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID42 e42 ( .InEdge(Out14), .OutEdge(In13[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID43 e43 ( .InEdge(Out12), .OutEdge(In13[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID44 e44 ( .InEdge(Out5), .OutEdge(In13[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID14_INDEGREE4 n14 ( .InEdges(In14), .OutEdge(Out14),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID45 e45 ( .InEdge(Out22), .OutEdge(In14[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID46 e46 ( .InEdge(Out15), .OutEdge(In14[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID47 e47 ( .InEdge(Out13), .OutEdge(In14[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID48 e48 ( .InEdge(Out6), .OutEdge(In14[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID15_INDEGREE3 n15 ( .InEdges(In15), .OutEdge(Out15),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID49 e49 ( .InEdge(Out23), .OutEdge(In15[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID50 e50 ( .InEdge(Out14), .OutEdge(In15[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID51 e51 ( .InEdge(Out7), .OutEdge(In15[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID16_INDEGREE3 n16 ( .InEdges(In16), .OutEdge(Out16),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID52 e52 ( .InEdge(Out24), .OutEdge(In16[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID53 e53 ( .InEdge(Out17), .OutEdge(In16[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID54 e54 ( .InEdge(Out8), .OutEdge(In16[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID17_INDEGREE4 n17 ( .InEdges(In17), .OutEdge(Out17),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID55 e55 ( .InEdge(Out25), .OutEdge(In17[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID56 e56 ( .InEdge(Out18), .OutEdge(In17[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID57 e57 ( .InEdge(Out16), .OutEdge(In17[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID58 e58 ( .InEdge(Out9), .OutEdge(In17[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID18_INDEGREE4 n18 ( .InEdges(In18), .OutEdge(Out18),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID59 e59 ( .InEdge(Out26), .OutEdge(In18[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID60 e60 ( .InEdge(Out19), .OutEdge(In18[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID61 e61 ( .InEdge(Out17), .OutEdge(In18[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID62 e62 ( .InEdge(Out10), .OutEdge(In18[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID19_INDEGREE4 n19 ( .InEdges(In19), .OutEdge(Out19),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID63 e63 ( .InEdge(Out27), .OutEdge(In19[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID64 e64 ( .InEdge(Out20), .OutEdge(In19[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID65 e65 ( .InEdge(Out18), .OutEdge(In19[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID66 e66 ( .InEdge(Out11), .OutEdge(In19[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID20_INDEGREE4 n20 ( .InEdges(In20), .OutEdge(Out20),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID67 e67 ( .InEdge(Out28), .OutEdge(In20[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID68 e68 ( .InEdge(Out21), .OutEdge(In20[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID69 e69 ( .InEdge(Out19), .OutEdge(In20[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID70 e70 ( .InEdge(Out12), .OutEdge(In20[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID21_INDEGREE4 n21 ( .InEdges(In21), .OutEdge(Out21),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID71 e71 ( .InEdge(Out29), .OutEdge(In21[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID72 e72 ( .InEdge(Out22), .OutEdge(In21[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID73 e73 ( .InEdge(Out20), .OutEdge(In21[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID74 e74 ( .InEdge(Out13), .OutEdge(In21[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID22_INDEGREE4 n22 ( .InEdges(In22), .OutEdge(Out22),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID75 e75 ( .InEdge(Out30), .OutEdge(In22[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID76 e76 ( .InEdge(Out23), .OutEdge(In22[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID77 e77 ( .InEdge(Out21), .OutEdge(In22[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID78 e78 ( .InEdge(Out14), .OutEdge(In22[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID23_INDEGREE3 n23 ( .InEdges(In23), .OutEdge(Out23),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID79 e79 ( .InEdge(Out31), .OutEdge(In23[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID80 e80 ( .InEdge(Out22), .OutEdge(In23[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID81 e81 ( .InEdge(Out15), .OutEdge(In23[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID24_INDEGREE3 n24 ( .InEdges(In24), .OutEdge(Out24),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID82 e82 ( .InEdge(Out32), .OutEdge(In24[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID83 e83 ( .InEdge(Out25), .OutEdge(In24[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID84 e84 ( .InEdge(Out16), .OutEdge(In24[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID25_INDEGREE4 n25 ( .InEdges(In25), .OutEdge(Out25),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID85 e85 ( .InEdge(Out33), .OutEdge(In25[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID86 e86 ( .InEdge(Out26), .OutEdge(In25[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID87 e87 ( .InEdge(Out24), .OutEdge(In25[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID88 e88 ( .InEdge(Out17), .OutEdge(In25[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID26_INDEGREE4 n26 ( .InEdges(In26), .OutEdge(Out26),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID89 e89 ( .InEdge(Out34), .OutEdge(In26[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID90 e90 ( .InEdge(Out27), .OutEdge(In26[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID91 e91 ( .InEdge(Out25), .OutEdge(In26[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID92 e92 ( .InEdge(Out18), .OutEdge(In26[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID27_INDEGREE4 n27 ( .InEdges(In27), .OutEdge(Out27),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID93 e93 ( .InEdge(Out35), .OutEdge(In27[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID94 e94 ( .InEdge(Out28), .OutEdge(In27[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID95 e95 ( .InEdge(Out26), .OutEdge(In27[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID96 e96 ( .InEdge(Out19), .OutEdge(In27[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID28_INDEGREE4 n28 ( .InEdges(In28), .OutEdge(Out28),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID97 e97 ( .InEdge(Out36), .OutEdge(In28[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID98 e98 ( .InEdge(Out29), .OutEdge(In28[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID99 e99 ( .InEdge(Out27), .OutEdge(In28[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID100 e100 ( .InEdge(Out20), .OutEdge(In28[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID29_INDEGREE4 n29 ( .InEdges(In29), .OutEdge(Out29),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID101 e101 ( .InEdge(Out37), .OutEdge(In29[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID102 e102 ( .InEdge(Out30), .OutEdge(In29[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID103 e103 ( .InEdge(Out28), .OutEdge(In29[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID104 e104 ( .InEdge(Out21), .OutEdge(In29[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID30_INDEGREE4 n30 ( .InEdges(In30), .OutEdge(Out30),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID105 e105 ( .InEdge(Out38), .OutEdge(In30[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID106 e106 ( .InEdge(Out31), .OutEdge(In30[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID107 e107 ( .InEdge(Out29), .OutEdge(In30[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID108 e108 ( .InEdge(Out22), .OutEdge(In30[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID31_INDEGREE3 n31 ( .InEdges(In31), .OutEdge(Out31),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID109 e109 ( .InEdge(Out39), .OutEdge(In31[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID110 e110 ( .InEdge(Out30), .OutEdge(In31[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID111 e111 ( .InEdge(Out23), .OutEdge(In31[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID32_INDEGREE3 n32 ( .InEdges(In32), .OutEdge(Out32),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID112 e112 ( .InEdge(Out40), .OutEdge(In32[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID113 e113 ( .InEdge(Out33), .OutEdge(In32[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID114 e114 ( .InEdge(Out24), .OutEdge(In32[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID33_INDEGREE4 n33 ( .InEdges(In33), .OutEdge(Out33),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID115 e115 ( .InEdge(Out41), .OutEdge(In33[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID116 e116 ( .InEdge(Out34), .OutEdge(In33[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID117 e117 ( .InEdge(Out32), .OutEdge(In33[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID118 e118 ( .InEdge(Out25), .OutEdge(In33[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID34_INDEGREE4 n34 ( .InEdges(In34), .OutEdge(Out34),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID119 e119 ( .InEdge(Out42), .OutEdge(In34[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID120 e120 ( .InEdge(Out35), .OutEdge(In34[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID121 e121 ( .InEdge(Out33), .OutEdge(In34[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID122 e122 ( .InEdge(Out26), .OutEdge(In34[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID35_INDEGREE4 n35 ( .InEdges(In35), .OutEdge(Out35),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID123 e123 ( .InEdge(Out43), .OutEdge(In35[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID124 e124 ( .InEdge(Out36), .OutEdge(In35[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID125 e125 ( .InEdge(Out34), .OutEdge(In35[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID126 e126 ( .InEdge(Out27), .OutEdge(In35[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID36_INDEGREE4 n36 ( .InEdges(In36), .OutEdge(Out36),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID127 e127 ( .InEdge(Out44), .OutEdge(In36[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID128 e128 ( .InEdge(Out37), .OutEdge(In36[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID129 e129 ( .InEdge(Out35), .OutEdge(In36[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID130 e130 ( .InEdge(Out28), .OutEdge(In36[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID37_INDEGREE4 n37 ( .InEdges(In37), .OutEdge(Out37),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID131 e131 ( .InEdge(Out45), .OutEdge(In37[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID132 e132 ( .InEdge(Out38), .OutEdge(In37[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID133 e133 ( .InEdge(Out36), .OutEdge(In37[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID134 e134 ( .InEdge(Out29), .OutEdge(In37[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID38_INDEGREE4 n38 ( .InEdges(In38), .OutEdge(Out38),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID135 e135 ( .InEdge(Out46), .OutEdge(In38[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID136 e136 ( .InEdge(Out39), .OutEdge(In38[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID137 e137 ( .InEdge(Out37), .OutEdge(In38[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID138 e138 ( .InEdge(Out30), .OutEdge(In38[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID39_INDEGREE3 n39 ( .InEdges(In39), .OutEdge(Out39),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID139 e139 ( .InEdge(Out47), .OutEdge(In39[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID140 e140 ( .InEdge(Out38), .OutEdge(In39[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID141 e141 ( .InEdge(Out31), .OutEdge(In39[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID40_INDEGREE3 n40 ( .InEdges(In40), .OutEdge(Out40),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID142 e142 ( .InEdge(Out48), .OutEdge(In40[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID143 e143 ( .InEdge(Out41), .OutEdge(In40[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID144 e144 ( .InEdge(Out32), .OutEdge(In40[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID41_INDEGREE4 n41 ( .InEdges(In41), .OutEdge(Out41),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID145 e145 ( .InEdge(Out49), .OutEdge(In41[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID146 e146 ( .InEdge(Out42), .OutEdge(In41[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID147 e147 ( .InEdge(Out40), .OutEdge(In41[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID148 e148 ( .InEdge(Out33), .OutEdge(In41[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID42_INDEGREE4 n42 ( .InEdges(In42), .OutEdge(Out42),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID149 e149 ( .InEdge(Out50), .OutEdge(In42[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID150 e150 ( .InEdge(Out43), .OutEdge(In42[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID151 e151 ( .InEdge(Out41), .OutEdge(In42[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID152 e152 ( .InEdge(Out34), .OutEdge(In42[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID43_INDEGREE4 n43 ( .InEdges(In43), .OutEdge(Out43),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID153 e153 ( .InEdge(Out51), .OutEdge(In43[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID154 e154 ( .InEdge(Out44), .OutEdge(In43[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID155 e155 ( .InEdge(Out42), .OutEdge(In43[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID156 e156 ( .InEdge(Out35), .OutEdge(In43[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID44_INDEGREE4 n44 ( .InEdges(In44), .OutEdge(Out44),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID157 e157 ( .InEdge(Out52), .OutEdge(In44[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID158 e158 ( .InEdge(Out45), .OutEdge(In44[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID159 e159 ( .InEdge(Out43), .OutEdge(In44[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID160 e160 ( .InEdge(Out36), .OutEdge(In44[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID45_INDEGREE4 n45 ( .InEdges(In45), .OutEdge(Out45),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID161 e161 ( .InEdge(Out53), .OutEdge(In45[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID162 e162 ( .InEdge(Out46), .OutEdge(In45[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID163 e163 ( .InEdge(Out44), .OutEdge(In45[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID164 e164 ( .InEdge(Out37), .OutEdge(In45[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID46_INDEGREE4 n46 ( .InEdges(In46), .OutEdge(Out46),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID165 e165 ( .InEdge(Out54), .OutEdge(In46[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID166 e166 ( .InEdge(Out47), .OutEdge(In46[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID167 e167 ( .InEdge(Out45), .OutEdge(In46[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID168 e168 ( .InEdge(Out38), .OutEdge(In46[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID47_INDEGREE3 n47 ( .InEdges(In47), .OutEdge(Out47),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID169 e169 ( .InEdge(Out55), .OutEdge(In47[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID170 e170 ( .InEdge(Out46), .OutEdge(In47[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID171 e171 ( .InEdge(Out39), .OutEdge(In47[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID48_INDEGREE3 n48 ( .InEdges(In48), .OutEdge(Out48),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID172 e172 ( .InEdge(Out56), .OutEdge(In48[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID173 e173 ( .InEdge(Out49), .OutEdge(In48[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID174 e174 ( .InEdge(Out40), .OutEdge(In48[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID49_INDEGREE4 n49 ( .InEdges(In49), .OutEdge(Out49),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID175 e175 ( .InEdge(Out57), .OutEdge(In49[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID176 e176 ( .InEdge(Out50), .OutEdge(In49[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID177 e177 ( .InEdge(Out48), .OutEdge(In49[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID178 e178 ( .InEdge(Out41), .OutEdge(In49[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID50_INDEGREE4 n50 ( .InEdges(In50), .OutEdge(Out50),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID179 e179 ( .InEdge(Out58), .OutEdge(In50[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID180 e180 ( .InEdge(Out51), .OutEdge(In50[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID181 e181 ( .InEdge(Out49), .OutEdge(In50[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID182 e182 ( .InEdge(Out42), .OutEdge(In50[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID51_INDEGREE4 n51 ( .InEdges(In51), .OutEdge(Out51),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID183 e183 ( .InEdge(Out59), .OutEdge(In51[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID184 e184 ( .InEdge(Out52), .OutEdge(In51[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID185 e185 ( .InEdge(Out50), .OutEdge(In51[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID186 e186 ( .InEdge(Out43), .OutEdge(In51[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID52_INDEGREE4 n52 ( .InEdges(In52), .OutEdge(Out52),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID187 e187 ( .InEdge(Out60), .OutEdge(In52[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID188 e188 ( .InEdge(Out53), .OutEdge(In52[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID189 e189 ( .InEdge(Out51), .OutEdge(In52[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID190 e190 ( .InEdge(Out44), .OutEdge(In52[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID53_INDEGREE4 n53 ( .InEdges(In53), .OutEdge(Out53),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID191 e191 ( .InEdge(Out61), .OutEdge(In53[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID192 e192 ( .InEdge(Out54), .OutEdge(In53[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID193 e193 ( .InEdge(Out52), .OutEdge(In53[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID194 e194 ( .InEdge(Out45), .OutEdge(In53[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID54_INDEGREE4 n54 ( .InEdges(In54), .OutEdge(Out54),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID195 e195 ( .InEdge(Out62), .OutEdge(In54[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID196 e196 ( .InEdge(Out55), .OutEdge(In54[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID197 e197 ( .InEdge(Out53), .OutEdge(In54[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID198 e198 ( .InEdge(Out46), .OutEdge(In54[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID55_INDEGREE3 n55 ( .InEdges(In55), .OutEdge(Out55),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID199 e199 ( .InEdge(Out63), .OutEdge(In55[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID200 e200 ( .InEdge(Out54), .OutEdge(In55[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID201 e201 ( .InEdge(Out47), .OutEdge(In55[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID56_INDEGREE2 n56 ( .InEdges(In56), .OutEdge(Out56),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID202 e202 ( .InEdge(Out57), .OutEdge(In56[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID203 e203 ( .InEdge(Out48), .OutEdge(In56[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID57_INDEGREE3 n57 ( .InEdges(In57), .OutEdge(Out57),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID204 e204 ( .InEdge(Out58), .OutEdge(In57[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID205 e205 ( .InEdge(Out56), .OutEdge(In57[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID206 e206 ( .InEdge(Out49), .OutEdge(In57[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID58_INDEGREE3 n58 ( .InEdges(In58), .OutEdge(Out58),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID207 e207 ( .InEdge(Out59), .OutEdge(In58[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID208 e208 ( .InEdge(Out57), .OutEdge(In58[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID209 e209 ( .InEdge(Out50), .OutEdge(In58[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID59_INDEGREE3 n59 ( .InEdges(In59), .OutEdge(Out59),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID210 e210 ( .InEdge(Out60), .OutEdge(In59[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID211 e211 ( .InEdge(Out58), .OutEdge(In59[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID212 e212 ( .InEdge(Out51), .OutEdge(In59[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID60_INDEGREE3 n60 ( .InEdges(In60), .OutEdge(Out60),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID213 e213 ( .InEdge(Out61), .OutEdge(In60[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID214 e214 ( .InEdge(Out59), .OutEdge(In60[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID215 e215 ( .InEdge(Out52), .OutEdge(In60[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID61_INDEGREE3 n61 ( .InEdges(In61), .OutEdge(Out61),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID216 e216 ( .InEdge(Out62), .OutEdge(In61[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID217 e217 ( .InEdge(Out60), .OutEdge(In61[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID218 e218 ( .InEdge(Out53), .OutEdge(In61[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID62_INDEGREE3 n62 ( .InEdges(In62), .OutEdge(Out62),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID219 e219 ( .InEdge(Out63), .OutEdge(In62[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID220 e220 ( .InEdge(Out61), .OutEdge(In62[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID221 e221 ( .InEdge(Out54), .OutEdge(In62[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID63_INDEGREE2 n63 ( .InEdges(In63), .OutEdge(Out63),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID222 e222 ( .InEdge(Out62), .OutEdge(In63[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID223 e223 ( .InEdge(Out55), .OutEdge(In63[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
endmodule
