
module EdgeAux_DW01_add_30_0 ( A, B, CI, SUM, CO );
input  [29:0] A;
input  [29:0] B;
output [29:0] SUM;
input  CI;
output CO;
    wire \SUM1[11] , \SUM1[2] , \SUM1[6] , \SUM1[4] , \SUM1[9] , \SUM1[0] , 
        \SUM1[13] , \SUM1[8] , \SUM1[1] , \SUM1[12] , \SUM1[5] , \SUM1[7] , 
        \SUM1[10] , \SUM1[3] ;
    assign \SUM1[13]  = A[13];
    assign \SUM1[12]  = A[12];
    assign \SUM1[11]  = A[11];
    assign \SUM1[10]  = A[10];
    assign \SUM1[9]  = A[9];
    assign \SUM1[8]  = A[8];
    assign \SUM1[7]  = A[7];
    assign \SUM1[6]  = A[6];
    assign \SUM1[5]  = A[5];
    assign \SUM1[4]  = A[4];
    assign \SUM1[3]  = A[3];
    assign \SUM1[2]  = A[2];
    assign \SUM1[1]  = A[1];
    assign \SUM1[0]  = A[0];
    assign SUM[13] = \SUM1[13] ;
    assign SUM[12] = \SUM1[12] ;
    assign SUM[11] = \SUM1[11] ;
    assign SUM[10] = \SUM1[10] ;
    assign SUM[9] = \SUM1[9] ;
    assign SUM[8] = \SUM1[8] ;
    assign SUM[7] = \SUM1[7] ;
    assign SUM[6] = \SUM1[6] ;
    assign SUM[5] = \SUM1[5] ;
    assign SUM[4] = \SUM1[4] ;
    assign SUM[3] = \SUM1[3] ;
    assign SUM[2] = \SUM1[2] ;
    assign SUM[1] = \SUM1[1] ;
    assign SUM[0] = \SUM1[0] ;
endmodule


module EdgeAux_DW02_mult_16_16_0 ( A, B, TC, PRODUCT );
input  [15:0] A;
input  [15:0] B;
output [31:0] PRODUCT;
input  TC;
    wire \ab[13][0] , \ab[9][1] , \A1[13] , \A1[6] , \A2[5] , \SUMB[12][1] , 
        \ab[3][7] , \SUMB[4][8] , \SUMB[5][2] , \CARRYB[6][3] , \CARRYB[2][1] , 
        \ab[7][5] , \ab[4][11] , \ab[12][3] , \ab[8][2] , \SUMB[13][2] , 
        \SUMB[3][11] , \CARRYB[9][4] , \ab[6][6] , \SUMB[1][9] , 
        \CARRYB[2][8] , \A1[29] , \CARRYB[3][2] , \ab[2][4] , \SUMB[4][1] , 
        \CARRYB[7][0] , \SUMB[1][4] , \CARRYB[2][5] , \ab[7][1] , \ab[3][3] , 
        \SUMB[5][6] , \CARRYB[6][7] , \ab[2][9] , \CARRYB[3][11] , \ab[9][5] , 
        \SUMB[2][13] , \A2[1] , \A1[2] , \CARRYB[8][3] , \ab[2][0] , 
        \SUMB[4][5] , \A2[8] , \CARRYB[7][4] , \ab[6][2] , \CARRYB[12][1] , 
        \CARRYB[3][6] , \ab[8][6] , \ab[7][8] , \CARRYB[9][0] , \ab[2][11] , 
        \CARRYB[9][2] , \ab[8][4] , \ab[3][8] , \ab[2][13] , \SUMB[4][7] , 
        \CARRYB[7][6] , \A1[9] , \ab[6][0] , \ab[2][2] , \CARRYB[3][4] , 
        \SUMB[2][11] , \A1[0] , \A2[3] , \CARRYB[8][1] , \ab[6][9] , 
        \ab[7][3] , \SUMB[1][6] , \CARRYB[13][0] , \CARRYB[2][7] , \ab[6][4] , 
        \ab[3][1] , \SUMB[5][4] , \CARRYB[6][5] , \CARRYB[2][11] , 
        \CARRYB[3][0] , \ab[2][6] , \SUMB[4][3] , \CARRYB[7][2] , \ab[12][1] , 
        \SUMB[5][9] , \CARRYB[6][8] , \ab[8][0] , \CARRYB[6][1] , \ab[3][5] , 
        \SUMB[1][2] , \CARRYB[2][3] , \ab[7][7] , \ab[13][2] , \ab[3][11] , 
        \CARRYB[3][9] , \SUMB[4][11] , \CARRYB[8][5] , \A1[11] , \A2[7] , 
        \A1[4] , \ab[9][3] , \SUMB[12][3] , \ab[11][4] , \SUMB[9][2] , 
        \SUMB[1][14] , \ab[1][3] , \ab[0][10] , \ab[0][9] , \SUMB[10][5] , 
        \ab[5][1] , \SUMB[7][6] , \CARRYB[4][7] , \SUMB[3][4] , 
        \CARRYB[11][2] , \SUMB[8][1] , \A2[14] , \ab[5][8] , \ab[4][2] , 
        \CARRYB[10][1] , \SUMB[2][7] , \CARRYB[1][6] , \SUMB[6][5] , 
        \CARRYB[5][4] , \CARRYB[1][10] , \ab[5][5] , \ab[1][7] , lsb_0, 
        \SUMB[7][2] , \CARRYB[4][3] , \ab[11][0] , \ab[0][14] , \SUMB[10][1] , 
        \SUMB[6][8] , \CARRYB[5][9] , \SUMB[9][6] , \SUMB[1][10] , \ab[0][4] , 
        \SUMB[6][1] , \CARRYB[5][0] , \ab[14][1] , \ab[4][6] , \ab[1][12] , 
        \SUMB[2][3] , \CARRYB[1][2] , \SUMB[3][9] , \ab[10][3] , \SUMB[8][5] , 
        \A2[10] , \SUMB[11][2] , \ab[1][10] , \ab[10][1] , \SUMB[8][7] , 
        \A2[12] , \ab[4][4] , \ab[0][6] , \CARRYB[4][8] , \SUMB[6][3] , 
        \CARRYB[5][2] , \SUMB[2][1] , \CARRYB[1][0] , \ab[15][0] , \ab[11][2] , 
        \SUMB[10][3] , \SUMB[14][1] , \SUMB[9][4] , \SUMB[1][12] , 
        \SUMB[2][8] , \CARRYB[1][9] , \ab[5][7] , \ab[1][5] , \SUMB[3][2] , 
        \CARRYB[4][1] , \ab[4][0] , \ab[0][2] , \SUMB[2][5] , \CARRYB[10][3] , 
        \CARRYB[1][4] , \SUMB[6][7] , \CARRYB[5][6] , \SUMB[11][4] , 
        \CARRYB[1][12] , \ab[10][5] , \ab[1][8] , \ab[1][14] , \SUMB[8][3] , 
        \ab[1][1] , \SUMB[7][4] , \CARRYB[4][5] , \ab[5][3] , \SUMB[3][6] , 
        \CARRYB[11][0] , \ab[4][9] , \ab[4][1] , \ab[0][12] , \ab[10][4] , 
        \SUMB[2][4] , \CARRYB[10][2] , \CARRYB[1][5] , \CARRYB[1][13] , 
        \ab[0][3] , \SUMB[6][6] , \CARRYB[14][0] , \CARRYB[5][7] , \ab[1][9] , 
        \SUMB[8][2] , \ab[1][0] , \CARRYB[4][4] , \SUMB[7][5] , \ab[5][2] , 
        \SUMB[3][7] , \CARRYB[11][1] , \ab[4][8] , \SUMB[9][1] , \ab[0][13] , 
        \ab[1][11] , \A2[13] , \SUMB[8][6] , \SUMB[11][1] , \SUMB[7][8] , 
        \ab[10][0] , \CARRYB[4][9] , \ab[0][7] , \CARRYB[5][3] , \SUMB[6][2] , 
        \ab[11][3] , \ab[4][5] , \CARRYB[1][1] , \SUMB[10][2] , \SUMB[2][9] , 
        \CARRYB[1][8] , \ab[5][6] , \SUMB[9][5] , \SUMB[1][13] , \SUMB[3][3] , 
        \ab[1][4] , \SUMB[7][1] , \ab[5][4] , \CARRYB[4][0] , \SUMB[3][1] , 
        \ab[1][6] , \CARRYB[4][2] , \ab[11][1] , \SUMB[7][3] , \SUMB[6][9] , 
        \ab[0][15] , \CARRYB[5][8] , \ab[0][5] , \SUMB[1][11] , \CARRYB[5][1] , 
        \ab[4][7] , \ab[14][0] , \CARRYB[10][4] , \CARRYB[1][3] , \SUMB[2][2] , 
        \ab[10][2] , \ab[1][13] , \SUMB[8][4] , \SUMB[3][8] , \A2[11] , 
        \SUMB[11][3] , \ab[0][11] , \SUMB[9][3] , \SUMB[10][4] , \ab[0][8] , 
        \ab[1][2] , \SUMB[7][7] , \CARRYB[4][6] , \ab[5][0] , \SUMB[3][5] , 
        \CARRYB[11][3] , \ab[5][9] , \ab[4][3] , \ab[12][0] , \SUMB[2][6] , 
        \CARRYB[10][0] , \CARRYB[1][7] , \ab[6][5] , \ab[0][1] , 
        \CARRYB[1][11] , \CARRYB[5][5] , \SUMB[6][4] , \CARRYB[3][1] , 
        \CARRYB[2][10] , \SUMB[4][2] , \CARRYB[7][3] , \ab[2][7] , \ab[8][1] , 
        \SUMB[13][1] , \SUMB[5][8] , \SUMB[5][1] , \SUMB[3][12] , 
        \CARRYB[6][0] , \ab[3][4] , \CARRYB[2][2] , \ab[7][6] , \SUMB[1][3] , 
        \CARRYB[8][4] , \A1[10] , \ab[3][10] , \SUMB[12][2] , \CARRYB[3][8] , 
        \SUMB[4][10] , \A1[5] , \A2[6] , \ab[9][2] , \CARRYB[9][3] , 
        \ab[3][9] , \ab[2][12] , \ab[8][5] , \ab[2][3] , \SUMB[4][6] , 
        \CARRYB[7][7] , \ab[6][1] , \A1[8] , \CARRYB[12][2] , \CARRYB[4][10] , 
        \CARRYB[3][5] , \SUMB[2][10] , \A2[2] , \A1[1] , \ab[9][6] , 
        \ab[6][8] , \ab[5][10] , \SUMB[1][7] , \CARRYB[8][0] , \CARRYB[13][1] , 
        \ab[7][2] , \CARRYB[2][6] , \ab[3][0] , \SUMB[5][5] , \CARRYB[6][4] , 
        \CARRYB[2][4] , \ab[9][4] , \ab[7][0] , \SUMB[1][5] , \ab[3][2] , 
        \CARRYB[3][10] , \SUMB[5][7] , \CARRYB[6][6] , \SUMB[2][12] , \A1[3] , 
        \ab[2][8] , \SUMB[4][4] , \CARRYB[8][2] , \CARRYB[7][5] , \ab[6][3] , 
        \ab[2][1] , \A2[9] , \CARRYB[12][0] , \CARRYB[3][7] , \SUMB[5][10] , 
        \CARRYB[9][1] , \ab[2][10] , \ab[8][7] , \ab[3][12] , \CARRYB[8][6] , 
        \A1[12] , \SUMB[4][9] , \ab[13][1] , \ab[9][0] , \A2[4] , \A1[7] , 
        \ab[3][6] , \SUMB[5][3] , \CARRYB[6][2] , \SUMB[1][1] , \ab[7][4] , 
        \CARRYB[2][0] , \ab[12][2] , \ab[8][3] , \ab[4][10] , \ab[6][7] , 
        \SUMB[1][8] , \CARRYB[9][5] , \CARRYB[2][9] , \SUMB[3][10] , 
        \CARRYB[3][3] , \CARRYB[2][12] , \ab[2][5] , \CARRYB[7][1] , n31, n32, 
        n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 , UNCONNECTED_23 , UNCONNECTED_24 , 
	UNCONNECTED_25 , UNCONNECTED_26 , UNCONNECTED_27 , UNCONNECTED_28 , 
	UNCONNECTED_29 , UNCONNECTED_30 , UNCONNECTED_31 , UNCONNECTED_32 , 
	UNCONNECTED_33 , UNCONNECTED_34 , UNCONNECTED_35 , UNCONNECTED_36 , 
	UNCONNECTED_37 , UNCONNECTED_38 , UNCONNECTED_39 , UNCONNECTED_40 , 
	UNCONNECTED_41 , UNCONNECTED_42 , UNCONNECTED_43 , UNCONNECTED_44 , 
	UNCONNECTED_45 , UNCONNECTED_46 ;
    VMW_PULLDOWN U3 ( .Z(n31) );
    VMW_PULLDOWN U4 ( .Z(n32) );
    VMW_PULLDOWN U5 ( .Z(n33) );
    VMW_PULLDOWN U6 ( .Z(n34) );
    VMW_PULLDOWN U7 ( .Z(n35) );
    VMW_PULLDOWN U8 ( .Z(n36) );
    VMW_PULLDOWN U9 ( .Z(n37) );
    VMW_PULLDOWN U10 ( .Z(n38) );
    VMW_PULLDOWN U11 ( .Z(n39) );
    VMW_PULLDOWN U12 ( .Z(n40) );
    VMW_PULLDOWN U13 ( .Z(n41) );
    VMW_PULLDOWN U14 ( .Z(n42) );
    VMW_PULLDOWN U15 ( .Z(n43) );
    VMW_PULLDOWN U16 ( .Z(n44) );
    VMW_PULLDOWN U17 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U18 ( .Z(\A2[9] ) );
    VMW_PULLDOWN U19 ( .Z(\A2[2] ) );
    VMW_PULLDOWN U20 ( .Z(\A2[6] ) );
    VMW_PULLDOWN U21 ( .Z(\A2[11] ) );
    VMW_PULLDOWN U22 ( .Z(\A2[13] ) );
    VMW_PULLDOWN U23 ( .Z(\A2[12] ) );
    VMW_PULLDOWN U24 ( .Z(\A2[10] ) );
    VMW_PULLDOWN U25 ( .Z(lsb_0) );
    VMW_PULLDOWN U26 ( .Z(\A2[14] ) );
    VMW_PULLDOWN U27 ( .Z(\A2[7] ) );
    VMW_PULLDOWN U28 ( .Z(\A2[3] ) );
    VMW_PULLDOWN U29 ( .Z(\A2[8] ) );
    VMW_PULLDOWN U30 ( .Z(\A2[1] ) );
    VMW_PULLDOWN U31 ( .Z(\A1[29] ) );
    VMW_PULLDOWN U32 ( .Z(\A2[5] ) );
    VMW_XOR2 U33 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
    VMW_FADD S0_13 ( .CI(n31), .A(\ab[0][14] ), .B(\ab[1][13] ), .S(
        \SUMB[1][13] ), .CO(\CARRYB[1][13] ) );
    VMW_FADD S0_12 ( .CI(n32), .A(\ab[0][13] ), .B(\ab[1][12] ), .S(
        \SUMB[1][12] ), .CO(\CARRYB[1][12] ) );
    VMW_FADD S0_11 ( .CI(n33), .A(\ab[0][12] ), .B(\ab[1][11] ), .S(
        \SUMB[1][11] ), .CO(\CARRYB[1][11] ) );
    VMW_FADD S0_10 ( .CI(n34), .A(\ab[0][11] ), .B(\ab[1][10] ), .S(
        \SUMB[1][10] ), .CO(\CARRYB[1][10] ) );
    VMW_FADD S0_9 ( .CI(n35), .A(\ab[0][10] ), .B(\ab[1][9] ), .S(\SUMB[1][9] 
        ), .CO(\CARRYB[1][9] ) );
    VMW_FADD S0_8 ( .CI(n36), .A(\ab[0][9] ), .B(\ab[1][8] ), .S(\SUMB[1][8] ), 
        .CO(\CARRYB[1][8] ) );
    VMW_FADD S0_7 ( .CI(n37), .A(\ab[0][8] ), .B(\ab[1][7] ), .S(\SUMB[1][7] ), 
        .CO(\CARRYB[1][7] ) );
    VMW_FADD S0_6 ( .CI(n38), .A(\ab[0][7] ), .B(\ab[1][6] ), .S(\SUMB[1][6] ), 
        .CO(\CARRYB[1][6] ) );
    VMW_FADD S0_5 ( .CI(n39), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_FADD S0_4 ( .CI(n40), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S0_3 ( .CI(n41), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_FADD S0_2 ( .CI(n42), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_FADD S0_1 ( .CI(n43), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_FADD S0_0 ( .CI(n44), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U34 ( .A(A[10]), .B(B[5]), .Z(\ab[10][5] ) );
    VMW_AND2 U35 ( .A(A[2]), .B(B[6]), .Z(\ab[2][6] ) );
    VMW_AND2 U36 ( .A(A[7]), .B(B[0]), .Z(\ab[7][0] ) );
    VMW_AND2 U37 ( .A(A[3]), .B(B[6]), .Z(\ab[3][6] ) );
    VMW_AND2 U38 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U39 ( .A(A[13]), .B(B[2]), .Z(\ab[13][2] ) );
    VMW_AND2 U40 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U41 ( .A(A[0]), .B(B[12]), .Z(\ab[0][12] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[5]), .Z(\ab[5][5] ) );
    VMW_AND2 U43 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U44 ( .A(A[12]), .B(B[0]), .Z(\ab[12][0] ) );
    VMW_AND2 U45 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[5]), .Z(\ab[4][5] ) );
    VMW_AND2 U47 ( .A(A[1]), .B(B[13]), .Z(\ab[1][13] ) );
    VMW_AND2 U48 ( .A(B[9]), .B(A[6]), .Z(\ab[6][9] ) );
    VMW_AND2 U49 ( .A(A[13]), .B(B[0]), .Z(\ab[13][0] ) );
    VMW_AND2 U50 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U51 ( .A(B[14]), .B(A[1]), .Z(\ab[1][14] ) );
    VMW_AND2 U52 ( .A(B[5]), .B(A[9]), .Z(\ab[9][5] ) );
    VMW_AND2 U53 ( .A(A[3]), .B(B[8]), .Z(\ab[3][8] ) );
    VMW_AND2 U54 ( .A(A[6]), .B(B[2]), .Z(\ab[6][2] ) );
    VMW_AND2 U55 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U56 ( .A(A[2]), .B(B[8]), .Z(\ab[2][8] ) );
    VMW_AND2 U57 ( .A(A[8]), .B(B[5]), .Z(\ab[8][5] ) );
    VMW_AND2 U58 ( .A(A[15]), .B(B[0]), .Z(\ab[15][0] ) );
    VMW_AND2 U59 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_AND2 U60 ( .A(A[3]), .B(B[10]), .Z(\ab[3][10] ) );
    VMW_AND2 U61 ( .A(A[6]), .B(B[7]), .Z(\ab[6][7] ) );
    VMW_AND2 U62 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U63 ( .A(A[7]), .B(B[7]), .Z(\ab[7][7] ) );
    VMW_AND2 U64 ( .A(A[8]), .B(B[2]), .Z(\ab[8][2] ) );
    VMW_AND2 U65 ( .A(A[2]), .B(B[11]), .Z(\ab[2][11] ) );
    VMW_AND2 U66 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_AND2 U67 ( .A(A[8]), .B(B[4]), .Z(\ab[8][4] ) );
    VMW_AND2 U68 ( .A(A[0]), .B(B[14]), .Z(\ab[0][14] ) );
    VMW_AND2 U69 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U70 ( .A(A[5]), .B(B[3]), .Z(\ab[5][3] ) );
    VMW_AND2 U71 ( .A(A[11]), .B(B[2]), .Z(\ab[11][2] ) );
    VMW_AND2 U72 ( .A(A[2]), .B(B[9]), .Z(\ab[2][9] ) );
    VMW_AND2 U73 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U74 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_AND2 U75 ( .A(A[3]), .B(B[9]), .Z(\ab[3][9] ) );
    VMW_AND2 U76 ( .A(B[4]), .B(A[9]), .Z(\ab[9][4] ) );
    VMW_AND2 U77 ( .A(A[2]), .B(B[10]), .Z(\ab[2][10] ) );
    VMW_AND2 U78 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
    VMW_AND2 U79 ( .A(A[7]), .B(B[6]), .Z(\ab[7][6] ) );
    VMW_AND2 U80 ( .A(A[10]), .B(B[3]), .Z(\ab[10][3] ) );
    VMW_AND2 U81 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U82 ( .A(A[3]), .B(B[11]), .Z(\ab[3][11] ) );
    VMW_AND2 U83 ( .A(A[6]), .B(B[6]), .Z(\ab[6][6] ) );
    VMW_AND2 U84 ( .A(A[11]), .B(B[3]), .Z(\ab[11][3] ) );
    VMW_AND2 U85 ( .A(A[11]), .B(B[4]), .Z(\ab[11][4] ) );
    VMW_AND2 U86 ( .A(A[3]), .B(B[7]), .Z(\ab[3][7] ) );
    VMW_AND2 U87 ( .A(A[6]), .B(B[1]), .Z(\ab[6][1] ) );
    VMW_AND2 U88 ( .A(A[10]), .B(B[4]), .Z(\ab[10][4] ) );
    VMW_AND2 U89 ( .A(A[2]), .B(B[7]), .Z(\ab[2][7] ) );
    VMW_AND2 U90 ( .A(A[7]), .B(B[1]), .Z(\ab[7][1] ) );
    VMW_AND2 U91 ( .A(A[1]), .B(B[12]), .Z(\ab[1][12] ) );
    VMW_AND2 U92 ( .A(B[3]), .B(A[9]), .Z(\ab[9][3] ) );
    VMW_AND2 U93 ( .A(A[4]), .B(B[4]), .Z(\ab[4][4] ) );
    VMW_AND2 U94 ( .A(A[6]), .B(B[8]), .Z(\ab[6][8] ) );
    VMW_AND2 U95 ( .A(A[13]), .B(B[1]), .Z(\ab[13][1] ) );
    VMW_AND2 U96 ( .A(A[0]), .B(B[13]), .Z(\ab[0][13] ) );
    VMW_AND2 U97 ( .A(A[5]), .B(B[4]), .Z(\ab[5][4] ) );
    VMW_AND2 U98 ( .A(B[8]), .B(A[7]), .Z(\ab[7][8] ) );
    VMW_AND2 U99 ( .A(A[8]), .B(B[3]), .Z(\ab[8][3] ) );
    VMW_AND2 U100 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U101 ( .A(A[2]), .B(B[5]), .Z(\ab[2][5] ) );
    VMW_AND2 U102 ( .A(A[4]), .B(B[10]), .Z(\ab[4][10] ) );
    VMW_AND2 U103 ( .A(A[7]), .B(B[3]), .Z(\ab[7][3] ) );
    VMW_AND2 U104 ( .A(A[10]), .B(B[2]), .Z(\ab[10][2] ) );
    VMW_AND2 U105 ( .A(A[0]), .B(B[9]), .Z(\ab[0][9] ) );
    VMW_AND2 U106 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_AND2 U107 ( .A(A[12]), .B(B[1]), .Z(\ab[12][1] ) );
    VMW_AND2 U108 ( .A(A[3]), .B(B[5]), .Z(\ab[3][5] ) );
    VMW_AND2 U109 ( .A(A[6]), .B(B[3]), .Z(\ab[6][3] ) );
    VMW_AND2 U110 ( .A(A[14]), .B(B[0]), .Z(\ab[14][0] ) );
    VMW_AND2 U111 ( .A(A[1]), .B(B[9]), .Z(\ab[1][9] ) );
    VMW_AND2 U112 ( .A(A[8]), .B(B[1]), .Z(\ab[8][1] ) );
    VMW_AND2 U113 ( .A(A[12]), .B(B[3]), .Z(\ab[12][3] ) );
    VMW_AND2 U114 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_AND2 U115 ( .A(A[0]), .B(B[11]), .Z(\ab[0][11] ) );
    VMW_AND2 U116 ( .A(A[5]), .B(B[6]), .Z(\ab[5][6] ) );
    VMW_AND2 U117 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VMW_AND2 U118 ( .A(A[4]), .B(B[6]), .Z(\ab[4][6] ) );
    VMW_AND2 U119 ( .A(A[1]), .B(B[10]), .Z(\ab[1][10] ) );
    VMW_AND2 U120 ( .A(B[1]), .B(A[9]), .Z(\ab[9][1] ) );
    VMW_AND2 U121 ( .A(A[9]), .B(B[6]), .Z(\ab[9][6] ) );
    VMW_AND2 U122 ( .A(B[15]), .B(A[0]), .Z(\ab[0][15] ) );
    VMW_AND2 U123 ( .A(A[1]), .B(B[7]), .Z(\ab[1][7] ) );
    VMW_AND2 U124 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U125 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U126 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U127 ( .A(A[8]), .B(B[6]), .Z(\ab[8][6] ) );
    VMW_AND2 U128 ( .A(A[6]), .B(B[4]), .Z(\ab[6][4] ) );
    VMW_AND2 U129 ( .A(A[11]), .B(B[1]), .Z(\ab[11][1] ) );
    VMW_AND2 U130 ( .A(A[4]), .B(B[8]), .Z(\ab[4][8] ) );
    VMW_AND2 U131 ( .A(A[7]), .B(B[4]), .Z(\ab[7][4] ) );
    VMW_AND2 U132 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U133 ( .A(A[5]), .B(B[8]), .Z(\ab[5][8] ) );
    VMW_AND2 U134 ( .A(A[2]), .B(B[12]), .Z(\ab[2][12] ) );
    VMW_AND2 U135 ( .A(A[10]), .B(B[1]), .Z(\ab[10][1] ) );
    VMW_AND2 U136 ( .A(B[7]), .B(A[8]), .Z(\ab[8][7] ) );
    VMW_AND2 U137 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U138 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_AND2 U139 ( .A(A[1]), .B(B[6]), .Z(\ab[1][6] ) );
    VMW_AND2 U140 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_AND2 U141 ( .A(B[13]), .B(A[2]), .Z(\ab[2][13] ) );
    VMW_AND2 U142 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_AND2 U143 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_AND2 U144 ( .A(A[5]), .B(B[9]), .Z(\ab[5][9] ) );
    VMW_AND2 U145 ( .A(A[7]), .B(B[5]), .Z(\ab[7][5] ) );
    VMW_AND2 U146 ( .A(B[12]), .B(A[3]), .Z(\ab[3][12] ) );
    VMW_AND2 U147 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_AND2 U148 ( .A(A[6]), .B(B[5]), .Z(\ab[6][5] ) );
    VMW_AND2 U149 ( .A(A[10]), .B(B[0]), .Z(\ab[10][0] ) );
    VMW_AND2 U150 ( .A(A[11]), .B(B[0]), .Z(\ab[11][0] ) );
    VMW_AND2 U151 ( .A(A[12]), .B(B[2]), .Z(\ab[12][2] ) );
    VMW_AND2 U152 ( .A(A[4]), .B(B[9]), .Z(\ab[4][9] ) );
    VMW_AND2 U153 ( .A(B[10]), .B(A[5]), .Z(\ab[5][10] ) );
    VMW_AND2 U154 ( .A(A[3]), .B(B[4]), .Z(\ab[3][4] ) );
    VMW_AND2 U155 ( .A(A[14]), .B(B[1]), .Z(\ab[14][1] ) );
    VMW_AND2 U156 ( .A(A[1]), .B(B[8]), .Z(\ab[1][8] ) );
    VMW_AND2 U157 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U158 ( .A(B[11]), .B(A[4]), .Z(\ab[4][11] ) );
    VMW_AND2 U159 ( .A(A[0]), .B(B[8]), .Z(\ab[0][8] ) );
    VMW_AND2 U160 ( .A(A[7]), .B(B[2]), .Z(\ab[7][2] ) );
    VMW_AND2 U161 ( .A(A[1]), .B(B[11]), .Z(\ab[1][11] ) );
    VMW_AND2 U162 ( .A(B[0]), .B(A[9]), .Z(\ab[9][0] ) );
    VMW_AND2 U163 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_AND2 U164 ( .A(A[4]), .B(B[7]), .Z(\ab[4][7] ) );
    VMW_AND2 U165 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_AND2 U166 ( .A(A[0]), .B(B[10]), .Z(\ab[0][10] ) );
    VMW_AND2 U167 ( .A(A[5]), .B(B[7]), .Z(\ab[5][7] ) );
    VMW_AND2 U168 ( .A(A[8]), .B(B[0]), .Z(\ab[8][0] ) );
    VMW_AND2 U169 ( .A(B[2]), .B(A[9]), .Z(\ab[9][2] ) );
    EdgeAux_DW01_add_30_0 FS ( .A({\A1[29] , UNCONNECTED_1, UNCONNECTED_2, 
        UNCONNECTED_3, UNCONNECTED_4, UNCONNECTED_5, UNCONNECTED_6, 
        UNCONNECTED_7, UNCONNECTED_8, UNCONNECTED_9, UNCONNECTED_10, 
        UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, UNCONNECTED_14, 
        UNCONNECTED_15, \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , 
        \A1[0] }), .B({UNCONNECTED_16, UNCONNECTED_17, UNCONNECTED_18, 
        UNCONNECTED_19, UNCONNECTED_20, UNCONNECTED_21, UNCONNECTED_22, 
        UNCONNECTED_23, UNCONNECTED_24, UNCONNECTED_25, UNCONNECTED_26, 
        UNCONNECTED_27, UNCONNECTED_28, UNCONNECTED_29, UNCONNECTED_30, 
        \A2[14] , \A2[13] , \A2[12] , \A2[11] , \A2[10] , \A2[9] , \A2[8] , 
        \A2[7] , \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , lsb_0}), 
        .CI(lsb_0), .SUM({UNCONNECTED_31, UNCONNECTED_32, UNCONNECTED_33, 
        UNCONNECTED_34, UNCONNECTED_35, UNCONNECTED_36, UNCONNECTED_37, 
        UNCONNECTED_38, UNCONNECTED_39, UNCONNECTED_40, UNCONNECTED_41, 
        UNCONNECTED_42, UNCONNECTED_43, UNCONNECTED_44, UNCONNECTED_45, 
        UNCONNECTED_46, PRODUCT[15], PRODUCT[14], PRODUCT[13], PRODUCT[12], 
        PRODUCT[11], PRODUCT[10], PRODUCT[9], PRODUCT[8], PRODUCT[7], 
        PRODUCT[6], PRODUCT[5], PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S2_7_4 ( .CI(\SUMB[6][5] ), .A(\ab[7][4] ), .B(\CARRYB[6][4] ), 
        .S(\SUMB[7][4] ), .CO(\CARRYB[7][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_FADD S2_5_8 ( .CI(\SUMB[4][9] ), .A(\ab[5][8] ), .B(\CARRYB[4][8] ), 
        .S(\SUMB[5][8] ), .CO(\CARRYB[5][8] ) );
    VMW_FADD S2_12_1 ( .CI(\SUMB[11][2] ), .A(\ab[12][1] ), .B(\CARRYB[11][1] 
        ), .S(\SUMB[12][1] ), .CO(\CARRYB[12][1] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_13_1 ( .CI(\SUMB[12][2] ), .A(\ab[13][1] ), .B(\CARRYB[12][1] 
        ), .S(\SUMB[13][1] ), .CO(\CARRYB[13][1] ) );
    VMW_FADD S2_4_8 ( .CI(\SUMB[3][9] ), .A(\ab[4][8] ), .B(\CARRYB[3][8] ), 
        .S(\SUMB[4][8] ), .CO(\CARRYB[4][8] ) );
    VMW_FADD S2_6_4 ( .CI(\SUMB[5][5] ), .A(\ab[6][4] ), .B(\CARRYB[5][4] ), 
        .S(\SUMB[6][4] ), .CO(\CARRYB[6][4] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_FADD S2_10_4 ( .CI(\SUMB[9][5] ), .A(\ab[10][4] ), .B(\CARRYB[9][4] ), 
        .S(\SUMB[10][4] ), .CO(\CARRYB[10][4] ) );
    VMW_FADD S2_8_6 ( .CI(\SUMB[7][7] ), .A(\ab[8][6] ), .B(\CARRYB[7][6] ), 
        .S(\SUMB[8][6] ), .CO(\CARRYB[8][6] ) );
    VMW_FADD S2_9_6 ( .CI(\SUMB[8][7] ), .A(\ab[9][6] ), .B(\CARRYB[8][6] ), 
        .S(\SUMB[9][6] ) );
    VMW_FADD S2_11_4 ( .CI(\SUMB[10][5] ), .A(\ab[11][4] ), .B(\CARRYB[10][4] 
        ), .S(\SUMB[11][4] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S2_4_6 ( .CI(\SUMB[3][7] ), .A(\ab[4][6] ), .B(\CARRYB[3][6] ), 
        .S(\SUMB[4][6] ), .CO(\CARRYB[4][6] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_FADD S1_10_0 ( .CI(\SUMB[9][1] ), .A(\ab[10][0] ), .B(\CARRYB[9][0] ), 
        .S(\A1[8] ), .CO(\CARRYB[10][0] ) );
    VMW_FADD S2_11_3 ( .CI(\SUMB[10][4] ), .A(\ab[11][3] ), .B(\CARRYB[10][3] 
        ), .S(\SUMB[11][3] ), .CO(\CARRYB[11][3] ) );
    VMW_FADD S2_3_11 ( .CI(\SUMB[2][12] ), .A(\ab[3][11] ), .B(\CARRYB[2][11] 
        ), .S(\SUMB[3][11] ), .CO(\CARRYB[3][11] ) );
    VMW_FADD S2_9_1 ( .CI(\SUMB[8][2] ), .A(\ab[9][1] ), .B(\CARRYB[8][1] ), 
        .S(\SUMB[9][1] ), .CO(\CARRYB[9][1] ) );
    VMW_FADD S1_11_0 ( .CI(\SUMB[10][1] ), .A(\ab[11][0] ), .B(\CARRYB[10][0] 
        ), .S(\A1[9] ), .CO(\CARRYB[11][0] ) );
    VMW_FADD S2_8_1 ( .CI(\SUMB[7][2] ), .A(\ab[8][1] ), .B(\CARRYB[7][1] ), 
        .S(\SUMB[8][1] ), .CO(\CARRYB[8][1] ) );
    VMW_FADD S2_10_3 ( .CI(\SUMB[9][4] ), .A(\ab[10][3] ), .B(\CARRYB[9][3] ), 
        .S(\SUMB[10][3] ), .CO(\CARRYB[10][3] ) );
    VMW_FADD S2_2_10 ( .CI(\SUMB[1][11] ), .A(\ab[2][10] ), .B(\CARRYB[1][10] 
        ), .S(\SUMB[2][10] ), .CO(\CARRYB[2][10] ) );
    VMW_FADD S2_5_6 ( .CI(\SUMB[4][7] ), .A(\ab[5][6] ), .B(\CARRYB[4][6] ), 
        .S(\SUMB[5][6] ), .CO(\CARRYB[5][6] ) );
    VMW_FADD S1_7_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), 
        .S(\A1[5] ), .CO(\CARRYB[7][0] ) );
    VMW_FADD S2_6_3 ( .CI(\SUMB[5][4] ), .A(\ab[6][3] ), .B(\CARRYB[5][3] ), 
        .S(\SUMB[6][3] ), .CO(\CARRYB[6][3] ) );
    VMW_FADD S2_3_5 ( .CI(\SUMB[2][6] ), .A(\ab[3][5] ), .B(\CARRYB[2][5] ), 
        .S(\SUMB[3][5] ), .CO(\CARRYB[3][5] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ), .CO(\CARRYB[2][5] ) );
    VMW_FADD S2_7_3 ( .CI(\SUMB[6][4] ), .A(\ab[7][3] ), .B(\CARRYB[6][3] ), 
        .S(\SUMB[7][3] ), .CO(\CARRYB[7][3] ) );
    VMW_FADD S2_2_11 ( .CI(\SUMB[1][12] ), .A(\ab[2][11] ), .B(\CARRYB[1][11] 
        ), .S(\SUMB[2][11] ), .CO(\CARRYB[2][11] ) );
    VMW_FADD S2_5_7 ( .CI(\SUMB[4][8] ), .A(\ab[5][7] ), .B(\CARRYB[4][7] ), 
        .S(\SUMB[5][7] ), .CO(\CARRYB[5][7] ) );
    VMW_FADD S2_10_2 ( .CI(\SUMB[9][3] ), .A(\ab[10][2] ), .B(\CARRYB[9][2] ), 
        .S(\SUMB[10][2] ), .CO(\CARRYB[10][2] ) );
    VMW_FADD S2_11_2 ( .CI(\SUMB[10][3] ), .A(\ab[11][2] ), .B(\CARRYB[10][2] 
        ), .S(\SUMB[11][2] ), .CO(\CARRYB[11][2] ) );
    VMW_FADD S2_3_10 ( .CI(\SUMB[2][11] ), .A(\ab[3][10] ), .B(\CARRYB[2][10] 
        ), .S(\SUMB[3][10] ), .CO(\CARRYB[3][10] ) );
    VMW_FADD S2_4_7 ( .CI(\SUMB[3][8] ), .A(\ab[4][7] ), .B(\CARRYB[3][7] ), 
        .S(\SUMB[4][7] ), .CO(\CARRYB[4][7] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_FADD S2_7_2 ( .CI(\SUMB[6][3] ), .A(\ab[7][2] ), .B(\CARRYB[6][2] ), 
        .S(\SUMB[7][2] ), .CO(\CARRYB[7][2] ) );
    VMW_FADD S2_6_2 ( .CI(\SUMB[5][3] ), .A(\ab[6][2] ), .B(\CARRYB[5][2] ), 
        .S(\SUMB[6][2] ), .CO(\CARRYB[6][2] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ), .CO(\CARRYB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_FADD S2_6_5 ( .CI(\SUMB[5][6] ), .A(\ab[6][5] ), .B(\CARRYB[5][5] ), 
        .S(\SUMB[6][5] ), .CO(\CARRYB[6][5] ) );
    VMW_FADD S2_4_9 ( .CI(\SUMB[3][10] ), .A(\ab[4][9] ), .B(\CARRYB[3][9] ), 
        .S(\SUMB[4][9] ), .CO(\CARRYB[4][9] ) );
    VMW_FADD S2_7_5 ( .CI(\SUMB[6][6] ), .A(\ab[7][5] ), .B(\CARRYB[6][5] ), 
        .S(\SUMB[7][5] ), .CO(\CARRYB[7][5] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S2_5_9 ( .CI(\SUMB[4][10] ), .A(\ab[5][9] ), .B(\CARRYB[4][9] ), 
        .S(\SUMB[5][9] ), .CO(\CARRYB[5][9] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_FADD S2_10_5 ( .CI(\SUMB[9][6] ), .A(\ab[10][5] ), .B(\CARRYB[9][5] ), 
        .S(\SUMB[10][5] ) );
    VMW_FADD S1_14_0 ( .CI(\SUMB[13][1] ), .A(\ab[14][0] ), .B(\CARRYB[13][0] 
        ), .S(\A1[12] ), .CO(\CARRYB[14][0] ) );
    VMW_FADD S2_8_7 ( .CI(\SUMB[7][8] ), .A(\ab[8][7] ), .B(\CARRYB[7][7] ), 
        .S(\SUMB[8][7] ) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_FADD S2_7_7 ( .CI(\SUMB[6][8] ), .A(\ab[7][7] ), .B(\CARRYB[6][7] ), 
        .S(\SUMB[7][7] ), .CO(\CARRYB[7][7] ) );
    VMW_FADD S2_12_2 ( .CI(\SUMB[11][3] ), .A(\ab[12][2] ), .B(\CARRYB[11][2] 
        ), .S(\SUMB[12][2] ), .CO(\CARRYB[12][2] ) );
    VMW_FADD S2_13_2 ( .CI(\SUMB[12][3] ), .A(\ab[13][2] ), .B(\CARRYB[12][2] 
        ), .S(\SUMB[13][2] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_6_7 ( .CI(\SUMB[5][8] ), .A(\ab[6][7] ), .B(\CARRYB[5][7] ), 
        .S(\SUMB[6][7] ), .CO(\CARRYB[6][7] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ), .CO(\CARRYB[5][2] ) );
    VMW_FADD S2_2_8 ( .CI(\SUMB[1][9] ), .A(\ab[2][8] ), .B(\CARRYB[1][8] ), 
        .S(\SUMB[2][8] ), .CO(\CARRYB[2][8] ) );
    VMW_FADD S2_4_11 ( .CI(\SUMB[3][12] ), .A(\ab[4][11] ), .B(\CARRYB[3][11] 
        ), .S(\SUMB[4][11] ) );
    VMW_FADD S2_8_5 ( .CI(\SUMB[7][6] ), .A(\ab[8][5] ), .B(\CARRYB[7][5] ), 
        .S(\SUMB[8][5] ), .CO(\CARRYB[8][5] ) );
    VMW_FADD S2_9_5 ( .CI(\SUMB[8][6] ), .A(\ab[9][5] ), .B(\CARRYB[8][5] ), 
        .S(\SUMB[9][5] ), .CO(\CARRYB[9][5] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_FADD S2_5_10 ( .CI(\SUMB[4][11] ), .A(\ab[5][10] ), .B(\CARRYB[4][10] 
        ), .S(\SUMB[5][10] ) );
    VMW_FADD S2_14_1 ( .CI(\SUMB[13][2] ), .A(\ab[14][1] ), .B(\CARRYB[13][1] 
        ), .S(\SUMB[14][1] ) );
    VMW_FADD S2_3_8 ( .CI(\SUMB[2][9] ), .A(\ab[3][8] ), .B(\CARRYB[2][8] ), 
        .S(\SUMB[3][8] ), .CO(\CARRYB[3][8] ) );
    VMW_FADD S2_4_5 ( .CI(\SUMB[3][6] ), .A(\ab[4][5] ), .B(\CARRYB[3][5] ), 
        .S(\SUMB[4][5] ), .CO(\CARRYB[4][5] ) );
    VMW_FADD S2_6_9 ( .CI(\SUMB[5][10] ), .A(\ab[6][9] ), .B(\CARRYB[5][9] ), 
        .S(\SUMB[6][9] ) );
    VMW_FADD S2_9_2 ( .CI(\SUMB[8][3] ), .A(\ab[9][2] ), .B(\CARRYB[8][2] ), 
        .S(\SUMB[9][2] ), .CO(\CARRYB[9][2] ) );
    VMW_FADD S2_3_12 ( .CI(\SUMB[2][13] ), .A(\ab[3][12] ), .B(\CARRYB[2][12] 
        ), .S(\SUMB[3][12] ) );
    VMW_FADD S2_8_2 ( .CI(\SUMB[7][3] ), .A(\ab[8][2] ), .B(\CARRYB[7][2] ), 
        .S(\SUMB[8][2] ), .CO(\CARRYB[8][2] ) );
    VMW_FADD S2_5_5 ( .CI(\SUMB[4][6] ), .A(\ab[5][5] ), .B(\CARRYB[4][5] ), 
        .S(\SUMB[5][5] ), .CO(\CARRYB[5][5] ) );
    VMW_FADD S2_2_13 ( .CI(\SUMB[1][14] ), .A(\ab[2][13] ), .B(\CARRYB[1][13] 
        ), .S(\SUMB[2][13] ) );
    VMW_FADD S2_3_6 ( .CI(\SUMB[2][7] ), .A(\ab[3][6] ), .B(\CARRYB[2][6] ), 
        .S(\SUMB[3][6] ), .CO(\CARRYB[3][6] ) );
    VMW_FADD S2_2_6 ( .CI(\SUMB[1][7] ), .A(\ab[2][6] ), .B(\CARRYB[1][6] ), 
        .S(\SUMB[2][6] ), .CO(\CARRYB[2][6] ) );
    VMW_FADD S2_5_4 ( .CI(\SUMB[4][5] ), .A(\ab[5][4] ), .B(\CARRYB[4][4] ), 
        .S(\SUMB[5][4] ), .CO(\CARRYB[5][4] ) );
    VMW_FADD S2_2_12 ( .CI(\SUMB[1][13] ), .A(\ab[2][12] ), .B(\CARRYB[1][12] 
        ), .S(\SUMB[2][12] ), .CO(\CARRYB[2][12] ) );
    VMW_FADD S2_7_8 ( .CI(\SUMB[6][9] ), .A(\ab[7][8] ), .B(\CARRYB[6][8] ), 
        .S(\SUMB[7][8] ) );
    VMW_FADD S2_8_3 ( .CI(\SUMB[7][4] ), .A(\ab[8][3] ), .B(\CARRYB[7][3] ), 
        .S(\SUMB[8][3] ), .CO(\CARRYB[8][3] ) );
    VMW_FADD S2_10_1 ( .CI(\SUMB[9][2] ), .A(\ab[10][1] ), .B(\CARRYB[9][1] ), 
        .S(\SUMB[10][1] ), .CO(\CARRYB[10][1] ) );
    VMW_FADD S2_9_3 ( .CI(\SUMB[8][4] ), .A(\ab[9][3] ), .B(\CARRYB[8][3] ), 
        .S(\SUMB[9][3] ), .CO(\CARRYB[9][3] ) );
    VMW_FADD S2_11_1 ( .CI(\SUMB[10][2] ), .A(\ab[11][1] ), .B(\CARRYB[10][1] 
        ), .S(\SUMB[11][1] ), .CO(\CARRYB[11][1] ) );
    VMW_FADD S2_4_4 ( .CI(\SUMB[3][5] ), .A(\ab[4][4] ), .B(\CARRYB[3][4] ), 
        .S(\SUMB[4][4] ), .CO(\CARRYB[4][4] ) );
    VMW_FADD S2_6_8 ( .CI(\SUMB[5][9] ), .A(\ab[6][8] ), .B(\CARRYB[5][8] ), 
        .S(\SUMB[6][8] ), .CO(\CARRYB[6][8] ) );
    VMW_FADD S2_7_1 ( .CI(\SUMB[6][2] ), .A(\ab[7][1] ), .B(\CARRYB[6][1] ), 
        .S(\SUMB[7][1] ), .CO(\CARRYB[7][1] ) );
    VMW_FADD S2_2_7 ( .CI(\SUMB[1][8] ), .A(\ab[2][7] ), .B(\CARRYB[1][7] ), 
        .S(\SUMB[2][7] ), .CO(\CARRYB[2][7] ) );
    VMW_FADD S1_8_0 ( .CI(\SUMB[7][1] ), .A(\ab[8][0] ), .B(\CARRYB[7][0] ), 
        .S(\A1[6] ), .CO(\CARRYB[8][0] ) );
    VMW_FADD S1_9_0 ( .CI(\SUMB[8][1] ), .A(\ab[9][0] ), .B(\CARRYB[8][0] ), 
        .S(\A1[7] ), .CO(\CARRYB[9][0] ) );
    VMW_FADD S2_3_7 ( .CI(\SUMB[2][8] ), .A(\ab[3][7] ), .B(\CARRYB[2][7] ), 
        .S(\SUMB[3][7] ), .CO(\CARRYB[3][7] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ), .CO(\CARRYB[6][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_6 ( .CI(\SUMB[5][7] ), .A(\ab[6][6] ), .B(\CARRYB[5][6] ), 
        .S(\SUMB[6][6] ), .CO(\CARRYB[6][6] ) );
    VMW_FADD S1_12_0 ( .CI(\SUMB[11][1] ), .A(\ab[12][0] ), .B(\CARRYB[11][0] 
        ), .S(\A1[10] ), .CO(\CARRYB[12][0] ) );
    VMW_FADD S4_0 ( .CI(\SUMB[14][1] ), .A(\ab[15][0] ), .B(\CARRYB[14][0] ), 
        .S(\A1[13] ) );
    VMW_FADD S2_12_3 ( .CI(\SUMB[11][4] ), .A(\ab[12][3] ), .B(\CARRYB[11][3] 
        ), .S(\SUMB[12][3] ) );
    VMW_FADD S1_13_0 ( .CI(\SUMB[12][1] ), .A(\ab[13][0] ), .B(\CARRYB[12][0] 
        ), .S(\A1[11] ), .CO(\CARRYB[13][0] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_FADD S2_7_6 ( .CI(\SUMB[6][7] ), .A(\ab[7][6] ), .B(\CARRYB[6][6] ), 
        .S(\SUMB[7][6] ), .CO(\CARRYB[7][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ), .CO(\CARRYB[4][3] ) );
    VMW_FADD S2_3_9 ( .CI(\SUMB[2][10] ), .A(\ab[3][9] ), .B(\CARRYB[2][9] ), 
        .S(\SUMB[3][9] ), .CO(\CARRYB[3][9] ) );
    VMW_FADD S2_9_4 ( .CI(\SUMB[8][5] ), .A(\ab[9][4] ), .B(\CARRYB[8][4] ), 
        .S(\SUMB[9][4] ), .CO(\CARRYB[9][4] ) );
    VMW_FADD S2_4_10 ( .CI(\SUMB[3][11] ), .A(\ab[4][10] ), .B(\CARRYB[3][10] 
        ), .S(\SUMB[4][10] ), .CO(\CARRYB[4][10] ) );
    VMW_FADD S2_8_4 ( .CI(\SUMB[7][5] ), .A(\ab[8][4] ), .B(\CARRYB[7][4] ), 
        .S(\SUMB[8][4] ), .CO(\CARRYB[8][4] ) );
    VMW_FADD S2_5_3 ( .CI(\SUMB[4][4] ), .A(\ab[5][3] ), .B(\CARRYB[4][3] ), 
        .S(\SUMB[5][3] ), .CO(\CARRYB[5][3] ) );
    VMW_FADD S2_2_9 ( .CI(\SUMB[1][10] ), .A(\ab[2][9] ), .B(\CARRYB[1][9] ), 
        .S(\SUMB[2][9] ), .CO(\CARRYB[2][9] ) );
endmodule


module EdgeAux ( Eid, InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [5:0] Eid;
input  [5:0] WeightAddr;
input  [15:0] InEdge;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire \Weight[11] , \Weight[6] , \Weight[15] , \Weight[2] , \Weight[0] , 
        \Weight[9] , \Weight[13] , \Weight[4] , \Weight[12] , \Weight[5] , 
        \Weight[1] , \Weight[8] , \Weight[14] , \Weight[3] , \Weight[10] , 
        \Weight[7] , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
        n101;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 ;
    VMW_PULLDOWN U15 ( .Z(n101) );
    VMW_AO22 U16 ( .A(\Weight[9] ), .B(n76), .C(WeightData[9]), .D(n77), .Z(
        n91) );
    VMW_AO22 U17 ( .A(\Weight[8] ), .B(n76), .C(WeightData[8]), .D(n77), .Z(
        n92) );
    VMW_AO22 U18 ( .A(\Weight[7] ), .B(n76), .C(WeightData[7]), .D(n77), .Z(
        n93) );
    VMW_AO22 U19 ( .A(\Weight[6] ), .B(n76), .C(WeightData[6]), .D(n77), .Z(
        n94) );
    VMW_AO22 U20 ( .A(\Weight[5] ), .B(n76), .C(WeightData[5]), .D(n77), .Z(
        n95) );
    VMW_AO22 U21 ( .A(\Weight[4] ), .B(n76), .C(WeightData[4]), .D(n77), .Z(
        n96) );
    VMW_AO22 U22 ( .A(\Weight[3] ), .B(n76), .C(WeightData[3]), .D(n77), .Z(
        n97) );
    VMW_AO22 U23 ( .A(\Weight[2] ), .B(n76), .C(WeightData[2]), .D(n77), .Z(
        n98) );
    VMW_AO22 U24 ( .A(\Weight[1] ), .B(n76), .C(WeightData[1]), .D(n77), .Z(
        n99) );
    VMW_AO22 U25 ( .A(\Weight[15] ), .B(n76), .C(WeightData[15]), .D(n77), .Z(
        n85) );
    VMW_AO22 U26 ( .A(\Weight[14] ), .B(n76), .C(WeightData[14]), .D(n77), .Z(
        n86) );
    VMW_AO22 U27 ( .A(\Weight[13] ), .B(n76), .C(WeightData[13]), .D(n77), .Z(
        n87) );
    VMW_AO22 U28 ( .A(\Weight[12] ), .B(n76), .C(WeightData[12]), .D(n77), .Z(
        n88) );
    VMW_AO22 U29 ( .A(\Weight[11] ), .B(n76), .C(WeightData[11]), .D(n77), .Z(
        n89) );
    VMW_AO22 U30 ( .A(\Weight[10] ), .B(n76), .C(WeightData[10]), .D(n77), .Z(
        n90) );
    VMW_AO22 U31 ( .A(\Weight[0] ), .B(n76), .C(WeightData[0]), .D(n77), .Z(
        n100) );
    VMW_AND3 U32 ( .A(n79), .B(n80), .C(n81), .Z(n78) );
    VMW_AND4 U33 ( .A(n82), .B(n83), .C(n84), .D(n78), .Z(n77) );
    VMW_XNOR2 U34 ( .A(WeightAddr[5]), .B(Eid[5]), .Z(n80) );
    VMW_XNOR2 U35 ( .A(WeightAddr[2]), .B(Eid[2]), .Z(n79) );
    VMW_XNOR2 U36 ( .A(WeightAddr[3]), .B(Eid[3]), .Z(n81) );
    VMW_XNOR2 U37 ( .A(WeightAddr[0]), .B(Eid[0]), .Z(n83) );
    VMW_XNOR2 U38 ( .A(WeightAddr[4]), .B(Eid[4]), .Z(n82) );
    VMW_XNOR2 U39 ( .A(WeightAddr[1]), .B(Eid[1]), .Z(n84) );
    VMW_INV U40 ( .A(n77), .Z(n76) );
    VMW_FD \Weight_reg[15]  ( .D(n85), .CP(Clk), .Q(\Weight[15] ) );
    VMW_FD \Weight_reg[14]  ( .D(n86), .CP(Clk), .Q(\Weight[14] ) );
    VMW_FD \Weight_reg[13]  ( .D(n87), .CP(Clk), .Q(\Weight[13] ) );
    VMW_FD \Weight_reg[12]  ( .D(n88), .CP(Clk), .Q(\Weight[12] ) );
    VMW_FD \Weight_reg[11]  ( .D(n89), .CP(Clk), .Q(\Weight[11] ) );
    VMW_FD \Weight_reg[10]  ( .D(n90), .CP(Clk), .Q(\Weight[10] ) );
    VMW_FD \Weight_reg[9]  ( .D(n91), .CP(Clk), .Q(\Weight[9] ) );
    VMW_FD \Weight_reg[8]  ( .D(n92), .CP(Clk), .Q(\Weight[8] ) );
    VMW_FD \Weight_reg[7]  ( .D(n93), .CP(Clk), .Q(\Weight[7] ) );
    VMW_FD \Weight_reg[6]  ( .D(n94), .CP(Clk), .Q(\Weight[6] ) );
    VMW_FD \Weight_reg[5]  ( .D(n95), .CP(Clk), .Q(\Weight[5] ) );
    VMW_FD \Weight_reg[4]  ( .D(n96), .CP(Clk), .Q(\Weight[4] ) );
    VMW_FD \Weight_reg[3]  ( .D(n97), .CP(Clk), .Q(\Weight[3] ) );
    VMW_FD \Weight_reg[2]  ( .D(n98), .CP(Clk), .Q(\Weight[2] ) );
    VMW_FD \Weight_reg[1]  ( .D(n99), .CP(Clk), .Q(\Weight[1] ) );
    VMW_FD \Weight_reg[0]  ( .D(n100), .CP(Clk), .Q(\Weight[0] ) );
    EdgeAux_DW02_mult_16_16_0 mul_92 ( .A({\Weight[15] , \Weight[14] , 
        \Weight[13] , \Weight[12] , \Weight[11] , \Weight[10] , \Weight[9] , 
        \Weight[8] , \Weight[7] , \Weight[6] , \Weight[5] , \Weight[4] , 
        \Weight[3] , \Weight[2] , \Weight[1] , \Weight[0] }), .B(InEdge), .TC(
        n101), .PRODUCT({UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, 
        UNCONNECTED_4, UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, 
        UNCONNECTED_8, UNCONNECTED_9, UNCONNECTED_10, UNCONNECTED_11, 
        UNCONNECTED_12, UNCONNECTED_13, UNCONNECTED_14, UNCONNECTED_15, 
        UNCONNECTED_16, OutEdge[15], OutEdge[14], OutEdge[13], OutEdge[12], 
        OutEdge[11], OutEdge[10], OutEdge[9], OutEdge[8], OutEdge[7], 
        OutEdge[6], OutEdge[5], OutEdge[4], OutEdge[3], OutEdge[2], OutEdge[1], 
        OutEdge[0]}) );
endmodule


module NodeAux_INDEGREE1_SOURCE1_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE1_SOURCE1 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [3:0] Nid;
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , n82, \OutEdge96[11] , \OutEdge96[5] , 
        \OutEdge96[15] , \OutEdge96[8] , \OutEdge96[1] , \OutEdge96[3] , 
        \OutEdge96[7] , \OutEdge96[13] , \OutEdge96[6] , \OutEdge96[12] , 
        \OutEdge96[2] , \OutEdge96[9] , \OutEdge96[14] , \OutEdge96[0] , 
        \OutEdge96[10] , \OutEdge96[4] , \path[1] , n267, n268, n269, n270, 
        n271, n272, n273, n274, n275, n276, n277, n278;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U46 ( .Z(n278) );
    VMW_AO22 U47 ( .A(OutEdge[15]), .B(n267), .C(InEdges[15]), .D(n268), .Z(
        \OutEdge96[15] ) );
    VMW_AO22 U48 ( .A(OutEdge[14]), .B(n267), .C(InEdges[14]), .D(n268), .Z(
        \OutEdge96[14] ) );
    VMW_AO22 U49 ( .A(OutEdge[13]), .B(n267), .C(InEdges[13]), .D(n268), .Z(
        \OutEdge96[13] ) );
    VMW_AO22 U50 ( .A(OutEdge[12]), .B(n267), .C(InEdges[12]), .D(n268), .Z(
        \OutEdge96[12] ) );
    VMW_AO22 U51 ( .A(OutEdge[11]), .B(n267), .C(InEdges[11]), .D(n268), .Z(
        \OutEdge96[11] ) );
    VMW_AO22 U52 ( .A(OutEdge[10]), .B(n267), .C(InEdges[10]), .D(n268), .Z(
        \OutEdge96[10] ) );
    VMW_AO22 U53 ( .A(OutEdge[9]), .B(n267), .C(InEdges[9]), .D(n268), .Z(
        \OutEdge96[9] ) );
    VMW_AO22 U54 ( .A(OutEdge[8]), .B(n267), .C(InEdges[8]), .D(n268), .Z(
        \OutEdge96[8] ) );
    VMW_AO22 U55 ( .A(OutEdge[7]), .B(n267), .C(InEdges[7]), .D(n268), .Z(
        \OutEdge96[7] ) );
    VMW_AO22 U56 ( .A(OutEdge[6]), .B(n267), .C(InEdges[6]), .D(n268), .Z(
        \OutEdge96[6] ) );
    VMW_AO22 U57 ( .A(OutEdge[5]), .B(n267), .C(InEdges[5]), .D(n268), .Z(
        \OutEdge96[5] ) );
    VMW_AO22 U58 ( .A(OutEdge[4]), .B(n267), .C(InEdges[4]), .D(n268), .Z(
        \OutEdge96[4] ) );
    VMW_AO22 U59 ( .A(OutEdge[3]), .B(n267), .C(InEdges[3]), .D(n268), .Z(
        \OutEdge96[3] ) );
    VMW_AO22 U60 ( .A(OutEdge[2]), .B(n267), .C(InEdges[2]), .D(n268), .Z(
        \OutEdge96[2] ) );
    VMW_AO22 U61 ( .A(OutEdge[1]), .B(n267), .C(InEdges[1]), .D(n268), .Z(
        \OutEdge96[1] ) );
    VMW_AO22 U62 ( .A(OutEdge[0]), .B(n267), .C(InEdges[0]), .D(n268), .Z(
        \OutEdge96[0] ) );
    VMW_AO21 U63 ( .A(Start), .B(\path[1] ), .C(n267), .Z(n277) );
    VMW_AO21 U64 ( .A(\path[2] ), .B(Start), .C(n267), .Z(n276) );
    VMW_AO21 U65 ( .A(Start), .B(\path[0] ), .C(n267), .Z(n275) );
    VMW_NOR2 U66 ( .A(n269), .B(Start), .Z(n268) );
    VMW_NOR2 U67 ( .A(Start), .B(n82), .Z(n267) );
    VMW_AND4 U68 ( .A(n270), .B(n271), .C(n272), .D(n273), .Z(n274) );
    VMW_XNOR2 U69 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n273) );
    VMW_XNOR2 U70 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n272) );
    VMW_XNOR2 U71 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n271) );
    VMW_XNOR2 U72 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n270) );
    VMW_INV U73 ( .A(n82), .Z(n269) );
    VMW_BUFIZ U74 ( .A(\path[1] ), .E(n274), .Z(\PathData[1] ) );
    VMW_BUFIZ U75 ( .A(\path[0] ), .E(n274), .Z(\PathData[0] ) );
    VMW_BUFIZ U76 ( .A(\path[2] ), .E(n274), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n275), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n276), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n277), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge96[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge96[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge96[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge96[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge96[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge96[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge96[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge96[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge96[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge96[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge96[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge96[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge96[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge96[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge96[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge96[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE1_SOURCE1_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges), 
        .LEQ(n278), .TC(n278), .GE_GT(n82) );
endmodule


module NodeAux_INDEGREE1_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE1_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [3:0] Nid;
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , n82, \OutEdge96[11] , \OutEdge96[5] , 
        \OutEdge96[15] , \OutEdge96[8] , \OutEdge96[1] , \OutEdge96[3] , 
        \OutEdge96[7] , \OutEdge96[13] , \OutEdge96[6] , \OutEdge96[12] , 
        \OutEdge96[2] , \OutEdge96[9] , \OutEdge96[14] , \OutEdge96[0] , 
        \OutEdge96[10] , \OutEdge96[4] , \path[1] , n267, n268, n269, n270, 
        n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
        n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U46 ( .Z(n293) );
    VMW_AO22 U47 ( .A(OutEdge[15]), .B(n267), .C(n268), .D(InEdges[15]), .Z(
        \OutEdge96[15] ) );
    VMW_OR2 U48 ( .A(n269), .B(Start), .Z(\OutEdge96[14] ) );
    VMW_OR2 U49 ( .A(n270), .B(Start), .Z(\OutEdge96[13] ) );
    VMW_OR2 U50 ( .A(n271), .B(Start), .Z(\OutEdge96[12] ) );
    VMW_OR2 U51 ( .A(n272), .B(Start), .Z(\OutEdge96[11] ) );
    VMW_OR2 U52 ( .A(n273), .B(Start), .Z(\OutEdge96[10] ) );
    VMW_OR2 U53 ( .A(n274), .B(Start), .Z(\OutEdge96[9] ) );
    VMW_OR2 U54 ( .A(n275), .B(Start), .Z(\OutEdge96[8] ) );
    VMW_OR2 U55 ( .A(n276), .B(Start), .Z(\OutEdge96[7] ) );
    VMW_OR2 U56 ( .A(n277), .B(Start), .Z(\OutEdge96[6] ) );
    VMW_OR2 U57 ( .A(n278), .B(Start), .Z(\OutEdge96[5] ) );
    VMW_OR2 U58 ( .A(n279), .B(Start), .Z(\OutEdge96[4] ) );
    VMW_OR2 U59 ( .A(n280), .B(Start), .Z(\OutEdge96[3] ) );
    VMW_OR2 U60 ( .A(n281), .B(Start), .Z(\OutEdge96[2] ) );
    VMW_OR2 U61 ( .A(n282), .B(Start), .Z(\OutEdge96[1] ) );
    VMW_OR2 U62 ( .A(n283), .B(Start), .Z(\OutEdge96[0] ) );
    VMW_AO21 U63 ( .A(\path[1] ), .B(Start), .C(n267), .Z(n292) );
    VMW_AO21 U64 ( .A(Start), .B(\path[2] ), .C(n267), .Z(n291) );
    VMW_AO21 U65 ( .A(\path[0] ), .B(Start), .C(n267), .Z(n290) );
    VMW_INV U66 ( .A(n82), .Z(n284) );
    VMW_NOR2 U67 ( .A(Start), .B(n82), .Z(n267) );
    VMW_NOR2 U68 ( .A(Start), .B(n284), .Z(n268) );
    VMW_AND4 U69 ( .A(n285), .B(n286), .C(n287), .D(n288), .Z(n289) );
    VMW_XNOR2 U70 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n288) );
    VMW_XNOR2 U71 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n287) );
    VMW_XNOR2 U72 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n286) );
    VMW_XNOR2 U73 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n285) );
    VMW_AO22 U74 ( .A(InEdges[9]), .B(n82), .C(OutEdge[9]), .D(n284), .Z(n274)
         );
    VMW_AO22 U75 ( .A(InEdges[8]), .B(n82), .C(OutEdge[8]), .D(n284), .Z(n275)
         );
    VMW_AO22 U76 ( .A(InEdges[7]), .B(n82), .C(OutEdge[7]), .D(n284), .Z(n276)
         );
    VMW_AO22 U77 ( .A(InEdges[6]), .B(n82), .C(OutEdge[6]), .D(n284), .Z(n277)
         );
    VMW_AO22 U78 ( .A(InEdges[5]), .B(n82), .C(OutEdge[5]), .D(n284), .Z(n278)
         );
    VMW_AO22 U79 ( .A(InEdges[4]), .B(n82), .C(OutEdge[4]), .D(n284), .Z(n279)
         );
    VMW_AO22 U80 ( .A(InEdges[3]), .B(n82), .C(OutEdge[3]), .D(n284), .Z(n280)
         );
    VMW_AO22 U81 ( .A(InEdges[2]), .B(n82), .C(OutEdge[2]), .D(n284), .Z(n281)
         );
    VMW_AO22 U82 ( .A(InEdges[1]), .B(n82), .C(OutEdge[1]), .D(n284), .Z(n282)
         );
    VMW_AO22 U83 ( .A(InEdges[14]), .B(n82), .C(OutEdge[14]), .D(n284), .Z(
        n269) );
    VMW_AO22 U84 ( .A(InEdges[13]), .B(n82), .C(OutEdge[13]), .D(n284), .Z(
        n270) );
    VMW_AO22 U85 ( .A(InEdges[12]), .B(n82), .C(OutEdge[12]), .D(n284), .Z(
        n271) );
    VMW_AO22 U86 ( .A(InEdges[11]), .B(n82), .C(OutEdge[11]), .D(n284), .Z(
        n272) );
    VMW_AO22 U87 ( .A(InEdges[10]), .B(n82), .C(OutEdge[10]), .D(n284), .Z(
        n273) );
    VMW_AO22 U88 ( .A(InEdges[0]), .B(n82), .C(OutEdge[0]), .D(n284), .Z(n283)
         );
    VMW_BUFIZ U89 ( .A(\path[1] ), .E(n289), .Z(\PathData[1] ) );
    VMW_BUFIZ U90 ( .A(\path[0] ), .E(n289), .Z(\PathData[0] ) );
    VMW_BUFIZ U91 ( .A(\path[2] ), .E(n289), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n290), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n291), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n292), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge96[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge96[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge96[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge96[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge96[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge96[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge96[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge96[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge96[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge96[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge96[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge96[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge96[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge96[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge96[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge96[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE1_SOURCE0_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges), 
        .LEQ(n293), .TC(n293), .GE_GT(n82) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n85) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n85), .D(n82), .Z(n86) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n86), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n93) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n93), .D(n90), .Z(n94) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n94), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n96), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n102), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n112) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n112), .D(n110), .Z(n113) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n114), .C(n113), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n114) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE2_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [3:0] Nid;
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp180[1] , \temp180[8] , \OutEdge106[5] , \temp180[5] , 
        \OutEdge106[8] , \OutEdge106[1] , \path[2] , \path[0] , 
        \OutEdge106[3] , \temp180[7] , \OutEdge106[7] , \temp180[3] , 
        \OutEdge106[13] , \temp180[12] , \temp180[10] , \OutEdge106[11] , 
        \OutEdge106[15] , \temp180[14] , n84, \OutEdge106[14] , \temp180[15] , 
        \temp180[11] , \OutEdge106[10] , \OutEdge106[12] , \temp180[13] , 
        \OutEdge106[6] , \temp180[2] , \path[1] , n92, \OutEdge106[2] , 
        \temp180[6] , \temp180[4] , \OutEdge106[9] , \OutEdge106[0] , 
        \temp180[0] , \temp180[9] , \OutEdge106[4] , n367, n368, n369, n370, 
        n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
        n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
        n395, n396, n397;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U55 ( .Z(n396) );
    VMW_PULLDOWN U56 ( .Z(n397) );
    VMW_NOR2 U57 ( .A(Start), .B(n367), .Z(\OutEdge106[15] ) );
    VMW_NAND2 U58 ( .A(n368), .B(n369), .Z(\OutEdge106[14] ) );
    VMW_NAND2 U59 ( .A(n370), .B(n369), .Z(\OutEdge106[13] ) );
    VMW_NAND2 U60 ( .A(n371), .B(n369), .Z(\OutEdge106[12] ) );
    VMW_NAND2 U61 ( .A(n372), .B(n369), .Z(\OutEdge106[11] ) );
    VMW_NAND2 U62 ( .A(n373), .B(n369), .Z(\OutEdge106[10] ) );
    VMW_NAND2 U63 ( .A(n374), .B(n369), .Z(\OutEdge106[9] ) );
    VMW_NAND2 U64 ( .A(n375), .B(n369), .Z(\OutEdge106[8] ) );
    VMW_NAND2 U65 ( .A(n376), .B(n369), .Z(\OutEdge106[7] ) );
    VMW_NAND2 U66 ( .A(n377), .B(n369), .Z(\OutEdge106[6] ) );
    VMW_NAND2 U67 ( .A(n378), .B(n369), .Z(\OutEdge106[5] ) );
    VMW_NAND2 U68 ( .A(n379), .B(n369), .Z(\OutEdge106[4] ) );
    VMW_NAND2 U69 ( .A(n380), .B(n369), .Z(\OutEdge106[3] ) );
    VMW_NAND2 U70 ( .A(n381), .B(n369), .Z(\OutEdge106[2] ) );
    VMW_NAND2 U71 ( .A(n382), .B(n369), .Z(\OutEdge106[1] ) );
    VMW_NAND2 U72 ( .A(n383), .B(n369), .Z(\OutEdge106[0] ) );
    VMW_AO21 U73 ( .A(Start), .B(\path[1] ), .C(n384), .Z(n395) );
    VMW_AO21 U74 ( .A(\path[2] ), .B(Start), .C(n384), .Z(n394) );
    VMW_OR2 U75 ( .A(n386), .B(n92), .Z(n385) );
    VMW_AO22 U76 ( .A(OutEdge[15]), .B(n386), .C(InEdges[15]), .D(n84), .Z(
        \temp180[15] ) );
    VMW_OAI22 U77 ( .A(\path[0] ), .B(n369), .C(n385), .D(Start), .Z(n387) );
    VMW_MUX2I U78 ( .A(\temp180[15] ), .B(InEdges[31]), .S(n92), .Z(n367) );
    VMW_NOR3 U79 ( .A(Start), .B(n84), .C(n92), .Z(n384) );
    VMW_AND4 U80 ( .A(n388), .B(n389), .C(n390), .D(n391), .Z(n392) );
    VMW_XNOR2 U81 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n391) );
    VMW_XNOR2 U82 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n390) );
    VMW_XNOR2 U83 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n389) );
    VMW_XNOR2 U84 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n388) );
    VMW_AO22 U85 ( .A(OutEdge[9]), .B(n386), .C(InEdges[9]), .D(n84), .Z(
        \temp180[9] ) );
    VMW_AO22 U86 ( .A(OutEdge[8]), .B(n386), .C(InEdges[8]), .D(n84), .Z(
        \temp180[8] ) );
    VMW_AO22 U87 ( .A(OutEdge[7]), .B(n386), .C(InEdges[7]), .D(n84), .Z(
        \temp180[7] ) );
    VMW_AO22 U88 ( .A(OutEdge[6]), .B(n386), .C(InEdges[6]), .D(n84), .Z(
        \temp180[6] ) );
    VMW_AO22 U89 ( .A(OutEdge[5]), .B(n386), .C(InEdges[5]), .D(n84), .Z(
        \temp180[5] ) );
    VMW_AO22 U90 ( .A(OutEdge[4]), .B(n386), .C(InEdges[4]), .D(n84), .Z(
        \temp180[4] ) );
    VMW_AO22 U91 ( .A(OutEdge[3]), .B(n386), .C(InEdges[3]), .D(n84), .Z(
        \temp180[3] ) );
    VMW_AO22 U92 ( .A(OutEdge[2]), .B(n386), .C(InEdges[2]), .D(n84), .Z(
        \temp180[2] ) );
    VMW_AO22 U93 ( .A(OutEdge[1]), .B(n386), .C(InEdges[1]), .D(n84), .Z(
        \temp180[1] ) );
    VMW_AO22 U94 ( .A(OutEdge[14]), .B(n386), .C(InEdges[14]), .D(n84), .Z(
        \temp180[14] ) );
    VMW_AO22 U95 ( .A(OutEdge[13]), .B(n386), .C(InEdges[13]), .D(n84), .Z(
        \temp180[13] ) );
    VMW_AO22 U96 ( .A(OutEdge[12]), .B(n386), .C(InEdges[12]), .D(n84), .Z(
        \temp180[12] ) );
    VMW_AO22 U97 ( .A(OutEdge[11]), .B(n386), .C(InEdges[11]), .D(n84), .Z(
        \temp180[11] ) );
    VMW_AO22 U98 ( .A(OutEdge[10]), .B(n386), .C(InEdges[10]), .D(n84), .Z(
        \temp180[10] ) );
    VMW_AO22 U99 ( .A(OutEdge[0]), .B(n386), .C(InEdges[0]), .D(n84), .Z(
        \temp180[0] ) );
    VMW_MUX2I U100 ( .A(\temp180[9] ), .B(InEdges[25]), .S(n92), .Z(n374) );
    VMW_MUX2I U101 ( .A(\temp180[8] ), .B(InEdges[24]), .S(n92), .Z(n375) );
    VMW_MUX2I U102 ( .A(\temp180[7] ), .B(InEdges[23]), .S(n92), .Z(n376) );
    VMW_MUX2I U103 ( .A(\temp180[6] ), .B(InEdges[22]), .S(n92), .Z(n377) );
    VMW_MUX2I U104 ( .A(\temp180[5] ), .B(InEdges[21]), .S(n92), .Z(n378) );
    VMW_MUX2I U105 ( .A(\temp180[4] ), .B(InEdges[20]), .S(n92), .Z(n379) );
    VMW_MUX2I U106 ( .A(\temp180[3] ), .B(InEdges[19]), .S(n92), .Z(n380) );
    VMW_MUX2I U107 ( .A(\temp180[2] ), .B(InEdges[18]), .S(n92), .Z(n381) );
    VMW_MUX2I U108 ( .A(\temp180[1] ), .B(InEdges[17]), .S(n92), .Z(n382) );
    VMW_MUX2I U109 ( .A(\temp180[14] ), .B(InEdges[30]), .S(n92), .Z(n368) );
    VMW_MUX2I U110 ( .A(\temp180[13] ), .B(InEdges[29]), .S(n92), .Z(n370) );
    VMW_MUX2I U111 ( .A(\temp180[12] ), .B(InEdges[28]), .S(n92), .Z(n371) );
    VMW_MUX2I U112 ( .A(\temp180[11] ), .B(InEdges[27]), .S(n92), .Z(n372) );
    VMW_MUX2I U113 ( .A(\temp180[10] ), .B(InEdges[26]), .S(n92), .Z(n373) );
    VMW_MUX2I U114 ( .A(\temp180[0] ), .B(InEdges[16]), .S(n92), .Z(n383) );
    VMW_INV U115 ( .A(n84), .Z(n386) );
    VMW_INV U116 ( .A(Start), .Z(n369) );
    VMW_INV U117 ( .A(n387), .Z(n393) );
    VMW_BUFIZ U118 ( .A(\path[1] ), .E(n392), .Z(\PathData[1] ) );
    VMW_BUFIZ U119 ( .A(\path[0] ), .E(n392), .Z(\PathData[0] ) );
    VMW_BUFIZ U120 ( .A(\path[2] ), .E(n392), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n393), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n394), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n395), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge106[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge106[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge106[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge106[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge106[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge106[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge106[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge106[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge106[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge106[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge106[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge106[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge106[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge106[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge106[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge106[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n397), .TC(n397), .GE_GT(n84) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 lte_55_1 ( .A({\temp180[15] , 
        \temp180[14] , \temp180[13] , \temp180[12] , \temp180[11] , 
        \temp180[10] , \temp180[9] , \temp180[8] , \temp180[7] , \temp180[6] , 
        \temp180[5] , \temp180[4] , \temp180[3] , \temp180[2] , \temp180[1] , 
        \temp180[0] }), .B(InEdges[31:16]), .LEQ(n396), .TC(n396), .GE_GT(n92)
         );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, 
        n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, n107, 
        n108, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n104), .B(B[12]), .Z(n103) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n96), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n104), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n103), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n104) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
        n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
        n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
        n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
        n163, n164;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n119), .B(B[2]), .Z(n118) );
    VMW_AO22 U5 ( .A(n121), .B(B[0]), .C(n122), .D(B[1]), .Z(n120) );
    VMW_OR2 U6 ( .A(B[2]), .B(n119), .Z(n123) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n122), .C(n123), .D(n120), .Z(n124) );
    VMW_NAND2 U8 ( .A(n126), .B(B[4]), .Z(n125) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n128), .C(n124), .D(n118), .Z(n127) );
    VMW_OR2 U10 ( .A(B[4]), .B(n126), .Z(n129) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n131), .C(n129), .D(n127), .Z(n130) );
    VMW_NAND2 U12 ( .A(n133), .B(B[6]), .Z(n132) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n135), .C(n130), .D(n125), .Z(n134) );
    VMW_OR2 U14 ( .A(B[6]), .B(n133), .Z(n136) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n138), .C(n136), .D(n134), .Z(n137) );
    VMW_NAND2 U16 ( .A(n140), .B(B[8]), .Z(n139) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n142), .C(n137), .D(n132), .Z(n141) );
    VMW_OR2 U18 ( .A(B[8]), .B(n140), .Z(n143) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n145), .C(n143), .D(n141), .Z(n144) );
    VMW_NAND2 U20 ( .A(n147), .B(B[10]), .Z(n146) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n149), .C(n144), .D(n139), .Z(n148) );
    VMW_NAND2 U22 ( .A(n149), .B(A[9]), .Z(n150) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n147), .C(n150), .D(n148), .Z(n151) );
    VMW_NAND2 U24 ( .A(n153), .B(B[12]), .Z(n152) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n155), .C(n151), .D(n146), .Z(n154) );
    VMW_NAND2 U26 ( .A(n155), .B(A[11]), .Z(n156) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n153), .C(n156), .D(n154), .Z(n157) );
    VMW_NAND2 U28 ( .A(n159), .B(B[14]), .Z(n158) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n161), .C(n157), .D(n152), .Z(n160) );
    VMW_NAND2 U30 ( .A(n161), .B(A[13]), .Z(n162) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n159), .C(n162), .D(n160), .Z(n163) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n164), .C(n163), .D(n158), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n153) );
    VMW_INV U34 ( .A(B[7]), .Z(n142) );
    VMW_INV U35 ( .A(A[7]), .Z(n145) );
    VMW_INV U36 ( .A(A[3]), .Z(n131) );
    VMW_INV U37 ( .A(B[3]), .Z(n128) );
    VMW_INV U38 ( .A(A[10]), .Z(n147) );
    VMW_INV U39 ( .A(B[9]), .Z(n149) );
    VMW_INV U40 ( .A(A[4]), .Z(n126) );
    VMW_INV U41 ( .A(A[8]), .Z(n140) );
    VMW_INV U42 ( .A(A[14]), .Z(n159) );
    VMW_INV U43 ( .A(B[11]), .Z(n155) );
    VMW_INV U44 ( .A(A[5]), .Z(n138) );
    VMW_INV U45 ( .A(B[5]), .Z(n135) );
    VMW_INV U46 ( .A(A[1]), .Z(n122) );
    VMW_INV U47 ( .A(B[15]), .Z(n164) );
    VMW_INV U48 ( .A(B[13]), .Z(n161) );
    VMW_INV U49 ( .A(A[6]), .Z(n133) );
    VMW_INV U50 ( .A(A[2]), .Z(n119) );
    VMW_INV U51 ( .A(A[0]), .Z(n121) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE3_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [3:0] Nid;
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp284[0] , \OutEdge116[6] , \temp284[9] , \temp284[11] , 
        \temp190[2] , \OutEdge116[2] , \temp284[4] , \temp190[6] , 
        \temp284[15] , \path[2] , \OutEdge116[9] , \path[0] , \temp190[4] , 
        \OutEdge116[0] , \temp284[6] , \temp284[13] , \temp190[0] , 
        \temp284[2] , \OutEdge116[4] , \temp190[9] , \temp190[10] , 
        \OutEdge116[11] , \OutEdge116[15] , \temp190[14] , \OutEdge116[13] , 
        \temp190[12] , n94, \OutEdge116[12] , \temp190[13] , n86, 
        \OutEdge116[14] , \temp190[15] , \temp190[11] , \OutEdge116[10] , 
        \temp284[12] , \temp190[1] , \temp284[3] , \OutEdge116[5] , 
        \temp190[8] , \path[1] , \OutEdge116[8] , \temp190[5] , 
        \OutEdge116[1] , \temp284[7] , n102, \OutEdge116[3] , \temp284[5] , 
        \temp190[7] , \temp284[14] , \temp284[1] , \OutEdge116[7] , 
        \temp284[8] , \temp284[10] , \temp190[3] , n467, n468, n469, n470, 
        n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
        n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U64 ( .Z(n500) );
    VMW_PULLDOWN U65 ( .Z(n502) );
    VMW_PULLDOWN U66 ( .Z(n501) );
    VMW_AND2 U67 ( .A(n467), .B(n468), .Z(\OutEdge116[15] ) );
    VMW_OR2 U68 ( .A(n469), .B(Start), .Z(\OutEdge116[14] ) );
    VMW_OR2 U69 ( .A(n470), .B(Start), .Z(\OutEdge116[13] ) );
    VMW_OR2 U70 ( .A(n471), .B(Start), .Z(\OutEdge116[12] ) );
    VMW_OR2 U71 ( .A(n472), .B(Start), .Z(\OutEdge116[11] ) );
    VMW_OR2 U72 ( .A(n473), .B(Start), .Z(\OutEdge116[10] ) );
    VMW_OR2 U73 ( .A(n474), .B(Start), .Z(\OutEdge116[9] ) );
    VMW_OR2 U74 ( .A(n475), .B(Start), .Z(\OutEdge116[8] ) );
    VMW_OR2 U75 ( .A(n476), .B(Start), .Z(\OutEdge116[7] ) );
    VMW_OR2 U76 ( .A(n477), .B(Start), .Z(\OutEdge116[6] ) );
    VMW_OR2 U77 ( .A(n478), .B(Start), .Z(\OutEdge116[5] ) );
    VMW_OR2 U78 ( .A(n479), .B(Start), .Z(\OutEdge116[4] ) );
    VMW_OR2 U79 ( .A(n480), .B(Start), .Z(\OutEdge116[3] ) );
    VMW_OR2 U80 ( .A(n481), .B(Start), .Z(\OutEdge116[2] ) );
    VMW_OR2 U81 ( .A(n482), .B(Start), .Z(\OutEdge116[1] ) );
    VMW_OR2 U82 ( .A(n483), .B(Start), .Z(\OutEdge116[0] ) );
    VMW_OR2 U83 ( .A(n484), .B(n485), .Z(n499) );
    VMW_AO22 U84 ( .A(\path[2] ), .B(Start), .C(n486), .D(n485), .Z(n498) );
    VMW_AO22 U85 ( .A(\temp190[15] ), .B(n487), .C(InEdges[31]), .D(n94), .Z(
        \temp284[15] ) );
    VMW_AND3 U86 ( .A(n467), .B(n488), .C(n487), .Z(n485) );
    VMW_INV U87 ( .A(Start), .Z(n467) );
    VMW_AO22 U88 ( .A(n490), .B(n467), .C(n491), .D(Start), .Z(n489) );
    VMW_AO22 U89 ( .A(\temp284[15] ), .B(n486), .C(InEdges[47]), .D(n102), .Z(
        n468) );
    VMW_INV U90 ( .A(n102), .Z(n486) );
    VMW_AND4 U91 ( .A(n492), .B(n493), .C(n494), .D(n495), .Z(n496) );
    VMW_XNOR2 U92 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n495) );
    VMW_XNOR2 U93 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n494) );
    VMW_XNOR2 U94 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n493) );
    VMW_XNOR2 U95 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n492) );
    VMW_AO22 U96 ( .A(InEdges[9]), .B(n86), .C(OutEdge[9]), .D(n488), .Z(
        \temp190[9] ) );
    VMW_AO22 U97 ( .A(\temp190[9] ), .B(n487), .C(InEdges[25]), .D(n94), .Z(
        \temp284[9] ) );
    VMW_AO22 U98 ( .A(InEdges[8]), .B(n86), .C(OutEdge[8]), .D(n488), .Z(
        \temp190[8] ) );
    VMW_AO22 U99 ( .A(\temp190[8] ), .B(n487), .C(InEdges[24]), .D(n94), .Z(
        \temp284[8] ) );
    VMW_AO22 U100 ( .A(InEdges[7]), .B(n86), .C(OutEdge[7]), .D(n488), .Z(
        \temp190[7] ) );
    VMW_AO22 U101 ( .A(\temp190[7] ), .B(n487), .C(InEdges[23]), .D(n94), .Z(
        \temp284[7] ) );
    VMW_AO22 U102 ( .A(InEdges[6]), .B(n86), .C(OutEdge[6]), .D(n488), .Z(
        \temp190[6] ) );
    VMW_AO22 U103 ( .A(\temp190[6] ), .B(n487), .C(InEdges[22]), .D(n94), .Z(
        \temp284[6] ) );
    VMW_AO22 U104 ( .A(InEdges[5]), .B(n86), .C(OutEdge[5]), .D(n488), .Z(
        \temp190[5] ) );
    VMW_AO22 U105 ( .A(\temp190[5] ), .B(n487), .C(InEdges[21]), .D(n94), .Z(
        \temp284[5] ) );
    VMW_AO22 U106 ( .A(InEdges[4]), .B(n86), .C(OutEdge[4]), .D(n488), .Z(
        \temp190[4] ) );
    VMW_AO22 U107 ( .A(\temp190[4] ), .B(n487), .C(InEdges[20]), .D(n94), .Z(
        \temp284[4] ) );
    VMW_AO22 U108 ( .A(InEdges[3]), .B(n86), .C(OutEdge[3]), .D(n488), .Z(
        \temp190[3] ) );
    VMW_AO22 U109 ( .A(\temp190[3] ), .B(n487), .C(InEdges[19]), .D(n94), .Z(
        \temp284[3] ) );
    VMW_AO22 U110 ( .A(InEdges[2]), .B(n86), .C(OutEdge[2]), .D(n488), .Z(
        \temp190[2] ) );
    VMW_AO22 U111 ( .A(\temp190[2] ), .B(n487), .C(InEdges[18]), .D(n94), .Z(
        \temp284[2] ) );
    VMW_AO22 U112 ( .A(InEdges[1]), .B(n86), .C(OutEdge[1]), .D(n488), .Z(
        \temp190[1] ) );
    VMW_AO22 U113 ( .A(\temp190[1] ), .B(n487), .C(InEdges[17]), .D(n94), .Z(
        \temp284[1] ) );
    VMW_AO22 U114 ( .A(InEdges[15]), .B(n86), .C(OutEdge[15]), .D(n488), .Z(
        \temp190[15] ) );
    VMW_AO22 U115 ( .A(InEdges[14]), .B(n86), .C(OutEdge[14]), .D(n488), .Z(
        \temp190[14] ) );
    VMW_AO22 U116 ( .A(\temp190[14] ), .B(n487), .C(InEdges[30]), .D(n94), .Z(
        \temp284[14] ) );
    VMW_AO22 U117 ( .A(InEdges[13]), .B(n86), .C(OutEdge[13]), .D(n488), .Z(
        \temp190[13] ) );
    VMW_AO22 U118 ( .A(\temp190[13] ), .B(n487), .C(InEdges[29]), .D(n94), .Z(
        \temp284[13] ) );
    VMW_AO22 U119 ( .A(InEdges[12]), .B(n86), .C(OutEdge[12]), .D(n488), .Z(
        \temp190[12] ) );
    VMW_AO22 U120 ( .A(\temp190[12] ), .B(n487), .C(InEdges[28]), .D(n94), .Z(
        \temp284[12] ) );
    VMW_AO22 U121 ( .A(InEdges[11]), .B(n86), .C(OutEdge[11]), .D(n488), .Z(
        \temp190[11] ) );
    VMW_AO22 U122 ( .A(\temp190[11] ), .B(n487), .C(InEdges[27]), .D(n94), .Z(
        \temp284[11] ) );
    VMW_AO22 U123 ( .A(InEdges[10]), .B(n86), .C(OutEdge[10]), .D(n488), .Z(
        \temp190[10] ) );
    VMW_AO22 U124 ( .A(\temp190[10] ), .B(n487), .C(InEdges[26]), .D(n94), .Z(
        \temp284[10] ) );
    VMW_AO22 U125 ( .A(InEdges[0]), .B(n86), .C(OutEdge[0]), .D(n488), .Z(
        \temp190[0] ) );
    VMW_AO22 U126 ( .A(\temp190[0] ), .B(n487), .C(InEdges[16]), .D(n94), .Z(
        \temp284[0] ) );
    VMW_AO22 U127 ( .A(\path[1] ), .B(Start), .C(n102), .D(n467), .Z(n484) );
    VMW_AO21 U128 ( .A(n487), .B(n86), .C(n102), .Z(n490) );
    VMW_AO22 U129 ( .A(\temp284[9] ), .B(n486), .C(InEdges[41]), .D(n102), .Z(
        n474) );
    VMW_AO22 U130 ( .A(\temp284[8] ), .B(n486), .C(InEdges[40]), .D(n102), .Z(
        n475) );
    VMW_AO22 U131 ( .A(\temp284[7] ), .B(n486), .C(InEdges[39]), .D(n102), .Z(
        n476) );
    VMW_AO22 U132 ( .A(\temp284[6] ), .B(n486), .C(InEdges[38]), .D(n102), .Z(
        n477) );
    VMW_AO22 U133 ( .A(\temp284[5] ), .B(n486), .C(InEdges[37]), .D(n102), .Z(
        n478) );
    VMW_AO22 U134 ( .A(\temp284[4] ), .B(n486), .C(InEdges[36]), .D(n102), .Z(
        n479) );
    VMW_AO22 U135 ( .A(\temp284[3] ), .B(n486), .C(InEdges[35]), .D(n102), .Z(
        n480) );
    VMW_AO22 U136 ( .A(\temp284[2] ), .B(n486), .C(InEdges[34]), .D(n102), .Z(
        n481) );
    VMW_AO22 U137 ( .A(\temp284[1] ), .B(n486), .C(InEdges[33]), .D(n102), .Z(
        n482) );
    VMW_AO22 U138 ( .A(\temp284[14] ), .B(n486), .C(InEdges[46]), .D(n102), 
        .Z(n469) );
    VMW_AO22 U139 ( .A(\temp284[13] ), .B(n486), .C(InEdges[45]), .D(n102), 
        .Z(n470) );
    VMW_AO22 U140 ( .A(\temp284[12] ), .B(n486), .C(InEdges[44]), .D(n102), 
        .Z(n471) );
    VMW_AO22 U141 ( .A(\temp284[11] ), .B(n486), .C(InEdges[43]), .D(n102), 
        .Z(n472) );
    VMW_AO22 U142 ( .A(\temp284[10] ), .B(n486), .C(InEdges[42]), .D(n102), 
        .Z(n473) );
    VMW_AO22 U143 ( .A(\temp284[0] ), .B(n486), .C(InEdges[32]), .D(n102), .Z(
        n483) );
    VMW_INV U144 ( .A(n86), .Z(n488) );
    VMW_INV U145 ( .A(n94), .Z(n487) );
    VMW_INV U146 ( .A(n489), .Z(n497) );
    VMW_INV U147 ( .A(\path[0] ), .Z(n491) );
    VMW_BUFIZ U148 ( .A(\path[1] ), .E(n496), .Z(\PathData[1] ) );
    VMW_BUFIZ U149 ( .A(\path[0] ), .E(n496), .Z(\PathData[0] ) );
    VMW_BUFIZ U150 ( .A(\path[2] ), .E(n496), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n497), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n498), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n499), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge116[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge116[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge116[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge116[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge116[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge116[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge116[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge116[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge116[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge116[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge116[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge116[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge116[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge116[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge116[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge116[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp190[15] , 
        \temp190[14] , \temp190[13] , \temp190[12] , \temp190[11] , 
        \temp190[10] , \temp190[9] , \temp190[8] , \temp190[7] , \temp190[6] , 
        \temp190[5] , \temp190[4] , \temp190[3] , \temp190[2] , \temp190[1] , 
        \temp190[0] }), .B(InEdges[31:16]), .LEQ(n502), .TC(n502), .GE_GT(n94)
         );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n501), .TC(n501), .GE_GT(n86) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 lte_55_2 ( .A({\temp284[15] , 
        \temp284[14] , \temp284[13] , \temp284[12] , \temp284[11] , 
        \temp284[10] , \temp284[9] , \temp284[8] , \temp284[7] , \temp284[6] , 
        \temp284[5] , \temp284[4] , \temp284[3] , \temp284[2] , \temp284[1] , 
        \temp284[0] }), .B(InEdges[47:32]), .LEQ(n500), .TC(n500), .GE_GT(n102
        ) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, 
        n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, 
        n108, n109, n110, n111, n113, n114, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n95), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n113), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n113), .B(A[13]), .Z(n114) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n114), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n113) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
        n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
        n164, n165;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n127), .B(B[4]), .Z(n126) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n129), .C(n125), .D(n119), .Z(n128) );
    VMW_OR2 U10 ( .A(B[4]), .B(n127), .Z(n130) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n132), .C(n130), .D(n128), .Z(n131) );
    VMW_NAND2 U12 ( .A(n134), .B(B[6]), .Z(n133) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n136), .C(n131), .D(n126), .Z(n135) );
    VMW_OR2 U14 ( .A(B[6]), .B(n134), .Z(n137) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n139), .C(n137), .D(n135), .Z(n138) );
    VMW_NAND2 U16 ( .A(n141), .B(B[8]), .Z(n140) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n143), .C(n138), .D(n133), .Z(n142) );
    VMW_OR2 U18 ( .A(B[8]), .B(n141), .Z(n144) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n146), .C(n144), .D(n142), .Z(n145) );
    VMW_NAND2 U20 ( .A(n148), .B(B[10]), .Z(n147) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n150), .C(n145), .D(n140), .Z(n149) );
    VMW_NAND2 U22 ( .A(n150), .B(A[9]), .Z(n151) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n148), .C(n151), .D(n149), .Z(n152) );
    VMW_NAND2 U24 ( .A(n154), .B(B[12]), .Z(n153) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n156), .C(n152), .D(n147), .Z(n155) );
    VMW_NAND2 U26 ( .A(n156), .B(A[11]), .Z(n157) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n154), .C(n157), .D(n155), .Z(n158) );
    VMW_NAND2 U28 ( .A(n160), .B(B[14]), .Z(n159) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n162), .C(n158), .D(n153), .Z(n161) );
    VMW_NAND2 U30 ( .A(n162), .B(A[13]), .Z(n163) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n160), .C(n163), .D(n161), .Z(n164) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n165), .C(n164), .D(n159), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n154) );
    VMW_INV U34 ( .A(B[7]), .Z(n143) );
    VMW_INV U35 ( .A(A[7]), .Z(n146) );
    VMW_INV U36 ( .A(A[3]), .Z(n132) );
    VMW_INV U37 ( .A(B[3]), .Z(n129) );
    VMW_INV U38 ( .A(A[10]), .Z(n148) );
    VMW_INV U39 ( .A(B[9]), .Z(n150) );
    VMW_INV U40 ( .A(A[4]), .Z(n127) );
    VMW_INV U41 ( .A(A[8]), .Z(n141) );
    VMW_INV U42 ( .A(A[14]), .Z(n160) );
    VMW_INV U43 ( .A(B[11]), .Z(n156) );
    VMW_INV U44 ( .A(A[5]), .Z(n139) );
    VMW_INV U45 ( .A(B[5]), .Z(n136) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n165) );
    VMW_INV U48 ( .A(B[13]), .Z(n162) );
    VMW_INV U49 ( .A(A[6]), .Z(n134) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
        n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
        n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
        n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
        n213, n214;
    VMW_OAI21 U3 ( .A(B[15]), .B(n166), .C(n167), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n169), .B(B[2]), .Z(n168) );
    VMW_AO22 U5 ( .A(n171), .B(B[0]), .C(n172), .D(B[1]), .Z(n170) );
    VMW_OR2 U6 ( .A(B[2]), .B(n169), .Z(n173) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n172), .C(n173), .D(n170), .Z(n174) );
    VMW_NAND2 U8 ( .A(n176), .B(B[4]), .Z(n175) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n178), .C(n174), .D(n168), .Z(n177) );
    VMW_OR2 U10 ( .A(B[4]), .B(n176), .Z(n179) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n181), .C(n179), .D(n177), .Z(n180) );
    VMW_NAND2 U12 ( .A(n183), .B(B[6]), .Z(n182) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n185), .C(n180), .D(n175), .Z(n184) );
    VMW_OR2 U14 ( .A(B[6]), .B(n183), .Z(n186) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n188), .C(n186), .D(n184), .Z(n187) );
    VMW_NAND2 U16 ( .A(n190), .B(B[8]), .Z(n189) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n192), .C(n187), .D(n182), .Z(n191) );
    VMW_OR2 U18 ( .A(B[8]), .B(n190), .Z(n193) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n195), .C(n193), .D(n191), .Z(n194) );
    VMW_NAND2 U20 ( .A(n197), .B(B[10]), .Z(n196) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n199), .C(n194), .D(n189), .Z(n198) );
    VMW_NAND2 U22 ( .A(n199), .B(A[9]), .Z(n200) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n197), .C(n200), .D(n198), .Z(n201) );
    VMW_NAND2 U24 ( .A(n203), .B(B[12]), .Z(n202) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n205), .C(n201), .D(n196), .Z(n204) );
    VMW_NAND2 U26 ( .A(n205), .B(A[11]), .Z(n206) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n203), .C(n206), .D(n204), .Z(n207) );
    VMW_NAND2 U28 ( .A(n209), .B(B[14]), .Z(n208) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n211), .C(n207), .D(n202), .Z(n210) );
    VMW_NAND2 U30 ( .A(n211), .B(A[13]), .Z(n212) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n209), .C(n212), .D(n210), .Z(n213) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n214), .C(n213), .D(n208), .Z(n167) );
    VMW_INV U33 ( .A(A[12]), .Z(n203) );
    VMW_INV U34 ( .A(B[7]), .Z(n192) );
    VMW_INV U35 ( .A(A[7]), .Z(n195) );
    VMW_INV U36 ( .A(A[3]), .Z(n181) );
    VMW_INV U37 ( .A(B[3]), .Z(n178) );
    VMW_INV U38 ( .A(A[10]), .Z(n197) );
    VMW_INV U39 ( .A(B[9]), .Z(n199) );
    VMW_INV U40 ( .A(A[4]), .Z(n176) );
    VMW_INV U41 ( .A(A[8]), .Z(n190) );
    VMW_INV U42 ( .A(A[14]), .Z(n209) );
    VMW_INV U43 ( .A(B[11]), .Z(n205) );
    VMW_INV U44 ( .A(A[5]), .Z(n188) );
    VMW_INV U45 ( .A(B[5]), .Z(n185) );
    VMW_INV U46 ( .A(A[1]), .Z(n172) );
    VMW_INV U47 ( .A(B[15]), .Z(n214) );
    VMW_INV U48 ( .A(B[13]), .Z(n211) );
    VMW_INV U49 ( .A(A[6]), .Z(n183) );
    VMW_INV U50 ( .A(A[2]), .Z(n169) );
    VMW_INV U51 ( .A(A[0]), .Z(n171) );
    VMW_INV U52 ( .A(A[15]), .Z(n166) );
endmodule


module NodeAux_INDEGREE4_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [3:0] Nid;
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp200[0] , \temp384[15] , \OutEdge126[12] , \temp200[15] , 
        \temp200[9] , \temp384[6] , \temp294[3] , n112, \temp294[13] , 
        \temp384[11] , \temp200[4] , \temp294[7] , \temp384[2] , \path[2] , 
        \temp200[11] , \temp200[13] , \path[0] , \temp294[5] , \temp384[0] , 
        \temp384[13] , \temp200[6] , \temp384[9] , \OutEdge126[14] , 
        \temp294[11] , \temp384[4] , \temp294[1] , \OutEdge126[10] , 
        \temp294[15] , \temp200[2] , \temp294[8] , \OutEdge126[8] , 
        \OutEdge126[1] , \OutEdge126[5] , n96, \OutEdge126[7] , 
        \OutEdge126[3] , \OutEdge126[2] , \OutEdge126[6] , \OutEdge126[4] , 
        n104, \OutEdge126[9] , n88, \OutEdge126[0] , \temp384[5] , 
        \temp294[0] , \OutEdge126[11] , \temp294[14] , \temp200[3] , 
        \temp294[9] , \path[1] , \temp200[12] , \temp294[4] , \temp384[1] , 
        \temp384[12] , \temp384[8] , \temp200[7] , \OutEdge126[15] , 
        \temp294[10] , \temp294[12] , \temp384[10] , \temp200[5] , 
        \temp294[6] , \temp384[3] , \temp200[10] , \temp200[1] , \temp384[14] , 
        \OutEdge126[13] , \temp200[14] , \temp384[7] , \temp200[8] , 
        \temp294[2] , n567, n568, n569, n570, n571, n572, n573, n574, n575, 
        n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
        n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
        n600, n601, n602, n603, n604, n605, n606;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U73 ( .Z(n603) );
    VMW_PULLDOWN U74 ( .Z(n604) );
    VMW_PULLDOWN U75 ( .Z(n605) );
    VMW_PULLDOWN U76 ( .Z(n606) );
    VMW_NOR2 U77 ( .A(Start), .B(n567), .Z(\OutEdge126[15] ) );
    VMW_NAND2 U78 ( .A(n568), .B(n569), .Z(\OutEdge126[14] ) );
    VMW_NAND2 U79 ( .A(n570), .B(n569), .Z(\OutEdge126[13] ) );
    VMW_NAND2 U80 ( .A(n571), .B(n569), .Z(\OutEdge126[12] ) );
    VMW_NAND2 U81 ( .A(n572), .B(n569), .Z(\OutEdge126[11] ) );
    VMW_NAND2 U82 ( .A(n573), .B(n569), .Z(\OutEdge126[10] ) );
    VMW_NAND2 U83 ( .A(n574), .B(n569), .Z(\OutEdge126[9] ) );
    VMW_NAND2 U84 ( .A(n575), .B(n569), .Z(\OutEdge126[8] ) );
    VMW_NAND2 U85 ( .A(n576), .B(n569), .Z(\OutEdge126[7] ) );
    VMW_NAND2 U86 ( .A(n577), .B(n569), .Z(\OutEdge126[6] ) );
    VMW_NAND2 U87 ( .A(n578), .B(n569), .Z(\OutEdge126[5] ) );
    VMW_NAND2 U88 ( .A(n579), .B(n569), .Z(\OutEdge126[4] ) );
    VMW_NAND2 U89 ( .A(n580), .B(n569), .Z(\OutEdge126[3] ) );
    VMW_NAND2 U90 ( .A(n581), .B(n569), .Z(\OutEdge126[2] ) );
    VMW_NAND2 U91 ( .A(n582), .B(n569), .Z(\OutEdge126[1] ) );
    VMW_NAND2 U92 ( .A(n583), .B(n569), .Z(\OutEdge126[0] ) );
    VMW_OAI211 U93 ( .A(n96), .B(n88), .C(n585), .D(n586), .Z(n584) );
    VMW_NAND2 U94 ( .A(n585), .B(n588), .Z(n587) );
    VMW_AO22 U95 ( .A(\temp294[15] ), .B(n586), .C(InEdges[47]), .D(n104), .Z(
        \temp384[15] ) );
    VMW_INV U96 ( .A(n88), .Z(n589) );
    VMW_OAI22 U97 ( .A(n591), .B(Start), .C(\path[2] ), .D(n569), .Z(n590) );
    VMW_OAI22 U98 ( .A(n584), .B(Start), .C(\path[1] ), .D(n569), .Z(n592) );
    VMW_OAI22 U99 ( .A(n587), .B(Start), .C(\path[0] ), .D(n569), .Z(n593) );
    VMW_MUX2I U100 ( .A(\temp384[15] ), .B(InEdges[63]), .S(n112), .Z(n567) );
    VMW_INV U101 ( .A(Start), .Z(n569) );
    VMW_INV U102 ( .A(n96), .Z(n594) );
    VMW_OAI21 U103 ( .A(n96), .B(n589), .C(n586), .Z(n588) );
    VMW_AND4 U104 ( .A(n595), .B(n596), .C(n597), .D(n598), .Z(n599) );
    VMW_XNOR2 U105 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n598) );
    VMW_XNOR2 U106 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n597) );
    VMW_XNOR2 U107 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n596) );
    VMW_XNOR2 U108 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n595) );
    VMW_AO22 U109 ( .A(InEdges[9]), .B(n88), .C(OutEdge[9]), .D(n589), .Z(
        \temp200[9] ) );
    VMW_AO22 U110 ( .A(InEdges[25]), .B(n96), .C(\temp200[9] ), .D(n594), .Z(
        \temp294[9] ) );
    VMW_AO22 U111 ( .A(\temp294[9] ), .B(n586), .C(InEdges[41]), .D(n104), .Z(
        \temp384[9] ) );
    VMW_AO22 U112 ( .A(InEdges[8]), .B(n88), .C(OutEdge[8]), .D(n589), .Z(
        \temp200[8] ) );
    VMW_AO22 U113 ( .A(InEdges[24]), .B(n96), .C(\temp200[8] ), .D(n594), .Z(
        \temp294[8] ) );
    VMW_AO22 U114 ( .A(\temp294[8] ), .B(n586), .C(InEdges[40]), .D(n104), .Z(
        \temp384[8] ) );
    VMW_AO22 U115 ( .A(InEdges[7]), .B(n88), .C(OutEdge[7]), .D(n589), .Z(
        \temp200[7] ) );
    VMW_AO22 U116 ( .A(InEdges[23]), .B(n96), .C(\temp200[7] ), .D(n594), .Z(
        \temp294[7] ) );
    VMW_AO22 U117 ( .A(\temp294[7] ), .B(n586), .C(InEdges[39]), .D(n104), .Z(
        \temp384[7] ) );
    VMW_AO22 U118 ( .A(InEdges[6]), .B(n88), .C(OutEdge[6]), .D(n589), .Z(
        \temp200[6] ) );
    VMW_AO22 U119 ( .A(InEdges[22]), .B(n96), .C(\temp200[6] ), .D(n594), .Z(
        \temp294[6] ) );
    VMW_AO22 U120 ( .A(\temp294[6] ), .B(n586), .C(InEdges[38]), .D(n104), .Z(
        \temp384[6] ) );
    VMW_AO22 U121 ( .A(InEdges[5]), .B(n88), .C(OutEdge[5]), .D(n589), .Z(
        \temp200[5] ) );
    VMW_AO22 U122 ( .A(InEdges[21]), .B(n96), .C(\temp200[5] ), .D(n594), .Z(
        \temp294[5] ) );
    VMW_AO22 U123 ( .A(\temp294[5] ), .B(n586), .C(InEdges[37]), .D(n104), .Z(
        \temp384[5] ) );
    VMW_AO22 U124 ( .A(InEdges[4]), .B(n88), .C(OutEdge[4]), .D(n589), .Z(
        \temp200[4] ) );
    VMW_AO22 U125 ( .A(InEdges[20]), .B(n96), .C(\temp200[4] ), .D(n594), .Z(
        \temp294[4] ) );
    VMW_AO22 U126 ( .A(\temp294[4] ), .B(n586), .C(InEdges[36]), .D(n104), .Z(
        \temp384[4] ) );
    VMW_AO22 U127 ( .A(InEdges[3]), .B(n88), .C(OutEdge[3]), .D(n589), .Z(
        \temp200[3] ) );
    VMW_AO22 U128 ( .A(InEdges[19]), .B(n96), .C(\temp200[3] ), .D(n594), .Z(
        \temp294[3] ) );
    VMW_AO22 U129 ( .A(\temp294[3] ), .B(n586), .C(InEdges[35]), .D(n104), .Z(
        \temp384[3] ) );
    VMW_AO22 U130 ( .A(InEdges[2]), .B(n88), .C(OutEdge[2]), .D(n589), .Z(
        \temp200[2] ) );
    VMW_AO22 U131 ( .A(InEdges[18]), .B(n96), .C(\temp200[2] ), .D(n594), .Z(
        \temp294[2] ) );
    VMW_AO22 U132 ( .A(\temp294[2] ), .B(n586), .C(InEdges[34]), .D(n104), .Z(
        \temp384[2] ) );
    VMW_AO22 U133 ( .A(InEdges[1]), .B(n88), .C(OutEdge[1]), .D(n589), .Z(
        \temp200[1] ) );
    VMW_AO22 U134 ( .A(InEdges[17]), .B(n96), .C(\temp200[1] ), .D(n594), .Z(
        \temp294[1] ) );
    VMW_AO22 U135 ( .A(\temp294[1] ), .B(n586), .C(InEdges[33]), .D(n104), .Z(
        \temp384[1] ) );
    VMW_AO22 U136 ( .A(InEdges[15]), .B(n88), .C(OutEdge[15]), .D(n589), .Z(
        \temp200[15] ) );
    VMW_AO22 U137 ( .A(InEdges[31]), .B(n96), .C(\temp200[15] ), .D(n594), .Z(
        \temp294[15] ) );
    VMW_AO22 U138 ( .A(InEdges[14]), .B(n88), .C(OutEdge[14]), .D(n589), .Z(
        \temp200[14] ) );
    VMW_AO22 U139 ( .A(InEdges[30]), .B(n96), .C(\temp200[14] ), .D(n594), .Z(
        \temp294[14] ) );
    VMW_AO22 U140 ( .A(\temp294[14] ), .B(n586), .C(InEdges[46]), .D(n104), 
        .Z(\temp384[14] ) );
    VMW_AO22 U141 ( .A(InEdges[13]), .B(n88), .C(OutEdge[13]), .D(n589), .Z(
        \temp200[13] ) );
    VMW_AO22 U142 ( .A(InEdges[29]), .B(n96), .C(\temp200[13] ), .D(n594), .Z(
        \temp294[13] ) );
    VMW_AO22 U143 ( .A(\temp294[13] ), .B(n586), .C(InEdges[45]), .D(n104), 
        .Z(\temp384[13] ) );
    VMW_AO22 U144 ( .A(InEdges[12]), .B(n88), .C(OutEdge[12]), .D(n589), .Z(
        \temp200[12] ) );
    VMW_AO22 U145 ( .A(InEdges[28]), .B(n96), .C(\temp200[12] ), .D(n594), .Z(
        \temp294[12] ) );
    VMW_AO22 U146 ( .A(\temp294[12] ), .B(n586), .C(InEdges[44]), .D(n104), 
        .Z(\temp384[12] ) );
    VMW_AO22 U147 ( .A(InEdges[11]), .B(n88), .C(OutEdge[11]), .D(n589), .Z(
        \temp200[11] ) );
    VMW_AO22 U148 ( .A(InEdges[27]), .B(n96), .C(\temp200[11] ), .D(n594), .Z(
        \temp294[11] ) );
    VMW_AO22 U149 ( .A(\temp294[11] ), .B(n586), .C(InEdges[43]), .D(n104), 
        .Z(\temp384[11] ) );
    VMW_AO22 U150 ( .A(InEdges[10]), .B(n88), .C(OutEdge[10]), .D(n589), .Z(
        \temp200[10] ) );
    VMW_AO22 U151 ( .A(InEdges[26]), .B(n96), .C(\temp200[10] ), .D(n594), .Z(
        \temp294[10] ) );
    VMW_AO22 U152 ( .A(\temp294[10] ), .B(n586), .C(InEdges[42]), .D(n104), 
        .Z(\temp384[10] ) );
    VMW_AO22 U153 ( .A(InEdges[0]), .B(n88), .C(OutEdge[0]), .D(n589), .Z(
        \temp200[0] ) );
    VMW_AO22 U154 ( .A(InEdges[16]), .B(n96), .C(\temp200[0] ), .D(n594), .Z(
        \temp294[0] ) );
    VMW_AO22 U155 ( .A(\temp294[0] ), .B(n586), .C(InEdges[32]), .D(n104), .Z(
        \temp384[0] ) );
    VMW_AND4 U156 ( .A(n594), .B(n586), .C(n589), .D(n585), .Z(n591) );
    VMW_MUX2I U157 ( .A(\temp384[9] ), .B(InEdges[57]), .S(n112), .Z(n574) );
    VMW_MUX2I U158 ( .A(\temp384[8] ), .B(InEdges[56]), .S(n112), .Z(n575) );
    VMW_MUX2I U159 ( .A(\temp384[7] ), .B(InEdges[55]), .S(n112), .Z(n576) );
    VMW_MUX2I U160 ( .A(\temp384[6] ), .B(InEdges[54]), .S(n112), .Z(n577) );
    VMW_MUX2I U161 ( .A(\temp384[5] ), .B(InEdges[53]), .S(n112), .Z(n578) );
    VMW_MUX2I U162 ( .A(\temp384[4] ), .B(InEdges[52]), .S(n112), .Z(n579) );
    VMW_MUX2I U163 ( .A(\temp384[3] ), .B(InEdges[51]), .S(n112), .Z(n580) );
    VMW_MUX2I U164 ( .A(\temp384[2] ), .B(InEdges[50]), .S(n112), .Z(n581) );
    VMW_MUX2I U165 ( .A(\temp384[1] ), .B(InEdges[49]), .S(n112), .Z(n582) );
    VMW_MUX2I U166 ( .A(\temp384[14] ), .B(InEdges[62]), .S(n112), .Z(n568) );
    VMW_MUX2I U167 ( .A(\temp384[13] ), .B(InEdges[61]), .S(n112), .Z(n570) );
    VMW_MUX2I U168 ( .A(\temp384[12] ), .B(InEdges[60]), .S(n112), .Z(n571) );
    VMW_MUX2I U169 ( .A(\temp384[11] ), .B(InEdges[59]), .S(n112), .Z(n572) );
    VMW_MUX2I U170 ( .A(\temp384[10] ), .B(InEdges[58]), .S(n112), .Z(n573) );
    VMW_MUX2I U171 ( .A(\temp384[0] ), .B(InEdges[48]), .S(n112), .Z(n583) );
    VMW_INV U172 ( .A(n104), .Z(n586) );
    VMW_INV U173 ( .A(n112), .Z(n585) );
    VMW_INV U174 ( .A(n590), .Z(n601) );
    VMW_INV U175 ( .A(n592), .Z(n602) );
    VMW_INV U176 ( .A(n593), .Z(n600) );
    VMW_BUFIZ U177 ( .A(\path[1] ), .E(n599), .Z(\PathData[1] ) );
    VMW_BUFIZ U178 ( .A(\path[0] ), .E(n599), .Z(\PathData[0] ) );
    VMW_BUFIZ U179 ( .A(\path[2] ), .E(n599), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n600), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n601), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n602), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge126[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge126[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge126[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge126[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge126[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge126[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge126[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge126[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge126[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge126[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge126[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge126[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge126[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge126[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge126[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge126[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n606), .TC(n606), .GE_GT(n88) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp200[15] , 
        \temp200[14] , \temp200[13] , \temp200[12] , \temp200[11] , 
        \temp200[10] , \temp200[9] , \temp200[8] , \temp200[7] , \temp200[6] , 
        \temp200[5] , \temp200[4] , \temp200[3] , \temp200[2] , \temp200[1] , 
        \temp200[0] }), .B(InEdges[31:16]), .LEQ(n605), .TC(n605), .GE_GT(n96)
         );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp294[15] , 
        \temp294[14] , \temp294[13] , \temp294[12] , \temp294[11] , 
        \temp294[10] , \temp294[9] , \temp294[8] , \temp294[7] , \temp294[6] , 
        \temp294[5] , \temp294[4] , \temp294[3] , \temp294[2] , \temp294[1] , 
        \temp294[0] }), .B(InEdges[47:32]), .LEQ(n604), .TC(n604), .GE_GT(n104
        ) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp384[15] , 
        \temp384[14] , \temp384[13] , \temp384[12] , \temp384[11] , 
        \temp384[10] , \temp384[9] , \temp384[8] , \temp384[7] , \temp384[6] , 
        \temp384[5] , \temp384[4] , \temp384[3] , \temp384[2] , \temp384[1] , 
        \temp384[0] }), .B(InEdges[63:48]), .LEQ(n603), .TC(n603), .GE_GT(n112
        ) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n91, n92, 
        n93, n94, n95, n96, n97, n99, n100, n101, n102, n103, n104, n105, n107, 
        n108, n109, n110, n111, n112, n113, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n100), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n104), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, 
        n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
        n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
        n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
        n165, n166;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n123), .B(B[0]), .C(n124), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n124), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n135), .B(B[6]), .Z(n134) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n137), .C(n132), .D(n127), .Z(n136) );
    VMW_OR2 U14 ( .A(B[6]), .B(n135), .Z(n138) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n140), .C(n138), .D(n136), .Z(n139) );
    VMW_NAND2 U16 ( .A(n142), .B(B[8]), .Z(n141) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n144), .C(n139), .D(n134), .Z(n143) );
    VMW_OR2 U18 ( .A(B[8]), .B(n142), .Z(n145) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n147), .C(n145), .D(n143), .Z(n146) );
    VMW_NAND2 U20 ( .A(n149), .B(B[10]), .Z(n148) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n151), .C(n146), .D(n141), .Z(n150) );
    VMW_NAND2 U22 ( .A(n151), .B(A[9]), .Z(n152) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n149), .C(n152), .D(n150), .Z(n153) );
    VMW_NAND2 U24 ( .A(n155), .B(B[12]), .Z(n154) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n157), .C(n153), .D(n148), .Z(n156) );
    VMW_NAND2 U26 ( .A(n157), .B(A[11]), .Z(n158) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n155), .C(n158), .D(n156), .Z(n159) );
    VMW_NAND2 U28 ( .A(n161), .B(B[14]), .Z(n160) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n163), .C(n159), .D(n154), .Z(n162) );
    VMW_NAND2 U30 ( .A(n163), .B(A[13]), .Z(n164) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n161), .C(n164), .D(n162), .Z(n165) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n166), .C(n165), .D(n160), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n155) );
    VMW_INV U34 ( .A(B[7]), .Z(n144) );
    VMW_INV U35 ( .A(A[7]), .Z(n147) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n149) );
    VMW_INV U39 ( .A(B[9]), .Z(n151) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n142) );
    VMW_INV U42 ( .A(A[14]), .Z(n161) );
    VMW_INV U43 ( .A(B[11]), .Z(n157) );
    VMW_INV U44 ( .A(A[5]), .Z(n140) );
    VMW_INV U45 ( .A(B[5]), .Z(n137) );
    VMW_INV U46 ( .A(A[1]), .Z(n124) );
    VMW_INV U47 ( .A(B[15]), .Z(n166) );
    VMW_INV U48 ( .A(B[13]), .Z(n163) );
    VMW_INV U49 ( .A(A[6]), .Z(n135) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n123) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
        n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
        n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
        n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
        n214, n215;
    VMW_OAI21 U3 ( .A(B[15]), .B(n167), .C(n168), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n170), .B(B[2]), .Z(n169) );
    VMW_AO22 U5 ( .A(n172), .B(B[0]), .C(n173), .D(B[1]), .Z(n171) );
    VMW_OR2 U6 ( .A(B[2]), .B(n170), .Z(n174) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n173), .C(n174), .D(n171), .Z(n175) );
    VMW_NAND2 U8 ( .A(n177), .B(B[4]), .Z(n176) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n179), .C(n175), .D(n169), .Z(n178) );
    VMW_OR2 U10 ( .A(B[4]), .B(n177), .Z(n180) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n182), .C(n180), .D(n178), .Z(n181) );
    VMW_NAND2 U12 ( .A(n184), .B(B[6]), .Z(n183) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n186), .C(n181), .D(n176), .Z(n185) );
    VMW_OR2 U14 ( .A(B[6]), .B(n184), .Z(n187) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n189), .C(n187), .D(n185), .Z(n188) );
    VMW_NAND2 U16 ( .A(n191), .B(B[8]), .Z(n190) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n193), .C(n188), .D(n183), .Z(n192) );
    VMW_OR2 U18 ( .A(B[8]), .B(n191), .Z(n194) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n196), .C(n194), .D(n192), .Z(n195) );
    VMW_NAND2 U20 ( .A(n198), .B(B[10]), .Z(n197) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n200), .C(n195), .D(n190), .Z(n199) );
    VMW_NAND2 U22 ( .A(n200), .B(A[9]), .Z(n201) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n198), .C(n201), .D(n199), .Z(n202) );
    VMW_NAND2 U24 ( .A(n204), .B(B[12]), .Z(n203) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n206), .C(n202), .D(n197), .Z(n205) );
    VMW_NAND2 U26 ( .A(n206), .B(A[11]), .Z(n207) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n204), .C(n207), .D(n205), .Z(n208) );
    VMW_NAND2 U28 ( .A(n210), .B(B[14]), .Z(n209) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n212), .C(n208), .D(n203), .Z(n211) );
    VMW_NAND2 U30 ( .A(n212), .B(A[13]), .Z(n213) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n210), .C(n213), .D(n211), .Z(n214) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n215), .C(n214), .D(n209), .Z(n168) );
    VMW_INV U33 ( .A(A[12]), .Z(n204) );
    VMW_INV U34 ( .A(B[7]), .Z(n193) );
    VMW_INV U35 ( .A(A[7]), .Z(n196) );
    VMW_INV U36 ( .A(A[3]), .Z(n182) );
    VMW_INV U37 ( .A(B[3]), .Z(n179) );
    VMW_INV U38 ( .A(A[10]), .Z(n198) );
    VMW_INV U39 ( .A(B[9]), .Z(n200) );
    VMW_INV U40 ( .A(A[4]), .Z(n177) );
    VMW_INV U41 ( .A(A[8]), .Z(n191) );
    VMW_INV U42 ( .A(A[14]), .Z(n210) );
    VMW_INV U43 ( .A(B[11]), .Z(n206) );
    VMW_INV U44 ( .A(A[5]), .Z(n189) );
    VMW_INV U45 ( .A(B[5]), .Z(n186) );
    VMW_INV U46 ( .A(A[1]), .Z(n173) );
    VMW_INV U47 ( .A(B[15]), .Z(n215) );
    VMW_INV U48 ( .A(B[13]), .Z(n212) );
    VMW_INV U49 ( .A(A[6]), .Z(n184) );
    VMW_INV U50 ( .A(A[2]), .Z(n170) );
    VMW_INV U51 ( .A(A[0]), .Z(n172) );
    VMW_INV U52 ( .A(A[15]), .Z(n167) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
        n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
        n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
        n263, n264;
    VMW_OAI21 U3 ( .A(B[15]), .B(n216), .C(n217), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n219), .B(B[2]), .Z(n218) );
    VMW_AO22 U5 ( .A(n221), .B(B[0]), .C(n222), .D(B[1]), .Z(n220) );
    VMW_OR2 U6 ( .A(B[2]), .B(n219), .Z(n223) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n222), .C(n223), .D(n220), .Z(n224) );
    VMW_NAND2 U8 ( .A(n226), .B(B[4]), .Z(n225) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n228), .C(n224), .D(n218), .Z(n227) );
    VMW_OR2 U10 ( .A(B[4]), .B(n226), .Z(n229) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n231), .C(n229), .D(n227), .Z(n230) );
    VMW_NAND2 U12 ( .A(n233), .B(B[6]), .Z(n232) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n235), .C(n230), .D(n225), .Z(n234) );
    VMW_OR2 U14 ( .A(B[6]), .B(n233), .Z(n236) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n238), .C(n236), .D(n234), .Z(n237) );
    VMW_NAND2 U16 ( .A(n240), .B(B[8]), .Z(n239) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n242), .C(n237), .D(n232), .Z(n241) );
    VMW_OR2 U18 ( .A(B[8]), .B(n240), .Z(n243) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n245), .C(n243), .D(n241), .Z(n244) );
    VMW_NAND2 U20 ( .A(n247), .B(B[10]), .Z(n246) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n249), .C(n244), .D(n239), .Z(n248) );
    VMW_NAND2 U22 ( .A(n249), .B(A[9]), .Z(n250) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n247), .C(n250), .D(n248), .Z(n251) );
    VMW_NAND2 U24 ( .A(n253), .B(B[12]), .Z(n252) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n255), .C(n251), .D(n246), .Z(n254) );
    VMW_NAND2 U26 ( .A(n255), .B(A[11]), .Z(n256) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n253), .C(n256), .D(n254), .Z(n257) );
    VMW_NAND2 U28 ( .A(n259), .B(B[14]), .Z(n258) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n261), .C(n257), .D(n252), .Z(n260) );
    VMW_NAND2 U30 ( .A(n261), .B(A[13]), .Z(n262) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n259), .C(n262), .D(n260), .Z(n263) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n264), .C(n263), .D(n258), .Z(n217) );
    VMW_INV U33 ( .A(A[12]), .Z(n253) );
    VMW_INV U34 ( .A(B[7]), .Z(n242) );
    VMW_INV U35 ( .A(A[7]), .Z(n245) );
    VMW_INV U36 ( .A(A[3]), .Z(n231) );
    VMW_INV U37 ( .A(B[3]), .Z(n228) );
    VMW_INV U38 ( .A(A[10]), .Z(n247) );
    VMW_INV U39 ( .A(B[9]), .Z(n249) );
    VMW_INV U40 ( .A(A[4]), .Z(n226) );
    VMW_INV U41 ( .A(A[8]), .Z(n240) );
    VMW_INV U42 ( .A(A[14]), .Z(n259) );
    VMW_INV U43 ( .A(B[11]), .Z(n255) );
    VMW_INV U44 ( .A(A[5]), .Z(n238) );
    VMW_INV U45 ( .A(B[5]), .Z(n235) );
    VMW_INV U46 ( .A(A[1]), .Z(n222) );
    VMW_INV U47 ( .A(B[15]), .Z(n264) );
    VMW_INV U48 ( .A(B[13]), .Z(n261) );
    VMW_INV U49 ( .A(A[6]), .Z(n233) );
    VMW_INV U50 ( .A(A[2]), .Z(n219) );
    VMW_INV U51 ( .A(A[0]), .Z(n221) );
    VMW_INV U52 ( .A(A[15]), .Z(n216) );
endmodule


module NodeAux_INDEGREE5_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [3:0] Nid;
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp210[13] , \temp484[4] , \temp394[5] , \temp304[13] , 
        \temp210[3] , \temp394[13] , \OutEdge136[14] , \temp394[1] , 
        \temp484[0] , \OutEdge136[10] , \path[2] , \temp394[8] , \temp210[7] , 
        \temp484[9] , \temp394[15] , \path[0] , \temp210[5] , \OutEdge136[12] , 
        \temp210[15] , \temp304[15] , \temp394[3] , \temp484[2] , \temp210[1] , 
        n90, \temp394[11] , \temp484[6] , \temp394[7] , \temp210[8] , 
        \temp304[11] , \temp210[11] , n98, n114, \OutEdge136[2] , \temp304[4] , 
        \OutEdge136[6] , \temp304[9] , \temp304[0] , \temp484[13] , n106, 
        \temp304[2] , \temp484[11] , \OutEdge136[4] , \temp484[15] , 
        \temp304[6] , \OutEdge136[9] , \OutEdge136[0] , \temp484[14] , 
        \OutEdge136[8] , \temp304[7] , \OutEdge136[1] , \temp304[3] , 
        \temp484[10] , \OutEdge136[5] , \OutEdge136[7] , \temp304[8] , 
        \temp304[1] , \temp484[12] , \OutEdge136[3] , \temp304[5] , 
        \temp394[10] , \temp210[0] , \temp484[7] , \temp210[9] , \temp304[10] , 
        \temp394[6] , \temp210[10] , \path[1] , \temp210[4] , \temp394[14] , 
        \OutEdge136[13] , \temp210[14] , n122, \temp394[2] , \temp304[14] , 
        \temp484[3] , \temp394[0] , \temp484[1] , \OutEdge136[11] , 
        \temp210[6] , \temp394[9] , \temp484[8] , \temp210[12] , \temp484[5] , 
        \temp304[12] , \temp394[4] , \OutEdge136[15] , \temp394[12] , 
        \temp210[2] , n667, n668, n669, n670, n671, n672, n673, n674, n675, 
        n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
        n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
        n700, n701, n702, n703, n704, n705, n706, n707, n708, n709;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U82 ( .Z(n708) );
    VMW_PULLDOWN U83 ( .Z(n705) );
    VMW_PULLDOWN U84 ( .Z(n707) );
    VMW_PULLDOWN U85 ( .Z(n706) );
    VMW_PULLDOWN U86 ( .Z(n709) );
    VMW_AO21 U87 ( .A(\temp484[15] ), .B(n667), .C(n668), .Z(\OutEdge136[15] )
         );
    VMW_NAND2 U88 ( .A(n669), .B(n670), .Z(\OutEdge136[14] ) );
    VMW_NAND2 U89 ( .A(n671), .B(n670), .Z(\OutEdge136[13] ) );
    VMW_NAND2 U90 ( .A(n672), .B(n670), .Z(\OutEdge136[12] ) );
    VMW_NAND2 U91 ( .A(n673), .B(n670), .Z(\OutEdge136[11] ) );
    VMW_NAND2 U92 ( .A(n674), .B(n670), .Z(\OutEdge136[10] ) );
    VMW_NAND2 U93 ( .A(n675), .B(n670), .Z(\OutEdge136[9] ) );
    VMW_NAND2 U94 ( .A(n676), .B(n670), .Z(\OutEdge136[8] ) );
    VMW_NAND2 U95 ( .A(n677), .B(n670), .Z(\OutEdge136[7] ) );
    VMW_NAND2 U96 ( .A(n678), .B(n670), .Z(\OutEdge136[6] ) );
    VMW_NAND2 U97 ( .A(n679), .B(n670), .Z(\OutEdge136[5] ) );
    VMW_NAND2 U98 ( .A(n680), .B(n670), .Z(\OutEdge136[4] ) );
    VMW_NAND2 U99 ( .A(n681), .B(n670), .Z(\OutEdge136[3] ) );
    VMW_NAND2 U100 ( .A(n682), .B(n670), .Z(\OutEdge136[2] ) );
    VMW_NAND2 U101 ( .A(n683), .B(n670), .Z(\OutEdge136[1] ) );
    VMW_NAND2 U102 ( .A(n684), .B(n670), .Z(\OutEdge136[0] ) );
    VMW_AO22 U103 ( .A(\path[1] ), .B(Start), .C(n667), .D(n685), .Z(n704) );
    VMW_OAI21 U104 ( .A(n670), .B(n686), .C(n687), .Z(n702) );
    VMW_OR2 U105 ( .A(n122), .B(n689), .Z(n688) );
    VMW_AO22 U106 ( .A(InEdges[63]), .B(n114), .C(\temp394[15] ), .D(n690), 
        .Z(\temp484[15] ) );
    VMW_INV U107 ( .A(Start), .Z(n670) );
    VMW_OR2 U108 ( .A(Start), .B(n122), .Z(n691) );
    VMW_OAI22 U109 ( .A(\path[2] ), .B(n670), .C(n688), .D(Start), .Z(n692) );
    VMW_INV U110 ( .A(n114), .Z(n690) );
    VMW_INV U111 ( .A(n106), .Z(n693) );
    VMW_NOR4 U112 ( .A(n98), .B(n106), .C(n90), .D(n114), .Z(n689) );
    VMW_OAI211 U113 ( .A(n90), .B(n98), .C(n693), .D(n690), .Z(n685) );
    VMW_OAI21 U114 ( .A(n98), .B(n695), .C(n693), .Z(n694) );
    VMW_AO21 U115 ( .A(n690), .B(n694), .C(n691), .Z(n687) );
    VMW_AND4 U116 ( .A(n696), .B(n697), .C(n698), .D(n699), .Z(n701) );
    VMW_AND3 U117 ( .A(n122), .B(n670), .C(InEdges[79]), .Z(n668) );
    VMW_XNOR2 U118 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n699) );
    VMW_XNOR2 U119 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n698) );
    VMW_XNOR2 U120 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n697) );
    VMW_XNOR2 U121 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n696) );
    VMW_AO22 U122 ( .A(OutEdge[9]), .B(n695), .C(InEdges[9]), .D(n90), .Z(
        \temp210[9] ) );
    VMW_AO22 U123 ( .A(\temp210[9] ), .B(n700), .C(InEdges[25]), .D(n98), .Z(
        \temp304[9] ) );
    VMW_AO22 U124 ( .A(\temp304[9] ), .B(n693), .C(InEdges[41]), .D(n106), .Z(
        \temp394[9] ) );
    VMW_AO22 U125 ( .A(\temp394[9] ), .B(n690), .C(InEdges[57]), .D(n114), .Z(
        \temp484[9] ) );
    VMW_AO22 U126 ( .A(OutEdge[8]), .B(n695), .C(InEdges[8]), .D(n90), .Z(
        \temp210[8] ) );
    VMW_AO22 U127 ( .A(\temp210[8] ), .B(n700), .C(InEdges[24]), .D(n98), .Z(
        \temp304[8] ) );
    VMW_AO22 U128 ( .A(\temp304[8] ), .B(n693), .C(InEdges[40]), .D(n106), .Z(
        \temp394[8] ) );
    VMW_AO22 U129 ( .A(\temp394[8] ), .B(n690), .C(InEdges[56]), .D(n114), .Z(
        \temp484[8] ) );
    VMW_AO22 U130 ( .A(OutEdge[7]), .B(n695), .C(InEdges[7]), .D(n90), .Z(
        \temp210[7] ) );
    VMW_AO22 U131 ( .A(\temp210[7] ), .B(n700), .C(InEdges[23]), .D(n98), .Z(
        \temp304[7] ) );
    VMW_AO22 U132 ( .A(\temp304[7] ), .B(n693), .C(InEdges[39]), .D(n106), .Z(
        \temp394[7] ) );
    VMW_AO22 U133 ( .A(\temp394[7] ), .B(n690), .C(InEdges[55]), .D(n114), .Z(
        \temp484[7] ) );
    VMW_AO22 U134 ( .A(OutEdge[6]), .B(n695), .C(InEdges[6]), .D(n90), .Z(
        \temp210[6] ) );
    VMW_AO22 U135 ( .A(\temp210[6] ), .B(n700), .C(InEdges[22]), .D(n98), .Z(
        \temp304[6] ) );
    VMW_AO22 U136 ( .A(\temp304[6] ), .B(n693), .C(InEdges[38]), .D(n106), .Z(
        \temp394[6] ) );
    VMW_AO22 U137 ( .A(\temp394[6] ), .B(n690), .C(InEdges[54]), .D(n114), .Z(
        \temp484[6] ) );
    VMW_AO22 U138 ( .A(OutEdge[5]), .B(n695), .C(InEdges[5]), .D(n90), .Z(
        \temp210[5] ) );
    VMW_AO22 U139 ( .A(\temp210[5] ), .B(n700), .C(InEdges[21]), .D(n98), .Z(
        \temp304[5] ) );
    VMW_AO22 U140 ( .A(\temp304[5] ), .B(n693), .C(InEdges[37]), .D(n106), .Z(
        \temp394[5] ) );
    VMW_AO22 U141 ( .A(\temp394[5] ), .B(n690), .C(InEdges[53]), .D(n114), .Z(
        \temp484[5] ) );
    VMW_AO22 U142 ( .A(OutEdge[4]), .B(n695), .C(InEdges[4]), .D(n90), .Z(
        \temp210[4] ) );
    VMW_AO22 U143 ( .A(\temp210[4] ), .B(n700), .C(InEdges[20]), .D(n98), .Z(
        \temp304[4] ) );
    VMW_AO22 U144 ( .A(\temp304[4] ), .B(n693), .C(InEdges[36]), .D(n106), .Z(
        \temp394[4] ) );
    VMW_AO22 U145 ( .A(\temp394[4] ), .B(n690), .C(InEdges[52]), .D(n114), .Z(
        \temp484[4] ) );
    VMW_AO22 U146 ( .A(OutEdge[3]), .B(n695), .C(InEdges[3]), .D(n90), .Z(
        \temp210[3] ) );
    VMW_AO22 U147 ( .A(\temp210[3] ), .B(n700), .C(InEdges[19]), .D(n98), .Z(
        \temp304[3] ) );
    VMW_AO22 U148 ( .A(\temp304[3] ), .B(n693), .C(InEdges[35]), .D(n106), .Z(
        \temp394[3] ) );
    VMW_AO22 U149 ( .A(\temp394[3] ), .B(n690), .C(InEdges[51]), .D(n114), .Z(
        \temp484[3] ) );
    VMW_AO22 U150 ( .A(OutEdge[2]), .B(n695), .C(InEdges[2]), .D(n90), .Z(
        \temp210[2] ) );
    VMW_AO22 U151 ( .A(\temp210[2] ), .B(n700), .C(InEdges[18]), .D(n98), .Z(
        \temp304[2] ) );
    VMW_AO22 U152 ( .A(\temp304[2] ), .B(n693), .C(InEdges[34]), .D(n106), .Z(
        \temp394[2] ) );
    VMW_AO22 U153 ( .A(\temp394[2] ), .B(n690), .C(InEdges[50]), .D(n114), .Z(
        \temp484[2] ) );
    VMW_AO22 U154 ( .A(OutEdge[1]), .B(n695), .C(InEdges[1]), .D(n90), .Z(
        \temp210[1] ) );
    VMW_AO22 U155 ( .A(\temp210[1] ), .B(n700), .C(InEdges[17]), .D(n98), .Z(
        \temp304[1] ) );
    VMW_AO22 U156 ( .A(\temp304[1] ), .B(n693), .C(InEdges[33]), .D(n106), .Z(
        \temp394[1] ) );
    VMW_AO22 U157 ( .A(\temp394[1] ), .B(n690), .C(InEdges[49]), .D(n114), .Z(
        \temp484[1] ) );
    VMW_AO22 U158 ( .A(OutEdge[15]), .B(n695), .C(InEdges[15]), .D(n90), .Z(
        \temp210[15] ) );
    VMW_AO22 U159 ( .A(\temp210[15] ), .B(n700), .C(InEdges[31]), .D(n98), .Z(
        \temp304[15] ) );
    VMW_AO22 U160 ( .A(\temp304[15] ), .B(n693), .C(InEdges[47]), .D(n106), 
        .Z(\temp394[15] ) );
    VMW_AO22 U161 ( .A(OutEdge[14]), .B(n695), .C(InEdges[14]), .D(n90), .Z(
        \temp210[14] ) );
    VMW_AO22 U162 ( .A(\temp210[14] ), .B(n700), .C(InEdges[30]), .D(n98), .Z(
        \temp304[14] ) );
    VMW_AO22 U163 ( .A(\temp304[14] ), .B(n693), .C(InEdges[46]), .D(n106), 
        .Z(\temp394[14] ) );
    VMW_AO22 U164 ( .A(\temp394[14] ), .B(n690), .C(InEdges[62]), .D(n114), 
        .Z(\temp484[14] ) );
    VMW_AO22 U165 ( .A(OutEdge[13]), .B(n695), .C(InEdges[13]), .D(n90), .Z(
        \temp210[13] ) );
    VMW_AO22 U166 ( .A(\temp210[13] ), .B(n700), .C(InEdges[29]), .D(n98), .Z(
        \temp304[13] ) );
    VMW_AO22 U167 ( .A(\temp304[13] ), .B(n693), .C(InEdges[45]), .D(n106), 
        .Z(\temp394[13] ) );
    VMW_AO22 U168 ( .A(\temp394[13] ), .B(n690), .C(InEdges[61]), .D(n114), 
        .Z(\temp484[13] ) );
    VMW_AO22 U169 ( .A(OutEdge[12]), .B(n695), .C(InEdges[12]), .D(n90), .Z(
        \temp210[12] ) );
    VMW_AO22 U170 ( .A(\temp210[12] ), .B(n700), .C(InEdges[28]), .D(n98), .Z(
        \temp304[12] ) );
    VMW_AO22 U171 ( .A(\temp304[12] ), .B(n693), .C(InEdges[44]), .D(n106), 
        .Z(\temp394[12] ) );
    VMW_AO22 U172 ( .A(\temp394[12] ), .B(n690), .C(InEdges[60]), .D(n114), 
        .Z(\temp484[12] ) );
    VMW_AO22 U173 ( .A(OutEdge[11]), .B(n695), .C(InEdges[11]), .D(n90), .Z(
        \temp210[11] ) );
    VMW_AO22 U174 ( .A(\temp210[11] ), .B(n700), .C(InEdges[27]), .D(n98), .Z(
        \temp304[11] ) );
    VMW_AO22 U175 ( .A(\temp304[11] ), .B(n693), .C(InEdges[43]), .D(n106), 
        .Z(\temp394[11] ) );
    VMW_AO22 U176 ( .A(\temp394[11] ), .B(n690), .C(InEdges[59]), .D(n114), 
        .Z(\temp484[11] ) );
    VMW_AO22 U177 ( .A(OutEdge[10]), .B(n695), .C(InEdges[10]), .D(n90), .Z(
        \temp210[10] ) );
    VMW_AO22 U178 ( .A(\temp210[10] ), .B(n700), .C(InEdges[26]), .D(n98), .Z(
        \temp304[10] ) );
    VMW_AO22 U179 ( .A(\temp304[10] ), .B(n693), .C(InEdges[42]), .D(n106), 
        .Z(\temp394[10] ) );
    VMW_AO22 U180 ( .A(\temp394[10] ), .B(n690), .C(InEdges[58]), .D(n114), 
        .Z(\temp484[10] ) );
    VMW_AO22 U181 ( .A(OutEdge[0]), .B(n695), .C(InEdges[0]), .D(n90), .Z(
        \temp210[0] ) );
    VMW_AO22 U182 ( .A(\temp210[0] ), .B(n700), .C(InEdges[16]), .D(n98), .Z(
        \temp304[0] ) );
    VMW_AO22 U183 ( .A(\temp304[0] ), .B(n693), .C(InEdges[32]), .D(n106), .Z(
        \temp394[0] ) );
    VMW_AO22 U184 ( .A(\temp394[0] ), .B(n690), .C(InEdges[48]), .D(n114), .Z(
        \temp484[0] ) );
    VMW_MUX2I U185 ( .A(\temp484[9] ), .B(InEdges[73]), .S(n122), .Z(n675) );
    VMW_MUX2I U186 ( .A(\temp484[8] ), .B(InEdges[72]), .S(n122), .Z(n676) );
    VMW_MUX2I U187 ( .A(\temp484[7] ), .B(InEdges[71]), .S(n122), .Z(n677) );
    VMW_MUX2I U188 ( .A(\temp484[6] ), .B(InEdges[70]), .S(n122), .Z(n678) );
    VMW_MUX2I U189 ( .A(\temp484[5] ), .B(InEdges[69]), .S(n122), .Z(n679) );
    VMW_MUX2I U190 ( .A(\temp484[4] ), .B(InEdges[68]), .S(n122), .Z(n680) );
    VMW_MUX2I U191 ( .A(\temp484[3] ), .B(InEdges[67]), .S(n122), .Z(n681) );
    VMW_MUX2I U192 ( .A(\temp484[2] ), .B(InEdges[66]), .S(n122), .Z(n682) );
    VMW_MUX2I U193 ( .A(\temp484[1] ), .B(InEdges[65]), .S(n122), .Z(n683) );
    VMW_MUX2I U194 ( .A(\temp484[14] ), .B(InEdges[78]), .S(n122), .Z(n669) );
    VMW_MUX2I U195 ( .A(\temp484[13] ), .B(InEdges[77]), .S(n122), .Z(n671) );
    VMW_MUX2I U196 ( .A(\temp484[12] ), .B(InEdges[76]), .S(n122), .Z(n672) );
    VMW_MUX2I U197 ( .A(\temp484[11] ), .B(InEdges[75]), .S(n122), .Z(n673) );
    VMW_MUX2I U198 ( .A(\temp484[10] ), .B(InEdges[74]), .S(n122), .Z(n674) );
    VMW_MUX2I U199 ( .A(\temp484[0] ), .B(InEdges[64]), .S(n122), .Z(n684) );
    VMW_INV U200 ( .A(n90), .Z(n695) );
    VMW_INV U201 ( .A(n98), .Z(n700) );
    VMW_INV U202 ( .A(n691), .Z(n667) );
    VMW_INV U203 ( .A(n692), .Z(n703) );
    VMW_INV U204 ( .A(\path[0] ), .Z(n686) );
    VMW_BUFIZ U205 ( .A(\path[1] ), .E(n701), .Z(\PathData[1] ) );
    VMW_BUFIZ U206 ( .A(\path[0] ), .E(n701), .Z(\PathData[0] ) );
    VMW_BUFIZ U207 ( .A(\path[2] ), .E(n701), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n702), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n703), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n704), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge136[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge136[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge136[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge136[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge136[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge136[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge136[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge136[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge136[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge136[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge136[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge136[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge136[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge136[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge136[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge136[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_4 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n709), .TC(n709), .GE_GT(n90) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_3 lte_55_4 ( .A({\temp484[15] , 
        \temp484[14] , \temp484[13] , \temp484[12] , \temp484[11] , 
        \temp484[10] , \temp484[9] , \temp484[8] , \temp484[7] , \temp484[6] , 
        \temp484[5] , \temp484[4] , \temp484[3] , \temp484[2] , \temp484[1] , 
        \temp484[0] }), .B(InEdges[79:64]), .LEQ(n708), .TC(n708), .GE_GT(n122
        ) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_2 lte_55_2 ( .A({\temp304[15] , 
        \temp304[14] , \temp304[13] , \temp304[12] , \temp304[11] , 
        \temp304[10] , \temp304[9] , \temp304[8] , \temp304[7] , \temp304[6] , 
        \temp304[5] , \temp304[4] , \temp304[3] , \temp304[2] , \temp304[1] , 
        \temp304[0] }), .B(InEdges[47:32]), .LEQ(n707), .TC(n707), .GE_GT(n106
        ) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_1 lte_55_1 ( .A({\temp210[15] , 
        \temp210[14] , \temp210[13] , \temp210[12] , \temp210[11] , 
        \temp210[10] , \temp210[9] , \temp210[8] , \temp210[7] , \temp210[6] , 
        \temp210[5] , \temp210[4] , \temp210[3] , \temp210[2] , \temp210[1] , 
        \temp210[0] }), .B(InEdges[31:16]), .LEQ(n706), .TC(n706), .GE_GT(n98)
         );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp394[15] , 
        \temp394[14] , \temp394[13] , \temp394[12] , \temp394[11] , 
        \temp394[10] , \temp394[9] , \temp394[8] , \temp394[7] , \temp394[6] , 
        \temp394[5] , \temp394[4] , \temp394[3] , \temp394[2] , \temp394[1] , 
        \temp394[0] }), .B(InEdges[63:48]), .LEQ(n705), .TC(n705), .GE_GT(n114
        ) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n93, n94, n95, n96, n97, n98, n99, n101, n102, n103, n104, n105, n106, 
        n107, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n91), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n99), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n107), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n125, n126, n127, n128, 
        n129, n130, n131, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
        n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
        n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
        n166, n167;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n134), .C(n131), .D(n129), .Z(n133) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n133), .D(n127), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n145), .C(n140), .D(n135), .Z(n144) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n146) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n148), .C(n146), .D(n144), .Z(n147) );
    VMW_NAND2 U20 ( .A(n150), .B(B[10]), .Z(n149) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n152), .C(n147), .D(n142), .Z(n151) );
    VMW_NAND2 U22 ( .A(n152), .B(A[9]), .Z(n153) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U24 ( .A(n156), .B(B[12]), .Z(n155) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_NAND2 U26 ( .A(n158), .B(A[11]), .Z(n159) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_NAND2 U28 ( .A(n162), .B(B[14]), .Z(n161) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_NAND2 U30 ( .A(n164), .B(A[13]), .Z(n165) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n162), .C(n165), .D(n163), .Z(n166) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n167), .C(n166), .D(n161), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n156) );
    VMW_INV U34 ( .A(B[7]), .Z(n145) );
    VMW_INV U35 ( .A(A[7]), .Z(n148) );
    VMW_INV U36 ( .A(A[3]), .Z(n134) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n150) );
    VMW_INV U39 ( .A(B[9]), .Z(n152) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n143) );
    VMW_INV U42 ( .A(A[14]), .Z(n162) );
    VMW_INV U43 ( .A(B[11]), .Z(n158) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n167) );
    VMW_INV U48 ( .A(B[13]), .Z(n164) );
    VMW_INV U49 ( .A(A[6]), .Z(n136) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
        n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216;
    VMW_OAI21 U3 ( .A(B[15]), .B(n168), .C(n169), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n171), .B(B[2]), .Z(n170) );
    VMW_AO22 U5 ( .A(n173), .B(B[0]), .C(n174), .D(B[1]), .Z(n172) );
    VMW_OR2 U6 ( .A(B[2]), .B(n171), .Z(n175) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n174), .C(n175), .D(n172), .Z(n176) );
    VMW_NAND2 U8 ( .A(n178), .B(B[4]), .Z(n177) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n180), .C(n176), .D(n170), .Z(n179) );
    VMW_OR2 U10 ( .A(B[4]), .B(n178), .Z(n181) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n183), .C(n181), .D(n179), .Z(n182) );
    VMW_NAND2 U12 ( .A(n185), .B(B[6]), .Z(n184) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n187), .C(n182), .D(n177), .Z(n186) );
    VMW_OR2 U14 ( .A(B[6]), .B(n185), .Z(n188) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n190), .C(n188), .D(n186), .Z(n189) );
    VMW_NAND2 U16 ( .A(n192), .B(B[8]), .Z(n191) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n194), .C(n189), .D(n184), .Z(n193) );
    VMW_OR2 U18 ( .A(B[8]), .B(n192), .Z(n195) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n197), .C(n195), .D(n193), .Z(n196) );
    VMW_NAND2 U20 ( .A(n199), .B(B[10]), .Z(n198) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n201), .C(n196), .D(n191), .Z(n200) );
    VMW_NAND2 U22 ( .A(n201), .B(A[9]), .Z(n202) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n199), .C(n202), .D(n200), .Z(n203) );
    VMW_NAND2 U24 ( .A(n205), .B(B[12]), .Z(n204) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n207), .C(n203), .D(n198), .Z(n206) );
    VMW_NAND2 U26 ( .A(n207), .B(A[11]), .Z(n208) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n205), .C(n208), .D(n206), .Z(n209) );
    VMW_NAND2 U28 ( .A(n211), .B(B[14]), .Z(n210) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n213), .C(n209), .D(n204), .Z(n212) );
    VMW_NAND2 U30 ( .A(n213), .B(A[13]), .Z(n214) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n211), .C(n214), .D(n212), .Z(n215) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n216), .C(n215), .D(n210), .Z(n169) );
    VMW_INV U33 ( .A(A[12]), .Z(n205) );
    VMW_INV U34 ( .A(B[7]), .Z(n194) );
    VMW_INV U35 ( .A(A[7]), .Z(n197) );
    VMW_INV U36 ( .A(A[3]), .Z(n183) );
    VMW_INV U37 ( .A(B[3]), .Z(n180) );
    VMW_INV U38 ( .A(A[10]), .Z(n199) );
    VMW_INV U39 ( .A(B[9]), .Z(n201) );
    VMW_INV U40 ( .A(A[4]), .Z(n178) );
    VMW_INV U41 ( .A(A[8]), .Z(n192) );
    VMW_INV U42 ( .A(A[14]), .Z(n211) );
    VMW_INV U43 ( .A(B[11]), .Z(n207) );
    VMW_INV U44 ( .A(A[5]), .Z(n190) );
    VMW_INV U45 ( .A(B[5]), .Z(n187) );
    VMW_INV U46 ( .A(A[1]), .Z(n174) );
    VMW_INV U47 ( .A(B[15]), .Z(n216) );
    VMW_INV U48 ( .A(B[13]), .Z(n213) );
    VMW_INV U49 ( .A(A[6]), .Z(n185) );
    VMW_INV U50 ( .A(A[2]), .Z(n171) );
    VMW_INV U51 ( .A(A[0]), .Z(n173) );
    VMW_INV U52 ( .A(A[15]), .Z(n168) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
        n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265;
    VMW_OAI21 U3 ( .A(B[15]), .B(n217), .C(n218), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n220), .B(B[2]), .Z(n219) );
    VMW_AO22 U5 ( .A(n222), .B(B[0]), .C(n223), .D(B[1]), .Z(n221) );
    VMW_OR2 U6 ( .A(B[2]), .B(n220), .Z(n224) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n223), .C(n224), .D(n221), .Z(n225) );
    VMW_NAND2 U8 ( .A(n227), .B(B[4]), .Z(n226) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n229), .C(n225), .D(n219), .Z(n228) );
    VMW_OR2 U10 ( .A(B[4]), .B(n227), .Z(n230) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n232), .C(n230), .D(n228), .Z(n231) );
    VMW_NAND2 U12 ( .A(n234), .B(B[6]), .Z(n233) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n236), .C(n231), .D(n226), .Z(n235) );
    VMW_OR2 U14 ( .A(B[6]), .B(n234), .Z(n237) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n239), .C(n237), .D(n235), .Z(n238) );
    VMW_NAND2 U16 ( .A(n241), .B(B[8]), .Z(n240) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n243), .C(n238), .D(n233), .Z(n242) );
    VMW_OR2 U18 ( .A(B[8]), .B(n241), .Z(n244) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n246), .C(n244), .D(n242), .Z(n245) );
    VMW_NAND2 U20 ( .A(n248), .B(B[10]), .Z(n247) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n250), .C(n245), .D(n240), .Z(n249) );
    VMW_NAND2 U22 ( .A(n250), .B(A[9]), .Z(n251) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n248), .C(n251), .D(n249), .Z(n252) );
    VMW_NAND2 U24 ( .A(n254), .B(B[12]), .Z(n253) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n256), .C(n252), .D(n247), .Z(n255) );
    VMW_NAND2 U26 ( .A(n256), .B(A[11]), .Z(n257) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n254), .C(n257), .D(n255), .Z(n258) );
    VMW_NAND2 U28 ( .A(n260), .B(B[14]), .Z(n259) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n262), .C(n258), .D(n253), .Z(n261) );
    VMW_NAND2 U30 ( .A(n262), .B(A[13]), .Z(n263) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n260), .C(n263), .D(n261), .Z(n264) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n265), .C(n264), .D(n259), .Z(n218) );
    VMW_INV U33 ( .A(A[12]), .Z(n254) );
    VMW_INV U34 ( .A(B[7]), .Z(n243) );
    VMW_INV U35 ( .A(A[7]), .Z(n246) );
    VMW_INV U36 ( .A(A[3]), .Z(n232) );
    VMW_INV U37 ( .A(B[3]), .Z(n229) );
    VMW_INV U38 ( .A(A[10]), .Z(n248) );
    VMW_INV U39 ( .A(B[9]), .Z(n250) );
    VMW_INV U40 ( .A(A[4]), .Z(n227) );
    VMW_INV U41 ( .A(A[8]), .Z(n241) );
    VMW_INV U42 ( .A(A[14]), .Z(n260) );
    VMW_INV U43 ( .A(B[11]), .Z(n256) );
    VMW_INV U44 ( .A(A[5]), .Z(n239) );
    VMW_INV U45 ( .A(B[5]), .Z(n236) );
    VMW_INV U46 ( .A(A[1]), .Z(n223) );
    VMW_INV U47 ( .A(B[15]), .Z(n265) );
    VMW_INV U48 ( .A(B[13]), .Z(n262) );
    VMW_INV U49 ( .A(A[6]), .Z(n234) );
    VMW_INV U50 ( .A(A[2]), .Z(n220) );
    VMW_INV U51 ( .A(A[0]), .Z(n222) );
    VMW_INV U52 ( .A(A[15]), .Z(n217) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
        n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
        n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
        n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
        n313, n314;
    VMW_OAI21 U3 ( .A(B[15]), .B(n266), .C(n267), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n269), .B(B[2]), .Z(n268) );
    VMW_AO22 U5 ( .A(n271), .B(B[0]), .C(n272), .D(B[1]), .Z(n270) );
    VMW_OR2 U6 ( .A(B[2]), .B(n269), .Z(n273) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n272), .C(n273), .D(n270), .Z(n274) );
    VMW_NAND2 U8 ( .A(n276), .B(B[4]), .Z(n275) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n278), .C(n274), .D(n268), .Z(n277) );
    VMW_OR2 U10 ( .A(B[4]), .B(n276), .Z(n279) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n281), .C(n279), .D(n277), .Z(n280) );
    VMW_NAND2 U12 ( .A(n283), .B(B[6]), .Z(n282) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n285), .C(n280), .D(n275), .Z(n284) );
    VMW_OR2 U14 ( .A(B[6]), .B(n283), .Z(n286) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n288), .C(n286), .D(n284), .Z(n287) );
    VMW_NAND2 U16 ( .A(n290), .B(B[8]), .Z(n289) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n292), .C(n287), .D(n282), .Z(n291) );
    VMW_OR2 U18 ( .A(B[8]), .B(n290), .Z(n293) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n295), .C(n293), .D(n291), .Z(n294) );
    VMW_NAND2 U20 ( .A(n297), .B(B[10]), .Z(n296) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n299), .C(n294), .D(n289), .Z(n298) );
    VMW_NAND2 U22 ( .A(n299), .B(A[9]), .Z(n300) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n297), .C(n300), .D(n298), .Z(n301) );
    VMW_NAND2 U24 ( .A(n303), .B(B[12]), .Z(n302) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n305), .C(n301), .D(n296), .Z(n304) );
    VMW_NAND2 U26 ( .A(n305), .B(A[11]), .Z(n306) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n303), .C(n306), .D(n304), .Z(n307) );
    VMW_NAND2 U28 ( .A(n309), .B(B[14]), .Z(n308) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n311), .C(n307), .D(n302), .Z(n310) );
    VMW_NAND2 U30 ( .A(n311), .B(A[13]), .Z(n312) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n309), .C(n312), .D(n310), .Z(n313) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n314), .C(n313), .D(n308), .Z(n267) );
    VMW_INV U33 ( .A(A[12]), .Z(n303) );
    VMW_INV U34 ( .A(B[7]), .Z(n292) );
    VMW_INV U35 ( .A(A[7]), .Z(n295) );
    VMW_INV U36 ( .A(A[3]), .Z(n281) );
    VMW_INV U37 ( .A(B[3]), .Z(n278) );
    VMW_INV U38 ( .A(A[10]), .Z(n297) );
    VMW_INV U39 ( .A(B[9]), .Z(n299) );
    VMW_INV U40 ( .A(A[4]), .Z(n276) );
    VMW_INV U41 ( .A(A[8]), .Z(n290) );
    VMW_INV U42 ( .A(A[14]), .Z(n309) );
    VMW_INV U43 ( .A(B[11]), .Z(n305) );
    VMW_INV U44 ( .A(A[5]), .Z(n288) );
    VMW_INV U45 ( .A(B[5]), .Z(n285) );
    VMW_INV U46 ( .A(A[1]), .Z(n272) );
    VMW_INV U47 ( .A(B[15]), .Z(n314) );
    VMW_INV U48 ( .A(B[13]), .Z(n311) );
    VMW_INV U49 ( .A(A[6]), .Z(n283) );
    VMW_INV U50 ( .A(A[2]), .Z(n269) );
    VMW_INV U51 ( .A(A[0]), .Z(n271) );
    VMW_INV U52 ( .A(A[15]), .Z(n266) );
endmodule


module NodeAux_INDEGREE6_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [3:0] Nid;
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp494[7] , \temp584[2] , n100, \OutEdge146[7] , \temp314[15] , 
        \OutEdge146[12] , \temp314[11] , \OutEdge146[3] , \temp494[3] , 
        \temp584[6] , \path[2] , \path[0] , \temp314[13] , \temp494[1] , 
        \OutEdge146[1] , \temp584[4] , \OutEdge146[8] , \temp494[8] , n132, 
        \OutEdge146[10] , \temp584[0] , \OutEdge146[5] , \temp494[5] , 
        \OutEdge146[14] , \temp584[9] , \temp220[10] , \temp220[4] , 
        \temp314[7] , \temp494[11] , \temp404[6] , \temp584[13] , 
        \temp404[11] , \temp404[2] , \temp220[0] , \temp314[3] , \temp494[15] , 
        \temp220[14] , \temp404[15] , \temp220[9] , \temp404[9] , \temp314[8] , 
        \temp220[2] , \temp404[0] , \temp314[1] , \temp584[15] , n108, 
        \temp404[13] , \temp584[11] , \temp220[12] , \temp220[6] , 
        \temp314[5] , \temp404[4] , \temp494[13] , \temp404[12] , 
        \temp584[10] , \temp220[7] , \temp314[4] , n124, \temp494[12] , 
        \temp220[13] , \temp404[5] , \temp404[8] , \temp314[9] , \temp404[1] , 
        \temp220[3] , \temp314[0] , \temp584[14] , \temp404[3] , \temp220[15] , 
        \temp220[1] , \temp314[2] , \temp494[14] , \temp220[8] , \temp404[14] , 
        n116, \temp220[5] , \temp314[6] , \temp494[10] , \temp220[11] , 
        \temp404[7] , \temp584[12] , \temp404[10] , \temp584[1] , 
        \OutEdge146[4] , \temp494[4] , \OutEdge146[15] , \temp584[8] , 
        \path[1] , \temp494[0] , \OutEdge146[0] , \temp314[12] , n92, 
        \temp584[5] , \OutEdge146[9] , \temp494[9] , \OutEdge146[11] , 
        \OutEdge146[13] , \temp494[2] , \OutEdge146[2] , \temp314[10] , 
        \temp584[7] , \temp584[3] , \temp314[14] , \temp494[6] , 
        \OutEdge146[6] , n767, n768, n769, n770, n771, n772, n773, n774, n775, 
        n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
        n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
        n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
        n812;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U91 ( .Z(n811) );
    VMW_PULLDOWN U92 ( .Z(n810) );
    VMW_PULLDOWN U93 ( .Z(n809) );
    VMW_PULLDOWN U94 ( .Z(n808) );
    VMW_PULLDOWN U95 ( .Z(n812) );
    VMW_PULLDOWN U96 ( .Z(n807) );
    VMW_NOR2 U97 ( .A(Start), .B(n767), .Z(\OutEdge146[15] ) );
    VMW_NAND2 U98 ( .A(n768), .B(n769), .Z(\OutEdge146[14] ) );
    VMW_NAND2 U99 ( .A(n770), .B(n769), .Z(\OutEdge146[13] ) );
    VMW_NAND2 U100 ( .A(n771), .B(n769), .Z(\OutEdge146[12] ) );
    VMW_NAND2 U101 ( .A(n772), .B(n769), .Z(\OutEdge146[11] ) );
    VMW_NAND2 U102 ( .A(n773), .B(n769), .Z(\OutEdge146[10] ) );
    VMW_NAND2 U103 ( .A(n774), .B(n769), .Z(\OutEdge146[9] ) );
    VMW_NAND2 U104 ( .A(n775), .B(n769), .Z(\OutEdge146[8] ) );
    VMW_NAND2 U105 ( .A(n776), .B(n769), .Z(\OutEdge146[7] ) );
    VMW_NAND2 U106 ( .A(n777), .B(n769), .Z(\OutEdge146[6] ) );
    VMW_NAND2 U107 ( .A(n778), .B(n769), .Z(\OutEdge146[5] ) );
    VMW_NAND2 U108 ( .A(n779), .B(n769), .Z(\OutEdge146[4] ) );
    VMW_NAND2 U109 ( .A(n780), .B(n769), .Z(\OutEdge146[3] ) );
    VMW_NAND2 U110 ( .A(n781), .B(n769), .Z(\OutEdge146[2] ) );
    VMW_NAND2 U111 ( .A(n782), .B(n769), .Z(\OutEdge146[1] ) );
    VMW_NAND2 U112 ( .A(n783), .B(n769), .Z(\OutEdge146[0] ) );
    VMW_AND4 U113 ( .A(n785), .B(n786), .C(n787), .D(n788), .Z(n784) );
    VMW_OR3 U114 ( .A(n784), .B(n124), .C(n132), .Z(n789) );
    VMW_OR2 U115 ( .A(n132), .B(n791), .Z(n790) );
    VMW_AO22 U116 ( .A(\temp494[15] ), .B(n792), .C(InEdges[79]), .D(n124), 
        .Z(\temp584[15] ) );
    VMW_OAI22 U117 ( .A(\path[2] ), .B(n769), .C(n789), .D(Start), .Z(n793) );
    VMW_OAI22 U118 ( .A(\path[1] ), .B(n769), .C(n795), .D(Start), .Z(n794) );
    VMW_OAI22 U119 ( .A(\path[0] ), .B(n769), .C(n790), .D(Start), .Z(n796) );
    VMW_MUX2I U120 ( .A(\temp584[15] ), .B(InEdges[95]), .S(n132), .Z(n767) );
    VMW_INV U121 ( .A(Start), .Z(n769) );
    VMW_INV U122 ( .A(n116), .Z(n786) );
    VMW_AOI211 U123 ( .A(n785), .B(n787), .C(n108), .D(n116), .Z(n797) );
    VMW_OAI21 U124 ( .A(n100), .B(n785), .C(n788), .Z(n798) );
    VMW_AOI21 U125 ( .A(n786), .B(n798), .C(n124), .Z(n791) );
    VMW_AND4 U126 ( .A(n799), .B(n800), .C(n801), .D(n802), .Z(n803) );
    VMW_XNOR2 U127 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n802) );
    VMW_XNOR2 U128 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n801) );
    VMW_XNOR2 U129 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n800) );
    VMW_XNOR2 U130 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n799) );
    VMW_AO22 U131 ( .A(OutEdge[9]), .B(n785), .C(InEdges[9]), .D(n92), .Z(
        \temp220[9] ) );
    VMW_AO22 U132 ( .A(\temp220[9] ), .B(n787), .C(InEdges[25]), .D(n100), .Z(
        \temp314[9] ) );
    VMW_AO22 U133 ( .A(\temp314[9] ), .B(n788), .C(InEdges[41]), .D(n108), .Z(
        \temp404[9] ) );
    VMW_AO22 U134 ( .A(\temp404[9] ), .B(n786), .C(InEdges[57]), .D(n116), .Z(
        \temp494[9] ) );
    VMW_AO22 U135 ( .A(\temp494[9] ), .B(n792), .C(InEdges[73]), .D(n124), .Z(
        \temp584[9] ) );
    VMW_AO22 U136 ( .A(OutEdge[8]), .B(n785), .C(InEdges[8]), .D(n92), .Z(
        \temp220[8] ) );
    VMW_AO22 U137 ( .A(\temp220[8] ), .B(n787), .C(InEdges[24]), .D(n100), .Z(
        \temp314[8] ) );
    VMW_AO22 U138 ( .A(\temp314[8] ), .B(n788), .C(InEdges[40]), .D(n108), .Z(
        \temp404[8] ) );
    VMW_AO22 U139 ( .A(\temp404[8] ), .B(n786), .C(InEdges[56]), .D(n116), .Z(
        \temp494[8] ) );
    VMW_AO22 U140 ( .A(\temp494[8] ), .B(n792), .C(InEdges[72]), .D(n124), .Z(
        \temp584[8] ) );
    VMW_AO22 U141 ( .A(OutEdge[7]), .B(n785), .C(InEdges[7]), .D(n92), .Z(
        \temp220[7] ) );
    VMW_AO22 U142 ( .A(\temp220[7] ), .B(n787), .C(InEdges[23]), .D(n100), .Z(
        \temp314[7] ) );
    VMW_AO22 U143 ( .A(\temp314[7] ), .B(n788), .C(InEdges[39]), .D(n108), .Z(
        \temp404[7] ) );
    VMW_AO22 U144 ( .A(\temp404[7] ), .B(n786), .C(InEdges[55]), .D(n116), .Z(
        \temp494[7] ) );
    VMW_AO22 U145 ( .A(\temp494[7] ), .B(n792), .C(InEdges[71]), .D(n124), .Z(
        \temp584[7] ) );
    VMW_AO22 U146 ( .A(OutEdge[6]), .B(n785), .C(InEdges[6]), .D(n92), .Z(
        \temp220[6] ) );
    VMW_AO22 U147 ( .A(\temp220[6] ), .B(n787), .C(InEdges[22]), .D(n100), .Z(
        \temp314[6] ) );
    VMW_AO22 U148 ( .A(\temp314[6] ), .B(n788), .C(InEdges[38]), .D(n108), .Z(
        \temp404[6] ) );
    VMW_AO22 U149 ( .A(\temp404[6] ), .B(n786), .C(InEdges[54]), .D(n116), .Z(
        \temp494[6] ) );
    VMW_AO22 U150 ( .A(\temp494[6] ), .B(n792), .C(InEdges[70]), .D(n124), .Z(
        \temp584[6] ) );
    VMW_AO22 U151 ( .A(OutEdge[5]), .B(n785), .C(InEdges[5]), .D(n92), .Z(
        \temp220[5] ) );
    VMW_AO22 U152 ( .A(\temp220[5] ), .B(n787), .C(InEdges[21]), .D(n100), .Z(
        \temp314[5] ) );
    VMW_AO22 U153 ( .A(\temp314[5] ), .B(n788), .C(InEdges[37]), .D(n108), .Z(
        \temp404[5] ) );
    VMW_AO22 U154 ( .A(\temp404[5] ), .B(n786), .C(InEdges[53]), .D(n116), .Z(
        \temp494[5] ) );
    VMW_AO22 U155 ( .A(\temp494[5] ), .B(n792), .C(InEdges[69]), .D(n124), .Z(
        \temp584[5] ) );
    VMW_AO22 U156 ( .A(OutEdge[4]), .B(n785), .C(InEdges[4]), .D(n92), .Z(
        \temp220[4] ) );
    VMW_AO22 U157 ( .A(\temp220[4] ), .B(n787), .C(InEdges[20]), .D(n100), .Z(
        \temp314[4] ) );
    VMW_AO22 U158 ( .A(\temp314[4] ), .B(n788), .C(InEdges[36]), .D(n108), .Z(
        \temp404[4] ) );
    VMW_AO22 U159 ( .A(\temp404[4] ), .B(n786), .C(InEdges[52]), .D(n116), .Z(
        \temp494[4] ) );
    VMW_AO22 U160 ( .A(\temp494[4] ), .B(n792), .C(InEdges[68]), .D(n124), .Z(
        \temp584[4] ) );
    VMW_AO22 U161 ( .A(OutEdge[3]), .B(n785), .C(InEdges[3]), .D(n92), .Z(
        \temp220[3] ) );
    VMW_AO22 U162 ( .A(\temp220[3] ), .B(n787), .C(InEdges[19]), .D(n100), .Z(
        \temp314[3] ) );
    VMW_AO22 U163 ( .A(\temp314[3] ), .B(n788), .C(InEdges[35]), .D(n108), .Z(
        \temp404[3] ) );
    VMW_AO22 U164 ( .A(\temp404[3] ), .B(n786), .C(InEdges[51]), .D(n116), .Z(
        \temp494[3] ) );
    VMW_AO22 U165 ( .A(\temp494[3] ), .B(n792), .C(InEdges[67]), .D(n124), .Z(
        \temp584[3] ) );
    VMW_AO22 U166 ( .A(OutEdge[2]), .B(n785), .C(InEdges[2]), .D(n92), .Z(
        \temp220[2] ) );
    VMW_AO22 U167 ( .A(\temp220[2] ), .B(n787), .C(InEdges[18]), .D(n100), .Z(
        \temp314[2] ) );
    VMW_AO22 U168 ( .A(\temp314[2] ), .B(n788), .C(InEdges[34]), .D(n108), .Z(
        \temp404[2] ) );
    VMW_AO22 U169 ( .A(\temp404[2] ), .B(n786), .C(InEdges[50]), .D(n116), .Z(
        \temp494[2] ) );
    VMW_AO22 U170 ( .A(\temp494[2] ), .B(n792), .C(InEdges[66]), .D(n124), .Z(
        \temp584[2] ) );
    VMW_AO22 U171 ( .A(OutEdge[1]), .B(n785), .C(InEdges[1]), .D(n92), .Z(
        \temp220[1] ) );
    VMW_AO22 U172 ( .A(\temp220[1] ), .B(n787), .C(InEdges[17]), .D(n100), .Z(
        \temp314[1] ) );
    VMW_AO22 U173 ( .A(\temp314[1] ), .B(n788), .C(InEdges[33]), .D(n108), .Z(
        \temp404[1] ) );
    VMW_AO22 U174 ( .A(\temp404[1] ), .B(n786), .C(InEdges[49]), .D(n116), .Z(
        \temp494[1] ) );
    VMW_AO22 U175 ( .A(\temp494[1] ), .B(n792), .C(InEdges[65]), .D(n124), .Z(
        \temp584[1] ) );
    VMW_AO22 U176 ( .A(OutEdge[15]), .B(n785), .C(InEdges[15]), .D(n92), .Z(
        \temp220[15] ) );
    VMW_AO22 U177 ( .A(\temp220[15] ), .B(n787), .C(InEdges[31]), .D(n100), 
        .Z(\temp314[15] ) );
    VMW_AO22 U178 ( .A(\temp314[15] ), .B(n788), .C(InEdges[47]), .D(n108), 
        .Z(\temp404[15] ) );
    VMW_AO22 U179 ( .A(\temp404[15] ), .B(n786), .C(InEdges[63]), .D(n116), 
        .Z(\temp494[15] ) );
    VMW_AO22 U180 ( .A(OutEdge[14]), .B(n785), .C(InEdges[14]), .D(n92), .Z(
        \temp220[14] ) );
    VMW_AO22 U181 ( .A(\temp220[14] ), .B(n787), .C(InEdges[30]), .D(n100), 
        .Z(\temp314[14] ) );
    VMW_AO22 U182 ( .A(\temp314[14] ), .B(n788), .C(InEdges[46]), .D(n108), 
        .Z(\temp404[14] ) );
    VMW_AO22 U183 ( .A(\temp404[14] ), .B(n786), .C(InEdges[62]), .D(n116), 
        .Z(\temp494[14] ) );
    VMW_AO22 U184 ( .A(\temp494[14] ), .B(n792), .C(InEdges[78]), .D(n124), 
        .Z(\temp584[14] ) );
    VMW_AO22 U185 ( .A(OutEdge[13]), .B(n785), .C(InEdges[13]), .D(n92), .Z(
        \temp220[13] ) );
    VMW_AO22 U186 ( .A(\temp220[13] ), .B(n787), .C(InEdges[29]), .D(n100), 
        .Z(\temp314[13] ) );
    VMW_AO22 U187 ( .A(\temp314[13] ), .B(n788), .C(InEdges[45]), .D(n108), 
        .Z(\temp404[13] ) );
    VMW_AO22 U188 ( .A(\temp404[13] ), .B(n786), .C(InEdges[61]), .D(n116), 
        .Z(\temp494[13] ) );
    VMW_AO22 U189 ( .A(\temp494[13] ), .B(n792), .C(InEdges[77]), .D(n124), 
        .Z(\temp584[13] ) );
    VMW_AO22 U190 ( .A(OutEdge[12]), .B(n785), .C(InEdges[12]), .D(n92), .Z(
        \temp220[12] ) );
    VMW_AO22 U191 ( .A(\temp220[12] ), .B(n787), .C(InEdges[28]), .D(n100), 
        .Z(\temp314[12] ) );
    VMW_AO22 U192 ( .A(\temp314[12] ), .B(n788), .C(InEdges[44]), .D(n108), 
        .Z(\temp404[12] ) );
    VMW_AO22 U193 ( .A(\temp404[12] ), .B(n786), .C(InEdges[60]), .D(n116), 
        .Z(\temp494[12] ) );
    VMW_AO22 U194 ( .A(\temp494[12] ), .B(n792), .C(InEdges[76]), .D(n124), 
        .Z(\temp584[12] ) );
    VMW_AO22 U195 ( .A(OutEdge[11]), .B(n785), .C(InEdges[11]), .D(n92), .Z(
        \temp220[11] ) );
    VMW_AO22 U196 ( .A(\temp220[11] ), .B(n787), .C(InEdges[27]), .D(n100), 
        .Z(\temp314[11] ) );
    VMW_AO22 U197 ( .A(\temp314[11] ), .B(n788), .C(InEdges[43]), .D(n108), 
        .Z(\temp404[11] ) );
    VMW_AO22 U198 ( .A(\temp404[11] ), .B(n786), .C(InEdges[59]), .D(n116), 
        .Z(\temp494[11] ) );
    VMW_AO22 U199 ( .A(\temp494[11] ), .B(n792), .C(InEdges[75]), .D(n124), 
        .Z(\temp584[11] ) );
    VMW_AO22 U200 ( .A(OutEdge[10]), .B(n785), .C(InEdges[10]), .D(n92), .Z(
        \temp220[10] ) );
    VMW_AO22 U201 ( .A(\temp220[10] ), .B(n787), .C(InEdges[26]), .D(n100), 
        .Z(\temp314[10] ) );
    VMW_AO22 U202 ( .A(\temp314[10] ), .B(n788), .C(InEdges[42]), .D(n108), 
        .Z(\temp404[10] ) );
    VMW_AO22 U203 ( .A(\temp404[10] ), .B(n786), .C(InEdges[58]), .D(n116), 
        .Z(\temp494[10] ) );
    VMW_AO22 U204 ( .A(\temp494[10] ), .B(n792), .C(InEdges[74]), .D(n124), 
        .Z(\temp584[10] ) );
    VMW_AO22 U205 ( .A(OutEdge[0]), .B(n785), .C(InEdges[0]), .D(n92), .Z(
        \temp220[0] ) );
    VMW_AO22 U206 ( .A(\temp220[0] ), .B(n787), .C(InEdges[16]), .D(n100), .Z(
        \temp314[0] ) );
    VMW_AO22 U207 ( .A(\temp314[0] ), .B(n788), .C(InEdges[32]), .D(n108), .Z(
        \temp404[0] ) );
    VMW_AO22 U208 ( .A(\temp404[0] ), .B(n786), .C(InEdges[48]), .D(n116), .Z(
        \temp494[0] ) );
    VMW_AO22 U209 ( .A(\temp494[0] ), .B(n792), .C(InEdges[64]), .D(n124), .Z(
        \temp584[0] ) );
    VMW_NOR3 U210 ( .A(n132), .B(n124), .C(n797), .Z(n795) );
    VMW_MUX2I U211 ( .A(\temp584[9] ), .B(InEdges[89]), .S(n132), .Z(n774) );
    VMW_MUX2I U212 ( .A(\temp584[8] ), .B(InEdges[88]), .S(n132), .Z(n775) );
    VMW_MUX2I U213 ( .A(\temp584[7] ), .B(InEdges[87]), .S(n132), .Z(n776) );
    VMW_MUX2I U214 ( .A(\temp584[6] ), .B(InEdges[86]), .S(n132), .Z(n777) );
    VMW_MUX2I U215 ( .A(\temp584[5] ), .B(InEdges[85]), .S(n132), .Z(n778) );
    VMW_MUX2I U216 ( .A(\temp584[4] ), .B(InEdges[84]), .S(n132), .Z(n779) );
    VMW_MUX2I U217 ( .A(\temp584[3] ), .B(InEdges[83]), .S(n132), .Z(n780) );
    VMW_MUX2I U218 ( .A(\temp584[2] ), .B(InEdges[82]), .S(n132), .Z(n781) );
    VMW_MUX2I U219 ( .A(\temp584[1] ), .B(InEdges[81]), .S(n132), .Z(n782) );
    VMW_MUX2I U220 ( .A(\temp584[14] ), .B(InEdges[94]), .S(n132), .Z(n768) );
    VMW_MUX2I U221 ( .A(\temp584[13] ), .B(InEdges[93]), .S(n132), .Z(n770) );
    VMW_MUX2I U222 ( .A(\temp584[12] ), .B(InEdges[92]), .S(n132), .Z(n771) );
    VMW_MUX2I U223 ( .A(\temp584[11] ), .B(InEdges[91]), .S(n132), .Z(n772) );
    VMW_MUX2I U224 ( .A(\temp584[10] ), .B(InEdges[90]), .S(n132), .Z(n773) );
    VMW_MUX2I U225 ( .A(\temp584[0] ), .B(InEdges[80]), .S(n132), .Z(n783) );
    VMW_INV U226 ( .A(n100), .Z(n787) );
    VMW_INV U227 ( .A(n92), .Z(n785) );
    VMW_INV U228 ( .A(n108), .Z(n788) );
    VMW_INV U229 ( .A(n124), .Z(n792) );
    VMW_INV U230 ( .A(n793), .Z(n805) );
    VMW_INV U231 ( .A(n794), .Z(n806) );
    VMW_INV U232 ( .A(n796), .Z(n804) );
    VMW_BUFIZ U233 ( .A(\path[1] ), .E(n803), .Z(\PathData[1] ) );
    VMW_BUFIZ U234 ( .A(\path[0] ), .E(n803), .Z(\PathData[0] ) );
    VMW_BUFIZ U235 ( .A(\path[2] ), .E(n803), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n804), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n805), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n806), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge146[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge146[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge146[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge146[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge146[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge146[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge146[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge146[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge146[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge146[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge146[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge146[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge146[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge146[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge146[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge146[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_5 lte_55_1 ( .A({\temp220[15] , 
        \temp220[14] , \temp220[13] , \temp220[12] , \temp220[11] , 
        \temp220[10] , \temp220[9] , \temp220[8] , \temp220[7] , \temp220[6] , 
        \temp220[5] , \temp220[4] , \temp220[3] , \temp220[2] , \temp220[1] , 
        \temp220[0] }), .B(InEdges[31:16]), .LEQ(n812), .TC(n812), .GE_GT(n100
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_4 lte_55_5 ( .A({\temp584[15] , 
        \temp584[14] , \temp584[13] , \temp584[12] , \temp584[11] , 
        \temp584[10] , \temp584[9] , \temp584[8] , \temp584[7] , \temp584[6] , 
        \temp584[5] , \temp584[4] , \temp584[3] , \temp584[2] , \temp584[1] , 
        \temp584[0] }), .B(InEdges[95:80]), .LEQ(n811), .TC(n811), .GE_GT(n132
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_3 lte_55_4 ( .A({\temp494[15] , 
        \temp494[14] , \temp494[13] , \temp494[12] , \temp494[11] , 
        \temp494[10] , \temp494[9] , \temp494[8] , \temp494[7] , \temp494[6] , 
        \temp494[5] , \temp494[4] , \temp494[3] , \temp494[2] , \temp494[1] , 
        \temp494[0] }), .B(InEdges[79:64]), .LEQ(n810), .TC(n810), .GE_GT(n124
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_2 lte_55_3 ( .A({\temp404[15] , 
        \temp404[14] , \temp404[13] , \temp404[12] , \temp404[11] , 
        \temp404[10] , \temp404[9] , \temp404[8] , \temp404[7] , \temp404[6] , 
        \temp404[5] , \temp404[4] , \temp404[3] , \temp404[2] , \temp404[1] , 
        \temp404[0] }), .B(InEdges[63:48]), .LEQ(n809), .TC(n809), .GE_GT(n116
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp314[15] , 
        \temp314[14] , \temp314[13] , \temp314[12] , \temp314[11] , 
        \temp314[10] , \temp314[9] , \temp314[8] , \temp314[7] , \temp314[6] , 
        \temp314[5] , \temp314[4] , \temp314[3] , \temp314[2] , \temp314[1] , 
        \temp314[0] }), .B(InEdges[47:32]), .LEQ(n808), .TC(n808), .GE_GT(n108
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n807), .TC(n807), .GE_GT(n92) );
endmodule


module library ( InEdges, OutEdge, PathAddr, PathData, WeightAddr, WeightData, 
    Nid, Eid, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
input  [5:0] WeightAddr;
input  [5:0] Eid;
output [2:0] PathData;
input  [15:0] WeightData;
input  [3:0] Nid;
input  Start, Clk;
    EdgeAux edgeAux ( .Eid(Eid), .InEdge(InEdges[15:0]), .OutEdge(OutEdge), 
        .WeightAddr(WeightAddr), .WeightData(WeightData), .Clk(Clk) );
    NodeAux_INDEGREE1_SOURCE1 n_1_1 ( .Nid(Nid), .InEdges(InEdges[15:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE1_SOURCE0 n_1_0 ( .Nid(Nid), .InEdges(InEdges[15:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE4_SOURCE0 n_4_0 ( .Nid(Nid), .InEdges(InEdges[63:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE5_SOURCE0 n_5_0 ( .Nid(Nid), .InEdges(InEdges[79:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE2_SOURCE0 n_2_0 ( .Nid(Nid), .InEdges(InEdges[31:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE6_SOURCE0 n_6_0 ( .Nid(Nid), .InEdges(InEdges), .OutEdge(
        OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(Start), 
        .Clk(Clk) );
    NodeAux_INDEGREE3_SOURCE0 n_3_0 ( .Nid(Nid), .InEdges(InEdges[47:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
endmodule



module Node_NID0_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE1 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID0 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID1_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID3 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID2_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID4 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID5 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID6 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID7 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID8 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID3_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID9 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID10 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID11 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID12 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID4_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID13 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID14 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID15 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID16 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID17 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID18 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID5_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID19 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID20 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID6_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID21 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID22 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID23 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID24 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID7_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID25 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID26 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID27 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID28 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID29 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID8_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID30 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID31 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID9_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID32 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID33 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID34 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID35 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID36 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID10_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID37 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID38 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID39 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID40 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID41 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID42 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID11_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID43 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID44 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID45 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID46 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID47 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID12_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID48 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID49 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID50 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID51 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID13_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID52 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID14_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID53 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID54 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID55 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID56 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID57 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID58 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID15_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [3:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID59 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID60 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID61 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID62 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID63 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [5:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module graph ( WeightAddr, WeightData, PathAddr, PathData, Start, Clk );
input  [5:0] WeightAddr;
input  [15:0] WeightData;
input  [3:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire [15:0] In0;
    wire [15:0] Out0;
    wire [47:0] In1;
    wire [15:0] Out1;
    wire [79:0] In2;
    wire [15:0] Out2;
    wire [63:0] In3;
    wire [15:0] Out3;
    wire [95:0] In4;
    wire [15:0] Out4;
    wire [31:0] In5;
    wire [15:0] Out5;
    wire [63:0] In6;
    wire [15:0] Out6;
    wire [79:0] In7;
    wire [15:0] Out7;
    wire [31:0] In8;
    wire [15:0] Out8;
    wire [79:0] In9;
    wire [15:0] Out9;
    wire [95:0] In10;
    wire [15:0] Out10;
    wire [79:0] In11;
    wire [15:0] Out11;
    wire [63:0] In12;
    wire [15:0] Out12;
    wire [15:0] In13;
    wire [15:0] Out13;
    wire [95:0] In14;
    wire [15:0] Out14;
    wire [79:0] In15;
    wire [15:0] Out15;

    Node_NID0_INDEGREE1 n0 ( .InEdges(In0), .OutEdge(Out0),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID0 e0 ( .InEdge(Out15), .OutEdge(In0[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID1_INDEGREE3 n1 ( .InEdges(In1), .OutEdge(Out1),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1 e1 ( .InEdge(Out10), .OutEdge(In1[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2 e2 ( .InEdge(Out8), .OutEdge(In1[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID3 e3 ( .InEdge(Out3), .OutEdge(In1[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID2_INDEGREE5 n2 ( .InEdges(In2), .OutEdge(Out2),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID4 e4 ( .InEdge(Out10), .OutEdge(In2[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID5 e5 ( .InEdge(Out14), .OutEdge(In2[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID6 e6 ( .InEdge(Out9), .OutEdge(In2[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID7 e7 ( .InEdge(Out7), .OutEdge(In2[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID8 e8 ( .InEdge(Out6), .OutEdge(In2[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID3_INDEGREE4 n3 ( .InEdges(In3), .OutEdge(Out3),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID9 e9 ( .InEdge(Out6), .OutEdge(In3[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID10 e10 ( .InEdge(Out1), .OutEdge(In3[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID11 e11 ( .InEdge(Out10), .OutEdge(In3[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID12 e12 ( .InEdge(Out7), .OutEdge(In3[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID4_INDEGREE6 n4 ( .InEdges(In4), .OutEdge(Out4),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID13 e13 ( .InEdge(Out3), .OutEdge(In4[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID14 e14 ( .InEdge(Out5), .OutEdge(In4[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID15 e15 ( .InEdge(Out15), .OutEdge(In4[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID16 e16 ( .InEdge(Out2), .OutEdge(In4[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID17 e17 ( .InEdge(Out7), .OutEdge(In4[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID18 e18 ( .InEdge(Out1), .OutEdge(In4[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID5_INDEGREE2 n5 ( .InEdges(In5), .OutEdge(Out5),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID19 e19 ( .InEdge(Out10), .OutEdge(In5[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID20 e20 ( .InEdge(Out1), .OutEdge(In5[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID6_INDEGREE4 n6 ( .InEdges(In6), .OutEdge(Out6),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID21 e21 ( .InEdge(Out13), .OutEdge(In6[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID22 e22 ( .InEdge(Out4), .OutEdge(In6[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID23 e23 ( .InEdge(Out0), .OutEdge(In6[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID24 e24 ( .InEdge(Out14), .OutEdge(In6[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID7_INDEGREE5 n7 ( .InEdges(In7), .OutEdge(Out7),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID25 e25 ( .InEdge(Out10), .OutEdge(In7[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID26 e26 ( .InEdge(Out13), .OutEdge(In7[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID27 e27 ( .InEdge(Out9), .OutEdge(In7[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID28 e28 ( .InEdge(Out6), .OutEdge(In7[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID29 e29 ( .InEdge(Out3), .OutEdge(In7[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID8_INDEGREE2 n8 ( .InEdges(In8), .OutEdge(Out8),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID30 e30 ( .InEdge(Out0), .OutEdge(In8[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID31 e31 ( .InEdge(Out4), .OutEdge(In8[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID9_INDEGREE5 n9 ( .InEdges(In9), .OutEdge(Out9),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID32 e32 ( .InEdge(Out3), .OutEdge(In9[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID33 e33 ( .InEdge(Out5), .OutEdge(In9[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID34 e34 ( .InEdge(Out1), .OutEdge(In9[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID35 e35 ( .InEdge(Out10), .OutEdge(In9[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID36 e36 ( .InEdge(Out4), .OutEdge(In9[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID10_INDEGREE6 n10 ( .InEdges(In10), .OutEdge(Out10),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID37 e37 ( .InEdge(Out4), .OutEdge(In10[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID38 e38 ( .InEdge(Out3), .OutEdge(In10[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID39 e39 ( .InEdge(Out7), .OutEdge(In10[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID40 e40 ( .InEdge(Out1), .OutEdge(In10[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID41 e41 ( .InEdge(Out11), .OutEdge(In10[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID42 e42 ( .InEdge(Out8), .OutEdge(In10[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID11_INDEGREE5 n11 ( .InEdges(In11), .OutEdge(Out11),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID43 e43 ( .InEdge(Out1), .OutEdge(In11[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID44 e44 ( .InEdge(Out3), .OutEdge(In11[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID45 e45 ( .InEdge(Out14), .OutEdge(In11[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID46 e46 ( .InEdge(Out8), .OutEdge(In11[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID47 e47 ( .InEdge(Out10), .OutEdge(In11[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID12_INDEGREE4 n12 ( .InEdges(In12), .OutEdge(Out12),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID48 e48 ( .InEdge(Out2), .OutEdge(In12[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID49 e49 ( .InEdge(Out6), .OutEdge(In12[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID50 e50 ( .InEdge(Out4), .OutEdge(In12[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID51 e51 ( .InEdge(Out9), .OutEdge(In12[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID13_INDEGREE1 n13 ( .InEdges(In13), .OutEdge(Out13),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID52 e52 ( .InEdge(Out9), .OutEdge(In13[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID14_INDEGREE6 n14 ( .InEdges(In14), .OutEdge(Out14),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID53 e53 ( .InEdge(Out1), .OutEdge(In14[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID54 e54 ( .InEdge(Out15), .OutEdge(In14[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID55 e55 ( .InEdge(Out9), .OutEdge(In14[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID56 e56 ( .InEdge(Out2), .OutEdge(In14[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID57 e57 ( .InEdge(Out4), .OutEdge(In14[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID58 e58 ( .InEdge(Out6), .OutEdge(In14[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID15_INDEGREE5 n15 ( .InEdges(In15), .OutEdge(Out15),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID59 e59 ( .InEdge(Out9), .OutEdge(In15[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID60 e60 ( .InEdge(Out1), .OutEdge(In15[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID61 e61 ( .InEdge(Out5), .OutEdge(In15[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID62 e62 ( .InEdge(Out4), .OutEdge(In15[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID63 e63 ( .InEdge(Out8), .OutEdge(In15[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
endmodule
