
module CELL_DUMMY0_DW01_add_5_0 ( A, B, CI, SUM, CO );
input  [4:0] A;
input  [4:0] B;
output [4:0] SUM;
input  CI;
output CO;
    wire n1, \carry[2] , n2, n3, \carry[1] ;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(n2), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_PULLDOWN U2 ( .Z(n2) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(n1), .S(SUM[2]), .CO(SUM[3])
         );
    VMW_FADD U1_0 ( .CI(n3), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_PULLDOWN U3 ( .Z(n3) );
endmodule


module CELL_DUMMY0_DW01_add_6_0 ( A, B, CI, SUM, CO );
input  [5:0] A;
input  [5:0] B;
output [5:0] SUM;
input  CI;
output CO;
    wire n4, n6, n7, \carry[2] , n5, \carry[3] , \carry[1] ;
    VMW_PULLDOWN U1 ( .Z(n4) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(n6), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_PULLDOWN U2 ( .Z(n5) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(n5), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_0 ( .CI(n7), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_PULLDOWN U3 ( .Z(n6) );
    VMW_PULLDOWN U4 ( .Z(n7) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(n4), .S(SUM[3]), .CO(SUM[4])
         );
endmodule


module CELL_DUMMY0_DW01_add_7_0 ( A, B, CI, SUM, CO );
input  [6:0] A;
input  [6:0] B;
output [6:0] SUM;
input  CI;
output CO;
    wire n8, n9, \carry[4] , n12, \carry[2] , n10, n11, \carry[3] , \carry[1] ;
    VMW_PULLDOWN U1 ( .Z(n8) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(n11), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_PULLDOWN U2 ( .Z(n9) );
    VMW_PULLDOWN U5 ( .Z(n12) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(n10), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_0 ( .CI(n12), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_PULLDOWN U3 ( .Z(n10) );
    VMW_PULLDOWN U4 ( .Z(n11) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(n8), .S(SUM[4]), .CO(SUM[5])
         );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(n9), .S(SUM[3]), .CO(
        \carry[4] ) );
endmodule


module CELL_DUMMY0_DW01_add_8_0 ( A, B, CI, SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n13, n15, \carry[4] , \carry[2] , n14, n16, n17, n18, \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n13) );
    VMW_PULLDOWN U6 ( .Z(n18) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(n17), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_PULLDOWN U2 ( .Z(n14) );
    VMW_PULLDOWN U5 ( .Z(n17) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(n16), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_0 ( .CI(n18), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_PULLDOWN U3 ( .Z(n15) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(n13), .S(SUM[5]), .CO(SUM[6]
        ) );
    VMW_PULLDOWN U4 ( .Z(n16) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(n14), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(n15), .S(SUM[3]), .CO(
        \carry[4] ) );
endmodule


module CELL_DUMMY0 ( DATA_IN, cell_value, Reset, WR, Enable, Clk, NEIGHBORS );
input  [7:0] NEIGHBORS;
input  DATA_IN, Reset, WR, Enable, Clk;
output cell_value;
    wire n759, n776, \count75[6] , n758, n764, \count358[3] , \count353[1] , 
        \count75[4] , \count75[0] , \count75[2] , n771, n757, \count358[1] , 
        n763, n762, n770, \count363[2] , \count368[4] , \count368[0] , 
        \count368[2] , n773, n775, \count363[5] , \count368[6] , n765, 
        \count363[0] , n767, \count363[4] , \count368[3] , n375, \count75[5] , 
        n769, n772, \count363[3] , \count363[1] , \count368[1] , n760, 
        \count368[5] , \count353[2] , n768, \count358[0] , n774, \count358[4] , 
        n761, \count75[1] , \count75[3] , n766, \count358[2] , \count353[0] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 ;
    VMW_PULLDOWN U123 ( .Z(n759) );
    VMW_PULLDOWN U125 ( .Z(n774) );
    VMW_PULLDOWN U126 ( .Z(n775) );
    VMW_AND2 U134 ( .A(NEIGHBORS[3]), .B(n758), .Z(n760) );
    VMW_XOR2 U141 ( .A(NEIGHBORS[3]), .B(n758), .Z(\count353[0] ) );
    VMW_INV U148 ( .A(\count75[1] ), .Z(n766) );
    VMW_PULLDOWN U127 ( .Z(n776) );
    VMW_PULLDOWN U128 ( .Z(n375) );
    CELL_DUMMY0_DW01_add_7_0 add_62_6 ( .A({n375, \count363[5] , \count363[4] , 
        \count363[3] , \count363[2] , \count363[1] , \count363[0] }), .B({n774, 
        n774, n774, n774, n774, n774, NEIGHBORS[6]}), .CI(n774), .SUM({
        UNCONNECTED_1, \count368[5] , \count368[4] , \count368[3] , 
        \count368[2] , \count368[1] , \count368[0] }) );
    VMW_PULLDOWN U129 ( .Z(\count358[4] ) );
    VMW_OR3 U132 ( .A(\count75[5] ), .B(\count75[4] ), .C(\count75[6] ), .Z(
        n767) );
    VMW_AND3 U133 ( .A(n757), .B(n758), .C(NEIGHBORS[3]), .Z(\count353[2] ) );
    VMW_MUX2I U146 ( .A(n768), .B(cell_value), .S(n761), .Z(n764) );
    CELL_DUMMY0_DW01_add_8_0 add_62_7 ( .A({n375, \count368[6] , \count368[5] , 
        \count368[4] , \count368[3] , \count368[2] , \count368[1] , 
        \count368[0] }), .B({n773, n773, n773, n773, n773, n773, n773, 
        NEIGHBORS[7]}), .CI(n773), .SUM({UNCONNECTED_2, \count75[6] , 
        \count75[5] , \count75[4] , \count75[3] , \count75[2] , \count75[1] , 
        \count75[0] }) );
    VMW_OR2 U147 ( .A(Reset), .B(n770), .Z(n771) );
    VMW_AND2 U135 ( .A(\count75[0] ), .B(n762), .Z(n761) );
    VMW_XOR2 U140 ( .A(n757), .B(n760), .Z(\count353[1] ) );
    VMW_XOR2 U137 ( .A(NEIGHBORS[1]), .B(NEIGHBORS[0]), .Z(n765) );
    VMW_INV U149 ( .A(cell_value), .Z(n769) );
    VMW_OR2 U142 ( .A(n762), .B(n769), .Z(n768) );
    VMW_FD cell_value_reg ( .D(n772), .CP(Clk), .Q(cell_value) );
    VMW_PULLDOWN U130 ( .Z(\count363[5] ) );
    VMW_NOR4 U139 ( .A(\count75[3] ), .B(\count75[2] ), .C(n766), .D(n767), 
        .Z(n762) );
    CELL_DUMMY0_DW01_add_6_0 add_62_5 ( .A({n375, \count358[4] , \count358[3] , 
        \count358[2] , \count358[1] , \count358[0] }), .B({n775, n775, n775, 
        n775, n775, NEIGHBORS[5]}), .CI(n775), .SUM({UNCONNECTED_3, 
        \count363[4] , \count363[3] , \count363[2] , \count363[1] , 
        \count363[0] }) );
    VMW_AO22 U145 ( .A(NEIGHBORS[1]), .B(NEIGHBORS[0]), .C(NEIGHBORS[2]), .D(
        n765), .Z(n757) );
    VMW_XOR2 U138 ( .A(NEIGHBORS[2]), .B(n765), .Z(n758) );
    VMW_PULLDOWN U124 ( .Z(n773) );
    VMW_PULLDOWN U131 ( .Z(\count368[6] ) );
    CELL_DUMMY0_DW01_add_5_0 add_62_4 ( .A({n375, n759, \count353[2] , 
        \count353[1] , \count353[0] }), .B({n776, n776, n776, n776, 
        NEIGHBORS[4]}), .CI(n776), .SUM({UNCONNECTED_4, \count358[3] , 
        \count358[2] , \count358[1] , \count358[0] }) );
    VMW_AOI211 U136 ( .A(n764), .B(Enable), .C(WR), .D(Reset), .Z(n763) );
    VMW_MUX2I U143 ( .A(n769), .B(DATA_IN), .S(WR), .Z(n770) );
    VMW_MUX2I U144 ( .A(n771), .B(n769), .S(n763), .Z(n772) );
endmodule


module Life_Block_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, 
    ScanIn, ScanOut, ScanEnable, Id, Enable, BLOCK_VALUE, NORTH_EDGE, 
    SOUTH_EDGE, EAST_EDGE, WEST_EDGE, NW_EDGE, SW_EDGE, NE_EDGE, SE_EDGE );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
output [31:0] BLOCK_VALUE;
input  [31:0] NORTH_EDGE;
input  [31:0] SOUTH_EDGE;
input  Clk, Reset, RD, WR, ScanEnable, Enable, EAST_EDGE, WEST_EDGE, NW_EDGE, 
    SW_EDGE, NE_EDGE, SE_EDGE;
    wire \BLOCK_VALUE[31] , \BLOCK_VALUE[5] , \BLOCK_VALUE[1] , 
        \BLOCK_VALUE[8] , \BLOCK_VALUE[7] , \BLOCK_VALUE[3] , 
        \BLOCK_VALUE[25] , \BLOCK_VALUE[16] , \BLOCK_VALUE[21] , 
        \BLOCK_VALUE[12] , \BLOCK_VALUE[28] , \BLOCK_VALUE[19] , 
        \BLOCK_VALUE[23] , \BLOCK_VALUE[10] , \BLOCK_VALUE[27] , 
        \BLOCK_VALUE[14] , \BLOCK_VALUE[26] , \BLOCK_VALUE[15] , 
        \BLOCK_VALUE[18] , \BLOCK_VALUE[22] , \BLOCK_VALUE[11] , 
        \BLOCK_VALUE[20] , \BLOCK_VALUE[13] , \BLOCK_VALUE[30] , 
        \BLOCK_VALUE[29] , \BLOCK_VALUE[24] , \BLOCK_VALUE[17] , 
        \BLOCK_VALUE[2] , \BLOCK_VALUE[6] , \BLOCK_VALUE[4] , \BLOCK_VALUE[0] , 
        \BLOCK_VALUE[9] ;
    assign ScanOut[31] = \BLOCK_VALUE[31] ;
    assign ScanOut[30] = \BLOCK_VALUE[30] ;
    assign ScanOut[29] = \BLOCK_VALUE[29] ;
    assign ScanOut[28] = \BLOCK_VALUE[28] ;
    assign ScanOut[27] = \BLOCK_VALUE[27] ;
    assign ScanOut[26] = \BLOCK_VALUE[26] ;
    assign ScanOut[25] = \BLOCK_VALUE[25] ;
    assign ScanOut[24] = \BLOCK_VALUE[24] ;
    assign ScanOut[23] = \BLOCK_VALUE[23] ;
    assign ScanOut[22] = \BLOCK_VALUE[22] ;
    assign ScanOut[21] = \BLOCK_VALUE[21] ;
    assign ScanOut[20] = \BLOCK_VALUE[20] ;
    assign ScanOut[19] = \BLOCK_VALUE[19] ;
    assign ScanOut[18] = \BLOCK_VALUE[18] ;
    assign ScanOut[17] = \BLOCK_VALUE[17] ;
    assign ScanOut[16] = \BLOCK_VALUE[16] ;
    assign ScanOut[15] = \BLOCK_VALUE[15] ;
    assign ScanOut[14] = \BLOCK_VALUE[14] ;
    assign ScanOut[13] = \BLOCK_VALUE[13] ;
    assign ScanOut[12] = \BLOCK_VALUE[12] ;
    assign ScanOut[11] = \BLOCK_VALUE[11] ;
    assign ScanOut[10] = \BLOCK_VALUE[10] ;
    assign ScanOut[9] = \BLOCK_VALUE[9] ;
    assign ScanOut[8] = \BLOCK_VALUE[8] ;
    assign ScanOut[7] = \BLOCK_VALUE[7] ;
    assign ScanOut[6] = \BLOCK_VALUE[6] ;
    assign ScanOut[5] = \BLOCK_VALUE[5] ;
    assign ScanOut[4] = \BLOCK_VALUE[4] ;
    assign ScanOut[3] = \BLOCK_VALUE[3] ;
    assign ScanOut[2] = \BLOCK_VALUE[2] ;
    assign ScanOut[1] = \BLOCK_VALUE[1] ;
    assign ScanOut[0] = \BLOCK_VALUE[0] ;
    assign BLOCK_VALUE[31] = \BLOCK_VALUE[31] ;
    assign BLOCK_VALUE[30] = \BLOCK_VALUE[30] ;
    assign BLOCK_VALUE[29] = \BLOCK_VALUE[29] ;
    assign BLOCK_VALUE[28] = \BLOCK_VALUE[28] ;
    assign BLOCK_VALUE[27] = \BLOCK_VALUE[27] ;
    assign BLOCK_VALUE[26] = \BLOCK_VALUE[26] ;
    assign BLOCK_VALUE[25] = \BLOCK_VALUE[25] ;
    assign BLOCK_VALUE[24] = \BLOCK_VALUE[24] ;
    assign BLOCK_VALUE[23] = \BLOCK_VALUE[23] ;
    assign BLOCK_VALUE[22] = \BLOCK_VALUE[22] ;
    assign BLOCK_VALUE[21] = \BLOCK_VALUE[21] ;
    assign BLOCK_VALUE[20] = \BLOCK_VALUE[20] ;
    assign BLOCK_VALUE[19] = \BLOCK_VALUE[19] ;
    assign BLOCK_VALUE[18] = \BLOCK_VALUE[18] ;
    assign BLOCK_VALUE[17] = \BLOCK_VALUE[17] ;
    assign BLOCK_VALUE[16] = \BLOCK_VALUE[16] ;
    assign BLOCK_VALUE[15] = \BLOCK_VALUE[15] ;
    assign BLOCK_VALUE[14] = \BLOCK_VALUE[14] ;
    assign BLOCK_VALUE[13] = \BLOCK_VALUE[13] ;
    assign BLOCK_VALUE[12] = \BLOCK_VALUE[12] ;
    assign BLOCK_VALUE[11] = \BLOCK_VALUE[11] ;
    assign BLOCK_VALUE[10] = \BLOCK_VALUE[10] ;
    assign BLOCK_VALUE[9] = \BLOCK_VALUE[9] ;
    assign BLOCK_VALUE[8] = \BLOCK_VALUE[8] ;
    assign BLOCK_VALUE[7] = \BLOCK_VALUE[7] ;
    assign BLOCK_VALUE[6] = \BLOCK_VALUE[6] ;
    assign BLOCK_VALUE[5] = \BLOCK_VALUE[5] ;
    assign BLOCK_VALUE[4] = \BLOCK_VALUE[4] ;
    assign BLOCK_VALUE[3] = \BLOCK_VALUE[3] ;
    assign BLOCK_VALUE[2] = \BLOCK_VALUE[2] ;
    assign BLOCK_VALUE[1] = \BLOCK_VALUE[1] ;
    assign BLOCK_VALUE[0] = \BLOCK_VALUE[0] ;
    CELL_DUMMY0 cell_4 ( .DATA_IN(ScanIn[4]), .cell_value(\BLOCK_VALUE[4] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[5], \BLOCK_VALUE[5] , SOUTH_EDGE[5], 
        SOUTH_EDGE[4], SOUTH_EDGE[3], \BLOCK_VALUE[3] , NORTH_EDGE[3], 
        NORTH_EDGE[4]}) );
    CELL_DUMMY0 cell_15 ( .DATA_IN(ScanIn[15]), .cell_value(\BLOCK_VALUE[15] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[16], \BLOCK_VALUE[16] , SOUTH_EDGE[16], 
        SOUTH_EDGE[15], SOUTH_EDGE[14], \BLOCK_VALUE[14] , NORTH_EDGE[14], 
        NORTH_EDGE[15]}) );
    CELL_DUMMY0 cell_29 ( .DATA_IN(ScanIn[29]), .cell_value(\BLOCK_VALUE[29] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[30], \BLOCK_VALUE[30] , SOUTH_EDGE[30], 
        SOUTH_EDGE[29], SOUTH_EDGE[28], \BLOCK_VALUE[28] , NORTH_EDGE[28], 
        NORTH_EDGE[29]}) );
    CELL_DUMMY0 cell_3 ( .DATA_IN(ScanIn[3]), .cell_value(\BLOCK_VALUE[3] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[4], \BLOCK_VALUE[4] , SOUTH_EDGE[4], 
        SOUTH_EDGE[3], SOUTH_EDGE[2], \BLOCK_VALUE[2] , NORTH_EDGE[2], 
        NORTH_EDGE[3]}) );
    CELL_DUMMY0 cell_20 ( .DATA_IN(ScanIn[20]), .cell_value(\BLOCK_VALUE[20] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[21], \BLOCK_VALUE[21] , SOUTH_EDGE[21], 
        SOUTH_EDGE[20], SOUTH_EDGE[19], \BLOCK_VALUE[19] , NORTH_EDGE[19], 
        NORTH_EDGE[20]}) );
    CELL_DUMMY0 cell_27 ( .DATA_IN(ScanIn[27]), .cell_value(\BLOCK_VALUE[27] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[28], \BLOCK_VALUE[28] , SOUTH_EDGE[28], 
        SOUTH_EDGE[27], SOUTH_EDGE[26], \BLOCK_VALUE[26] , NORTH_EDGE[26], 
        NORTH_EDGE[27]}) );
    CELL_DUMMY0 cell_12 ( .DATA_IN(ScanIn[12]), .cell_value(\BLOCK_VALUE[12] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[13], \BLOCK_VALUE[13] , SOUTH_EDGE[13], 
        SOUTH_EDGE[12], SOUTH_EDGE[11], \BLOCK_VALUE[11] , NORTH_EDGE[11], 
        NORTH_EDGE[12]}) );
    CELL_DUMMY0 cell_26 ( .DATA_IN(ScanIn[26]), .cell_value(\BLOCK_VALUE[26] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[27], \BLOCK_VALUE[27] , SOUTH_EDGE[27], 
        SOUTH_EDGE[26], SOUTH_EDGE[25], \BLOCK_VALUE[25] , NORTH_EDGE[25], 
        NORTH_EDGE[26]}) );
    CELL_DUMMY0 cell_2 ( .DATA_IN(ScanIn[2]), .cell_value(\BLOCK_VALUE[2] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[3], \BLOCK_VALUE[3] , SOUTH_EDGE[3], 
        SOUTH_EDGE[2], SOUTH_EDGE[1], \BLOCK_VALUE[1] , NORTH_EDGE[1], 
        NORTH_EDGE[2]}) );
    CELL_DUMMY0 cell_5 ( .DATA_IN(ScanIn[5]), .cell_value(\BLOCK_VALUE[5] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[6], \BLOCK_VALUE[6] , SOUTH_EDGE[6], 
        SOUTH_EDGE[5], SOUTH_EDGE[4], \BLOCK_VALUE[4] , NORTH_EDGE[4], 
        NORTH_EDGE[5]}) );
    CELL_DUMMY0 cell_13 ( .DATA_IN(ScanIn[13]), .cell_value(\BLOCK_VALUE[13] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[14], \BLOCK_VALUE[14] , SOUTH_EDGE[14], 
        SOUTH_EDGE[13], SOUTH_EDGE[12], \BLOCK_VALUE[12] , NORTH_EDGE[12], 
        NORTH_EDGE[13]}) );
    CELL_DUMMY0 cell_14 ( .DATA_IN(ScanIn[14]), .cell_value(\BLOCK_VALUE[14] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[15], \BLOCK_VALUE[15] , SOUTH_EDGE[15], 
        SOUTH_EDGE[14], SOUTH_EDGE[13], \BLOCK_VALUE[13] , NORTH_EDGE[13], 
        NORTH_EDGE[14]}) );
    CELL_DUMMY0 cell_21 ( .DATA_IN(ScanIn[21]), .cell_value(\BLOCK_VALUE[21] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[22], \BLOCK_VALUE[22] , SOUTH_EDGE[22], 
        SOUTH_EDGE[21], SOUTH_EDGE[20], \BLOCK_VALUE[20] , NORTH_EDGE[20], 
        NORTH_EDGE[21]}) );
    CELL_DUMMY0 cell_28 ( .DATA_IN(ScanIn[28]), .cell_value(\BLOCK_VALUE[28] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[29], \BLOCK_VALUE[29] , SOUTH_EDGE[29], 
        SOUTH_EDGE[28], SOUTH_EDGE[27], \BLOCK_VALUE[27] , NORTH_EDGE[27], 
        NORTH_EDGE[28]}) );
    CELL_DUMMY0 cell_0 ( .DATA_IN(ScanIn[0]), .cell_value(\BLOCK_VALUE[0] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[1], \BLOCK_VALUE[1] , SOUTH_EDGE[1], 
        SOUTH_EDGE[0], SE_EDGE, EAST_EDGE, NE_EDGE, NORTH_EDGE[0]}) );
    CELL_DUMMY0 cell_7 ( .DATA_IN(ScanIn[7]), .cell_value(\BLOCK_VALUE[7] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[8], \BLOCK_VALUE[8] , SOUTH_EDGE[8], 
        SOUTH_EDGE[7], SOUTH_EDGE[6], \BLOCK_VALUE[6] , NORTH_EDGE[6], 
        NORTH_EDGE[7]}) );
    CELL_DUMMY0 cell_16 ( .DATA_IN(ScanIn[16]), .cell_value(\BLOCK_VALUE[16] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[17], \BLOCK_VALUE[17] , SOUTH_EDGE[17], 
        SOUTH_EDGE[16], SOUTH_EDGE[15], \BLOCK_VALUE[15] , NORTH_EDGE[15], 
        NORTH_EDGE[16]}) );
    CELL_DUMMY0 cell_31 ( .DATA_IN(ScanIn[31]), .cell_value(\BLOCK_VALUE[31] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NW_EDGE, WEST_EDGE, SW_EDGE, SOUTH_EDGE[31], 
        SOUTH_EDGE[30], \BLOCK_VALUE[30] , NORTH_EDGE[30], NORTH_EDGE[31]}) );
    CELL_DUMMY0 cell_9 ( .DATA_IN(ScanIn[9]), .cell_value(\BLOCK_VALUE[9] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[10], \BLOCK_VALUE[10] , SOUTH_EDGE[10], 
        SOUTH_EDGE[9], SOUTH_EDGE[8], \BLOCK_VALUE[8] , NORTH_EDGE[8], 
        NORTH_EDGE[9]}) );
    CELL_DUMMY0 cell_18 ( .DATA_IN(ScanIn[18]), .cell_value(\BLOCK_VALUE[18] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[19], \BLOCK_VALUE[19] , SOUTH_EDGE[19], 
        SOUTH_EDGE[18], SOUTH_EDGE[17], \BLOCK_VALUE[17] , NORTH_EDGE[17], 
        NORTH_EDGE[18]}) );
    CELL_DUMMY0 cell_23 ( .DATA_IN(ScanIn[23]), .cell_value(\BLOCK_VALUE[23] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[24], \BLOCK_VALUE[24] , SOUTH_EDGE[24], 
        SOUTH_EDGE[23], SOUTH_EDGE[22], \BLOCK_VALUE[22] , NORTH_EDGE[22], 
        NORTH_EDGE[23]}) );
    CELL_DUMMY0 cell_24 ( .DATA_IN(ScanIn[24]), .cell_value(\BLOCK_VALUE[24] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[25], \BLOCK_VALUE[25] , SOUTH_EDGE[25], 
        SOUTH_EDGE[24], SOUTH_EDGE[23], \BLOCK_VALUE[23] , NORTH_EDGE[23], 
        NORTH_EDGE[24]}) );
    CELL_DUMMY0 cell_1 ( .DATA_IN(ScanIn[1]), .cell_value(\BLOCK_VALUE[1] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[2], \BLOCK_VALUE[2] , SOUTH_EDGE[2], 
        SOUTH_EDGE[1], SOUTH_EDGE[0], \BLOCK_VALUE[0] , NORTH_EDGE[0], 
        NORTH_EDGE[1]}) );
    CELL_DUMMY0 cell_8 ( .DATA_IN(ScanIn[8]), .cell_value(\BLOCK_VALUE[8] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[9], \BLOCK_VALUE[9] , SOUTH_EDGE[9], 
        SOUTH_EDGE[8], SOUTH_EDGE[7], \BLOCK_VALUE[7] , NORTH_EDGE[7], 
        NORTH_EDGE[8]}) );
    CELL_DUMMY0 cell_11 ( .DATA_IN(ScanIn[11]), .cell_value(\BLOCK_VALUE[11] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[12], \BLOCK_VALUE[12] , SOUTH_EDGE[12], 
        SOUTH_EDGE[11], SOUTH_EDGE[10], \BLOCK_VALUE[10] , NORTH_EDGE[10], 
        NORTH_EDGE[11]}) );
    CELL_DUMMY0 cell_19 ( .DATA_IN(ScanIn[19]), .cell_value(\BLOCK_VALUE[19] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[20], \BLOCK_VALUE[20] , SOUTH_EDGE[20], 
        SOUTH_EDGE[19], SOUTH_EDGE[18], \BLOCK_VALUE[18] , NORTH_EDGE[18], 
        NORTH_EDGE[19]}) );
    CELL_DUMMY0 cell_25 ( .DATA_IN(ScanIn[25]), .cell_value(\BLOCK_VALUE[25] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[26], \BLOCK_VALUE[26] , SOUTH_EDGE[26], 
        SOUTH_EDGE[25], SOUTH_EDGE[24], \BLOCK_VALUE[24] , NORTH_EDGE[24], 
        NORTH_EDGE[25]}) );
    CELL_DUMMY0 cell_6 ( .DATA_IN(ScanIn[6]), .cell_value(\BLOCK_VALUE[6] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[7], \BLOCK_VALUE[7] , SOUTH_EDGE[7], 
        SOUTH_EDGE[6], SOUTH_EDGE[5], \BLOCK_VALUE[5] , NORTH_EDGE[5], 
        NORTH_EDGE[6]}) );
    CELL_DUMMY0 cell_10 ( .DATA_IN(ScanIn[10]), .cell_value(\BLOCK_VALUE[10] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[11], \BLOCK_VALUE[11] , SOUTH_EDGE[11], 
        SOUTH_EDGE[10], SOUTH_EDGE[9], \BLOCK_VALUE[9] , NORTH_EDGE[9], 
        NORTH_EDGE[10]}) );
    CELL_DUMMY0 cell_17 ( .DATA_IN(ScanIn[17]), .cell_value(\BLOCK_VALUE[17] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[18], \BLOCK_VALUE[18] , SOUTH_EDGE[18], 
        SOUTH_EDGE[17], SOUTH_EDGE[16], \BLOCK_VALUE[16] , NORTH_EDGE[16], 
        NORTH_EDGE[17]}) );
    CELL_DUMMY0 cell_30 ( .DATA_IN(ScanIn[30]), .cell_value(\BLOCK_VALUE[30] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[31], \BLOCK_VALUE[31] , SOUTH_EDGE[31], 
        SOUTH_EDGE[30], SOUTH_EDGE[29], \BLOCK_VALUE[29] , NORTH_EDGE[29], 
        NORTH_EDGE[30]}) );
    CELL_DUMMY0 cell_22 ( .DATA_IN(ScanIn[22]), .cell_value(\BLOCK_VALUE[22] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[23], \BLOCK_VALUE[23] , SOUTH_EDGE[23], 
        SOUTH_EDGE[22], SOUTH_EDGE[21], \BLOCK_VALUE[21] , NORTH_EDGE[21], 
        NORTH_EDGE[22]}) );
endmodule


module Life_Control_WIDTH32_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 ( A, SUM );
input  [6:0] A;
output [6:0] SUM;
    wire n5, n9, n7, n12, n6, n13, n8, n10, n11;
    VMW_AO21 U3 ( .A(n5), .B(A[2]), .C(n6), .Z(SUM[2]) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(n9), .Z(SUM[1]) );
    VMW_INV U6 ( .A(A[0]), .Z(SUM[0]) );
    VMW_AO22 U14 ( .A(A[5]), .B(n13), .C(n12), .D(n10), .Z(SUM[5]) );
    VMW_AO21 U7 ( .A(n8), .B(A[4]), .C(n10), .Z(SUM[4]) );
    VMW_AND2 U8 ( .A(n10), .B(n12), .Z(n11) );
    VMW_XOR2 U13 ( .A(A[6]), .B(n11), .Z(SUM[6]) );
    VMW_OR2 U9 ( .A(A[0]), .B(A[1]), .Z(n5) );
    VMW_NOR2 U12 ( .A(n8), .B(A[4]), .Z(n10) );
    VMW_INV U15 ( .A(A[5]), .Z(n12) );
    VMW_INV U17 ( .A(A[3]), .Z(n7) );
    VMW_NOR2 U10 ( .A(n5), .B(A[2]), .Z(n6) );
    VMW_NAND2 U11 ( .A(n6), .B(n7), .Z(n8) );
    VMW_OAI21 U4 ( .A(n6), .B(n7), .C(n8), .Z(SUM[3]) );
    VMW_INV U18 ( .A(n5), .Z(n9) );
    VMW_INV U16 ( .A(n10), .Z(n13) );
endmodule


module Life_Control_WIDTH32_CWIDTH7_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, ScanId, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire n330, n317, \count[2] , n362, n345, \count[6] , n339, n357, n322, 
        n325, n350, n319, \count[4] , n342, \count[0] , n359, n356, n337, n318, 
        n351, \ScanReg[15] , \ScanReg[26] , \ScanReg[2] , \count260[3] , n324, 
        \ScanReg[18] , n336, n358, n343, \ScanReg[22] , \ScanReg[11] , 
        \ScanReg[6] , \count260[5] , \ScanReg[20] , \ScanReg[13] , 
        \ScanReg[4] , n344, \count260[1] , n316, \ScanReg[29] , \ScanReg[30] , 
        n331, n323, \ScanReg[17] , \ScanReg[24] , \ScanReg[0] , \ScanReg[9] , 
        n338, n314, \count260[0] , n333, \ScanReg[16] , \ScanReg[25] , n361, 
        n346, \ScanReg[1] , \ScanReg[8] , \ScanReg[7] , n328, \ScanReg[5] , 
        \count260[4] , \ScanReg[21] , \ScanReg[12] , n354, \ScanReg[28] , 
        \ScanReg[31] , n321, n326, \ScanReg[19] , n348, \count260[6] , n353, 
        \ScanReg[10] , \ScanReg[23] , n341, \ScanReg[14] , \ScanReg[27] , n313, 
        \ScanReg[3] , \count260[2] , n334, \count[1] , n352, n349, n327, n335, 
        n360, n340, \count[5] , n347, n329, n332, n315, n320, \count[3] , n355;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U54 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U73 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_NOR2 U113 ( .A(n318), .B(n316), .Z(n314) );
    VMW_INV U134 ( .A(n321), .Z(ScanEnable) );
    VMW_AND2 U68 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_AND2 U96 ( .A(\ScanReg[13] ), .B(n316), .Z(n340) );
    VMW_AO21 U108 ( .A(RD), .B(ScanEnable), .C(n317), .Z(n328) );
    VMW_BUFIZ U141 ( .A(n330), .E(n328), .Z(\arr[27] ) );
    VMW_BUFIZ U166 ( .A(n355), .E(n328), .Z(\arr[8] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \count_reg[6]  ( .D(n356), .CP(Clk), .Q(\count[6] ) );
    VMW_AND2 U53 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U61 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_AND2 U84 ( .A(\ScanReg[8] ), .B(n316), .Z(n355) );
    VMW_BUFIZ U148 ( .A(n337), .E(n328), .Z(\arr[21] ) );
    VMW_BUFIZ U153 ( .A(n342), .E(n328), .Z(\arr[29] ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    Life_Control_WIDTH32_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 sub_281 ( .A({
        \count[6] , \count[5] , \count[4] , \count[3] , \count[2] , \count[1] , 
        \count[0] }), .SUM({\count260[6] , \count260[5] , \count260[4] , 
        \count260[3] , \count260[2] , \count260[1] , \count260[0] }) );
    VMW_FD \count_reg[2]  ( .D(n360), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U66 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AND2 U101 ( .A(\ScanReg[16] ), .B(n316), .Z(n333) );
    VMW_AND2 U106 ( .A(\ScanReg[10] ), .B(n316), .Z(n326) );
    VMW_OAI21 U121 ( .A(RD), .B(WR), .C(n322), .Z(n321) );
    VMW_AO22 U126 ( .A(\count[2] ), .B(n317), .C(\ScanReg[2] ), .D(n316), .Z(
        n339) );
    VMW_AO22 U83 ( .A(ScanOut[6]), .B(n314), .C(\count260[6] ), .D(n315), .Z(
        n356) );
    VMW_FD \count_reg[0]  ( .D(n362), .CP(Clk), .Q(\count[0] ) );
    VMW_AND2 U91 ( .A(\ScanReg[17] ), .B(n316), .Z(n346) );
    VMW_AND2 U98 ( .A(\ScanReg[21] ), .B(n316), .Z(n337) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(\count[0] ), .B(n317), .C(\ScanReg[0] ), .D(n316), .Z(
        n324) );
    VMW_BUFIZ U154 ( .A(n343), .E(n328), .Z(\arr[20] ) );
    VMW_FD \count_reg[4]  ( .D(n358), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U146 ( .A(n335), .E(n328), .Z(\arr[6] ) );
    VMW_BUFIZ U161 ( .A(n350), .E(n328), .Z(\arr[15] ) );
    VMW_AND2 U74 ( .A(DataIn[9]), .B(WR), .Z(ScanOut[9]) );
    VMW_AND2 U114 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_INV U133 ( .A(Reset), .Z(n320) );
    VMW_AND2 U99 ( .A(\ScanReg[31] ), .B(n316), .Z(n336) );
    VMW_BUFIZ U155 ( .A(n344), .E(n328), .Z(\arr[3] ) );
    VMW_AND2 U52 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U67 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_AO22 U82 ( .A(ScanOut[5]), .B(n314), .C(\count260[5] ), .D(n315), .Z(
        n357) );
    VMW_AND2 U107 ( .A(\ScanReg[23] ), .B(n316), .Z(n325) );
    VMW_AND2 U120 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U55 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U69 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U75 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U115 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_XNOR2 U132 ( .A(Addr[0]), .B(ScanId), .Z(n322) );
    VMW_AND2 U90 ( .A(\ScanReg[7] ), .B(n316), .Z(n347) );
    VMW_AND2 U109 ( .A(\ScanReg[19] ), .B(n316), .Z(n323) );
    VMW_OR4 U129 ( .A(\count[3] ), .B(\count[4] ), .C(\count[5] ), .D(
        \count[6] ), .Z(n313) );
    VMW_BUFIZ U147 ( .A(n336), .E(n328), .Z(\arr[31] ) );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_BUFIZ U160 ( .A(n349), .E(n328), .Z(\arr[26] ) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_AND2 U72 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_AND2 U97 ( .A(\ScanReg[28] ), .B(n316), .Z(n338) );
    VMW_BUFIZ U140 ( .A(n329), .E(n328), .Z(\arr[4] ) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_NOR2 U112 ( .A(n318), .B(n319), .Z(n315) );
    VMW_BUFIZ U135 ( .A(n323), .E(n328), .Z(\arr[19] ) );
    VMW_AND2 U60 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U85 ( .A(\ScanReg[11] ), .B(n316), .Z(n353) );
    VMW_AND2 U100 ( .A(\ScanReg[12] ), .B(n316), .Z(n334) );
    VMW_AO22 U127 ( .A(\count[1] ), .B(n317), .C(\ScanReg[1] ), .D(n316), .Z(
        n354) );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_BUFIZ U149 ( .A(n338), .E(n328), .Z(\arr[28] ) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_BUFIZ U152 ( .A(n341), .E(n328), .Z(\arr[30] ) );
    VMW_OR4 U51 ( .A(\count[1] ), .B(\count[2] ), .C(\count[0] ), .D(n313), 
        .Z(Enable) );
    VMW_AND2 U57 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_BUFIZ U137 ( .A(n325), .E(n328), .Z(\arr[23] ) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_AND2 U58 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U59 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_AND2 U62 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_AND2 U70 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AO22 U79 ( .A(ScanOut[2]), .B(n314), .C(\count260[2] ), .D(n315), .Z(
        n360) );
    VMW_AND2 U95 ( .A(\ScanReg[30] ), .B(n316), .Z(n341) );
    VMW_XOR2 U110 ( .A(Addr[0]), .B(Id), .Z(n316) );
    VMW_BUFIZ U159 ( .A(n348), .E(n328), .Z(\arr[5] ) );
    VMW_AND2 U119 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_BUFIZ U142 ( .A(n331), .E(n328), .Z(\arr[14] ) );
    VMW_BUFIZ U165 ( .A(n354), .E(n328), .Z(\arr[1] ) );
    VMW_AND2 U87 ( .A(\ScanReg[18] ), .B(n316), .Z(n351) );
    VMW_BUFIZ U150 ( .A(n339), .E(n328), .Z(\arr[2] ) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(\count[3] ), .B(n317), .C(\ScanReg[3] ), .D(n316), .Z(
        n344) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U65 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AND2 U102 ( .A(\ScanReg[25] ), .B(n316), .Z(n332) );
    VMW_AND2 U105 ( .A(\ScanReg[9] ), .B(n316), .Z(n327) );
    VMW_AO22 U80 ( .A(ScanOut[3]), .B(n314), .C(\count260[3] ), .D(n315), .Z(
        n359) );
    VMW_AO22 U122 ( .A(\count[6] ), .B(n317), .C(\ScanReg[6] ), .D(n316), .Z(
        n335) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_BUFIZ U139 ( .A(n327), .E(n328), .Z(\arr[9] ) );
    VMW_BUFIZ U157 ( .A(n346), .E(n328), .Z(\arr[17] ) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO22 U77 ( .A(ScanOut[0]), .B(n314), .C(\count260[0] ), .D(n315), .Z(
        n362) );
    VMW_AND2 U89 ( .A(\ScanReg[26] ), .B(n316), .Z(n349) );
    VMW_AND2 U92 ( .A(\ScanReg[24] ), .B(n316), .Z(n345) );
    VMW_BUFIZ U145 ( .A(n334), .E(n328), .Z(\arr[12] ) );
    VMW_BUFIZ U162 ( .A(n351), .E(n328), .Z(\arr[18] ) );
    VMW_AND2 U117 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AND2 U130 ( .A(n317), .B(WR), .Z(n319) );
    VMW_BUFIZ U138 ( .A(n326), .E(n328), .Z(\arr[10] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n357), .CP(Clk), .Q(\count[5] ) );
    VMW_AND2 U64 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AO22 U81 ( .A(ScanOut[4]), .B(n314), .C(\count260[4] ), .D(n315), .Z(
        n358) );
    VMW_BUFIZ U156 ( .A(n345), .E(n328), .Z(\arr[24] ) );
    VMW_AND2 U104 ( .A(\ScanReg[27] ), .B(n316), .Z(n330) );
    VMW_AND2 U76 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_AND2 U116 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AO22 U123 ( .A(\count[5] ), .B(n317), .C(\ScanReg[5] ), .D(n316), .Z(
        n348) );
    VMW_AND2 U56 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U88 ( .A(\ScanReg[15] ), .B(n316), .Z(n350) );
    VMW_AND2 U93 ( .A(\ScanReg[20] ), .B(n316), .Z(n343) );
    VMW_INV U131 ( .A(n316), .Z(n317) );
    VMW_FD \count_reg[1]  ( .D(n361), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(\ScanReg[29] ), .B(n316), .Z(n342) );
    VMW_BUFIZ U143 ( .A(n332), .E(n328), .Z(\arr[25] ) );
    VMW_BUFIZ U144 ( .A(n333), .E(n328), .Z(\arr[16] ) );
    VMW_BUFIZ U163 ( .A(n352), .E(n328), .Z(\arr[22] ) );
    VMW_BUFIZ U158 ( .A(n347), .E(n328), .Z(\arr[7] ) );
    VMW_BUFIZ U164 ( .A(n353), .E(n328), .Z(\arr[11] ) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_FD \count_reg[3]  ( .D(n359), .CP(Clk), .Q(\count[3] ) );
    VMW_BUFIZ U136 ( .A(n324), .E(n328), .Z(\arr[0] ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AND2 U63 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U71 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_OAI21 U111 ( .A(n319), .B(Enable), .C(n320), .Z(n318) );
    VMW_AO22 U124 ( .A(\count[4] ), .B(n317), .C(\ScanReg[4] ), .D(n316), .Z(
        n329) );
    VMW_AO22 U78 ( .A(ScanOut[1]), .B(n314), .C(\count260[1] ), .D(n315), .Z(
        n361) );
    VMW_AND2 U86 ( .A(\ScanReg[22] ), .B(n316), .Z(n352) );
    VMW_AND2 U103 ( .A(\ScanReg[14] ), .B(n316), .Z(n331) );
    VMW_AND2 U118 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_BUFIZ U151 ( .A(n340), .E(n328), .Z(\arr[13] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \nOut1_20[5] , \nScanOut2[20] , \nOut0_18[15] , \nOut1_20[20] , 
        \nOut1_55[10] , \nScanOut103[25] , \nScanOut91[17] , \nScanOut120[14] , 
        \nOut1_63[15] , \nScanOut2[13] , \nOut1_16[25] , \nScanOut84[23] , 
        \nOut1_16[16] , \nOut1_23[6] , \nScanOut29[23] , \nOut1_35[14] , 
        \nOut1_40[24] , \nScanOut116[11] , \nScanOut49[27] , \nScanOut84[10] , 
        \nScanOut108[0] , \nOut0_18[26] , \nOut1_63[26] , \nOut1_20[13] , 
        \nOut1_35[27] , \nOut1_40[17] , \nScanOut116[22] , \nOut1_44[1] , 
        \nOut1_55[23] , \nScanOut91[24] , \nScanOut103[16] , \nScanOut120[27] , 
        \nOut0_1[1] , \nOut0_2[2] , \nOut0_3[22] , \nScanOut11[1] , 
        \nScanOut29[10] , \nOut1_47[2] , \nScanOut70[8] , \nScanOut49[14] , 
        \nScanOut110[2] , \nOut0_3[11] , \nOut1_9[6] , \nScanOut12[2] , 
        \nOut0_19[1] , \nOut1_38[7] , \nOut1_25[8] , \nScanOut113[1] , 
        \nScanOut14[19] , \nScanOut37[31] , \nScanOut37[28] , \nScanOut61[29] , 
        \nScanOut42[18] , \nScanOut61[30] , \nScanOut4[1] , \nScanOut7[2] , 
        \nOut1_8[23] , \nOut0_13[19] , \nOut0_63[9] , \nScanOut108[29] , 
        \nScanOut75[5] , \nScanOut108[30] , \nOut0_30[31] , \nOut0_30[28] , 
        \nOut0_45[18] , \nScanOut76[6] , \nScanOut52[0] , \nOut0_59[3] , 
        \nScanOut80[6] , \nScanOut6[22] , \nOut0_7[20] , \nOut0_7[13] , 
        \nOut1_8[10] , \nOut0_17[31] , \nOut0_17[28] , \nOut1_19[18] , 
        \nOut0_41[30] , \nOut0_62[18] , \nScanOut83[5] , \nOut0_34[19] , 
        \nOut0_41[29] , \nScanOut51[3] , \nScanOut65[18] , \nScanOut10[31] , 
        \nScanOut10[28] , \nScanOut46[30] , \nOut0_20[8] , \nScanOut33[19] , 
        \nScanOut36[4] , \nScanOut46[29] , \nScanOut28[8] , \nScanOut35[7] , 
        \nScanOut38[15] , \nOut0_42[2] , \nOut1_63[4] , \nScanOut58[11] , 
        \nScanOut86[8] , \nScanOut49[1] , \nOut1_12[27] , \nScanOut80[21] , 
        \nOut1_24[22] , \nOut1_31[16] , \nOut1_44[26] , \nScanOut112[13] , 
        \nOut1_51[12] , \nScanOut107[27] , \nScanOut38[26] , \nOut0_41[1] , 
        \nOut1_60[7] , \nScanOut95[15] , \nScanOut124[16] , \nScanOut98[4] , 
        \nScanOut58[22] , \nOut1_12[14] , \nOut1_24[11] , \nOut0_25[5] , 
        \nOut0_26[6] , \nScanOut33[9] , \nOut1_51[21] , \nScanOut80[12] , 
        \nScanOut95[26] , \nScanOut107[14] , \nScanOut124[25] , \nOut1_2[25] , 
        \nOut0_6[19] , \nScanOut6[11] , \nOut1_31[25] , \nOut1_44[15] , 
        \nScanOut112[20] , \nOut0_9[9] , \nOut1_11[4] , \nOut1_12[7] , 
        \nOut0_16[11] , \nOut0_35[20] , \nScanOut38[2] , \nOut0_40[10] , 
        \nScanOut118[15] , \nOut1_18[21] , \nOut0_63[21] , \nOut0_20[14] , 
        \nOut0_33[1] , \nScanOut27[27] , \nScanOut52[17] , \nOut0_55[24] , 
        \nScanOut71[26] , \nOut0_30[2] , \nScanOut32[13] , \nScanOut47[23] , 
        \nOut1_9[30] , \nScanOut9[4] , \nScanOut11[22] , \nScanOut64[12] , 
        \nOut0_16[22] , \nOut1_18[12] , \nOut0_20[27] , \nOut0_55[17] , 
        \nOut0_35[13] , \nOut0_40[23] , \nScanOut41[9] , \nOut0_57[5] , 
        \nOut0_63[12] , \nScanOut118[26] , \nScanOut32[20] , \nOut0_49[9] , 
        \nOut1_9[29] , \nScanOut11[11] , \nScanOut47[10] , \nOut1_14[9] , 
        \nScanOut27[14] , \nScanOut64[21] , \nScanOut71[15] , \nOut0_28[0] , 
        \nScanOut52[24] , \nOut0_54[6] , \nScanOut122[0] , \nScanOut81[18] , 
        \nScanOut20[0] , \nScanOut23[3] , \nScanOut121[3] , \nOut1_2[16] , 
        \nScanOut7[31] , \nScanOut47[7] , \nScanOut59[31] , \nScanOut59[28] , 
        \nScanOut113[19] , \nScanOut7[28] , \nOut1_25[31] , \nOut1_25[28] , 
        \nOut1_50[18] , \nScanOut95[1] , \nScanOut96[2] , \nScanOut3[19] , 
        \nOut1_6[27] , \nScanOut44[4] , \nOut0_52[8] , \nOut0_9[24] , 
        \nOut1_57[8] , \nScanOut60[2] , \nScanOut63[1] , \nOut1_49[4] , 
        \nScanOut117[31] , \nScanOut117[28] , \nOut1_4[3] , \nOut1_6[14] , 
        \nScanOut19[9] , \nOut1_21[19] , \nOut1_54[30] , \nOut1_54[29] , 
        \nScanOut8[26] , \nOut0_9[17] , \nScanOut28[30] , \nScanOut28[29] , 
        \nScanOut105[5] , \nScanOut85[30] , \nScanOut106[6] , \nScanOut85[29] , 
        \nOut0_11[9] , \nOut0_12[13] , \nScanOut15[20] , \nScanOut36[11] , 
        \nScanOut43[21] , \nOut1_51[6] , \nScanOut60[10] , \nScanOut23[25] , 
        \nScanOut56[15] , \nScanOut75[24] , \nOut0_24[16] , \nOut1_52[5] , 
        \nOut0_31[22] , \nOut0_51[26] , \nScanOut109[23] , \nOut0_44[12] , 
        \nOut0_14[4] , \nScanOut23[16] , \nScanOut75[17] , \nScanOut78[0] , 
        \nOut1_35[2] , \nScanOut15[13] , \nScanOut36[22] , \nScanOut56[26] , 
        \nScanOut43[12] , \nScanOut60[23] , \nOut0_1[8] , \nOut1_1[7] , 
        \nOut0_2[31] , \nOut0_2[28] , \nOut1_7[0] , \nScanOut100[8] , 
        \nOut0_2[21] , \nOut0_6[23] , \nScanOut7[21] , \nScanOut8[15] , 
        \nOut0_12[20] , \nOut0_17[7] , \nOut1_36[1] , \nOut0_44[21] , 
        \nOut0_31[11] , \nOut0_24[25] , \nOut0_51[15] , \nOut1_25[21] , 
        \nOut1_50[11] , \nOut0_51[2] , \nScanOut109[10] , \nScanOut88[7] , 
        \nScanOut94[16] , \nScanOut125[15] , \nScanOut106[24] , \nOut1_30[15] , 
        \nOut1_45[25] , \nScanOut95[8] , \nScanOut113[10] , \nScanOut7[12] , 
        \nOut1_13[24] , \nScanOut81[22] , \nOut1_13[17] , \nOut0_28[9] , 
        \nScanOut39[16] , \nOut0_52[1] , \nScanOut59[12] , \nScanOut59[2] , 
        \nOut1_30[26] , \nOut1_45[16] , \nScanOut113[23] , \nScanOut81[11] , 
        \nOut1_14[0] , \nOut1_25[12] , \nScanOut94[25] , \nScanOut125[26] , 
        \nOut0_35[6] , \nOut1_50[22] , \nScanOut122[9] , \nScanOut106[17] , 
        \nOut1_17[3] , \nOut0_36[5] , \nScanOut20[9] , \nScanOut39[25] , 
        \nScanOut59[21] , \nScanOut41[0] , \nScanOut93[6] , \nOut0_6[10] , 
        \nOut1_9[20] , \nScanOut11[18] , \nScanOut32[29] , \nScanOut42[3] , 
        \nOut0_49[0] , \nScanOut90[5] , \nScanOut47[19] , \nScanOut64[31] , 
        \nScanOut32[30] , \nScanOut64[28] , \nOut0_9[0] , \nOut0_16[18] , 
        \nOut1_18[31] , \nScanOut25[4] , \nOut0_33[8] , \nScanOut124[7] , 
        \nOut0_35[29] , \nOut0_40[19] , \nOut0_63[31] , \nOut1_18[28] , 
        \nOut0_35[30] , \nOut0_63[28] , \nScanOut26[7] , \nOut1_9[13] , 
        \nOut1_28[4] , \nScanOut103[2] , \nScanOut127[4] , \nOut0_2[12] , 
        \nOut1_7[9] , \nScanOut100[1] , \nOut0_12[30] , \nOut0_31[18] , 
        \nOut1_36[8] , \nScanOut109[19] , \nOut0_44[28] , \nOut0_12[29] , 
        \nOut0_44[31] , \nScanOut15[30] , \nScanOut36[18] , \nScanOut43[28] , 
        \nScanOut66[5] , \nScanOut15[29] , \nScanOut43[31] , \nScanOut60[19] , 
        \nScanOut65[6] , \nOut1_2[4] , \nOut0_12[3] , \nOut1_33[5] , 
        \nScanOut78[9] , \nScanOut118[3] , \nScanOut19[0] , \nScanOut28[20] , 
        \nScanOut48[24] , \nScanOut3[23] , \nOut0_19[16] , \nOut1_34[17] , 
        \nOut1_41[27] , \nScanOut117[12] , \nOut1_62[16] , \nOut1_17[26] , 
        \nScanOut85[20] , \nScanOut121[17] , \nScanOut2[30] , \nScanOut2[29] , 
        \nOut0_3[18] , \nScanOut3[10] , \nOut0_11[0] , \nOut1_21[23] , 
        \nOut1_54[13] , \nScanOut90[14] , \nScanOut102[26] , \nOut1_30[6] , 
        \nOut1_17[15] , \nOut1_21[10] , \nScanOut28[13] , \nScanOut48[17] , 
        \nOut1_54[2] , \nOut1_57[1] , \nScanOut63[8] , \nScanOut90[27] , 
        \nScanOut121[24] , \nOut1_34[24] , \nOut1_54[20] , \nScanOut102[15] , 
        \nOut1_41[14] , \nScanOut117[21] , \nScanOut85[13] , \nOut0_19[25] , 
        \nOut1_62[25] , \nScanOut68[3] , \nOut1_7[24] , \nOut0_8[27] , 
        \nScanOut9[25] , \nOut0_13[10] , \nScanOut9[16] , \nOut0_13[23] , 
        \nScanOut14[23] , \nScanOut22[26] , \nOut0_25[15] , \nOut0_30[21] , 
        \nOut1_42[6] , \nOut0_45[11] , \nOut0_63[0] , \nOut0_50[25] , 
        \nScanOut108[20] , \nScanOut57[16] , \nScanOut61[13] , 
        \nScanOut74[27] , \nOut0_25[26] , \nScanOut37[12] , \nOut1_41[5] , 
        \nOut0_60[3] , \nScanOut42[22] , \nOut0_50[16] , \nScanOut108[13] , 
        \nScanOut11[8] , \nOut1_26[2] , \nOut0_45[22] , \nScanOut14[10] , 
        \nOut0_19[8] , \nOut0_30[12] , \nScanOut113[8] , \nScanOut22[15] , 
        \nScanOut37[21] , \nScanOut61[20] , \nScanOut42[11] , \nOut1_25[1] , 
        \nScanOut57[25] , \nOut1_59[7] , \nScanOut74[14] , \nScanOut84[19] , 
        \nOut1_44[8] , \nScanOut70[1] , \nScanOut73[2] , \nOut0_8[14] , 
        \nScanOut17[6] , \nScanOut29[19] , \nScanOut116[18] , \nScanOut116[5] , 
        \nOut1_3[26] , \nOut1_7[17] , \nOut1_20[30] , \nOut1_20[29] , 
        \nOut1_55[19] , \nScanOut115[6] , \nScanOut14[5] , \nScanOut108[9] , 
        \nScanOut30[3] , \nScanOut33[0] , \nOut1_3[15] , \nScanOut6[18] , 
        \nScanOut112[30] , \nOut1_19[5] , \nOut0_38[3] , \nOut1_24[18] , 
        \nScanOut112[29] , \nOut1_51[31] , \nOut1_51[28] , \nScanOut54[7] , 
        \nScanOut1[5] , \nScanOut49[8] , \nScanOut86[1] , \nScanOut58[18] , 
        \nScanOut2[6] , \nScanOut80[28] , \nScanOut85[2] , \nOut0_4[5] , 
        \nOut0_41[8] , \nScanOut80[31] , \nScanOut57[4] , \nScanOut4[8] , 
        \nOut0_7[6] , \nOut1_8[19] , \nScanOut10[21] , \nScanOut65[11] , 
        \nOut0_17[12] , \nOut0_20[1] , \nOut0_21[17] , \nOut0_23[2] , 
        \nScanOut26[24] , \nScanOut33[10] , \nScanOut46[20] , \nScanOut53[14] , 
        \nScanOut70[25] , \nOut0_54[27] , \nOut1_19[22] , \nOut0_62[22] , 
        \nScanOut28[1] , \nOut0_34[23] , \nOut0_41[13] , \nScanOut119[16] , 
        \nScanOut10[12] , \nScanOut26[17] , \nOut0_44[5] , \nScanOut52[9] , 
        \nScanOut53[27] , \nScanOut70[16] , \nScanOut33[23] , \nScanOut65[22] , 
        \nScanOut46[13] , \nOut0_7[30] , \nOut0_7[29] , \nOut1_7[4] , 
        \nScanOut8[22] , \nOut0_12[17] , \nOut0_17[21] , \nOut1_19[11] , 
        \nOut0_62[11] , \nOut0_21[24] , \nOut0_34[10] , \nOut0_41[20] , 
        \nOut0_47[6] , \nOut0_54[14] , \nScanOut119[25] , \nScanOut78[4] , 
        \nScanOut8[11] , \nOut0_12[24] , \nScanOut15[24] , \nScanOut23[21] , 
        \nOut0_24[12] , \nOut0_31[26] , \nOut0_44[16] , \nOut0_51[22] , 
        \nOut1_52[1] , \nScanOut109[27] , \nScanOut56[11] , \nScanOut60[14] , 
        \nScanOut75[20] , \nOut0_24[21] , \nScanOut36[15] , \nScanOut43[25] , 
        \nOut1_51[2] , \nScanOut66[8] , \nOut0_51[11] , \nScanOut109[14] , 
        \nOut0_17[3] , \nOut1_36[5] , \nOut0_44[25] , \nOut0_31[15] , 
        \nOut1_4[7] , \nOut1_28[9] , \nOut0_14[0] , \nScanOut15[17] , 
        \nScanOut23[12] , \nScanOut36[26] , \nScanOut60[27] , \nScanOut43[16] , 
        \nOut1_35[6] , \nScanOut56[22] , \nScanOut75[13] , \nOut0_1[5] , 
        \nScanOut1[8] , \nOut1_2[21] , \nOut1_2[9] , \nOut1_6[23] , 
        \nOut0_9[20] , \nOut1_17[18] , \nOut1_34[30] , \nScanOut102[18] , 
        \nScanOut121[30] , \nScanOut121[29] , \nOut0_19[31] , \nOut0_19[28] , 
        \nOut1_34[29] , \nOut1_62[28] , \nOut1_49[0] , \nOut1_41[19] , 
        \nOut1_62[31] , \nScanOut60[6] , \nScanOut63[5] , \nOut1_6[10] , 
        \nOut0_9[13] , \nScanOut48[30] , \nScanOut90[19] , \nScanOut106[2] , 
        \nScanOut105[1] , \nOut1_33[8] , \nScanOut48[29] , \nScanOut39[31] , 
        \nOut1_2[12] , \nScanOut20[4] , \nOut0_36[8] , \nScanOut39[28] , 
        \nScanOut121[7] , \nScanOut23[7] , \nOut0_28[4] , \nScanOut44[0] , 
        \nScanOut94[31] , \nScanOut94[28] , \nScanOut122[4] , \nOut1_3[18] , 
        \nScanOut6[26] , \nScanOut9[0] , \nOut1_11[0] , \nScanOut11[26] , 
        \nOut1_13[30] , \nOut1_13[29] , \nOut1_45[31] , \nScanOut95[5] , 
        \nScanOut96[6] , \nScanOut106[29] , \nScanOut106[30] , 
        \nScanOut125[18] , \nOut1_45[28] , \nOut1_30[18] , \nScanOut47[3] , 
        \nScanOut64[16] , \nScanOut127[9] , \nOut0_30[6] , \nScanOut11[15] , 
        \nOut1_12[3] , \nScanOut27[23] , \nScanOut32[17] , \nScanOut47[27] , 
        \nScanOut52[13] , \nOut0_33[5] , \nScanOut71[22] , \nOut0_16[15] , 
        \nOut0_20[10] , \nScanOut25[9] , \nOut0_55[20] , \nOut1_18[25] , 
        \nOut0_63[25] , \nScanOut27[10] , \nOut0_35[24] , \nScanOut38[6] , 
        \nOut0_40[14] , \nScanOut118[11] , \nScanOut52[20] , \nOut0_54[2] , 
        \nScanOut71[11] , \nOut0_16[26] , \nOut1_18[16] , \nScanOut32[24] , 
        \nScanOut64[25] , \nScanOut47[14] , \nOut0_63[16] , \nScanOut90[8] , 
        \nOut0_35[17] , \nOut0_40[27] , \nOut0_57[1] , \nScanOut118[22] , 
        \nOut0_20[23] , \nOut0_55[13] , \nOut1_24[26] , \nOut0_41[5] , 
        \nOut1_60[3] , \nOut1_51[16] , \nScanOut57[9] , \nScanOut95[11] , 
        \nScanOut98[0] , \nScanOut124[12] , \nScanOut107[23] , \nOut1_31[12] , 
        \nOut1_44[22] , \nScanOut112[17] , \nOut1_12[23] , \nScanOut80[25] , 
        \nScanOut38[11] , \nScanOut49[5] , \nScanOut58[15] , \nOut1_19[8] , 
        \nOut0_42[6] , \nOut1_63[0] , \nOut1_31[21] , \nOut1_44[11] , 
        \nScanOut112[24] , \nScanOut80[16] , \nOut0_2[6] , \nScanOut6[15] , 
        \nOut1_12[10] , \nOut1_24[15] , \nScanOut95[22] , \nScanOut124[21] , 
        \nOut0_25[1] , \nOut1_51[25] , \nScanOut107[10] , \nOut0_26[2] , 
        \nScanOut2[24] , \nOut0_3[26] , \nOut0_4[8] , \nScanOut4[5] , 
        \nOut0_7[24] , \nOut0_21[30] , \nScanOut38[22] , \nScanOut58[26] , 
        \nScanOut51[7] , \nScanOut119[28] , \nScanOut119[31] , \nOut0_21[29] , 
        \nOut0_54[19] , \nScanOut83[1] , \nOut0_7[17] , \nScanOut7[6] , 
        \nOut0_59[7] , \nScanOut80[2] , \nOut1_8[27] , \nOut0_44[8] , 
        \nScanOut52[4] , \nOut1_8[14] , \nScanOut35[3] , \nScanOut36[0] , 
        \nScanOut26[30] , \nScanOut70[28] , \nScanOut26[29] , \nScanOut53[19] , 
        \nScanOut70[31] , \nOut1_9[2] , \nScanOut57[31] , \nScanOut74[19] , 
        \nScanOut12[6] , \nScanOut22[18] , \nScanOut57[28] , \nOut0_19[5] , 
        \nOut1_38[3] , \nScanOut113[5] , \nOut0_3[15] , \nScanOut9[31] , 
        \nScanOut11[5] , \nScanOut110[6] , \nOut1_41[8] , \nScanOut76[2] , 
        \nScanOut9[28] , \nOut0_25[18] , \nOut0_50[31] , \nOut0_50[28] , 
        \nScanOut75[1] , \nScanOut14[8] , \nOut1_23[2] , \nScanOut108[4] , 
        \nOut0_18[11] , \nScanOut29[27] , \nOut1_35[10] , \nOut1_40[20] , 
        \nScanOut49[23] , \nScanOut116[15] , \nScanOut116[8] , \nOut1_16[21] , 
        \nOut1_63[11] , \nScanOut84[27] , \nOut1_20[24] , \nOut1_55[14] , 
        \nScanOut91[13] , \nScanOut120[10] , \nScanOut103[21] , \nOut1_7[30] , 
        \nOut0_8[19] , \nOut1_20[1] , \nScanOut49[10] , \nOut1_7[29] , 
        \nScanOut29[14] , \nOut1_44[5] , \nOut1_47[6] , \nScanOut1[1] , 
        \nScanOut2[17] , \nOut1_16[12] , \nOut1_20[17] , \nScanOut91[20] , 
        \nScanOut120[23] , \nOut1_35[23] , \nOut1_55[27] , \nScanOut103[12] , 
        \nOut1_40[13] , \nScanOut116[26] , \nScanOut84[14] , \nOut0_18[22] , 
        \nScanOut2[2] , \nOut1_3[22] , \nOut0_4[1] , \nOut0_7[2] , 
        \nOut1_63[22] , \nScanOut10[25] , \nOut0_17[16] , \nScanOut28[5] , 
        \nOut0_34[27] , \nOut0_41[17] , \nScanOut119[12] , \nOut1_19[26] , 
        \nOut0_62[26] , \nOut0_20[5] , \nOut0_21[13] , \nOut0_23[6] , 
        \nScanOut26[20] , \nScanOut53[10] , \nOut0_54[23] , \nScanOut70[21] , 
        \nScanOut33[14] , \nScanOut36[9] , \nScanOut46[24] , \nScanOut65[15] , 
        \nScanOut10[16] , \nOut0_17[25] , \nOut1_19[15] , \nOut0_21[20] , 
        \nOut0_54[10] , \nOut0_34[14] , \nOut0_41[24] , \nOut0_47[2] , 
        \nOut0_62[15] , \nScanOut119[21] , \nScanOut33[27] , \nScanOut83[8] , 
        \nScanOut46[17] , \nOut1_12[19] , \nOut1_19[1] , \nScanOut26[13] , 
        \nScanOut65[26] , \nScanOut70[12] , \nOut1_31[28] , \nOut0_38[7] , 
        \nOut0_44[1] , \nScanOut53[23] , \nScanOut107[19] , \nScanOut124[28] , 
        \nScanOut124[31] , \nOut1_31[31] , \nOut1_44[18] , \nOut0_25[8] , 
        \nScanOut30[7] , \nScanOut33[4] , \nScanOut57[0] , \nScanOut98[9] , 
        \nScanOut85[6] , \nScanOut95[18] , \nOut1_3[11] , \nScanOut38[18] , 
        \nScanOut86[5] , \nOut1_7[20] , \nScanOut49[19] , \nScanOut54[3] , 
        \nOut1_63[9] , \nScanOut70[5] , \nScanOut73[6] , \nOut1_1[3] , 
        \nOut1_7[13] , \nOut0_8[23] , \nScanOut14[1] , \nOut1_59[3] , 
        \nScanOut91[30] , \nScanOut91[29] , \nOut0_8[10] , \nOut1_16[31] , 
        \nOut1_40[29] , \nScanOut103[31] , \nScanOut115[2] , \nScanOut120[19] , 
        \nScanOut103[28] , \nScanOut116[1] , \nOut1_16[28] , \nOut0_18[18] , 
        \nOut1_35[19] , \nOut1_40[30] , \nOut1_63[18] , \nScanOut9[21] , 
        \nOut0_13[14] , \nScanOut14[27] , \nScanOut17[2] , \nOut1_20[8] , 
        \nScanOut37[16] , \nOut1_41[1] , \nOut0_60[7] , \nScanOut42[26] , 
        \nScanOut61[17] , \nScanOut22[22] , \nScanOut57[12] , \nScanOut74[23] , 
        \nOut0_25[11] , \nOut0_63[4] , \nOut0_30[25] , \nOut1_42[2] , 
        \nScanOut108[24] , \nOut0_50[21] , \nScanOut75[8] , \nOut0_45[15] , 
        \nScanOut9[12] , \nOut0_13[27] , \nScanOut14[14] , \nScanOut22[11] , 
        \nScanOut68[7] , \nScanOut74[10] , \nOut1_25[5] , \nScanOut37[25] , 
        \nScanOut57[21] , \nScanOut42[15] , \nOut1_26[6] , \nScanOut61[24] , 
        \nOut0_30[16] , \nOut0_45[26] , \nOut0_11[4] , \nOut0_25[22] , 
        \nOut0_50[12] , \nOut1_30[2] , \nScanOut108[17] , \nOut1_21[27] , 
        \nOut1_54[17] , \nScanOut102[22] , \nScanOut121[13] , \nOut0_2[25] , 
        \nOut1_2[0] , \nScanOut3[27] , \nOut0_19[12] , \nScanOut90[10] , 
        \nOut1_6[19] , \nOut1_17[22] , \nOut1_62[12] , \nScanOut85[24] , 
        \nOut1_34[13] , \nOut1_41[23] , \nScanOut117[16] , \nScanOut3[14] , 
        \nOut0_12[7] , \nScanOut19[4] , \nScanOut48[20] , \nScanOut28[24] , 
        \nScanOut105[8] , \nOut1_33[1] , \nOut1_17[11] , \nScanOut85[17] , 
        \nScanOut118[7] , \nOut0_19[21] , \nScanOut8[18] , \nOut0_9[30] , 
        \nOut1_21[14] , \nOut1_34[20] , \nOut1_49[9] , \nOut1_62[21] , 
        \nOut1_41[10] , \nScanOut117[25] , \nOut1_54[24] , \nOut1_54[6] , 
        \nScanOut90[23] , \nScanOut102[11] , \nScanOut121[20] , \nOut0_9[29] , 
        \nScanOut28[17] , \nOut1_57[5] , \nScanOut48[13] , \nOut0_24[31] , 
        \nOut0_24[28] , \nOut0_51[18] , \nScanOut100[5] , \nOut1_1[1] , 
        \nOut0_2[16] , \nOut0_14[9] , \nOut1_28[0] , \nScanOut103[6] , 
        \nOut1_2[31] , \nOut1_2[28] , \nOut0_6[27] , \nOut1_9[24] , 
        \nScanOut23[31] , \nScanOut23[28] , \nOut1_52[8] , \nScanOut56[18] , 
        \nScanOut65[2] , \nScanOut66[1] , \nScanOut75[30] , \nScanOut75[29] , 
        \nScanOut27[19] , \nScanOut42[7] , \nScanOut52[29] , \nOut0_49[4] , 
        \nScanOut52[30] , \nScanOut71[18] , \nScanOut90[1] , \nOut0_6[14] , 
        \nOut0_9[4] , \nScanOut9[9] , \nScanOut93[2] , \nScanOut41[4] , 
        \nOut0_57[8] , \nScanOut127[0] , \nOut1_9[17] , \nOut1_11[9] , 
        \nOut0_20[19] , \nScanOut26[3] , \nScanOut118[18] , \nScanOut25[0] , 
        \nOut0_55[30] , \nOut0_55[29] , \nScanOut124[3] , \nScanOut7[25] , 
        \nScanOut39[12] , \nScanOut44[9] , \nOut0_52[5] , \nScanOut59[16] , 
        \nScanOut59[6] , \nOut1_13[20] , \nScanOut81[26] , \nOut1_25[25] , 
        \nOut1_30[11] , \nOut1_45[21] , \nScanOut113[14] , \nOut1_50[15] , 
        \nScanOut106[20] , \nOut0_51[6] , \nScanOut94[12] , \nScanOut125[11] , 
        \nScanOut88[3] , \nScanOut39[21] , \nOut1_2[2] , \nScanOut7[16] , 
        \nOut1_13[13] , \nOut1_14[4] , \nOut1_17[7] , \nOut0_36[1] , 
        \nScanOut59[25] , \nOut0_35[2] , \nOut1_25[16] , \nOut1_50[26] , 
        \nScanOut81[15] , \nScanOut94[21] , \nScanOut106[13] , 
        \nScanOut125[22] , \nOut0_12[5] , \nOut1_30[22] , \nOut1_45[12] , 
        \nScanOut113[27] , \nScanOut118[5] , \nScanOut28[26] , \nOut1_33[3] , 
        \nScanOut3[25] , \nOut1_17[20] , \nScanOut19[6] , \nScanOut48[22] , 
        \nScanOut85[26] , \nOut0_19[10] , \nOut1_62[10] , \nOut1_21[25] , 
        \nOut1_34[11] , \nOut1_41[21] , \nScanOut106[9] , \nScanOut117[14] , 
        \nOut1_54[15] , \nScanOut102[20] , \nScanOut1[3] , \nOut0_2[27] , 
        \nScanOut3[16] , \nOut1_6[31] , \nOut1_6[28] , \nOut0_9[18] , 
        \nOut0_11[6] , \nScanOut90[12] , \nScanOut121[11] , \nOut1_30[0] , 
        \nOut0_19[23] , \nOut1_21[16] , \nScanOut28[15] , \nScanOut48[11] , 
        \nOut1_54[26] , \nOut1_54[4] , \nOut1_57[7] , \nScanOut102[13] , 
        \nScanOut90[21] , \nScanOut121[22] , \nOut1_62[23] , \nOut1_17[13] , 
        \nScanOut85[15] , \nScanOut23[19] , \nOut1_34[22] , \nOut1_41[12] , 
        \nScanOut117[27] , \nScanOut56[29] , \nOut1_28[2] , \nScanOut56[30] , 
        \nScanOut75[18] , \nScanOut103[4] , \nScanOut100[7] , \nOut0_2[14] , 
        \nScanOut8[30] , \nScanOut8[29] , \nOut0_17[8] , \nOut1_51[9] , 
        \nScanOut66[3] , \nOut0_24[19] , \nOut0_51[29] , \nScanOut65[0] , 
        \nOut0_51[30] , \nOut1_2[19] , \nOut0_6[25] , \nOut0_20[31] , 
        \nOut0_20[28] , \nScanOut41[6] , \nScanOut118[30] , \nScanOut118[29] , 
        \nOut0_55[18] , \nScanOut93[0] , \nOut0_6[16] , \nOut1_9[26] , 
        \nScanOut42[5] , \nOut0_49[6] , \nScanOut90[3] , \nOut0_54[9] , 
        \nScanOut7[27] , \nOut0_9[6] , \nOut1_12[8] , \nScanOut25[2] , 
        \nScanOut124[1] , \nOut1_9[15] , \nOut1_13[22] , \nOut1_25[27] , 
        \nScanOut26[1] , \nScanOut27[31] , \nScanOut27[28] , \nScanOut52[18] , 
        \nScanOut71[30] , \nScanOut47[8] , \nScanOut71[29] , \nScanOut127[2] , 
        \nOut0_51[4] , \nScanOut88[1] , \nOut1_50[17] , \nScanOut81[24] , 
        \nScanOut94[10] , \nScanOut106[22] , \nScanOut125[13] , \nOut1_30[13] , 
        \nOut1_45[23] , \nScanOut113[16] , \nOut1_3[20] , \nOut0_4[3] , 
        \nScanOut7[14] , \nScanOut39[10] , \nScanOut59[4] , \nOut0_52[7] , 
        \nScanOut59[14] , \nOut1_13[11] , \nScanOut81[17] , \nOut1_14[6] , 
        \nOut1_25[14] , \nOut1_30[20] , \nOut1_45[10] , \nScanOut113[25] , 
        \nOut1_50[24] , \nScanOut106[11] , \nScanOut94[23] , \nScanOut125[20] , 
        \nOut1_17[5] , \nOut0_35[0] , \nOut0_36[3] , \nScanOut39[23] , 
        \nScanOut59[27] , \nOut0_7[0] , \nScanOut10[27] , \nOut0_20[7] , 
        \nScanOut33[16] , \nScanOut46[26] , \nOut0_17[14] , \nOut1_19[24] , 
        \nOut0_21[11] , \nScanOut26[22] , \nScanOut65[17] , \nScanOut70[23] , 
        \nScanOut35[8] , \nScanOut53[12] , \nOut0_54[21] , \nOut0_23[4] , 
        \nOut0_34[25] , \nOut0_41[15] , \nScanOut119[10] , \nOut0_62[24] , 
        \nScanOut10[14] , \nScanOut26[11] , \nScanOut28[7] , \nScanOut53[21] , 
        \nScanOut70[10] , \nScanOut33[25] , \nOut0_44[3] , \nScanOut46[15] , 
        \nScanOut65[24] , \nOut0_17[27] , \nOut0_34[16] , \nScanOut80[9] , 
        \nScanOut119[23] , \nOut0_41[26] , \nOut0_47[0] , \nOut1_19[17] , 
        \nOut0_62[17] , \nOut0_21[22] , \nScanOut38[29] , \nOut0_54[12] , 
        \nOut1_3[13] , \nOut1_19[3] , \nOut0_26[9] , \nScanOut30[5] , 
        \nScanOut38[30] , \nScanOut33[6] , \nOut0_38[5] , \nScanOut54[1] , 
        \nScanOut95[30] , \nScanOut95[29] , \nScanOut86[7] , \nScanOut2[0] , 
        \nOut1_12[31] , \nOut1_31[19] , \nScanOut85[4] , \nScanOut107[31] , 
        \nScanOut124[19] , \nScanOut107[28] , \nOut1_7[22] , \nOut0_8[21] , 
        \nOut1_12[28] , \nOut1_44[29] , \nOut1_16[19] , \nOut0_18[30] , 
        \nOut1_44[30] , \nScanOut57[2] , \nOut1_60[8] , \nScanOut103[19] , 
        \nScanOut120[31] , \nScanOut120[28] , \nOut0_18[29] , \nOut1_35[28] , 
        \nOut1_40[18] , \nOut1_59[1] , \nOut1_63[30] , \nOut1_63[29] , 
        \nOut1_35[31] , \nScanOut70[7] , \nScanOut73[4] , \nOut0_1[7] , 
        \nScanEnable[0] , \nScanOut2[9] , \nOut1_7[11] , \nOut0_8[12] , 
        \nScanOut17[0] , \nScanOut49[28] , \nScanOut91[18] , \nScanOut116[3] , 
        \nScanOut115[0] , \nOut1_9[9] , \nScanOut9[23] , \nOut0_13[16] , 
        \nScanOut14[3] , \nScanOut49[31] , \nOut1_23[9] , \nOut0_30[27] , 
        \nOut0_45[17] , \nScanOut68[5] , \nScanOut9[10] , \nOut0_13[25] , 
        \nScanOut14[25] , \nScanOut22[20] , \nOut0_25[13] , \nOut1_42[0] , 
        \nOut0_50[23] , \nScanOut108[26] , \nOut0_63[6] , \nScanOut74[21] , 
        \nScanOut37[14] , \nScanOut57[10] , \nScanOut76[9] , \nOut1_41[3] , 
        \nScanOut42[24] , \nOut0_60[5] , \nOut0_25[20] , \nScanOut61[15] , 
        \nScanOut108[15] , \nOut1_26[4] , \nOut0_30[14] , \nOut0_50[10] , 
        \nOut0_45[24] , \nScanOut14[16] , \nScanOut37[27] , \nOut1_38[8] , 
        \nScanOut42[17] , \nScanOut61[26] , \nScanOut74[12] , \nScanOut22[13] , 
        \nScanOut57[23] , \nOut1_25[7] , \nOut1_31[10] , \nScanOut38[13] , 
        \nOut0_42[4] , \nScanOut54[8] , \nScanOut49[7] , \nScanOut58[17] , 
        \nOut1_63[2] , \nScanOut112[15] , \nScanOut6[24] , \nOut1_12[21] , 
        \nOut1_44[20] , \nScanOut80[27] , \nScanOut95[13] , \nScanOut124[10] , 
        \nOut0_2[4] , \nOut1_3[30] , \nOut1_24[24] , \nOut0_41[7] , 
        \nOut1_51[14] , \nScanOut98[2] , \nScanOut107[21] , \nOut1_60[1] , 
        \nOut1_3[29] , \nScanOut38[20] , \nScanOut6[17] , \nOut1_24[17] , 
        \nOut0_25[3] , \nOut0_26[0] , \nScanOut58[24] , \nOut1_51[27] , 
        \nScanOut95[20] , \nScanOut124[23] , \nScanOut107[12] , \nOut1_31[23] , 
        \nOut1_44[13] , \nScanOut112[26] , \nOut1_12[12] , \nScanOut80[14] , 
        \nOut0_3[24] , \nScanOut4[7] , \nOut0_7[26] , \nScanOut7[4] , 
        \nOut1_8[25] , \nScanOut26[18] , \nScanOut52[6] , \nScanOut53[31] , 
        \nScanOut53[28] , \nScanOut70[19] , \nOut0_59[5] , \nScanOut80[0] , 
        \nOut0_7[15] , \nOut0_7[9] , \nOut1_8[16] , \nScanOut36[2] , 
        \nOut0_47[9] , \nScanOut51[5] , \nScanOut83[3] , \nOut0_21[18] , 
        \nScanOut35[1] , \nOut0_54[31] , \nScanOut119[19] , \nOut0_54[28] , 
        \nScanOut9[19] , \nScanOut11[7] , \nOut0_25[30] , \nOut0_25[29] , 
        \nOut0_50[19] , \nOut0_3[17] , \nOut1_9[0] , \nOut0_19[7] , 
        \nScanOut110[4] , \nOut1_38[1] , \nScanOut113[7] , \nScanOut12[4] , 
        \nScanOut17[9] , \nScanOut22[30] , \nOut1_42[9] , \nScanOut75[3] , 
        \nScanOut76[0] , \nScanOut22[29] , \nScanOut74[28] , \nScanOut57[19] , 
        \nScanOut74[31] , \nOut1_20[3] , \nScanOut2[26] , \nOut1_16[23] , 
        \nOut1_20[26] , \nScanOut91[11] , \nScanOut120[12] , \nOut1_35[12] , 
        \nOut1_55[16] , \nScanOut103[23] , \nOut1_40[22] , \nScanOut116[17] , 
        \nScanOut84[25] , \nOut0_18[13] , \nOut1_63[13] , \nScanOut2[15] , 
        \nOut1_7[18] , \nScanOut49[21] , \nOut0_18[20] , \nOut1_23[0] , 
        \nScanOut29[25] , \nScanOut115[9] , \nOut1_35[21] , \nOut1_40[11] , 
        \nScanOut108[6] , \nScanOut116[24] , \nOut1_59[8] , \nOut1_63[20] , 
        \nOut1_16[10] , \nScanOut84[16] , \nOut1_20[15] , \nOut1_55[25] , 
        \nScanOut91[22] , \nScanOut120[21] , \nScanOut103[10] , \nOut0_8[31] , 
        \nOut0_8[28] , \nOut1_44[7] , \nScanOut8[20] , \nOut0_12[15] , 
        \nScanOut15[26] , \nScanOut29[16] , \nOut1_47[4] , \nScanOut49[12] , 
        \nScanOut23[23] , \nScanOut36[17] , \nScanOut60[16] , \nScanOut43[27] , 
        \nOut1_51[0] , \nOut0_24[10] , \nOut0_51[20] , \nScanOut56[13] , 
        \nScanOut65[9] , \nScanOut75[22] , \nOut1_52[3] , \nScanOut109[25] , 
        \nOut0_14[2] , \nScanOut23[10] , \nOut0_31[24] , \nOut0_44[14] , 
        \nScanOut56[20] , \nScanOut78[6] , \nScanOut15[15] , \nOut1_35[4] , 
        \nScanOut60[25] , \nScanOut75[11] , \nScanOut36[24] , \nScanOut43[14] , 
        \nOut1_1[8] , \nOut1_4[5] , \nOut1_6[21] , \nOut1_7[6] , 
        \nScanOut8[13] , \nOut0_12[26] , \nOut0_17[1] , \nOut0_31[17] , 
        \nOut0_24[23] , \nOut1_36[7] , \nOut0_44[27] , \nScanOut109[16] , 
        \nOut0_51[13] , \nOut1_6[12] , \nOut0_9[22] , \nScanOut48[18] , 
        \nScanOut60[4] , \nScanOut63[7] , \nOut1_49[2] , \nScanOut90[31] , 
        \nScanOut90[28] , \nScanOut102[29] , \nScanOut105[3] , \nScanOut1[7] , 
        \nOut0_2[9] , \nOut1_2[23] , \nOut0_9[11] , \nOut1_17[30] , 
        \nOut1_17[29] , \nScanOut102[30] , \nScanOut121[18] , \nOut0_19[19] , 
        \nOut1_34[18] , \nOut1_41[31] , \nOut1_62[19] , \nOut1_30[9] , 
        \nOut1_41[28] , \nScanOut106[0] , \nOut1_13[18] , \nScanOut106[18] , 
        \nScanOut125[30] , \nScanOut122[6] , \nScanOut125[29] , 
        \nScanOut20[6] , \nScanOut23[5] , \nOut0_28[6] , \nOut1_30[30] , 
        \nOut1_45[19] , \nOut1_30[29] , \nOut0_35[9] , \nOut1_2[10] , 
        \nScanOut47[1] , \nScanOut121[5] , \nScanOut88[8] , \nScanOut94[19] , 
        \nScanOut95[7] , \nScanOut2[18] , \nOut0_3[30] , \nScanOut9[27] , 
        \nScanOut9[2] , \nOut1_11[2] , \nScanOut11[24] , \nOut1_12[1] , 
        \nOut0_16[17] , \nOut1_18[27] , \nScanOut38[4] , \nScanOut39[19] , 
        \nScanOut96[4] , \nScanOut44[2] , \nScanOut124[8] , \nOut0_63[27] , 
        \nOut0_20[12] , \nOut0_35[26] , \nOut0_40[16] , \nScanOut118[13] , 
        \nOut0_55[22] , \nScanOut27[21] , \nOut0_33[7] , \nScanOut52[11] , 
        \nScanOut71[20] , \nScanOut26[8] , \nScanOut64[14] , \nScanOut32[15] , 
        \nOut0_20[21] , \nOut0_30[4] , \nScanOut47[25] , \nScanOut11[17] , 
        \nOut0_16[24] , \nOut0_55[11] , \nOut1_18[14] , \nOut0_63[14] , 
        \nOut0_35[15] , \nScanOut118[20] , \nOut0_40[25] , \nOut0_57[3] , 
        \nScanOut64[27] , \nScanOut93[9] , \nOut0_13[12] , \nScanOut14[21] , 
        \nScanOut27[12] , \nScanOut32[26] , \nScanOut47[16] , \nScanOut52[22] , 
        \nOut0_54[0] , \nScanOut71[13] , \nScanOut22[24] , \nScanOut37[10] , 
        \nScanOut61[11] , \nOut1_41[7] , \nScanOut42[20] , \nOut0_60[1] , 
        \nOut0_25[17] , \nOut0_50[27] , \nScanOut57[14] , \nScanOut74[25] , 
        \nScanOut108[22] , \nOut1_42[4] , \nOut0_63[2] , \nScanOut12[9] , 
        \nOut0_30[23] , \nOut0_45[13] , \nScanOut57[27] , \nScanOut68[1] , 
        \nScanOut14[12] , \nScanOut22[17] , \nOut1_25[3] , \nScanOut61[22] , 
        \nScanOut74[16] , \nScanOut37[23] , \nScanOut42[13] , \nOut0_3[29] , 
        \nScanOut110[9] , \nOut1_7[26] , \nScanOut9[14] , \nOut0_13[21] , 
        \nOut0_25[24] , \nOut1_26[0] , \nOut0_30[10] , \nOut0_45[20] , 
        \nScanOut108[11] , \nOut0_50[14] , \nOut0_8[25] , \nOut1_47[9] , 
        \nScanOut70[3] , \nScanOut73[0] , \nScanOut116[30] , \nOut1_3[24] , 
        \nOut1_7[15] , \nScanOut14[7] , \nOut1_20[18] , \nOut1_55[28] , 
        \nOut1_59[5] , \nScanOut116[29] , \nOut1_55[31] , \nOut0_8[16] , 
        \nScanOut17[4] , \nScanOut29[31] , \nScanOut29[28] , \nScanOut115[4] , 
        \nScanOut84[31] , \nScanOut84[28] , \nScanOut116[7] , \nOut1_19[7] , 
        \nScanOut80[19] , \nScanOut30[1] , \nScanOut33[2] , \nOut0_38[1] , 
        \nScanOut58[30] , \nScanOut58[29] , \nScanOut2[4] , \nScanOut6[29] , 
        \nScanOut57[6] , \nScanOut112[18] , \nScanOut6[30] , \nOut1_24[30] , 
        \nOut1_24[29] , \nOut1_51[19] , \nScanOut85[0] , \nOut1_1[5] , 
        \nOut0_2[23] , \nOut1_3[17] , \nOut0_4[7] , \nOut0_7[18] , 
        \nOut0_7[4] , \nScanOut28[3] , \nOut0_42[9] , \nScanOut54[5] , 
        \nScanOut86[3] , \nScanOut10[23] , \nOut0_17[10] , \nOut1_19[20] , 
        \nOut0_62[20] , \nOut0_21[15] , \nOut0_34[21] , \nOut0_41[11] , 
        \nScanOut119[14] , \nOut0_54[25] , \nOut0_23[0] , \nScanOut26[26] , 
        \nScanOut53[16] , \nScanOut70[27] , \nOut0_20[3] , \nScanOut33[12] , 
        \nScanOut65[13] , \nScanOut46[22] , \nOut0_6[21] , \nScanOut7[23] , 
        \nScanOut7[9] , \nOut0_17[23] , \nOut0_21[26] , \nOut0_54[16] , 
        \nOut1_19[13] , \nOut0_62[13] , \nOut0_34[12] , \nScanOut119[27] , 
        \nOut0_41[22] , \nOut0_47[4] , \nScanOut51[8] , \nOut1_8[31] , 
        \nOut1_8[28] , \nOut0_59[8] , \nScanOut65[20] , \nScanOut10[10] , 
        \nScanOut46[11] , \nOut1_13[26] , \nScanOut26[15] , \nScanOut33[21] , 
        \nScanOut53[25] , \nOut1_30[17] , \nScanOut39[14] , \nOut0_44[7] , 
        \nOut0_52[3] , \nScanOut70[14] , \nScanOut59[10] , \nScanOut59[0] , 
        \nScanOut96[9] , \nOut1_45[27] , \nScanOut113[12] , \nScanOut81[20] , 
        \nScanOut7[10] , \nOut1_14[2] , \nOut1_17[1] , \nOut1_25[23] , 
        \nScanOut94[14] , \nScanOut125[17] , \nScanOut39[27] , \nOut1_50[13] , 
        \nOut0_51[0] , \nScanOut88[5] , \nScanOut106[26] , \nScanOut121[8] , 
        \nScanOut59[23] , \nScanOut23[8] , \nOut0_36[7] , \nOut1_25[10] , 
        \nOut0_35[4] , \nOut1_50[20] , \nScanOut94[27] , \nScanOut125[24] , 
        \nScanOut106[15] , \nOut1_30[24] , \nOut1_45[14] , \nScanOut113[21] , 
        \nOut1_9[22] , \nOut1_13[15] , \nScanOut81[13] , \nScanOut42[1] , 
        \nOut0_49[2] , \nScanOut90[7] , \nOut0_6[12] , \nOut0_9[2] , 
        \nScanOut11[30] , \nOut0_16[30] , \nScanOut41[2] , \nScanOut93[4] , 
        \nOut0_16[29] , \nOut0_35[18] , \nOut0_40[28] , \nOut1_18[19] , 
        \nOut0_40[31] , \nOut0_63[19] , \nScanOut26[5] , \nScanOut127[6] , 
        \nScanOut11[29] , \nOut0_30[9] , \nScanOut32[18] , \nScanOut47[28] , 
        \nOut1_9[11] , \nScanOut47[31] , \nScanOut25[6] , \nScanOut64[19] , 
        \nScanOut124[5] , \nScanOut38[9] , \nOut0_2[10] , \nOut1_4[8] , 
        \nScanOut100[3] , \nScanOut15[18] , \nOut1_28[6] , \nOut1_35[9] , 
        \nScanOut103[0] , \nScanOut36[30] , \nScanOut36[29] , \nScanOut43[19] , 
        \nScanOut60[31] , \nScanOut60[28] , \nOut0_11[2] , \nOut0_12[18] , 
        \nOut0_31[30] , \nOut0_31[29] , \nOut0_44[19] , \nScanOut65[4] , 
        \nScanOut109[31] , \nScanOut109[28] , \nScanOut66[7] , \nOut1_30[4] , 
        \nOut0_2[19] , \nOut1_2[27] , \nOut1_2[6] , \nScanOut3[21] , 
        \nOut1_17[24] , \nOut1_21[21] , \nScanOut90[16] , \nScanOut121[15] , 
        \nOut1_34[15] , \nOut1_54[11] , \nScanOut102[24] , \nOut1_41[25] , 
        \nScanOut117[10] , \nScanOut85[22] , \nOut0_19[14] , \nScanOut19[2] , 
        \nOut1_62[14] , \nScanOut48[26] , \nScanOut3[12] , \nOut0_12[1] , 
        \nScanOut28[22] , \nOut0_19[27] , \nOut1_33[7] , \nOut1_34[26] , 
        \nOut1_41[16] , \nScanOut117[23] , \nScanOut118[1] , \nOut0_6[31] , 
        \nOut0_6[28] , \nOut1_9[18] , \nOut1_11[6] , \nOut1_17[17] , 
        \nOut1_62[27] , \nScanOut85[11] , \nOut1_21[12] , \nOut1_54[22] , 
        \nScanOut90[25] , \nScanOut121[26] , \nScanOut102[17] , 
        \nScanOut28[11] , \nOut1_54[0] , \nOut1_57[3] , \nScanOut60[9] , 
        \nScanOut32[11] , \nScanOut48[15] , \nScanOut11[20] , \nOut0_30[0] , 
        \nScanOut47[21] , \nScanOut64[10] , \nScanOut11[13] , \nOut1_12[5] , 
        \nScanOut27[25] , \nScanOut71[24] , \nScanOut52[15] , \nOut0_55[26] , 
        \nOut0_16[13] , \nOut1_18[23] , \nOut0_20[16] , \nOut0_33[3] , 
        \nOut0_35[22] , \nOut0_40[12] , \nScanOut118[17] , \nOut0_63[23] , 
        \nScanOut27[16] , \nScanOut38[0] , \nScanOut42[8] , \nScanOut52[26] , 
        \nScanOut71[17] , \nScanOut32[22] , \nScanOut47[12] , \nOut0_54[4] , 
        \nScanOut64[23] , \nScanOut9[6] , \nOut0_16[20] , \nOut0_35[11] , 
        \nScanOut118[24] , \nOut0_40[21] , \nOut0_57[7] , \nOut1_18[10] , 
        \nOut0_63[10] , \nOut0_20[25] , \nOut0_55[15] , \nScanOut121[1] , 
        \nOut1_2[14] , \nScanOut7[19] , \nOut1_17[8] , \nScanOut20[2] , 
        \nScanOut23[1] , \nOut0_28[2] , \nScanOut113[28] , \nScanOut113[31] , 
        \nOut1_25[19] , \nOut1_50[30] , \nOut1_50[29] , \nScanOut44[6] , 
        \nScanOut122[2] , \nScanOut59[9] , \nScanOut96[0] , \nScanOut3[31] , 
        \nOut1_6[25] , \nOut0_9[26] , \nScanOut47[5] , \nScanOut59[19] , 
        \nScanOut81[30] , \nScanOut95[3] , \nScanOut81[29] , \nOut1_49[6] , 
        \nOut0_51[9] , \nScanOut85[18] , \nOut1_54[9] , \nScanOut63[3] , 
        \nScanOut60[0] , \nOut0_9[15] , \nScanOut28[18] , \nScanOut106[4] , 
        \nScanOut117[19] , \nScanOut3[28] , \nOut1_6[16] , \nOut1_21[31] , 
        \nOut1_21[28] , \nOut1_54[18] , \nScanOut105[7] , \nOut0_12[8] , 
        \nScanOut118[8] , \nOut1_4[1] , \nOut1_7[2] , \nScanOut8[24] , 
        \nOut0_12[11] , \nOut0_31[20] , \nOut0_44[10] , \nScanOut78[2] , 
        \nScanOut8[17] , \nOut0_12[22] , \nScanOut15[22] , \nScanOut23[27] , 
        \nOut0_24[14] , \nOut0_51[24] , \nScanOut109[21] , \nOut1_52[7] , 
        \nScanOut75[26] , \nScanOut36[13] , \nScanOut56[17] , \nScanOut43[23] , 
        \nOut1_51[4] , \nOut0_17[5] , \nOut0_24[27] , \nScanOut60[12] , 
        \nScanOut109[12] , \nOut0_31[13] , \nOut0_51[17] , \nOut1_36[3] , 
        \nOut0_44[23] , \nScanOut103[9] , \nScanOut2[22] , \nOut0_14[6] , 
        \nScanOut15[11] , \nScanOut36[20] , \nScanOut43[10] , \nScanOut60[21] , 
        \nScanOut23[14] , \nScanOut56[24] , \nScanOut75[15] , \nOut1_16[27] , 
        \nOut1_23[4] , \nOut1_35[0] , \nScanOut108[2] , \nScanOut29[21] , 
        \nScanOut49[25] , \nScanOut84[21] , \nOut0_18[17] , \nOut1_20[22] , 
        \nOut1_35[16] , \nOut1_63[17] , \nOut1_40[26] , \nScanOut116[13] , 
        \nOut1_55[12] , \nScanOut91[15] , \nScanOut103[27] , \nScanOut120[16] , 
        \nOut1_20[7] , \nScanOut29[12] , \nScanOut49[16] , \nOut1_47[0] , 
        \nScanOut73[9] , \nOut0_1[26] , \nOut0_1[15] , \nOut0_1[3] , 
        \nScanOut2[11] , \nOut0_18[24] , \nOut1_20[11] , \nOut1_44[3] , 
        \nOut1_55[21] , \nScanOut103[14] , \nScanOut91[26] , \nScanOut120[25] , 
        \nOut0_3[20] , \nOut1_9[4] , \nScanOut12[0] , \nOut1_16[14] , 
        \nOut1_63[24] , \nScanOut84[12] , \nOut1_35[25] , \nOut1_40[15] , 
        \nScanOut116[20] , \nOut0_19[3] , \nScanOut113[3] , \nOut1_38[5] , 
        \nScanOut110[0] , \nOut0_3[13] , \nScanOut11[3] , \nOut0_13[31] , 
        \nOut0_13[28] , \nScanOut108[18] , \nOut0_45[30] , \nScanOut14[31] , 
        \nScanOut14[28] , \nOut1_26[9] , \nOut0_30[19] , \nOut0_45[29] , 
        \nScanOut42[30] , \nScanOut61[18] , \nScanOut76[4] , \nScanOut37[19] , 
        \nScanOut42[29] , \nOut0_60[8] , \nScanOut68[8] , \nScanOut75[7] , 
        \nScanOut4[3] , \nScanOut51[1] , \nScanOut83[7] , \nScanOut6[20] , 
        \nOut0_7[22] , \nOut0_7[11] , \nScanOut7[0] , \nOut0_59[1] , 
        \nScanOut80[4] , \nOut1_8[21] , \nScanOut52[2] , \nScanOut10[19] , 
        \nScanOut33[31] , \nScanOut65[29] , \nScanOut33[28] , \nScanOut46[18] , 
        \nScanOut65[30] , \nOut1_8[12] , \nOut0_17[19] , \nOut1_19[29] , 
        \nOut0_23[9] , \nScanOut35[5] , \nOut0_62[29] , \nOut0_34[31] , 
        \nOut1_19[30] , \nOut0_41[18] , \nOut0_62[30] , \nOut0_34[28] , 
        \nOut1_12[25] , \nOut1_24[20] , \nScanOut36[6] , \nOut0_41[3] , 
        \nScanOut98[6] , \nOut1_60[5] , \nOut1_51[10] , \nScanOut85[9] , 
        \nScanOut80[23] , \nScanOut95[17] , \nScanOut107[25] , 
        \nScanOut124[14] , \nScanOut6[13] , \nOut1_31[14] , \nScanOut38[17] , 
        \nOut1_44[24] , \nScanOut112[11] , \nScanOut49[3] , \nOut0_42[0] , 
        \nScanOut58[13] , \nOut1_63[6] , \nScanOut80[10] , \nScanOut0[24] , 
        \nScanOut0[17] , \nOut0_2[0] , \nOut1_12[16] , \nOut1_24[13] , 
        \nOut1_31[27] , \nOut0_38[8] , \nOut1_44[17] , \nScanOut112[22] , 
        \nOut1_51[23] , \nScanOut107[16] , \nOut0_25[7] , \nScanOut95[24] , 
        \nScanOut124[27] , \nOut0_26[4] , \nScanOut30[8] , \nScanOut58[20] , 
        \nOut1_5[30] , \nOut1_5[29] , \nScanOut38[24] , \nScanOut68[21] , 
        \nOut0_45[3] , \nOut0_46[0] , \nOut0_5[3] , \nOut0_6[0] , 
        \nOut1_14[12] , \nOut1_61[22] , \nOut0_22[4] , \nOut1_22[17] , 
        \nOut1_37[23] , \nOut0_39[13] , \nOut1_42[13] , \nScanOut86[14] , 
        \nScanOut81[9] , \nScanOut114[26] , \nOut1_57[27] , \nScanOut101[12] , 
        \nOut0_59[17] , \nScanOut34[8] , \nScanOut93[20] , \nScanOut122[23] , 
        \nScanOut68[12] , \nScanOut128[4] , \nOut1_22[24] , \nScanOut29[7] , 
        \nOut0_59[24] , \nOut1_57[14] , \nScanOut101[21] , \nScanOut93[13] , 
        \nScanOut122[10] , \nOut1_14[21] , \nScanOut86[27] , \nScanOut3[0] , 
        \nOut0_21[7] , \nOut1_37[10] , \nOut1_61[11] , \nOut0_39[20] , 
        \nOut1_42[20] , \nScanOut114[15] , \nScanOut84[4] , \nOut0_27[18] , 
        \nOut1_29[28] , \nOut0_52[28] , \nScanOut55[1] , \nScanOut56[2] , 
        \nOut1_61[8] , \nOut1_29[31] , \nOut0_52[31] , \nScanOut87[7] , 
        \nScanOut0[3] , \nOut1_18[3] , \nScanOut20[18] , \nScanOut32[6] , 
        \nScanOut55[28] , \nScanOut55[31] , \nScanOut76[19] , \nOut0_39[5] , 
        \nScanOut4[26] , \nScanOut4[15] , \nOut0_5[24] , \nOut0_5[17] , 
        \nOut0_27[9] , \nScanOut31[5] , \nScanOut114[0] , \nScanOut15[3] , 
        \nScanOut89[30] , \nScanOut89[29] , \nScanOut16[0] , \nOut1_22[9] , 
        \nScanOut24[30] , \nScanOut24[29] , \nScanOut51[19] , \nScanOut72[31] , 
        \nScanOut72[28] , \nOut0_23[30] , \nOut0_23[29] , \nScanOut117[3] , 
        \nOut0_56[19] , \nOut1_58[29] , \nOut1_58[30] , \nScanOut71[7] , 
        \nOut1_26[15] , \nOut0_28[25] , \nOut1_58[1] , \nScanOut72[4] , 
        \nOut1_53[25] , \nScanOut105[10] , \nScanOut97[22] , \nScanOut126[21] , 
        \nOut1_8[9] , \nOut1_10[10] , \nOut1_33[21] , \nOut1_39[8] , 
        \nOut1_46[11] , \nScanOut82[16] , \nScanOut110[24] , \nOut0_48[21] , 
        \nOut1_10[23] , \nScanOut19[13] , \nOut1_24[7] , \nOut1_27[4] , 
        \nOut1_40[3] , \nScanOut77[9] , \nScanOut79[17] , \nOut0_61[5] , 
        \nScanOut82[25] , \nOut1_26[26] , \nOut1_33[12] , \nOut1_46[22] , 
        \nOut0_48[12] , \nScanOut110[17] , \nOut0_28[16] , \nOut1_53[16] , 
        \nScanOut105[23] , \nScanOut97[11] , \nOut1_0[21] , \nOut1_0[12] , 
        \nOut1_0[1] , \nOut1_1[18] , \nScanOut19[20] , \nScanOut79[24] , 
        \nScanOut126[12] , \nScanOut13[15] , \nScanOut30[24] , \nOut1_43[0] , 
        \nScanOut69[5] , \nScanOut45[14] , \nOut0_62[6] , \nScanOut66[25] , 
        \nOut0_14[26] , \nOut0_22[23] , \nScanOut25[10] , \nScanOut50[20] , 
        \nScanOut73[11] , \nOut1_55[4] , \nOut0_37[17] , \nOut0_57[13] , 
        \nOut1_59[23] , \nOut1_39[27] , \nOut0_42[27] , \nOut1_56[7] , 
        \nOut0_61[16] , \nScanOut88[10] , \nScanOut107[9] , \nOut1_3[2] , 
        \nOut0_10[6] , \nScanOut25[23] , \nScanOut73[22] , \nScanOut30[17] , 
        \nScanOut50[13] , \nScanOut45[27] , \nOut0_13[5] , \nScanOut13[26] , 
        \nOut1_31[0] , \nOut0_14[15] , \nOut0_37[24] , \nOut1_39[14] , 
        \nScanOut66[16] , \nOut0_42[14] , \nScanOut119[5] , \nOut0_61[25] , 
        \nScanOut88[23] , \nOut0_57[20] , \nOut0_22[10] , \nOut1_32[3] , 
        \nOut1_59[10] , \nScanOut18[6] , \nScanOut64[0] , \nOut1_11[30] , 
        \nOut1_11[29] , \nOut1_32[18] , \nOut1_47[28] , \nOut0_49[18] , 
        \nOut1_47[31] , \nOut1_50[9] , \nScanOut67[3] , \nScanOut104[30] , 
        \nScanOut127[18] , \nScanOut104[29] , \nScanOut101[7] , 
        \nScanOut18[19] , \nOut0_8[6] , \nOut0_16[8] , \nOut1_29[2] , 
        \nScanOut96[31] , \nScanOut96[28] , \nScanOut102[4] , \nScanOut27[1] , 
        \nOut1_4[10] , \nScanOut69[18] , \nScanOut92[19] , \nScanOut126[2] , 
        \nOut1_13[8] , \nScanOut24[2] , \nScanOut125[1] , \nOut1_15[18] , 
        \nOut1_36[30] , \nOut1_36[29] , \nOut0_38[19] , \nOut1_43[19] , 
        \nOut1_60[31] , \nScanOut91[3] , \nOut0_48[6] , \nOut1_60[28] , 
        \nScanOut43[5] , \nScanOut100[18] , \nScanOut123[29] , 
        \nScanOut123[30] , \nOut0_55[9] , \nOut0_0[25] , \nOut0_0[16] , 
        \nOut1_0[31] , \nOut1_4[23] , \nScanOut40[6] , \nScanOut92[0] , 
        \nOut1_6[6] , \nOut0_10[24] , \nOut1_16[5] , \nOut0_33[15] , 
        \nOut1_48[15] , \nOut0_37[3] , \nOut0_46[25] , \nOut0_10[17] , 
        \nOut1_15[6] , \nOut0_26[21] , \nScanOut99[26] , \nScanOut128[25] , 
        \nOut1_28[11] , \nOut0_53[11] , \nScanOut54[22] , \nScanOut77[13] , 
        \nScanOut17[17] , \nScanOut21[12] , \nOut0_34[0] , \nScanOut34[26] , 
        \nScanOut41[16] , \nScanOut62[27] , \nOut0_26[12] , \nOut1_28[22] , 
        \nOut0_53[22] , \nScanOut58[4] , \nScanOut99[15] , \nScanOut128[16] , 
        \nOut0_53[7] , \nOut0_33[26] , \nOut0_46[16] , \nOut1_48[26] , 
        \nScanOut17[24] , \nScanOut34[15] , \nScanOut89[1] , \nScanOut41[25] , 
        \nScanOut46[8] , \nOut0_50[4] , \nScanOut21[21] , \nScanOut62[14] , 
        \nScanOut77[20] , \nScanOut54[11] , \nScanOut78[14] , \nOut1_0[28] , 
        \nOut1_0[8] , \nOut1_5[5] , \nScanOut5[16] , \nOut0_15[2] , 
        \nOut0_16[1] , \nScanOut18[10] , \nOut1_37[7] , \nOut1_32[22] , 
        \nOut1_34[4] , \nOut1_47[12] , \nScanOut111[27] , \nOut0_49[22] , 
        \nScanOut5[25] , \nOut1_11[20] , \nOut1_11[13] , \nScanOut18[23] , 
        \nOut1_27[16] , \nOut0_29[26] , \nScanOut83[15] , \nScanOut96[21] , 
        \nScanOut127[22] , \nOut1_52[26] , \nScanOut104[13] , \nOut1_53[3] , 
        \nScanOut64[9] , \nScanOut79[6] , \nOut1_27[25] , \nScanOut78[27] , 
        \nScanOut96[12] , \nScanOut127[11] , \nOut0_29[15] , \nOut1_32[11] , 
        \nOut1_52[15] , \nScanOut104[20] , \nOut1_47[21] , \nOut0_49[11] , 
        \nScanOut111[14] , \nScanOut83[26] , \nOut1_50[0] , \nOut0_4[27] , 
        \nOut0_4[14] , \nOut0_22[19] , \nOut1_31[9] , \nScanOut107[0] , 
        \nOut0_57[30] , \nOut0_57[29] , \nOut1_59[19] , \nScanOut25[19] , 
        \nScanOut50[30] , \nScanOut73[18] , \nScanOut104[3] , \nScanOut50[29] , 
        \nScanOut62[7] , \nOut1_48[2] , \nScanOut61[4] , \nScanOut88[19] , 
        \nScanOut21[31] , \nScanOut45[2] , \nScanOut97[4] , \nScanOut21[28] , 
        \nScanOut77[29] , \nScanOut21[6] , \nOut0_26[31] , \nScanOut46[1] , 
        \nScanOut54[18] , \nScanOut77[30] , \nScanOut89[8] , \nScanOut94[7] , 
        \nOut0_26[28] , \nOut1_28[18] , \nOut0_53[18] , \nScanOut1[14] , 
        \nScanOut22[5] , \nOut0_29[6] , \nScanOut120[5] , \nScanOut123[6] , 
        \nOut1_23[14] , \nOut0_34[9] , \nOut1_56[24] , \nScanOut92[23] , 
        \nScanOut123[20] , \nScanOut100[11] , \nOut0_58[14] , \nOut1_36[20] , 
        \nOut0_38[10] , \nOut1_43[10] , \nScanOut115[25] , \nOut1_15[11] , 
        \nOut1_60[21] , \nOut0_55[0] , \nScanOut87[17] , \nScanOut1[27] , 
        \nScanOut8[2] , \nOut1_10[2] , \nScanOut27[8] , \nOut0_56[3] , 
        \nScanOut69[22] , \nScanOut92[9] , \nOut1_15[22] , \nOut0_31[4] , 
        \nOut1_36[13] , \nOut0_38[23] , \nOut1_43[23] , \nScanOut115[16] , 
        \nScanOut87[24] , \nOut1_23[27] , \nOut0_58[27] , \nOut1_60[12] , 
        \nScanOut92[10] , \nScanOut123[13] , \nOut1_56[17] , \nScanOut100[22] , 
        \nOut0_0[31] , \nOut0_0[7] , \nOut1_4[19] , \nScanOut39[4] , 
        \nScanOut125[8] , \nOut1_13[1] , \nScanOut69[11] , \nScanOut16[14] , 
        \nOut0_32[7] , \nScanOut63[24] , \nScanOut20[11] , \nOut0_24[3] , 
        \nScanOut35[25] , \nScanOut40[15] , \nScanOut55[21] , \nScanOut76[10] , 
        \nOut1_1[22] , \nOut1_1[11] , \nOut0_3[4] , \nScanOut3[9] , 
        \nOut0_11[27] , \nOut0_27[22] , \nOut1_29[12] , \nOut0_52[12] , 
        \nScanOut98[25] , \nOut0_27[0] , \nOut0_32[16] , \nOut1_49[16] , 
        \nOut0_47[26] , \nOut1_5[20] , \nOut1_5[13] , \nOut0_6[9] , 
        \nOut0_11[14] , \nScanOut16[27] , \nScanOut20[22] , \nScanOut55[12] , 
        \nScanOut76[23] , \nScanOut35[16] , \nScanOut63[17] , \nScanOut99[2] , 
        \nOut0_40[7] , \nScanOut40[26] , \nOut1_61[1] , \nOut0_27[11] , 
        \nOut1_29[21] , \nOut0_32[25] , \nOut0_47[15] , \nOut1_49[25] , 
        \nOut0_52[21] , \nScanOut55[8] , \nOut0_43[4] , \nScanOut34[1] , 
        \nScanOut48[7] , \nOut1_62[2] , \nScanOut98[16] , \nOut1_14[31] , 
        \nOut1_14[28] , \nOut0_39[30] , \nOut1_42[30] , \nOut1_61[18] , 
        \nOut1_37[19] , \nScanOut37[2] , \nOut0_39[29] , \nOut1_42[29] , 
        \nScanOut101[31] , \nScanOut101[28] , \nScanOut122[19] , 
        \nScanOut68[28] , \nScanOut5[7] , \nScanOut68[31] , \nScanOut6[4] , 
        \nOut0_46[9] , \nScanOut50[5] , \nScanOut82[3] , \nScanOut53[6] , 
        \nScanOut93[30] , \nScanOut19[29] , \nOut0_58[5] , \nScanOut81[0] , 
        \nScanOut93[29] , \nScanOut77[0] , \nScanOut97[18] , \nOut1_8[0] , 
        \nOut1_10[19] , \nScanOut19[30] , \nOut1_33[31] , \nOut1_43[9] , 
        \nScanOut74[3] , \nOut0_18[7] , \nOut1_33[28] , \nOut1_46[18] , 
        \nOut0_48[31] , \nOut1_39[1] , \nOut0_48[28] , \nScanOut105[19] , 
        \nScanOut112[7] , \nScanOut126[31] , \nScanOut126[28] , 
        \nScanOut10[7] , \nScanOut13[4] , \nScanOut12[25] , \nScanOut12[16] , 
        \nOut0_15[25] , \nScanOut111[4] , \nOut0_23[20] , \nOut0_36[14] , 
        \nOut0_60[15] , \nScanOut89[13] , \nOut1_38[24] , \nOut0_43[24] , 
        \nOut1_46[4] , \nScanOut24[13] , \nOut1_45[7] , \nScanOut51[23] , 
        \nOut0_56[10] , \nOut1_58[20] , \nOut1_58[8] , \nScanOut67[26] , 
        \nScanOut72[12] , \nOut0_15[16] , \nOut1_22[0] , \nScanOut31[27] , 
        \nScanOut44[17] , \nOut0_56[23] , \nScanOut114[9] , \nOut0_23[13] , 
        \nOut1_58[13] , \nOut0_60[26] , \nScanOut89[20] , \nOut0_36[27] , 
        \nOut1_38[17] , \nOut0_43[17] , \nScanOut109[6] , \nOut1_15[2] , 
        \nScanOut16[9] , \nScanOut31[14] , \nScanOut67[15] , \nScanOut17[13] , 
        \nOut1_21[3] , \nScanOut44[24] , \nScanOut24[20] , \nScanOut51[10] , 
        \nScanOut62[23] , \nScanOut72[21] , \nScanOut22[8] , \nScanOut34[22] , 
        \nScanOut41[12] , \nScanOut54[26] , \nScanOut21[16] , \nOut0_34[4] , 
        \nScanOut77[17] , \nOut0_0[28] , \nScanOut120[8] , \nOut1_4[14] , 
        \nOut0_10[20] , \nOut0_26[25] , \nOut1_28[15] , \nOut0_53[15] , 
        \nScanOut99[22] , \nScanOut128[21] , \nOut0_10[13] , \nOut1_16[1] , 
        \nOut0_33[11] , \nOut1_48[11] , \nOut0_46[21] , \nScanOut17[20] , 
        \nScanOut21[25] , \nOut0_37[7] , \nScanOut54[15] , \nScanOut77[24] , 
        \nScanOut34[11] , \nScanOut62[10] , \nScanOut89[5] , \nScanOut41[21] , 
        \nOut0_50[0] , \nScanOut24[6] , \nOut0_26[16] , \nOut1_28[26] , 
        \nOut0_33[22] , \nOut0_46[12] , \nOut1_48[22] , \nOut0_53[26] , 
        \nOut0_53[3] , \nScanOut58[0] , \nScanOut99[11] , \nScanOut128[12] , 
        \nScanOut97[9] , \nScanOut125[5] , \nScanOut39[9] , \nScanOut87[30] , 
        \nScanOut87[29] , \nScanOut126[6] , \nOut1_4[27] , \nOut0_8[2] , 
        \nScanOut27[5] , \nOut0_31[9] , \nScanOut40[2] , \nScanOut92[4] , 
        \nOut1_0[25] , \nOut1_0[16] , \nScanOut1[19] , \nOut1_23[19] , 
        \nScanOut43[1] , \nOut1_56[29] , \nOut0_58[19] , \nOut1_56[30] , 
        \nScanOut5[31] , \nScanOut5[28] , \nOut1_27[31] , \nOut1_27[28] , 
        \nOut0_48[2] , \nScanOut91[7] , \nScanOut115[31] , \nScanOut115[28] , 
        \nScanOut67[7] , \nOut0_29[18] , \nOut1_52[18] , \nScanOut111[19] , 
        \nOut1_5[8] , \nScanOut64[4] , \nOut1_29[6] , \nScanOut83[18] , 
        \nOut1_34[9] , \nScanOut102[0] , \nScanOut78[19] , \nOut1_0[5] , 
        \nOut1_3[6] , \nScanOut13[11] , \nOut0_14[22] , \nScanOut101[3] , 
        \nOut0_22[27] , \nOut0_37[13] , \nOut0_61[12] , \nScanOut61[9] , 
        \nScanOut88[14] , \nOut1_39[23] , \nOut0_42[23] , \nOut1_56[3] , 
        \nScanOut25[14] , \nScanOut50[24] , \nOut0_57[17] , \nOut1_59[27] , 
        \nOut1_55[0] , \nScanOut66[21] , \nScanOut73[15] , \nScanOut18[2] , 
        \nScanOut30[20] , \nScanOut45[10] , \nOut0_4[19] , \nOut0_10[2] , 
        \nOut0_13[1] , \nOut0_57[24] , \nScanOut13[22] , \nOut0_14[11] , 
        \nOut0_22[14] , \nOut1_32[7] , \nOut1_59[14] , \nOut0_61[21] , 
        \nScanOut88[27] , \nOut0_37[20] , \nOut1_39[10] , \nOut0_42[10] , 
        \nScanOut119[1] , \nScanOut30[13] , \nScanOut66[12] , \nScanOut45[23] , 
        \nScanOut25[27] , \nOut1_31[4] , \nScanOut50[17] , \nScanOut73[26] , 
        \nScanOut4[11] , \nScanOut13[9] , \nScanOut19[17] , \nScanOut79[13] , 
        \nScanOut111[9] , \nOut1_27[0] , \nOut1_24[3] , \nOut1_33[25] , 
        \nOut1_46[15] , \nScanOut110[20] , \nOut0_48[25] , \nOut1_10[14] , 
        \nScanOut19[24] , \nOut1_26[11] , \nOut0_28[21] , \nScanOut82[12] , 
        \nScanOut97[26] , \nScanOut126[25] , \nOut1_53[21] , \nScanOut105[14] , 
        \nOut1_43[4] , \nOut0_62[2] , \nScanOut69[1] , \nScanOut79[20] , 
        \nScanOut97[15] , \nOut0_0[3] , \nOut0_1[22] , \nOut0_1[11] , 
        \nScanOut0[7] , \nScanOut4[22] , \nOut1_10[27] , \nOut1_26[22] , 
        \nScanOut126[16] , \nOut0_28[12] , \nOut1_33[16] , \nOut1_53[12] , 
        \nScanOut105[27] , \nOut1_46[26] , \nOut0_48[16] , \nScanOut110[13] , 
        \nScanOut82[21] , \nOut0_5[20] , \nOut0_5[13] , \nScanOut12[31] , 
        \nScanOut31[19] , \nOut1_40[7] , \nOut0_61[1] , \nScanOut117[7] , 
        \nScanOut12[28] , \nScanOut16[4] , \nScanOut44[29] , \nScanOut15[7] , 
        \nScanOut44[30] , \nScanOut67[18] , \nOut1_58[5] , \nScanOut72[0] , 
        \nScanOut114[4] , \nOut0_15[31] , \nOut0_36[19] , \nOut0_15[28] , 
        \nOut1_38[29] , \nScanOut71[3] , \nOut0_43[29] , \nOut1_46[9] , 
        \nOut1_38[30] , \nOut0_43[30] , \nOut0_60[18] , \nScanOut3[4] , 
        \nOut0_11[19] , \nOut0_32[28] , \nOut0_47[18] , \nScanOut87[3] , 
        \nOut1_49[28] , \nOut1_49[31] , \nOut0_32[31] , \nOut0_43[9] , 
        \nScanOut55[5] , \nScanOut56[6] , \nScanOut31[1] , \nScanOut84[0] , 
        \nScanOut98[31] , \nScanOut98[28] , \nOut1_1[26] , \nOut1_1[15] , 
        \nScanOut0[20] , \nScanOut0[13] , \nOut0_3[9] , \nScanOut6[9] , 
        \nScanOut16[19] , \nOut1_18[7] , \nScanOut35[28] , \nOut0_39[1] , 
        \nScanOut40[18] , \nScanOut63[30] , \nScanOut63[29] , \nScanOut32[2] , 
        \nScanOut35[31] , \nOut1_57[23] , \nScanOut93[24] , \nScanOut122[27] , 
        \nScanOut101[16] , \nOut0_59[13] , \nOut1_22[13] , \nOut1_37[27] , 
        \nOut0_39[17] , \nOut1_42[17] , \nOut0_58[8] , \nScanOut114[22] , 
        \nOut1_61[26] , \nOut1_14[25] , \nOut1_14[16] , \nOut0_21[3] , 
        \nOut0_45[7] , \nScanOut86[10] , \nOut0_46[4] , \nScanOut50[8] , 
        \nScanOut68[25] , \nOut1_37[14] , \nOut0_39[24] , \nOut1_42[24] , 
        \nScanOut114[11] , \nOut1_61[15] , \nScanOut86[23] , \nOut0_5[30] , 
        \nOut0_5[29] , \nOut0_5[7] , \nScanOut93[17] , \nScanOut122[14] , 
        \nOut0_6[4] , \nOut1_22[20] , \nOut0_59[20] , \nScanOut29[3] , 
        \nOut1_57[10] , \nScanOut101[25] , \nScanOut68[16] , \nScanOut12[12] , 
        \nOut0_22[0] , \nScanOut128[0] , \nScanOut31[23] , \nScanOut44[13] , 
        \nScanOut67[22] , \nScanOut24[17] , \nOut1_45[3] , \nScanOut51[27] , 
        \nScanOut72[16] , \nScanOut72[9] , \nScanOut12[21] , \nOut0_15[21] , 
        \nOut0_23[24] , \nOut0_36[10] , \nOut0_56[14] , \nOut1_58[24] , 
        \nOut1_38[20] , \nOut0_43[20] , \nOut1_46[0] , \nOut1_21[7] , 
        \nScanOut24[24] , \nOut0_60[11] , \nScanOut72[25] , \nScanOut89[17] , 
        \nScanOut31[10] , \nScanOut51[14] , \nScanOut44[20] , \nOut0_15[12] , 
        \nOut0_36[23] , \nOut1_38[13] , \nScanOut67[11] , \nOut0_43[13] , 
        \nScanOut109[2] , \nOut0_60[22] , \nScanOut89[24] , \nOut1_22[4] , 
        \nOut0_23[17] , \nOut0_56[27] , \nOut1_58[17] , \nScanOut69[8] , 
        \nScanOut74[7] , \nScanOut79[30] , \nScanOut79[29] , \nOut0_61[8] , 
        \nScanOut77[4] , \nScanOut82[31] , \nScanOut82[28] , \nScanOut111[0] , 
        \nScanOut0[30] , \nScanOut4[18] , \nOut1_8[4] , \nScanOut10[3] , 
        \nScanOut13[0] , \nOut1_27[9] , \nOut0_18[3] , \nOut1_26[18] , 
        \nOut0_28[31] , \nOut0_28[28] , \nOut1_53[31] , \nOut1_53[28] , 
        \nScanOut112[3] , \nScanOut110[29] , \nOut1_39[5] , \nOut1_22[30] , 
        \nScanOut37[6] , \nScanOut110[30] , \nOut0_59[30] , \nOut1_22[29] , 
        \nOut0_59[29] , \nOut1_57[19] , \nScanOut0[29] , \nScanOut114[18] , 
        \nOut0_3[0] , \nOut1_5[24] , \nOut1_5[17] , \nScanOut5[3] , 
        \nScanOut6[0] , \nOut0_22[9] , \nScanOut34[5] , \nOut0_58[1] , 
        \nScanOut81[4] , \nScanOut128[9] , \nScanOut86[19] , \nScanOut50[1] , 
        \nScanOut53[2] , \nScanOut82[7] , \nOut0_11[23] , \nOut0_27[4] , 
        \nScanOut31[8] , \nOut1_49[12] , \nOut0_32[12] , \nOut0_47[22] , 
        \nOut0_27[26] , \nScanOut98[21] , \nOut1_29[16] , \nOut0_52[16] , 
        \nOut0_1[18] , \nScanOut16[10] , \nScanOut20[15] , \nOut0_24[7] , 
        \nOut0_39[8] , \nScanOut55[25] , \nScanOut76[14] , \nScanOut35[21] , 
        \nScanOut40[11] , \nScanOut63[20] , \nScanOut1[10] , \nScanOut8[6] , 
        \nOut0_11[10] , \nOut0_27[15] , \nOut1_29[25] , \nScanOut48[3] , 
        \nOut0_52[25] , \nScanOut98[12] , \nOut0_43[0] , \nOut1_62[6] , 
        \nOut0_32[21] , \nOut0_47[11] , \nOut1_49[21] , \nScanOut16[23] , 
        \nScanOut35[12] , \nScanOut99[6] , \nOut0_40[3] , \nScanOut40[22] , 
        \nOut1_61[5] , \nScanOut20[26] , \nScanOut63[13] , \nScanOut76[27] , 
        \nScanOut55[16] , \nOut0_56[7] , \nScanOut69[26] , \nScanOut84[9] , 
        \nScanOut43[8] , \nOut0_55[4] , \nOut1_60[25] , \nOut1_13[5] , 
        \nOut1_15[15] , \nOut1_23[10] , \nOut1_36[24] , \nOut0_38[14] , 
        \nOut1_43[14] , \nScanOut87[13] , \nScanOut115[21] , \nOut1_56[20] , 
        \nScanOut100[15] , \nOut0_58[10] , \nScanOut92[27] , \nScanOut123[24] , 
        \nOut0_32[3] , \nScanOut39[0] , \nScanOut69[15] , \nOut0_0[21] , 
        \nOut0_0[12] , \nScanOut1[23] , \nOut1_15[26] , \nOut1_23[23] , 
        \nOut0_58[23] , \nOut1_56[13] , \nScanOut100[26] , \nScanOut92[14] , 
        \nScanOut123[17] , \nOut1_60[16] , \nScanOut87[20] , \nOut1_10[6] , 
        \nOut1_36[17] , \nOut0_38[27] , \nOut1_43[27] , \nScanOut115[12] , 
        \nScanOut17[30] , \nScanOut17[29] , \nOut0_31[0] , \nScanOut94[3] , 
        \nScanOut34[18] , \nScanOut41[31] , \nScanOut62[19] , \nScanOut41[28] , 
        \nScanOut46[5] , \nScanOut45[6] , \nOut0_50[9] , \nScanOut58[9] , 
        \nScanOut99[18] , \nScanOut97[0] , \nScanOut22[1] , \nOut0_29[2] , 
        \nScanOut120[1] , \nScanOut123[2] , \nOut0_4[10] , \nOut0_10[30] , 
        \nOut0_10[29] , \nScanOut21[2] , \nOut0_33[18] , \nOut0_46[31] , 
        \nOut1_48[18] , \nOut1_16[8] , \nOut0_46[28] , \nScanOut104[7] , 
        \nScanOut128[31] , \nScanOut128[28] , \nOut0_14[18] , \nOut0_61[28] , 
        \nOut0_37[30] , \nOut1_39[19] , \nScanOut1[21] , \nScanOut1[12] , 
        \nOut0_4[23] , \nOut0_13[8] , \nOut0_37[29] , \nOut0_42[19] , 
        \nOut0_61[31] , \nScanOut119[8] , \nScanOut61[0] , \nScanOut107[4] , 
        \nOut1_5[1] , \nScanOut5[12] , \nScanOut13[18] , \nOut1_48[6] , 
        \nScanOut66[28] , \nOut1_27[12] , \nOut0_29[22] , \nScanOut30[30] , 
        \nScanOut30[29] , \nScanOut45[19] , \nScanOut66[31] , \nOut1_55[9] , 
        \nScanOut62[3] , \nOut1_52[22] , \nScanOut104[17] , \nScanOut102[9] , 
        \nScanOut96[25] , \nScanOut127[26] , \nScanOut5[21] , \nOut1_6[2] , 
        \nOut1_11[17] , \nOut0_15[6] , \nOut1_32[26] , \nOut1_47[16] , 
        \nScanOut83[11] , \nScanOut111[23] , \nOut0_49[26] , \nOut0_16[5] , 
        \nOut1_34[0] , \nScanOut18[14] , \nOut1_37[3] , \nScanOut78[10] , 
        \nOut1_11[24] , \nOut1_50[4] , \nScanOut83[22] , \nOut1_15[17] , 
        \nScanOut18[27] , \nOut1_27[21] , \nOut1_32[15] , \nOut1_47[25] , 
        \nOut0_49[15] , \nScanOut111[10] , \nOut0_29[11] , \nOut1_52[11] , 
        \nScanOut104[24] , \nScanOut78[23] , \nScanOut96[16] , 
        \nScanOut127[15] , \nOut1_23[12] , \nOut1_53[7] , \nScanOut79[2] , 
        \nOut0_58[12] , \nOut1_56[22] , \nScanOut100[17] , \nScanOut92[25] , 
        \nScanOut123[26] , \nScanOut87[11] , \nOut0_8[9] , \nScanOut8[4] , 
        \nOut1_36[26] , \nOut0_48[9] , \nOut1_60[27] , \nOut0_38[16] , 
        \nOut1_43[16] , \nScanOut115[23] , \nOut0_55[6] , \nOut1_10[4] , 
        \nOut0_31[2] , \nScanOut40[9] , \nOut0_56[5] , \nScanOut69[24] , 
        \nOut1_15[24] , \nOut1_60[14] , \nOut1_23[21] , \nOut1_36[15] , 
        \nOut0_38[25] , \nOut1_43[25] , \nScanOut87[22] , \nScanOut115[10] , 
        \nOut1_56[11] , \nScanOut100[24] , \nOut0_58[21] , \nScanOut92[16] , 
        \nScanOut123[15] , \nOut0_0[23] , \nOut0_0[10] , \nOut1_13[7] , 
        \nOut0_32[1] , \nScanOut39[2] , \nScanOut69[17] , \nScanOut97[2] , 
        \nOut0_10[18] , \nOut0_33[30] , \nOut1_48[30] , \nScanOut21[0] , 
        \nOut0_33[29] , \nOut1_48[29] , \nScanOut45[4] , \nOut0_46[19] , 
        \nOut0_53[8] , \nScanOut46[7] , \nScanOut128[19] , \nScanOut94[1] , 
        \nScanOut99[30] , \nScanOut99[29] , \nScanOut120[3] , \nOut0_4[21] , 
        \nOut0_4[12] , \nOut0_10[9] , \nScanOut13[29] , \nOut1_15[9] , 
        \nScanOut17[18] , \nOut0_29[0] , \nScanOut123[0] , \nScanOut34[30] , 
        \nScanOut34[29] , \nScanOut62[28] , \nScanOut41[19] , \nScanOut62[31] , 
        \nScanOut22[3] , \nScanOut45[31] , \nScanOut107[6] , \nScanOut66[19] , 
        \nScanOut45[28] , \nScanOut13[30] , \nScanOut18[9] , \nScanOut30[18] , 
        \nOut1_48[4] , \nScanOut62[1] , \nScanOut104[5] , \nOut0_5[18] , 
        \nOut1_5[3] , \nOut1_6[0] , \nOut0_14[30] , \nOut0_14[29] , 
        \nOut1_39[31] , \nOut0_42[31] , \nOut0_61[19] , \nOut1_39[28] , 
        \nOut0_42[28] , \nOut1_56[8] , \nScanOut61[2] , \nOut0_37[18] , 
        \nOut1_11[15] , \nOut0_15[4] , \nOut0_16[7] , \nScanOut18[16] , 
        \nScanOut78[12] , \nOut1_37[1] , \nScanOut101[8] , \nOut1_34[2] , 
        \nScanOut83[13] , \nScanOut5[23] , \nScanOut5[10] , \nScanOut18[25] , 
        \nOut1_27[10] , \nOut1_32[24] , \nOut1_47[14] , \nOut0_49[24] , 
        \nScanOut111[21] , \nOut0_29[20] , \nScanOut104[15] , \nOut1_52[20] , 
        \nOut1_53[5] , \nScanOut96[27] , \nScanOut127[24] , \nOut1_27[23] , 
        \nOut0_29[13] , \nScanOut78[21] , \nScanOut79[0] , \nScanOut104[26] , 
        \nOut1_52[13] , \nScanOut96[14] , \nScanOut127[17] , \nOut1_11[26] , 
        \nScanOut12[10] , \nOut0_15[23] , \nOut1_32[17] , \nOut1_47[27] , 
        \nScanOut83[20] , \nScanOut111[12] , \nOut0_36[12] , \nOut1_38[22] , 
        \nOut0_49[17] , \nOut1_50[6] , \nOut0_43[22] , \nOut1_46[2] , 
        \nOut0_60[13] , \nScanOut71[8] , \nScanOut89[15] , \nOut0_23[26] , 
        \nOut0_56[16] , \nScanOut24[15] , \nOut1_45[1] , \nOut1_58[26] , 
        \nScanOut72[14] , \nScanOut31[21] , \nScanOut51[25] , \nScanOut44[11] , 
        \nScanOut67[20] , \nScanOut12[23] , \nOut0_15[10] , \nOut1_22[6] , 
        \nOut0_23[15] , \nOut0_36[21] , \nOut0_56[25] , \nOut1_58[15] , 
        \nScanOut109[0] , \nOut1_38[11] , \nOut0_43[11] , \nOut1_21[5] , 
        \nScanOut44[22] , \nOut0_60[20] , \nScanOut89[26] , \nScanOut31[12] , 
        \nScanOut67[13] , \nScanOut24[26] , \nScanOut51[16] , \nScanOut72[27] , 
        \nScanOut77[6] , \nOut0_0[1] , \nOut1_1[24] , \nOut1_1[17] , 
        \nScanOut4[30] , \nOut1_26[30] , \nOut1_26[29] , \nOut0_28[19] , 
        \nOut1_53[19] , \nScanOut4[29] , \nScanOut110[18] , \nOut1_8[6] , 
        \nScanOut13[2] , \nOut0_18[1] , \nOut1_39[7] , \nOut0_62[9] , 
        \nScanOut74[5] , \nOut1_24[8] , \nScanOut82[19] , \nScanOut112[1] , 
        \nScanOut10[1] , \nScanOut79[18] , \nScanOut111[2] , \nScanOut0[18] , 
        \nOut1_5[26] , \nOut1_5[15] , \nScanOut29[8] , \nScanOut34[7] , 
        \nScanOut5[1] , \nOut0_21[8] , \nScanOut86[31] , \nScanOut86[28] , 
        \nScanOut37[4] , \nScanOut6[2] , \nScanOut50[3] , \nScanOut82[5] , 
        \nScanOut53[0] , \nOut1_57[31] , \nOut0_59[18] , \nOut1_22[18] , 
        \nOut1_57[28] , \nOut0_58[3] , \nScanOut81[6] , \nScanOut114[29] , 
        \nScanOut16[12] , \nScanOut35[23] , \nScanOut114[30] , 
        \nScanOut40[13] , \nScanOut20[17] , \nOut0_24[5] , \nScanOut63[22] , 
        \nScanOut76[16] , \nScanOut32[9] , \nScanOut55[27] , \nOut0_1[30] , 
        \nOut0_1[29] , \nOut0_3[2] , \nScanOut4[20] , \nScanOut4[13] , 
        \nOut1_10[16] , \nOut0_11[21] , \nOut0_27[24] , \nOut1_29[14] , 
        \nOut0_52[14] , \nScanOut98[23] , \nOut0_27[6] , \nOut0_32[10] , 
        \nOut0_47[20] , \nOut1_49[10] , \nOut0_11[12] , \nScanOut16[21] , 
        \nScanOut20[24] , \nScanOut55[14] , \nScanOut76[25] , \nScanOut35[10] , 
        \nOut0_40[1] , \nScanOut40[20] , \nOut1_61[7] , \nScanOut63[11] , 
        \nScanOut99[4] , \nOut0_32[23] , \nOut1_49[23] , \nOut0_47[13] , 
        \nOut0_18[8] , \nOut1_26[13] , \nOut0_27[17] , \nScanOut98[10] , 
        \nOut1_29[27] , \nOut0_43[2] , \nOut1_62[4] , \nOut0_52[27] , 
        \nScanOut48[1] , \nScanOut87[8] , \nScanOut97[24] , \nScanOut112[8] , 
        \nScanOut126[27] , \nOut0_28[23] , \nScanOut105[16] , \nOut1_33[27] , 
        \nOut1_53[23] , \nOut1_46[17] , \nOut0_48[27] , \nScanOut110[22] , 
        \nScanOut82[10] , \nScanOut10[8] , \nOut1_24[1] , \nOut1_27[2] , 
        \nScanOut19[15] , \nOut1_33[14] , \nOut1_40[5] , \nOut0_61[3] , 
        \nScanOut79[11] , \nOut1_46[24] , \nScanOut110[11] , \nOut0_48[14] , 
        \nOut1_10[25] , \nScanOut82[23] , \nScanOut126[14] , \nOut0_5[11] , 
        \nScanOut19[26] , \nOut1_26[20] , \nOut0_28[10] , \nScanOut97[17] , 
        \nScanOut105[25] , \nOut1_53[10] , \nScanOut69[3] , \nScanOut79[22] , 
        \nOut1_43[6] , \nOut0_62[0] , \nScanOut114[6] , \nOut0_15[19] , 
        \nOut0_36[31] , \nOut0_36[28] , \nScanOut109[9] , \nOut1_38[18] , 
        \nOut0_43[18] , \nOut0_60[30] , \nScanOut15[5] , \nOut0_60[29] , 
        \nScanOut16[6] , \nScanOut117[5] , \nOut0_0[19] , \nOut0_0[8] , 
        \nOut0_1[13] , \nScanOut3[6] , \nOut0_5[22] , \nScanOut71[1] , 
        \nScanOut12[19] , \nScanOut31[31] , \nScanOut31[28] , \nOut1_58[7] , 
        \nScanOut44[18] , \nScanOut67[30] , \nOut1_45[8] , \nScanOut67[29] , 
        \nScanOut72[2] , \nScanOut84[2] , \nScanOut16[31] , \nOut0_40[8] , 
        \nScanOut40[29] , \nScanOut16[28] , \nScanOut35[19] , \nScanOut40[30] , 
        \nScanOut56[4] , \nScanOut63[18] , \nScanOut55[7] , \nScanOut98[19] , 
        \nScanOut0[5] , \nScanOut48[8] , \nScanOut87[1] , \nScanOut32[0] , 
        \nOut0_1[20] , \nOut1_18[5] , \nOut0_39[3] , \nScanOut0[22] , 
        \nScanOut0[11] , \nScanOut5[8] , \nOut0_11[31] , \nOut0_47[29] , 
        \nOut1_49[19] , \nOut0_11[28] , \nScanOut31[3] , \nOut0_32[19] , 
        \nOut0_47[30] , \nOut1_14[14] , \nOut1_37[25] , \nOut0_45[5] , 
        \nOut0_46[6] , \nScanOut68[27] , \nScanOut53[9] , \nOut0_39[15] , 
        \nOut1_42[15] , \nScanOut114[20] , \nScanOut86[12] , \nOut0_5[5] , 
        \nOut0_6[6] , \nOut0_22[2] , \nOut1_22[11] , \nOut0_59[11] , 
        \nOut1_61[24] , \nScanOut93[26] , \nScanOut122[25] , \nOut1_57[21] , 
        \nScanOut101[14] , \nScanOut29[1] , \nScanOut128[2] , \nScanOut68[14] , 
        \nScanOut122[16] , \nOut1_22[22] , \nOut1_57[12] , \nScanOut93[15] , 
        \nScanOut101[27] , \nOut0_59[22] , \nOut1_37[16] , \nOut0_39[26] , 
        \nOut1_42[26] , \nScanOut114[13] , \nOut0_10[22] , \nOut1_14[27] , 
        \nOut1_61[17] , \nOut0_21[1] , \nScanOut86[21] , \nOut1_15[0] , 
        \nOut1_16[3] , \nOut0_37[5] , \nScanOut21[9] , \nOut0_33[13] , 
        \nOut0_46[23] , \nOut1_48[13] , \nOut0_26[27] , \nOut1_28[17] , 
        \nOut0_53[17] , \nOut0_29[9] , \nScanOut99[20] , \nScanOut128[23] , 
        \nOut0_34[6] , \nScanOut123[9] , \nScanOut17[11] , \nScanOut21[14] , 
        \nScanOut54[24] , \nScanOut77[15] , \nScanOut34[20] , \nScanOut62[21] , 
        \nScanOut41[10] , \nScanOut58[2] , \nOut0_8[0] , \nOut0_10[11] , 
        \nOut0_26[14] , \nOut1_28[24] , \nOut0_53[24] , \nOut0_53[1] , 
        \nScanOut99[13] , \nScanOut128[10] , \nScanOut17[22] , \nOut0_33[20] , 
        \nOut1_48[20] , \nOut0_46[10] , \nScanOut62[12] , \nScanOut21[27] , 
        \nScanOut34[13] , \nScanOut41[23] , \nOut0_50[2] , \nScanOut54[17] , 
        \nScanOut89[7] , \nScanOut27[7] , \nScanOut77[26] , \nScanOut94[8] , 
        \nScanOut1[31] , \nScanOut1[28] , \nOut1_23[31] , \nOut1_23[28] , 
        \nOut1_56[18] , \nOut0_58[28] , \nOut0_58[31] , \nOut1_4[16] , 
        \nScanOut115[19] , \nScanOut126[4] , \nScanOut24[4] , \nOut0_32[8] , 
        \nScanOut125[7] , \nOut0_48[0] , \nScanOut87[18] , \nScanOut91[5] , 
        \nOut0_0[27] , \nOut0_0[14] , \nOut0_0[5] , \nOut1_0[27] , 
        \nOut1_0[14] , \nOut1_4[25] , \nScanOut40[0] , \nScanOut43[3] , 
        \nScanOut92[6] , \nScanOut64[6] , \nScanOut78[31] , \nScanOut78[28] , 
        \nScanOut67[5] , \nScanOut79[9] , \nScanOut83[30] , \nScanOut83[29] , 
        \nOut1_0[7] , \nOut0_4[31] , \nScanOut5[19] , \nOut1_6[9] , 
        \nScanOut101[1] , \nOut1_27[19] , \nOut1_37[8] , \nScanOut102[2] , 
        \nOut0_29[30] , \nOut0_29[29] , \nOut1_52[29] , \nOut1_52[30] , 
        \nScanOut13[13] , \nOut1_29[4] , \nScanOut111[31] , \nScanOut111[28] , 
        \nScanOut25[16] , \nScanOut30[22] , \nScanOut66[23] , \nScanOut45[12] , 
        \nOut1_55[2] , \nScanOut50[26] , \nScanOut62[8] , \nScanOut73[17] , 
        \nOut0_4[28] , \nOut0_14[20] , \nOut0_22[25] , \nOut0_57[15] , 
        \nOut1_59[25] , \nOut0_61[10] , \nScanOut88[16] , \nOut0_37[11] , 
        \nOut1_39[21] , \nOut0_42[21] , \nOut1_56[1] , \nOut0_3[6] , 
        \nOut1_3[4] , \nOut0_10[0] , \nScanOut13[20] , \nScanOut25[25] , 
        \nScanOut50[15] , \nScanOut66[10] , \nScanOut73[24] , \nOut1_31[6] , 
        \nScanOut45[21] , \nOut0_13[3] , \nOut0_14[13] , \nScanOut30[11] , 
        \nOut0_22[16] , \nOut1_32[5] , \nOut0_37[22] , \nOut0_61[23] , 
        \nScanOut88[25] , \nScanOut119[3] , \nOut1_39[12] , \nOut0_42[12] , 
        \nScanOut18[0] , \nOut0_57[26] , \nOut1_59[16] , \nOut0_11[25] , 
        \nOut0_27[20] , \nOut0_27[2] , \nOut1_29[10] , \nOut0_32[14] , 
        \nOut0_47[24] , \nOut1_49[14] , \nOut0_52[10] , \nScanOut98[27] , 
        \nOut1_18[8] , \nOut1_0[19] , \nOut1_1[20] , \nOut1_1[13] , 
        \nScanOut0[8] , \nScanOut16[16] , \nScanOut20[13] , \nOut0_24[1] , 
        \nScanOut55[23] , \nScanOut76[12] , \nScanOut35[27] , \nScanOut63[26] , 
        \nScanOut40[17] , \nScanOut48[5] , \nOut0_5[8] , \nOut0_11[16] , 
        \nOut0_27[13] , \nOut1_62[0] , \nOut1_29[23] , \nOut0_43[6] , 
        \nOut0_52[23] , \nScanOut98[14] , \nScanOut16[25] , \nOut0_32[27] , 
        \nOut1_49[27] , \nOut0_47[17] , \nScanOut63[15] , \nScanOut20[20] , 
        \nScanOut35[14] , \nOut0_40[5] , \nScanOut40[24] , \nOut1_61[3] , 
        \nScanOut55[10] , \nScanOut56[9] , \nScanOut99[0] , \nScanOut37[0] , 
        \nScanOut76[21] , \nOut1_5[22] , \nOut1_5[11] , \nScanOut93[18] , 
        \nScanOut6[6] , \nOut1_14[19] , \nScanOut34[3] , \nScanOut68[19] , 
        \nOut1_37[31] , \nOut1_37[28] , \nOut0_58[7] , \nOut1_61[29] , 
        \nOut0_39[18] , \nOut1_42[18] , \nOut1_61[30] , \nScanOut81[2] , 
        \nOut0_45[8] , \nScanOut101[19] , \nScanOut122[31] , \nScanOut122[28] , 
        \nScanOut50[7] , \nScanOut53[4] , \nScanOut82[1] , \nScanOut5[5] , 
        \nScanOut74[1] , \nOut1_10[31] , \nOut1_10[28] , \nOut1_46[30] , 
        \nOut1_33[19] , \nOut1_46[29] , \nScanOut19[18] , \nOut1_40[8] , 
        \nOut0_48[19] , \nScanOut105[31] , \nScanOut105[28] , 
        \nScanOut126[19] , \nScanOut77[2] , \nOut1_5[7] , \nOut1_8[2] , 
        \nScanOut10[5] , \nScanOut111[6] , \nOut1_11[11] , \nScanOut12[27] , 
        \nScanOut12[14] , \nScanOut13[6] , \nOut0_18[5] , \nOut1_39[3] , 
        \nScanOut97[30] , \nScanOut112[5] , \nScanOut97[29] , \nOut0_15[27] , 
        \nOut0_23[22] , \nScanOut24[11] , \nScanOut31[25] , \nScanOut67[24] , 
        \nScanOut44[15] , \nOut1_45[5] , \nScanOut51[21] , \nOut0_56[12] , 
        \nScanOut72[10] , \nOut1_58[22] , \nOut0_60[17] , \nScanOut89[11] , 
        \nScanOut24[22] , \nOut0_36[16] , \nOut1_38[26] , \nOut0_43[26] , 
        \nOut1_46[6] , \nScanOut51[12] , \nScanOut117[8] , \nScanOut67[17] , 
        \nScanOut72[23] , \nOut0_15[14] , \nOut1_21[1] , \nScanOut44[26] , 
        \nScanOut31[16] , \nScanOut15[8] , \nOut1_22[2] , \nOut0_23[11] , 
        \nOut0_36[25] , \nOut0_60[24] , \nScanOut89[22] , \nScanOut109[4] , 
        \nOut1_38[15] , \nOut0_43[15] , \nOut1_58[11] , \nOut1_27[14] , 
        \nOut0_56[21] , \nScanOut96[23] , \nScanOut127[20] , \nOut0_29[24] , 
        \nScanOut104[11] , \nOut1_29[9] , \nOut1_32[20] , \nOut1_52[24] , 
        \nOut1_47[10] , \nOut0_49[20] , \nScanOut111[25] , \nScanOut83[17] , 
        \nScanOut5[27] , \nScanOut5[14] , \nOut1_6[4] , \nOut0_15[0] , 
        \nOut1_34[6] , \nOut0_16[3] , \nOut1_37[5] , \nScanOut18[12] , 
        \nOut1_32[13] , \nOut1_47[23] , \nOut1_50[2] , \nScanOut78[16] , 
        \nScanOut67[8] , \nScanOut111[16] , \nOut0_49[13] , \nOut1_11[22] , 
        \nOut1_27[27] , \nOut0_29[17] , \nScanOut83[24] , \nScanOut96[10] , 
        \nScanOut127[13] , \nScanOut104[22] , \nOut1_52[17] , \nScanOut78[25] , 
        \nScanOut79[4] , \nOut1_3[9] , \nOut0_4[16] , \nScanOut18[21] , 
        \nOut1_53[1] , \nScanOut104[1] , \nOut0_4[25] , \nOut0_22[31] , 
        \nScanOut25[31] , \nOut1_32[8] , \nScanOut88[31] , \nScanOut88[28] , 
        \nScanOut73[29] , \nScanOut25[28] , \nScanOut50[18] , \nScanOut73[30] , 
        \nScanOut107[2] , \nOut0_22[28] , \nOut0_57[18] , \nOut1_59[31] , 
        \nOut1_59[28] , \nScanOut61[6] , \nOut0_26[19] , \nOut1_28[30] , 
        \nScanOut46[3] , \nOut1_48[0] , \nScanOut62[5] , \nScanOut94[5] , 
        \nOut0_53[30] , \nOut1_28[29] , \nScanOut45[0] , \nOut0_53[29] , 
        \nScanOut21[19] , \nScanOut54[30] , \nScanOut97[6] , \nScanOut77[18] , 
        \nScanOut22[7] , \nOut0_29[4] , \nScanOut54[29] , \nScanOut123[4] , 
        \nScanOut1[16] , \nOut1_4[31] , \nScanOut21[4] , \nOut0_37[8] , 
        \nScanOut120[7] , \nOut1_4[28] , \nScanOut69[20] , \nScanOut8[0] , 
        \nOut0_56[1] , \nOut1_15[13] , \nOut1_36[22] , \nOut0_55[2] , 
        \nOut0_38[12] , \nOut1_43[12] , \nScanOut91[8] , \nScanOut115[27] , 
        \nOut1_60[23] , \nScanOut87[15] , \nOut1_13[3] , \nOut1_23[16] , 
        \nOut0_58[16] , \nScanOut92[21] , \nScanOut123[22] , \nOut0_32[5] , 
        \nOut1_56[26] , \nScanOut100[13] , \nScanOut24[9] , \nScanOut39[6] , 
        \nScanOut69[13] , \nScanOut1[25] , \nOut1_23[25] , \nOut1_56[15] , 
        \nScanOut92[12] , \nScanOut123[11] , \nScanOut100[20] , \nOut0_58[25] , 
        \nOut1_36[11] , \nOut0_38[21] , \nOut1_43[21] , \nScanOut115[14] , 
        \nScanOut126[9] , \nOut1_60[10] , \nOut1_10[0] , \nOut1_15[20] , 
        \nOut0_31[6] , \nScanOut87[26] , \nOut1_0[23] , \nOut1_0[10] , 
        \nOut1_0[3] , \nOut1_3[0] , \nScanOut13[17] , \nOut0_14[24] , 
        \nOut0_37[15] , \nOut1_39[25] , \nOut0_42[25] , \nOut1_56[5] , 
        \nOut0_61[14] , \nScanOut88[12] , \nOut0_22[21] , \nOut0_57[11] , 
        \nScanOut25[12] , \nOut1_48[9] , \nOut1_59[21] , \nOut1_55[6] , 
        \nScanOut73[13] , \nScanOut30[26] , \nScanOut50[22] , \nScanOut45[16] , 
        \nScanOut66[27] , \nOut0_10[4] , \nOut0_13[7] , \nScanOut18[4] , 
        \nOut0_22[12] , \nScanOut104[8] , \nOut1_32[1] , \nOut0_14[17] , 
        \nOut0_37[26] , \nOut0_57[22] , \nOut1_59[12] , \nScanOut119[7] , 
        \nOut1_39[16] , \nOut0_42[16] , \nOut1_31[2] , \nScanOut45[25] , 
        \nOut0_61[27] , \nScanOut88[21] , \nScanOut13[24] , \nScanOut30[15] , 
        \nScanOut66[14] , \nScanOut25[21] , \nScanOut50[11] , \nScanOut73[20] , 
        \nScanOut18[31] , \nScanOut67[1] , \nScanOut96[19] , \nOut1_11[18] , 
        \nScanOut18[28] , \nOut1_29[0] , \nOut1_53[8] , \nScanOut64[2] , 
        \nOut1_32[29] , \nOut1_47[19] , \nOut0_49[29] , \nOut0_15[9] , 
        \nOut1_32[30] , \nOut0_49[30] , \nScanOut102[6] , \nScanOut127[29] , 
        \nScanOut104[18] , \nScanOut127[30] , \nScanOut101[5] , 
        \nScanOut24[0] , \nScanOut125[3] , \nOut1_4[12] , \nOut1_15[30] , 
        \nOut1_36[18] , \nOut0_38[28] , \nOut1_43[28] , \nScanOut126[0] , 
        \nOut1_15[29] , \nOut0_38[31] , \nOut1_43[31] , \nOut1_60[19] , 
        \nScanOut100[30] , \nScanOut100[29] , \nScanOut123[18] , \nOut1_4[21] , 
        \nOut0_8[4] , \nOut1_10[9] , \nScanOut27[3] , \nScanOut69[30] , 
        \nScanOut8[9] , \nScanOut69[29] , \nScanOut92[2] , \nScanOut40[4] , 
        \nOut0_56[8] , \nScanOut43[7] , \nOut0_1[24] , \nOut0_1[17] , 
        \nScanOut0[26] , \nScanOut0[15] , \nOut0_10[26] , \nOut1_15[4] , 
        \nScanOut17[15] , \nScanOut34[24] , \nOut0_48[4] , \nScanOut92[31] , 
        \nScanOut92[28] , \nScanOut91[1] , \nScanOut41[14] , \nOut0_34[2] , 
        \nScanOut62[25] , \nScanOut77[11] , \nOut1_16[7] , \nScanOut21[10] , 
        \nOut0_26[23] , \nOut1_28[13] , \nOut0_53[13] , \nScanOut54[20] , 
        \nScanOut99[24] , \nScanOut128[27] , \nOut0_37[1] , \nOut0_46[27] , 
        \nOut0_33[17] , \nOut1_48[17] , \nOut0_10[15] , \nScanOut17[26] , 
        \nScanOut21[23] , \nScanOut54[13] , \nScanOut77[22] , \nScanOut34[17] , 
        \nScanOut41[27] , \nOut0_50[6] , \nScanOut62[16] , \nScanOut89[3] , 
        \nOut0_33[24] , \nOut1_48[24] , \nOut0_46[14] , \nOut1_14[10] , 
        \nOut1_22[15] , \nOut0_26[10] , \nScanOut99[17] , \nScanOut128[14] , 
        \nOut1_28[20] , \nScanOut45[9] , \nOut0_53[5] , \nOut0_53[20] , 
        \nScanOut58[6] , \nOut0_59[15] , \nOut1_57[25] , \nScanOut101[10] , 
        \nScanOut93[22] , \nScanOut122[21] , \nOut1_61[20] , \nScanOut86[16] , 
        \nOut0_21[5] , \nOut1_37[21] , \nOut0_39[11] , \nOut1_42[11] , 
        \nScanOut114[24] , \nOut0_45[1] , \nOut0_46[2] , \nScanOut68[23] , 
        \nScanOut82[8] , \nScanOut37[9] , \nOut1_61[13] , \nScanOut0[1] , 
        \nOut0_5[1] , \nOut1_14[23] , \nOut1_22[26] , \nOut1_37[12] , 
        \nOut0_39[22] , \nOut1_42[22] , \nScanOut86[25] , \nScanOut114[17] , 
        \nOut1_57[16] , \nScanOut101[23] , \nOut0_59[26] , \nScanOut122[12] , 
        \nOut1_5[18] , \nOut0_6[2] , \nScanOut93[11] , \nScanOut68[10] , 
        \nOut0_22[6] , \nScanOut29[5] , \nScanOut128[6] , \nScanOut87[5] , 
        \nScanOut3[2] , \nScanOut20[30] , \nScanOut20[29] , \nScanOut55[19] , 
        \nScanOut55[3] , \nOut1_62[9] , \nScanOut76[31] , \nScanOut76[28] , 
        \nScanOut56[0] , \nScanOut99[9] , \nOut0_27[30] , \nOut0_27[29] , 
        \nOut1_29[19] , \nOut0_52[19] , \nScanOut84[6] , \nScanOut31[7] , 
        \nOut1_1[30] , \nOut1_1[29] , \nOut0_5[26] , \nOut0_5[15] , 
        \nScanOut15[1] , \nScanOut16[2] , \nOut1_18[1] , \nOut0_39[7] , 
        \nOut1_21[8] , \nOut0_24[8] , \nScanOut32[4] , \nScanOut117[1] , 
        \nOut0_23[18] , \nOut0_56[28] , \nOut1_58[18] , \nOut0_56[31] , 
        \nScanOut24[18] , \nScanOut114[2] , \nScanOut51[31] , \nScanOut51[28] , 
        \nScanOut72[6] , \nOut1_58[3] , \nScanOut72[19] , \nScanOut19[11] , 
        \nScanOut71[5] , \nScanOut89[18] , \nScanOut79[15] , \nScanOut4[17] , 
        \nOut1_10[12] , \nOut1_24[5] , \nOut1_27[6] , \nScanOut82[14] , 
        \nScanOut19[22] , \nOut1_26[17] , \nOut1_33[23] , \nOut1_46[13] , 
        \nOut0_48[23] , \nScanOut110[26] , \nOut0_28[27] , \nScanOut105[12] , 
        \nOut1_43[2] , \nOut1_53[27] , \nOut0_62[4] , \nScanOut97[20] , 
        \nScanOut126[23] , \nScanOut74[8] , \nOut1_26[24] , \nOut0_28[14] , 
        \nScanOut69[7] , \nScanOut79[26] , \nScanOut105[21] , \nOut1_53[14] , 
        \nScanOut126[10] , \nOut0_0[4] , \nScanOut4[24] , \nScanOut97[13] , 
        \nOut0_5[9] , \nOut1_5[10] , \nOut1_10[21] , \nOut1_33[10] , 
        \nOut1_46[20] , \nScanOut82[27] , \nScanOut110[15] , \nOut1_40[1] , 
        \nOut0_48[10] , \nOut0_61[7] , \nScanOut68[18] , \nScanOut34[2] , 
        \nScanOut37[1] , \nOut1_5[23] , \nScanOut5[4] , \nScanOut50[6] , 
        \nScanOut93[19] , \nScanOut6[7] , \nScanOut82[0] , \nScanOut122[29] , 
        \nOut1_14[18] , \nOut1_37[29] , \nScanOut101[18] , \nScanOut122[30] , 
        \nOut0_39[19] , \nOut0_58[6] , \nOut1_42[19] , \nScanOut81[3] , 
        \nOut1_61[31] , \nOut1_37[30] , \nOut0_45[9] , \nOut1_61[28] , 
        \nScanOut53[5] , \nOut1_0[18] , \nOut1_1[21] , \nOut1_1[12] , 
        \nScanOut0[9] , \nOut0_3[7] , \nOut0_11[24] , \nScanOut16[17] , 
        \nOut1_18[9] , \nScanOut35[26] , \nScanOut40[16] , \nScanOut20[12] , 
        \nScanOut63[27] , \nScanOut76[13] , \nOut0_24[0] , \nOut0_27[21] , 
        \nOut1_29[11] , \nScanOut55[22] , \nScanOut98[26] , \nOut0_52[11] , 
        \nOut0_27[3] , \nOut0_32[15] , \nOut0_47[25] , \nOut1_49[15] , 
        \nScanOut16[24] , \nScanOut20[21] , \nScanOut55[11] , \nScanOut76[20] , 
        \nScanOut35[15] , \nOut0_40[4] , \nOut1_61[2] , \nScanOut40[25] , 
        \nScanOut56[8] , \nScanOut63[14] , \nScanOut99[1] , \nOut1_10[30] , 
        \nOut0_11[17] , \nOut0_32[26] , \nScanOut48[4] , \nOut0_47[16] , 
        \nOut1_49[26] , \nScanOut12[26] , \nScanOut12[15] , \nOut0_15[26] , 
        \nOut0_27[12] , \nScanOut98[15] , \nOut1_29[22] , \nOut0_43[7] , 
        \nOut1_62[1] , \nOut0_36[17] , \nOut1_38[27] , \nOut0_43[27] , 
        \nOut0_52[22] , \nOut1_46[7] , \nOut0_60[16] , \nScanOut89[10] , 
        \nOut0_23[23] , \nOut0_56[13] , \nOut1_58[23] , \nScanOut24[10] , 
        \nScanOut72[11] , \nScanOut31[24] , \nOut1_45[4] , \nScanOut51[20] , 
        \nScanOut44[14] , \nOut0_15[15] , \nScanOut15[9] , \nOut1_22[3] , 
        \nOut1_58[10] , \nScanOut67[25] , \nOut0_23[10] , \nOut0_36[24] , 
        \nOut0_56[20] , \nOut1_38[14] , \nOut0_43[14] , \nScanOut109[5] , 
        \nOut1_21[0] , \nOut0_60[25] , \nScanOut89[23] , \nScanOut117[9] , 
        \nScanOut31[17] , \nScanOut44[27] , \nScanOut67[16] , \nScanOut24[23] , 
        \nScanOut51[13] , \nScanOut72[22] , \nOut1_33[18] , \nOut1_46[28] , 
        \nScanOut105[30] , \nScanOut105[29] , \nScanOut126[18] , 
        \nOut0_48[18] , \nOut1_10[29] , \nOut1_46[31] , \nOut1_40[9] , 
        \nScanOut74[0] , \nScanOut77[3] , \nOut1_8[3] , \nScanOut13[7] , 
        \nOut0_18[4] , \nOut1_39[2] , \nScanOut19[19] , \nScanOut97[31] , 
        \nScanOut97[28] , \nScanOut112[4] , \nScanOut111[7] , \nOut1_3[8] , 
        \nOut0_4[17] , \nScanOut10[4] , \nScanOut25[30] , \nScanOut25[29] , 
        \nScanOut50[19] , \nScanOut73[31] , \nScanOut73[28] , \nScanOut107[3] , 
        \nOut0_4[24] , \nOut0_22[30] , \nOut0_22[29] , \nOut1_32[9] , 
        \nScanOut104[0] , \nOut1_48[1] , \nScanOut88[30] , \nScanOut88[29] , 
        \nOut0_57[19] , \nScanOut61[7] , \nScanOut62[4] , \nOut1_59[29] , 
        \nOut1_59[30] , \nOut1_5[6] , \nScanOut5[15] , \nOut1_6[5] , 
        \nOut0_16[2] , \nOut1_37[4] , \nOut1_11[10] , \nScanOut18[13] , 
        \nScanOut78[17] , \nScanOut83[16] , \nOut0_15[1] , \nOut1_27[15] , 
        \nOut1_29[8] , \nOut1_32[21] , \nOut0_49[21] , \nOut1_47[11] , 
        \nScanOut111[24] , \nOut0_29[25] , \nOut1_52[25] , \nOut1_34[7] , 
        \nScanOut96[22] , \nScanOut104[10] , \nScanOut127[21] , 
        \nScanOut1[24] , \nScanOut1[17] , \nScanOut5[26] , \nScanOut18[20] , 
        \nOut1_27[26] , \nOut0_29[16] , \nOut1_50[3] , \nOut1_53[0] , 
        \nScanOut78[24] , \nScanOut79[5] , \nOut1_52[16] , \nScanOut67[9] , 
        \nScanOut104[23] , \nScanOut96[11] , \nScanOut127[12] , \nOut1_11[23] , 
        \nScanOut83[25] , \nOut1_15[12] , \nOut1_23[17] , \nOut1_32[12] , 
        \nOut1_47[22] , \nScanOut111[17] , \nOut0_49[12] , \nOut0_55[3] , 
        \nOut1_56[27] , \nOut0_58[17] , \nScanOut87[14] , \nScanOut92[20] , 
        \nScanOut100[12] , \nScanOut123[23] , \nOut1_4[30] , \nOut1_4[29] , 
        \nOut1_36[23] , \nOut1_60[22] , \nOut0_38[13] , \nScanOut91[9] , 
        \nOut1_43[13] , \nScanOut115[26] , \nScanOut69[21] , \nScanOut8[1] , 
        \nOut0_56[0] , \nOut1_15[21] , \nOut1_60[11] , \nScanOut87[27] , 
        \nOut1_23[24] , \nOut1_36[10] , \nOut0_38[20] , \nOut1_43[20] , 
        \nScanOut115[15] , \nScanOut126[8] , \nOut1_56[14] , \nScanOut100[21] , 
        \nOut0_58[24] , \nScanOut92[13] , \nScanOut123[10] , \nOut1_10[1] , 
        \nOut0_31[7] , \nOut1_13[2] , \nOut0_32[4] , \nScanOut24[8] , 
        \nOut0_0[26] , \nOut0_0[15] , \nOut0_26[18] , \nScanOut39[7] , 
        \nScanOut69[12] , \nOut1_28[31] , \nOut1_28[28] , \nScanOut45[1] , 
        \nOut0_53[28] , \nOut0_53[31] , \nScanOut97[7] , \nScanOut46[2] , 
        \nScanOut94[4] , \nScanOut120[6] , \nOut1_0[22] , \nOut1_0[11] , 
        \nScanOut21[18] , \nScanOut21[5] , \nOut0_37[9] , \nScanOut22[6] , 
        \nScanOut54[28] , \nOut0_29[5] , \nScanOut54[31] , \nScanOut77[19] , 
        \nScanOut123[5] , \nScanOut18[30] , \nScanOut18[29] , \nOut1_53[9] , 
        \nScanOut64[3] , \nScanOut67[0] , \nScanOut96[18] , \nOut1_0[2] , 
        \nOut0_10[5] , \nOut1_11[19] , \nOut0_49[31] , \nScanOut101[4] , 
        \nScanOut102[7] , \nScanOut104[19] , \nScanOut127[31] , 
        \nScanOut127[28] , \nScanOut13[25] , \nScanOut13[16] , \nOut0_15[8] , 
        \nOut1_29[1] , \nOut1_32[31] , \nOut0_49[28] , \nOut1_32[28] , 
        \nOut1_47[18] , \nOut1_48[8] , \nOut0_14[25] , \nOut0_22[20] , 
        \nScanOut25[13] , \nScanOut30[27] , \nScanOut66[26] , \nScanOut45[17] , 
        \nScanOut50[23] , \nOut1_55[7] , \nOut0_57[10] , \nScanOut73[12] , 
        \nOut1_59[20] , \nOut0_61[15] , \nScanOut88[13] , \nScanOut25[20] , 
        \nOut0_37[14] , \nOut1_39[24] , \nOut0_42[24] , \nOut1_56[4] , 
        \nScanOut50[10] , \nScanOut66[15] , \nScanOut73[21] , \nOut1_31[3] , 
        \nScanOut30[14] , \nScanOut45[24] , \nOut1_3[1] , \nScanOut18[5] , 
        \nScanOut104[9] , \nOut0_8[5] , \nOut0_10[27] , \nOut0_13[6] , 
        \nOut0_14[16] , \nOut0_22[13] , \nOut1_32[0] , \nOut0_37[27] , 
        \nOut0_61[26] , \nScanOut88[20] , \nOut1_39[17] , \nOut0_42[17] , 
        \nScanOut119[6] , \nOut1_59[13] , \nOut0_57[23] , \nOut0_10[14] , 
        \nOut1_15[5] , \nOut1_16[6] , \nOut0_37[0] , \nScanOut21[11] , 
        \nOut0_26[22] , \nOut1_28[12] , \nOut0_33[16] , \nOut0_46[26] , 
        \nOut1_48[16] , \nOut0_53[12] , \nScanOut99[25] , \nScanOut128[26] , 
        \nOut0_34[3] , \nScanOut17[14] , \nScanOut54[21] , \nScanOut77[10] , 
        \nOut0_26[11] , \nScanOut34[25] , \nScanOut62[24] , \nScanOut41[15] , 
        \nOut1_28[21] , \nOut0_53[4] , \nScanOut45[8] , \nOut0_53[21] , 
        \nScanOut99[16] , \nScanOut128[15] , \nOut1_10[8] , \nOut1_15[31] , 
        \nOut1_15[28] , \nScanOut17[27] , \nOut0_33[25] , \nOut0_46[15] , 
        \nOut1_48[25] , \nScanOut58[7] , \nScanOut62[17] , \nScanOut21[22] , 
        \nScanOut34[16] , \nScanOut41[26] , \nOut0_50[7] , \nScanOut54[12] , 
        \nScanOut89[2] , \nOut0_38[30] , \nScanOut77[23] , \nScanOut100[31] , 
        \nScanOut100[28] , \nScanOut123[19] , \nOut1_43[30] , \nOut1_60[18] , 
        \nOut1_36[19] , \nOut0_38[29] , \nScanOut126[1] , \nOut1_43[29] , 
        \nScanOut27[2] , \nOut1_4[13] , \nScanOut24[1] , \nScanOut125[2] , 
        \nOut0_1[25] , \nOut0_1[16] , \nScanOut3[3] , \nOut1_4[20] , 
        \nScanOut43[6] , \nOut0_48[5] , \nScanOut69[28] , \nScanOut91[0] , 
        \nScanOut92[30] , \nScanOut92[29] , \nScanOut92[3] , \nScanOut8[8] , 
        \nScanOut40[5] , \nOut0_56[9] , \nScanOut69[31] , \nScanOut20[31] , 
        \nScanOut56[1] , \nScanOut76[29] , \nScanOut99[8] , \nScanOut20[28] , 
        \nScanOut55[18] , \nScanOut76[30] , \nScanOut84[7] , \nScanOut0[0] , 
        \nScanOut87[4] , \nOut1_18[0] , \nOut0_39[6] , \nScanOut55[2] , 
        \nOut1_62[8] , \nOut0_24[9] , \nOut0_27[31] , \nScanOut31[6] , 
        \nScanOut32[5] , \nOut0_27[28] , \nOut1_29[18] , \nOut0_52[18] , 
        \nOut1_1[31] , \nScanOut0[27] , \nScanOut0[14] , \nOut1_14[11] , 
        \nOut1_37[20] , \nOut0_46[3] , \nScanOut68[22] , \nScanOut82[9] , 
        \nOut0_39[10] , \nOut1_42[10] , \nScanOut114[25] , \nScanOut86[17] , 
        \nOut0_5[0] , \nOut1_5[19] , \nOut0_6[3] , \nOut1_22[14] , 
        \nOut1_61[21] , \nScanOut93[23] , \nScanOut122[20] , \nScanOut29[4] , 
        \nOut0_45[0] , \nOut1_57[24] , \nOut0_59[14] , \nScanOut101[11] , 
        \nOut0_21[4] , \nOut0_22[7] , \nScanOut68[11] , \nScanOut128[7] , 
        \nScanOut37[8] , \nOut1_22[27] , \nOut1_57[17] , \nScanOut93[10] , 
        \nScanOut122[13] , \nScanOut101[22] , \nOut1_37[13] , \nOut0_39[23] , 
        \nOut0_59[27] , \nOut1_42[23] , \nScanOut114[16] , \nScanOut4[16] , 
        \nOut1_10[13] , \nOut1_14[22] , \nOut1_61[12] , \nScanOut86[24] , 
        \nOut1_24[4] , \nOut1_26[16] , \nScanOut97[21] , \nScanOut126[22] , 
        \nOut0_28[26] , \nOut1_53[26] , \nOut1_33[22] , \nOut0_48[22] , 
        \nScanOut105[13] , \nOut1_46[12] , \nScanOut110[27] , \nScanOut82[15] , 
        \nOut1_1[28] , \nScanOut19[10] , \nScanOut4[25] , \nOut1_27[7] , 
        \nScanOut79[14] , \nOut1_33[11] , \nOut1_46[21] , \nScanOut110[14] , 
        \nOut0_48[11] , \nOut1_10[20] , \nScanOut82[26] , \nScanOut126[11] , 
        \nOut0_0[22] , \nOut0_0[11] , \nOut0_5[27] , \nOut0_5[14] , 
        \nScanOut15[0] , \nScanOut19[23] , \nOut1_26[25] , \nOut0_28[15] , 
        \nOut1_53[15] , \nScanOut97[12] , \nScanOut105[20] , \nOut1_40[0] , 
        \nOut0_61[6] , \nOut1_43[3] , \nOut0_62[5] , \nScanOut69[6] , 
        \nScanOut74[9] , \nScanOut79[27] , \nOut0_23[19] , \nOut0_56[30] , 
        \nOut1_58[19] , \nOut0_56[29] , \nScanOut114[3] , \nScanOut16[3] , 
        \nOut1_21[9] , \nScanOut117[0] , \nScanOut24[19] , \nScanOut51[30] , 
        \nScanOut71[4] , \nScanOut89[19] , \nScanOut72[18] , \nScanOut46[6] , 
        \nScanOut51[29] , \nOut1_58[2] , \nScanOut72[7] , \nScanOut94[0] , 
        \nOut0_10[19] , \nOut0_33[31] , \nOut0_33[28] , \nScanOut45[5] , 
        \nOut0_53[9] , \nScanOut97[3] , \nScanOut128[18] , \nOut0_46[18] , 
        \nOut1_48[28] , \nOut1_15[8] , \nOut0_29[1] , \nOut1_48[31] , 
        \nScanOut123[1] , \nScanOut17[19] , \nScanOut22[2] , \nScanOut34[31] , 
        \nScanOut34[28] , \nScanOut41[18] , \nScanOut62[30] , \nScanOut21[1] , 
        \nScanOut62[29] , \nScanOut99[31] , \nScanOut99[28] , \nScanOut1[13] , 
        \nScanOut8[5] , \nScanOut40[8] , \nOut0_56[4] , \nScanOut120[2] , 
        \nOut1_15[16] , \nOut1_36[27] , \nScanOut69[25] , \nOut0_38[17] , 
        \nOut0_48[8] , \nOut1_43[17] , \nScanOut115[22] , \nScanOut87[10] , 
        \nOut1_60[26] , \nOut1_23[13] , \nScanOut92[24] , \nScanOut123[27] , 
        \nScanOut39[3] , \nOut0_55[7] , \nOut1_56[23] , \nOut0_58[13] , 
        \nScanOut100[16] , \nScanOut69[16] , \nOut1_1[16] , \nScanOut1[20] , 
        \nOut0_8[8] , \nOut1_13[6] , \nOut0_32[0] , \nOut1_10[5] , 
        \nOut0_31[3] , \nOut1_23[20] , \nOut1_56[10] , \nScanOut92[17] , 
        \nScanOut123[14] , \nScanOut100[25] , \nOut1_36[14] , \nOut0_38[24] , 
        \nOut0_58[20] , \nOut1_43[24] , \nScanOut115[11] , \nOut1_60[15] , 
        \nOut0_4[20] , \nOut0_4[13] , \nOut1_5[2] , \nScanOut5[11] , 
        \nOut1_11[14] , \nOut0_15[5] , \nOut1_15[25] , \nScanOut87[23] , 
        \nOut1_34[3] , \nOut1_27[11] , \nScanOut96[26] , \nScanOut127[25] , 
        \nOut0_29[21] , \nOut1_52[21] , \nOut1_32[25] , \nOut0_49[25] , 
        \nScanOut104[14] , \nOut1_47[15] , \nScanOut111[20] , \nScanOut83[12] , 
        \nScanOut5[22] , \nOut1_6[1] , \nScanOut18[17] , \nScanOut101[9] , 
        \nOut0_16[6] , \nOut1_37[0] , \nScanOut78[13] , \nOut1_32[16] , 
        \nOut1_47[26] , \nScanOut111[13] , \nOut0_49[16] , \nOut1_11[27] , 
        \nScanOut83[21] , \nScanOut18[24] , \nOut1_27[22] , \nOut0_29[12] , 
        \nOut1_52[12] , \nScanOut96[15] , \nScanOut127[16] , \nScanOut104[27] , 
        \nOut1_50[7] , \nOut1_53[4] , \nScanOut78[20] , \nScanOut79[1] , 
        \nScanOut104[4] , \nOut0_10[8] , \nScanOut18[8] , \nScanOut107[7] , 
        \nScanOut13[31] , \nScanOut45[29] , \nScanOut13[28] , \nScanOut30[19] , 
        \nScanOut45[30] , \nScanOut66[18] , \nOut0_14[31] , \nOut1_39[29] , 
        \nOut0_42[29] , \nOut1_56[9] , \nOut0_14[28] , \nOut0_37[19] , 
        \nScanOut61[3] , \nOut1_39[30] , \nOut0_42[30] , \nOut0_61[18] , 
        \nOut1_48[5] , \nScanOut62[0] , \nScanOut4[31] , \nScanOut4[28] , 
        \nOut0_62[8] , \nScanOut74[4] , \nScanOut77[7] , \nScanOut110[19] , 
        \nOut1_26[28] , \nOut0_28[18] , \nOut1_53[18] , \nOut0_0[0] , 
        \nOut0_1[31] , \nOut1_1[25] , \nScanOut10[0] , \nOut1_26[31] , 
        \nOut0_3[3] , \nOut0_5[19] , \nOut1_8[7] , \nOut0_18[0] , 
        \nOut1_39[6] , \nScanOut79[19] , \nScanOut111[3] , \nScanOut82[18] , 
        \nScanOut112[0] , \nScanOut12[22] , \nScanOut12[11] , \nScanOut13[3] , 
        \nOut1_24[9] , \nOut0_15[22] , \nOut0_23[27] , \nScanOut24[14] , 
        \nScanOut31[20] , \nScanOut67[21] , \nScanOut44[10] , \nOut1_45[0] , 
        \nScanOut51[24] , \nOut0_56[17] , \nScanOut72[15] , \nOut1_58[27] , 
        \nOut0_60[12] , \nScanOut89[14] , \nScanOut24[27] , \nOut0_36[13] , 
        \nOut1_38[23] , \nOut0_43[23] , \nOut1_46[3] , \nScanOut51[17] , 
        \nScanOut71[9] , \nScanOut67[12] , \nScanOut72[26] , \nOut1_21[4] , 
        \nScanOut31[13] , \nScanOut44[23] , \nOut0_15[11] , \nOut1_22[7] , 
        \nOut0_23[14] , \nOut0_36[20] , \nOut0_60[21] , \nScanOut89[27] , 
        \nOut1_38[10] , \nOut0_43[10] , \nScanOut109[1] , \nOut1_58[14] , 
        \nOut0_56[24] , \nOut0_1[28] , \nOut0_11[20] , \nScanOut16[13] , 
        \nScanOut20[16] , \nOut0_27[25] , \nOut0_27[7] , \nOut1_29[15] , 
        \nOut0_32[11] , \nOut0_47[21] , \nOut1_49[11] , \nOut0_52[15] , 
        \nScanOut98[22] , \nOut0_24[4] , \nScanOut32[8] , \nScanOut55[26] , 
        \nScanOut76[17] , \nScanOut35[22] , \nScanOut63[23] , \nScanOut40[12] , 
        \nScanOut0[19] , \nOut1_5[14] , \nOut0_11[13] , \nOut0_27[16] , 
        \nOut1_62[5] , \nOut1_29[26] , \nOut0_43[3] , \nOut0_52[26] , 
        \nScanOut98[11] , \nScanOut16[20] , \nOut0_32[22] , \nOut0_47[12] , 
        \nOut1_49[22] , \nScanOut48[0] , \nScanOut87[9] , \nScanOut63[10] , 
        \nScanOut20[25] , \nScanOut35[11] , \nOut0_40[0] , \nOut1_61[6] , 
        \nScanOut40[21] , \nScanOut55[15] , \nScanOut99[5] , \nOut0_21[9] , 
        \nScanOut76[24] , \nScanOut86[30] , \nScanOut86[29] , \nScanOut34[6] , 
        \nScanOut37[5] , \nScanOut29[9] , \nScanOut53[1] , \nScanOut114[31] , 
        \nScanOut4[12] , \nOut0_5[23] , \nOut0_5[10] , \nOut1_5[27] , 
        \nScanOut6[3] , \nOut1_22[19] , \nOut0_58[2] , \nScanOut81[7] , 
        \nScanOut114[28] , \nOut1_57[30] , \nOut1_57[29] , \nOut0_59[19] , 
        \nScanOut82[4] , \nScanOut5[0] , \nScanOut16[7] , \nScanOut50[2] , 
        \nScanOut117[4] , \nScanOut12[18] , \nOut0_15[18] , \nScanOut15[4] , 
        \nScanOut114[7] , \nOut0_36[30] , \nScanOut31[30] , \nOut0_36[29] , 
        \nOut0_60[28] , \nOut1_38[19] , \nOut0_43[19] , \nOut0_60[31] , 
        \nScanOut109[8] , \nOut1_45[9] , \nOut1_58[6] , \nScanOut72[3] , 
        \nScanOut31[29] , \nScanOut67[28] , \nScanOut44[19] , \nScanOut67[31] , 
        \nScanOut71[0] , \nOut1_10[17] , \nScanOut10[9] , \nOut1_27[3] , 
        \nScanOut19[14] , \nScanOut79[10] , \nScanOut82[11] , \nOut0_18[9] , 
        \nOut0_48[26] , \nScanOut19[27] , \nOut1_24[0] , \nOut1_26[12] , 
        \nOut1_33[26] , \nOut1_46[16] , \nScanOut110[23] , \nOut0_28[22] , 
        \nOut1_53[22] , \nScanOut112[9] , \nScanOut97[25] , \nScanOut105[17] , 
        \nScanOut126[26] , \nOut1_26[21] , \nOut0_28[11] , \nOut1_40[4] , 
        \nOut1_43[7] , \nOut0_62[1] , \nScanOut69[2] , \nScanOut79[23] , 
        \nOut0_61[2] , \nOut1_53[11] , \nScanOut105[24] , \nScanOut126[15] , 
        \nOut0_0[9] , \nOut0_1[21] , \nOut0_1[12] , \nScanOut0[23] , 
        \nScanOut0[10] , \nScanOut4[21] , \nScanOut97[16] , \nOut1_10[24] , 
        \nScanOut82[22] , \nOut1_14[15] , \nOut1_22[10] , \nOut1_33[15] , 
        \nOut1_46[25] , \nScanOut110[10] , \nOut0_48[15] , \nOut0_45[4] , 
        \nScanOut53[8] , \nOut1_57[20] , \nOut0_59[10] , \nScanOut86[13] , 
        \nScanOut93[27] , \nScanOut101[15] , \nScanOut122[24] , \nOut1_61[25] , 
        \nScanOut5[9] , \nOut1_37[24] , \nOut0_39[14] , \nOut1_42[14] , 
        \nScanOut114[21] , \nScanOut68[26] , \nOut0_46[7] , \nOut1_61[16] , 
        \nScanOut0[4] , \nOut0_5[4] , \nOut1_14[26] , \nScanOut86[20] , 
        \nOut1_22[23] , \nOut1_37[17] , \nOut0_39[27] , \nOut1_42[27] , 
        \nScanOut114[12] , \nOut1_57[13] , \nScanOut101[26] , \nOut0_59[23] , 
        \nOut0_6[7] , \nOut0_21[0] , \nScanOut93[14] , \nScanOut122[17] , 
        \nOut0_22[3] , \nScanOut128[3] , \nScanOut29[0] , \nScanOut68[15] , 
        \nScanOut55[6] , \nScanOut98[18] , \nScanOut48[9] , \nScanOut87[0] , 
        \nScanOut3[7] , \nScanOut16[30] , \nScanOut16[29] , \nScanOut40[31] , 
        \nScanOut84[3] , \nScanOut63[19] , \nOut0_40[9] , \nScanOut40[28] , 
        \nScanOut56[5] , \nScanOut35[18] , \nOut0_11[30] , \nOut0_11[29] , 
        \nOut0_47[31] , \nScanOut31[2] , \nOut0_47[28] , \nOut1_18[4] , 
        \nOut0_32[18] , \nScanOut32[1] , \nOut1_49[18] , \nOut0_39[2] , 
        \nOut1_4[17] , \nScanOut125[6] , \nScanOut24[5] , \nOut0_32[9] , 
        \nScanOut1[30] , \nOut0_8[1] , \nScanOut27[6] , \nScanOut115[18] , 
        \nScanOut126[5] , \nScanOut1[29] , \nOut1_4[24] , \nOut1_23[30] , 
        \nOut1_23[29] , \nOut1_56[19] , \nOut0_58[30] , \nScanOut40[1] , 
        \nOut0_58[29] , \nScanOut43[2] , \nOut0_48[1] , \nScanOut92[7] , 
        \nScanOut87[19] , \nScanOut91[4] , \nOut0_0[18] , \nOut0_10[23] , 
        \nOut1_15[1] , \nScanOut17[10] , \nOut0_29[8] , \nScanOut123[8] , 
        \nScanOut34[21] , \nScanOut41[11] , \nScanOut21[15] , \nScanOut62[20] , 
        \nScanOut77[14] , \nOut0_34[7] , \nOut1_16[2] , \nOut0_26[26] , 
        \nOut1_28[16] , \nScanOut54[25] , \nScanOut99[21] , \nScanOut128[22] , 
        \nOut0_53[16] , \nOut0_37[4] , \nOut0_46[22] , \nScanOut21[8] , 
        \nOut0_33[12] , \nOut1_48[12] , \nScanOut17[23] , \nScanOut21[26] , 
        \nScanOut54[16] , \nScanOut77[27] , \nScanOut34[12] , \nScanOut41[22] , 
        \nOut0_50[3] , \nScanOut62[13] , \nScanOut89[6] , \nScanOut94[9] , 
        \nOut1_0[26] , \nOut1_0[15] , \nOut1_0[6] , \nOut1_3[5] , 
        \nOut0_4[30] , \nOut0_4[29] , \nOut0_10[10] , \nOut0_33[21] , 
        \nScanOut58[3] , \nOut0_46[11] , \nOut1_48[21] , \nOut0_26[15] , 
        \nScanOut99[12] , \nScanOut128[11] , \nOut1_28[25] , \nOut0_53[0] , 
        \nOut0_53[25] , \nOut0_13[2] , \nScanOut13[12] , \nOut0_14[21] , 
        \nOut0_37[10] , \nOut1_39[20] , \nOut0_42[20] , \nOut1_56[0] , 
        \nOut0_61[11] , \nScanOut88[17] , \nOut0_22[24] , \nOut0_57[14] , 
        \nOut1_59[24] , \nScanOut25[17] , \nScanOut73[16] , \nScanOut30[23] , 
        \nScanOut50[27] , \nOut1_55[3] , \nScanOut62[9] , \nScanOut45[13] , 
        \nOut0_22[17] , \nOut1_59[17] , \nScanOut66[22] , \nOut1_32[4] , 
        \nOut0_14[12] , \nOut0_37[23] , \nOut0_57[27] , \nOut1_39[13] , 
        \nOut0_42[13] , \nScanOut119[2] , \nOut0_61[22] , \nScanOut88[24] , 
        \nScanOut18[1] , \nOut0_10[1] , \nOut1_31[7] , \nScanOut13[21] , 
        \nScanOut30[10] , \nScanOut45[20] , \nScanOut66[11] , \nScanOut25[24] , 
        \nScanOut50[14] , \nScanOut73[25] , \nScanOut64[7] , \nScanOut67[4] , 
        \nScanOut83[31] , \nScanOut83[28] , \nScanOut79[8] , \nScanOut5[18] , 
        \nOut1_29[5] , \nScanOut78[30] , \nScanOut78[29] , \nScanOut111[30] , 
        \nScanOut111[29] , \nOut1_6[8] , \nOut1_27[18] , \nOut0_29[31] , 
        \nOut1_52[31] , \nOut0_29[28] , \nOut1_52[28] , \nScanOut102[3] , 
        \nScanOut101[0] , \nOut0_8[3] , \nOut1_37[9] , \nScanOut87[31] , 
        \nScanOut87[28] , \nScanOut126[7] , \nScanOut27[4] , \nOut0_31[8] , 
        \nOut1_4[15] , \nScanOut24[7] , \nScanOut39[8] , \nScanOut43[0] , 
        \nScanOut125[4] , \nOut0_0[30] , \nOut0_0[29] , \nScanOut1[18] , 
        \nOut0_48[3] , \nScanOut91[6] , \nScanOut115[29] , \nScanOut115[30] , 
        \nOut1_4[26] , \nOut1_23[18] , \nOut1_56[31] , \nOut1_56[28] , 
        \nOut0_58[18] , \nScanOut92[5] , \nScanOut40[3] , \nOut1_0[24] , 
        \nOut1_0[17] , \nOut1_0[4] , \nOut0_10[21] , \nOut1_16[0] , 
        \nOut0_33[10] , \nScanOut120[9] , \nOut1_48[10] , \nOut0_37[6] , 
        \nOut0_46[20] , \nOut0_10[12] , \nOut1_15[3] , \nScanOut21[17] , 
        \nScanOut22[9] , \nOut0_26[24] , \nScanOut99[23] , \nScanOut128[20] , 
        \nOut1_28[14] , \nOut0_53[14] , \nScanOut54[27] , \nScanOut77[16] , 
        \nScanOut17[12] , \nOut0_34[5] , \nScanOut34[23] , \nScanOut41[13] , 
        \nScanOut62[22] , \nOut0_26[17] , \nOut1_28[27] , \nScanOut99[10] , 
        \nScanOut128[13] , \nOut0_53[27] , \nOut0_53[2] , \nOut0_33[23] , 
        \nOut0_46[13] , \nOut1_48[23] , \nOut0_10[3] , \nScanOut13[10] , 
        \nScanOut17[21] , \nScanOut34[10] , \nScanOut58[1] , \nScanOut97[8] , 
        \nScanOut89[4] , \nScanOut41[20] , \nOut0_50[1] , \nScanOut21[24] , 
        \nScanOut62[11] , \nScanOut77[25] , \nScanOut30[21] , \nScanOut45[11] , 
        \nScanOut54[14] , \nScanOut66[20] , \nOut0_14[23] , \nOut0_22[26] , 
        \nScanOut25[15] , \nScanOut50[25] , \nScanOut73[14] , \nOut1_55[1] , 
        \nOut1_59[26] , \nOut0_37[12] , \nOut0_57[16] , \nScanOut61[8] , 
        \nOut1_39[22] , \nOut0_42[22] , \nOut1_56[2] , \nScanOut25[26] , 
        \nOut0_61[13] , \nScanOut88[15] , \nScanOut73[27] , \nScanOut30[12] , 
        \nScanOut50[16] , \nScanOut13[23] , \nOut1_31[5] , \nScanOut45[22] , 
        \nScanOut66[13] , \nOut1_3[7] , \nOut0_4[18] , \nOut0_13[0] , 
        \nOut0_14[10] , \nScanOut18[3] , \nOut0_37[21] , \nOut1_39[11] , 
        \nOut0_42[11] , \nOut0_61[20] , \nScanOut88[26] , \nScanOut119[0] , 
        \nOut0_57[25] , \nOut1_59[15] , \nOut0_22[15] , \nOut1_32[6] , 
        \nScanOut5[30] , \nScanOut64[5] , \nScanOut67[6] , \nScanOut111[18] , 
        \nScanOut5[29] , \nOut1_27[30] , \nOut1_27[29] , \nOut0_29[19] , 
        \nOut1_52[19] , \nScanOut101[2] , \nScanOut4[23] , \nScanOut4[10] , 
        \nOut0_5[21] , \nOut0_5[12] , \nOut1_5[9] , \nOut1_29[7] , 
        \nScanOut78[18] , \nScanOut102[1] , \nScanOut15[6] , \nOut1_34[8] , 
        \nScanOut83[19] , \nScanOut114[5] , \nScanOut12[30] , \nScanOut12[29] , 
        \nScanOut117[6] , \nScanOut16[5] , \nScanOut44[31] , \nScanOut67[19] , 
        \nScanOut31[18] , \nScanOut44[28] , \nScanOut13[8] , \nOut0_15[30] , 
        \nOut0_15[29] , \nOut0_36[18] , \nOut1_38[31] , \nOut0_43[31] , 
        \nOut0_60[19] , \nScanOut71[2] , \nOut1_38[28] , \nOut0_43[28] , 
        \nOut1_46[8] , \nOut1_58[4] , \nScanOut72[1] , \nOut1_24[2] , 
        \nOut1_26[10] , \nOut0_28[20] , \nOut1_53[20] , \nScanOut105[15] , 
        \nScanOut97[27] , \nScanOut126[24] , \nOut1_10[26] , \nOut1_10[15] , 
        \nScanOut82[13] , \nScanOut19[16] , \nOut1_33[24] , \nOut1_46[14] , 
        \nScanOut110[21] , \nOut0_48[24] , \nOut1_27[1] , \nScanOut79[12] , 
        \nScanOut111[8] , \nScanOut82[20] , \nOut1_26[23] , \nOut1_33[17] , 
        \nOut0_48[17] , \nOut1_46[27] , \nScanOut110[12] , \nOut0_28[13] , 
        \nOut1_53[13] , \nScanOut105[26] , \nScanOut97[14] , \nOut0_0[13] , 
        \nOut0_0[2] , \nOut0_1[23] , \nOut0_1[10] , \nScanOut0[21] , 
        \nScanOut0[12] , \nScanOut19[25] , \nOut1_40[6] , \nScanOut126[17] , 
        \nOut1_43[5] , \nOut0_61[0] , \nOut0_62[3] , \nScanOut79[21] , 
        \nOut0_46[5] , \nScanOut50[9] , \nScanOut69[0] , \nScanOut68[24] , 
        \nOut0_5[6] , \nOut0_6[5] , \nScanOut6[8] , \nOut1_14[17] , 
        \nOut1_61[27] , \nScanOut86[11] , \nOut1_22[12] , \nOut1_37[26] , 
        \nOut0_39[16] , \nScanOut114[23] , \nOut1_42[16] , \nOut1_57[22] , 
        \nOut0_58[9] , \nScanOut101[17] , \nOut0_45[6] , \nOut0_59[12] , 
        \nScanOut93[25] , \nScanOut122[26] , \nScanOut68[17] , \nOut0_21[2] , 
        \nOut0_22[1] , \nScanOut29[2] , \nScanOut128[1] , \nOut1_22[21] , 
        \nOut1_57[11] , \nOut0_59[21] , \nScanOut93[16] , \nScanOut101[24] , 
        \nOut1_14[24] , \nScanOut86[22] , \nScanOut122[15] , \nScanOut3[5] , 
        \nOut1_37[15] , \nOut1_61[14] , \nOut0_39[25] , \nScanOut114[10] , 
        \nOut1_42[25] , \nScanOut56[7] , \nScanOut84[1] , \nScanOut87[2] , 
        \nScanOut0[6] , \nOut0_3[8] , \nOut0_11[18] , \nOut0_43[8] , 
        \nScanOut55[4] , \nScanOut16[18] , \nOut1_18[6] , \nOut0_32[30] , 
        \nOut0_32[29] , \nOut0_47[19] , \nOut1_49[30] , \nOut1_49[29] , 
        \nScanOut32[3] , \nOut0_39[0] , \nScanOut63[28] , \nScanOut31[0] , 
        \nScanOut35[30] , \nScanOut35[29] , \nScanOut40[19] , \nScanOut63[31] , 
        \nScanOut98[30] , \nScanOut98[29] , \nOut1_1[27] , \nOut1_1[14] , 
        \nOut0_61[9] , \nScanOut77[5] , \nScanOut82[30] , \nScanOut82[29] , 
        \nScanOut74[6] , \nScanOut4[19] , \nOut1_8[5] , \nScanOut69[9] , 
        \nScanOut79[31] , \nScanOut79[28] , \nScanOut13[1] , \nScanOut110[31] , 
        \nOut0_18[2] , \nScanOut110[28] , \nOut1_26[19] , \nOut0_28[29] , 
        \nOut1_39[4] , \nOut1_53[29] , \nOut0_28[30] , \nOut1_53[30] , 
        \nScanOut112[2] , \nOut0_5[31] , \nScanOut10[2] , \nScanOut111[1] , 
        \nOut1_27[8] , \nOut0_5[28] , \nScanOut12[20] , \nScanOut12[13] , 
        \nOut0_15[20] , \nOut0_23[25] , \nOut0_36[11] , \nOut0_60[10] , 
        \nScanOut89[16] , \nOut1_38[21] , \nOut0_43[21] , \nOut1_46[1] , 
        \nOut1_58[25] , \nScanOut24[16] , \nScanOut51[26] , \nOut0_56[15] , 
        \nScanOut72[8] , \nOut1_45[2] , \nScanOut67[23] , \nScanOut72[17] , 
        \nOut0_15[13] , \nOut1_22[5] , \nScanOut31[22] , \nScanOut44[12] , 
        \nOut0_56[26] , \nOut1_58[16] , \nOut0_23[16] , \nOut0_60[23] , 
        \nScanOut89[25] , \nOut0_36[22] , \nOut1_38[12] , \nOut0_43[12] , 
        \nScanOut109[3] , \nOut1_21[6] , \nScanOut31[11] , \nScanOut67[10] , 
        \nScanOut24[25] , \nScanOut44[21] , \nOut0_39[9] , \nScanOut51[15] , 
        \nScanOut72[24] , \nOut0_1[19] , \nOut0_3[1] , \nOut0_11[22] , 
        \nScanOut16[11] , \nScanOut63[21] , \nScanOut20[14] , \nScanOut35[20] , 
        \nScanOut40[10] , \nScanOut55[24] , \nOut0_24[6] , \nOut0_27[27] , 
        \nScanOut76[15] , \nOut1_29[17] , \nOut0_52[17] , \nScanOut98[20] , 
        \nOut0_27[5] , \nScanOut31[9] , \nOut0_32[13] , \nOut0_47[23] , 
        \nOut1_49[13] , \nScanOut16[22] , \nScanOut20[27] , \nScanOut55[17] , 
        \nScanOut76[26] , \nScanOut35[13] , \nScanOut63[12] , \nScanOut99[7] , 
        \nOut0_40[2] , \nScanOut40[23] , \nOut1_61[4] , \nScanOut48[2] , 
        \nScanOut84[8] , \nScanOut0[31] , \nScanOut0[28] , \nOut1_5[16] , 
        \nOut0_11[11] , \nOut0_27[14] , \nOut1_29[24] , \nOut0_32[20] , 
        \nOut0_47[10] , \nOut1_49[20] , \nOut0_43[1] , \nOut0_52[24] , 
        \nOut1_62[7] , \nScanOut98[13] , \nOut0_22[8] , \nScanOut34[4] , 
        \nScanOut128[8] , \nScanOut37[7] , \nScanOut114[19] , \nOut1_5[25] , 
        \nOut1_22[31] , \nOut1_22[28] , \nOut1_57[18] , \nOut0_59[28] , 
        \nScanOut50[0] , \nOut0_59[31] , \nScanOut5[2] , \nScanOut6[1] , 
        \nScanOut82[6] , \nScanOut45[7] , \nScanOut53[3] , \nOut0_58[0] , 
        \nScanOut81[5] , \nScanOut86[18] , \nScanOut99[19] , \nScanOut58[8] , 
        \nScanOut97[1] , \nScanOut94[2] , \nOut0_0[20] , \nScanOut17[31] , 
        \nScanOut34[19] , \nScanOut46[4] , \nScanOut17[28] , \nScanOut41[29] , 
        \nOut0_50[8] , \nScanOut41[30] , \nScanOut62[18] , \nScanOut1[22] , 
        \nScanOut1[11] , \nOut0_10[31] , \nOut0_33[19] , \nScanOut120[0] , 
        \nScanOut128[30] , \nScanOut128[29] , \nOut0_10[28] , \nOut1_16[9] , 
        \nScanOut21[3] , \nOut0_46[29] , \nOut1_48[19] , \nScanOut22[0] , 
        \nOut0_46[30] , \nOut1_23[11] , \nOut0_29[3] , \nScanOut123[3] , 
        \nScanOut43[9] , \nOut0_55[5] , \nOut1_56[21] , \nScanOut92[26] , 
        \nScanOut123[25] , \nScanOut100[14] , \nOut1_36[25] , \nOut0_38[15] , 
        \nOut0_58[11] , \nScanOut115[20] , \nOut1_43[15] , \nScanOut8[7] , 
        \nOut1_15[14] , \nOut1_60[24] , \nScanOut87[12] , \nScanOut69[27] , 
        \nOut1_15[27] , \nOut1_36[16] , \nOut0_56[6] , \nOut0_38[26] , 
        \nScanOut115[13] , \nOut1_43[26] , \nScanOut87[21] , \nOut1_10[7] , 
        \nOut1_23[22] , \nOut1_60[17] , \nScanOut92[15] , \nScanOut123[16] , 
        \nOut1_56[12] , \nOut0_58[22] , \nScanOut100[27] , \nOut1_13[4] , 
        \nOut0_31[1] , \nOut0_32[2] , \nOut0_1[27] , \nOut0_1[14] , 
        \nScanOut0[2] , \nOut0_4[22] , \nOut0_4[11] , \nOut1_5[0] , 
        \nOut1_6[3] , \nOut0_16[4] , \nScanOut39[1] , \nScanOut69[14] , 
        \nOut1_37[2] , \nScanOut78[11] , \nScanOut18[15] , \nOut1_32[27] , 
        \nOut1_47[17] , \nScanOut111[22] , \nOut0_49[27] , \nScanOut5[20] , 
        \nScanOut5[13] , \nOut1_11[25] , \nOut1_11[16] , \nScanOut83[10] , 
        \nOut0_15[7] , \nOut1_27[13] , \nOut0_29[23] , \nOut1_52[23] , 
        \nScanOut96[24] , \nScanOut127[27] , \nScanOut104[16] , 
        \nScanOut102[8] , \nScanOut18[26] , \nOut1_34[1] , \nScanOut79[3] , 
        \nOut1_27[20] , \nOut1_50[5] , \nOut1_53[6] , \nScanOut78[22] , 
        \nScanOut96[17] , \nScanOut127[14] , \nOut0_29[10] , \nOut1_52[10] , 
        \nScanOut104[25] , \nOut1_32[14] , \nOut0_49[14] , \nOut1_47[24] , 
        \nScanOut111[11] , \nScanOut83[23] , \nScanOut107[5] , \nOut0_13[9] , 
        \nScanOut104[6] , \nScanOut13[19] , \nOut0_14[19] , \nOut0_37[28] , 
        \nOut1_39[18] , \nOut0_42[18] , \nOut0_61[30] , \nOut0_61[29] , 
        \nScanOut119[9] , \nScanOut30[28] , \nOut0_37[31] , \nScanOut45[18] , 
        \nOut1_48[7] , \nOut1_55[8] , \nScanOut62[2] , \nScanOut66[30] , 
        \nScanOut66[29] , \nScanOut30[31] , \nScanOut61[1] , \nOut0_27[19] , 
        \nOut1_29[30] , \nOut1_29[29] , \nOut0_52[30] , \nOut0_52[29] , 
        \nScanOut55[0] , \nScanOut3[1] , \nScanOut87[6] , \nScanOut56[3] , 
        \nScanOut84[5] , \nOut1_61[9] , \nOut1_1[19] , \nScanOut0[25] , 
        \nScanOut0[16] , \nOut1_18[2] , \nScanOut20[19] , \nOut0_27[8] , 
        \nScanOut31[4] , \nScanOut32[7] , \nScanOut55[30] , \nScanOut76[18] , 
        \nScanOut55[29] , \nOut1_22[16] , \nOut0_39[4] , \nOut0_45[2] , 
        \nOut1_57[26] , \nScanOut93[21] , \nScanOut122[22] , \nScanOut101[13] , 
        \nOut1_37[22] , \nOut0_39[12] , \nOut0_59[16] , \nScanOut114[27] , 
        \nOut1_42[12] , \nScanOut81[8] , \nOut1_61[23] , \nOut1_5[31] , 
        \nOut1_14[13] , \nScanOut86[15] , \nOut1_5[28] , \nScanOut68[20] , 
        \nOut1_14[20] , \nOut1_37[11] , \nOut0_46[1] , \nOut0_39[21] , 
        \nScanOut114[14] , \nOut1_42[21] , \nScanOut86[26] , \nOut1_61[10] , 
        \nScanOut4[14] , \nOut0_5[2] , \nScanOut93[12] , \nOut0_6[1] , 
        \nOut0_21[6] , \nOut1_22[25] , \nScanOut122[11] , \nOut1_57[15] , 
        \nOut0_59[25] , \nScanOut101[20] , \nOut0_22[5] , \nScanOut34[9] , 
        \nScanOut128[5] , \nScanOut29[6] , \nScanOut68[13] , \nScanOut19[12] , 
        \nOut1_27[5] , \nScanOut79[16] , \nOut1_33[20] , \nOut1_39[9] , 
        \nOut1_46[10] , \nScanOut110[25] , \nOut0_48[20] , \nOut1_8[8] , 
        \nOut1_10[11] , \nScanOut82[17] , \nOut1_24[6] , \nOut1_26[14] , 
        \nOut0_28[24] , \nOut1_53[24] , \nScanOut97[23] , \nScanOut126[20] , 
        \nScanOut105[11] , \nScanOut19[21] , \nScanOut69[4] , \nOut1_40[2] , 
        \nOut1_43[1] , \nScanOut79[25] , \nOut0_62[7] , \nScanOut77[8] , 
        \nOut0_61[4] , \nScanOut97[10] , \nOut1_0[20] , \nOut1_0[13] , 
        \nScanOut4[27] , \nOut1_10[22] , \nOut1_26[27] , \nScanOut126[13] , 
        \nOut0_28[17] , \nOut1_53[17] , \nScanOut105[22] , \nOut1_33[13] , 
        \nOut0_48[13] , \nOut1_46[23] , \nScanOut110[16] , \nScanOut82[24] , 
        \nOut0_5[25] , \nOut0_5[16] , \nScanOut16[1] , \nScanOut24[31] , 
        \nScanOut24[28] , \nScanOut72[29] , \nScanOut51[18] , \nScanOut72[30] , 
        \nScanOut117[2] , \nScanOut15[2] , \nScanOut114[1] , \nOut1_22[8] , 
        \nOut0_23[31] , \nOut1_58[31] , \nOut1_58[0] , \nScanOut89[31] , 
        \nScanOut89[28] , \nScanOut71[6] , \nScanOut72[5] , \nOut0_23[28] , 
        \nOut1_58[28] , \nOut0_56[18] , \nOut1_11[31] , \nOut1_11[28] , 
        \nScanOut104[31] , \nScanOut104[28] , \nScanOut127[19] , 
        \nOut1_47[30] , \nOut0_49[19] , \nOut1_32[19] , \nOut1_47[29] , 
        \nOut1_50[8] , \nScanOut67[2] , \nScanOut64[1] , \nOut1_29[3] , 
        \nScanOut96[30] , \nScanOut96[29] , \nScanOut102[5] , \nOut1_0[0] , 
        \nOut1_3[3] , \nOut0_13[4] , \nScanOut13[14] , \nOut0_14[27] , 
        \nOut0_16[9] , \nScanOut18[18] , \nScanOut101[6] , \nOut0_22[22] , 
        \nOut0_37[16] , \nOut0_61[17] , \nScanOut88[11] , \nOut1_39[26] , 
        \nOut0_42[26] , \nOut1_56[6] , \nOut1_59[22] , \nScanOut25[11] , 
        \nScanOut50[21] , \nOut0_57[12] , \nOut1_55[5] , \nScanOut66[24] , 
        \nScanOut73[10] , \nScanOut30[25] , \nScanOut45[15] , \nOut0_57[21] , 
        \nOut1_59[11] , \nOut0_14[14] , \nOut0_22[11] , \nOut1_32[2] , 
        \nOut0_61[24] , \nScanOut88[22] , \nScanOut18[7] , \nOut0_37[25] , 
        \nOut1_39[15] , \nOut0_42[15] , \nScanOut119[4] , \nOut1_4[11] , 
        \nOut0_10[25] , \nOut0_10[7] , \nScanOut13[27] , \nScanOut107[8] , 
        \nScanOut30[16] , \nScanOut66[17] , \nOut1_15[7] , \nScanOut17[16] , 
        \nScanOut25[22] , \nOut1_31[1] , \nScanOut45[26] , \nScanOut50[12] , 
        \nScanOut62[26] , \nScanOut73[23] , \nScanOut21[13] , \nScanOut34[27] , 
        \nScanOut41[17] , \nScanOut54[23] , \nOut0_26[20] , \nOut0_34[1] , 
        \nScanOut77[12] , \nOut1_28[10] , \nOut0_53[10] , \nScanOut99[27] , 
        \nScanOut128[24] , \nOut0_10[16] , \nOut1_16[4] , \nOut0_33[14] , 
        \nOut0_46[24] , \nOut1_48[14] , \nScanOut17[25] , \nScanOut21[20] , 
        \nOut0_37[2] , \nScanOut54[10] , \nScanOut77[21] , \nScanOut34[14] , 
        \nScanOut46[9] , \nScanOut62[15] , \nScanOut89[0] , \nScanOut41[24] , 
        \nOut0_50[5] , \nScanOut58[5] , \nOut0_26[13] , \nOut1_28[23] , 
        \nOut0_33[27] , \nOut0_46[17] , \nOut1_48[27] , \nOut0_53[23] , 
        \nOut0_53[6] , \nScanOut99[14] , \nScanOut125[0] , \nScanOut128[17] , 
        \nOut1_13[9] , \nScanOut24[3] , \nScanOut69[19] , \nOut1_4[22] , 
        \nOut0_8[7] , \nScanOut27[0] , \nScanOut40[7] , \nScanOut92[18] , 
        \nScanOut126[3] , \nOut1_15[19] , \nOut1_36[31] , \nOut1_60[29] , 
        \nScanOut92[1] , \nScanOut100[19] , \nScanOut123[31] , 
        \nScanOut123[28] , \nOut1_36[28] , \nOut0_38[18] , \nScanOut91[2] , 
        \nOut1_43[18] , \nOut1_60[30] , \nOut0_48[7] , \nOut1_0[30] , 
        \nOut1_0[29] , \nOut1_0[9] , \nOut0_4[15] , \nOut0_22[18] , 
        \nScanOut43[4] , \nOut0_55[8] , \nOut0_57[28] , \nOut1_59[18] , 
        \nOut0_57[31] , \nScanOut104[2] , \nScanOut107[1] , \nOut0_4[26] , 
        \nOut1_31[8] , \nOut1_5[4] , \nOut0_15[3] , \nScanOut25[18] , 
        \nScanOut50[28] , \nScanOut61[5] , \nScanOut88[18] , \nScanOut62[6] , 
        \nOut1_48[3] , \nScanOut50[31] , \nScanOut73[19] , \nOut1_27[17] , 
        \nOut0_29[27] , \nOut1_34[5] , \nOut1_52[27] , \nScanOut104[12] , 
        \nScanOut96[20] , \nScanOut127[23] , \nScanOut5[17] , \nOut1_11[12] , 
        \nScanOut83[14] , \nOut1_32[23] , \nOut1_47[13] , \nScanOut111[26] , 
        \nOut0_49[23] , \nScanOut18[11] , \nScanOut1[15] , \nScanOut5[24] , 
        \nOut1_6[7] , \nScanOut78[15] , \nOut1_11[21] , \nOut0_16[0] , 
        \nOut1_37[6] , \nScanOut83[27] , \nScanOut8[3] , \nScanOut18[22] , 
        \nOut1_27[24] , \nOut1_32[10] , \nOut0_49[10] , \nOut1_47[20] , 
        \nScanOut111[15] , \nOut0_29[14] , \nOut1_52[14] , \nScanOut104[21] , 
        \nOut1_50[1] , \nScanOut96[13] , \nScanOut127[10] , \nOut1_53[2] , 
        \nScanOut64[8] , \nScanOut78[26] , \nOut0_56[2] , \nScanOut79[7] , 
        \nOut1_60[20] , \nScanOut69[23] , \nScanOut92[8] , \nOut1_15[10] , 
        \nScanOut87[16] , \nOut1_23[15] , \nOut1_36[21] , \nOut0_38[11] , 
        \nScanOut115[24] , \nOut1_43[11] , \nOut1_56[25] , \nScanOut100[10] , 
        \nOut0_58[15] , \nScanOut92[22] , \nScanOut123[21] , \nOut1_4[18] , 
        \nOut0_55[1] , \nScanOut69[10] , \nScanOut39[5] , \nOut0_0[24] , 
        \nOut0_0[17] , \nScanOut1[26] , \nOut1_10[3] , \nOut1_13[0] , 
        \nScanOut125[9] , \nScanOut27[9] , \nOut0_32[6] , \nOut1_15[23] , 
        \nOut1_23[26] , \nOut0_31[5] , \nOut1_56[16] , \nOut0_58[26] , 
        \nScanOut87[25] , \nScanOut92[11] , \nScanOut100[23] , 
        \nScanOut123[12] , \nOut1_60[13] , \nScanOut21[30] , \nScanOut21[29] , 
        \nOut1_36[12] , \nOut0_38[22] , \nScanOut115[17] , \nOut1_43[22] , 
        \nScanOut46[0] , \nScanOut89[9] , \nScanOut54[19] , \nScanOut77[31] , 
        \nScanOut77[28] , \nScanOut94[6] , \nScanOut97[5] , \nScanOut21[7] , 
        \nScanOut22[4] , \nOut0_29[7] , \nScanOut45[3] , \nScanOut123[7] , 
        \nOut0_34[8] , \nOut0_26[30] , \nOut0_26[29] , \nOut1_28[19] , 
        \nOut0_53[19] , \nScanOut120[4] , \nOut0_0[6] , \nOut0_3[5] , 
        \nOut1_5[21] , \nOut1_5[12] , \nOut0_6[8] , \nOut1_14[30] , 
        \nScanOut101[30] , \nScanOut122[18] , \nScanOut101[29] , 
        \nOut1_14[29] , \nOut1_37[18] , \nOut0_39[28] , \nOut1_42[28] , 
        \nScanOut34[0] , \nScanOut37[3] , \nOut0_39[31] , \nOut1_42[31] , 
        \nOut1_61[19] , \nScanOut5[6] , \nScanOut6[5] , \nScanOut53[7] , 
        \nOut0_58[4] , \nScanOut81[1] , \nScanOut93[31] , \nScanOut93[28] , 
        \nScanOut68[30] , \nScanOut82[2] , \nOut0_46[8] , \nScanOut50[4] , 
        \nScanOut68[29] , \nOut0_11[26] , \nOut0_27[1] , \nOut0_32[17] , 
        \nOut0_47[27] , \nOut1_49[17] , \nScanOut16[15] , \nScanOut20[10] , 
        \nOut0_27[23] , \nScanOut98[24] , \nOut1_29[13] , \nOut0_52[13] , 
        \nScanOut55[20] , \nScanOut76[11] , \nOut0_24[2] , \nScanOut35[24] , 
        \nScanOut40[14] , \nScanOut63[25] , \nOut1_1[23] , \nOut1_1[10] , 
        \nScanOut3[8] , \nOut0_11[15] , \nOut0_27[10] , \nOut1_29[20] , 
        \nScanOut98[17] , \nOut0_43[5] , \nOut0_52[20] , \nScanOut55[9] , 
        \nOut1_62[3] , \nOut0_32[24] , \nOut0_47[14] , \nOut1_49[24] , 
        \nScanOut48[6] , \nScanOut12[24] , \nScanOut12[17] , \nScanOut16[26] , 
        \nScanOut35[17] , \nScanOut99[3] , \nOut0_40[6] , \nScanOut40[27] , 
        \nOut1_61[0] , \nScanOut20[23] , \nScanOut63[16] , \nScanOut76[22] , 
        \nScanOut31[26] , \nScanOut44[16] , \nScanOut55[13] , \nOut1_58[9] , 
        \nScanOut67[27] , \nOut0_15[24] , \nOut0_23[21] , \nScanOut24[12] , 
        \nScanOut51[22] , \nScanOut72[13] , \nOut1_45[6] , \nOut1_58[21] , 
        \nOut0_36[15] , \nOut0_56[11] , \nOut1_38[25] , \nOut0_43[25] , 
        \nOut1_46[5] , \nScanOut16[8] , \nScanOut24[21] , \nOut0_60[14] , 
        \nScanOut72[20] , \nScanOut89[12] , \nScanOut51[11] , \nOut1_21[2] , 
        \nScanOut31[15] , \nScanOut44[25] , \nOut0_15[17] , \nOut0_36[26] , 
        \nOut1_38[16] , \nOut0_43[16] , \nScanOut67[14] , \nScanOut114[8] , 
        \nOut0_60[27] , \nScanOut109[7] , \nScanOut89[21] , \nScanOut19[31] , 
        \nOut1_22[1] , \nOut0_23[12] , \nOut0_56[22] , \nOut1_58[12] , 
        \nScanOut19[28] , \nScanOut10[6] , \nOut1_43[8] , \nScanOut74[2] , 
        \nScanOut77[1] , \nScanOut97[19] , \nScanOut111[5] , \nOut0_2[8] , 
        \nScanOut2[19] , \nOut0_8[24] , \nOut1_8[1] , \nOut1_10[18] , 
        \nOut0_18[6] , \nOut1_46[19] , \nScanOut105[18] , \nScanOut126[29] , 
        \nScanOut112[6] , \nScanOut126[30] , \nOut0_48[29] , \nOut1_33[30] , 
        \nOut1_33[29] , \nOut1_39[0] , \nOut0_48[30] , \nScanOut13[5] , 
        \nOut1_20[19] , \nOut1_55[30] , \nScanOut73[1] , \nOut1_55[29] , 
        \nOut1_59[4] , \nScanOut116[28] , \nOut0_3[31] , \nOut0_3[28] , 
        \nOut1_7[27] , \nScanOut116[31] , \nOut1_7[14] , \nOut0_8[17] , 
        \nOut1_47[8] , \nScanOut70[2] , \nScanOut84[30] , \nScanOut84[29] , 
        \nScanOut116[6] , \nScanOut14[6] , \nScanOut17[5] , \nScanOut29[30] , 
        \nScanOut29[29] , \nScanOut115[5] , \nScanOut9[26] , \nOut0_30[22] , 
        \nOut0_45[12] , \nOut0_13[13] , \nScanOut14[20] , \nScanOut22[25] , 
        \nOut0_25[16] , \nOut1_42[5] , \nOut0_50[26] , \nOut0_63[3] , 
        \nScanOut108[23] , \nScanOut68[0] , \nScanOut74[24] , \nScanOut37[11] , 
        \nScanOut57[15] , \nOut1_41[6] , \nScanOut42[21] , \nOut0_60[0] , 
        \nScanOut61[10] , \nOut0_4[6] , \nScanOut9[15] , \nOut0_25[25] , 
        \nScanOut110[8] , \nOut1_26[1] , \nOut0_30[11] , \nOut0_50[15] , 
        \nScanOut108[10] , \nOut0_45[21] , \nScanOut10[22] , \nScanOut12[8] , 
        \nOut0_13[20] , \nScanOut14[13] , \nScanOut37[22] , \nScanOut42[12] , 
        \nScanOut61[23] , \nScanOut74[17] , \nOut0_20[2] , \nScanOut22[16] , 
        \nOut1_25[2] , \nScanOut57[26] , \nScanOut33[13] , \nScanOut46[23] , 
        \nScanOut26[27] , \nScanOut65[12] , \nScanOut70[26] , \nScanOut53[17] , 
        \nOut0_7[19] , \nOut0_7[5] , \nScanOut7[8] , \nOut0_17[11] , 
        \nOut1_19[21] , \nOut0_21[14] , \nScanOut28[2] , \nOut0_54[24] , 
        \nOut0_23[1] , \nOut0_34[20] , \nOut0_41[10] , \nScanOut119[15] , 
        \nOut0_62[21] , \nOut0_59[9] , \nOut1_8[30] , \nScanOut26[14] , 
        \nOut0_44[6] , \nScanOut53[24] , \nScanOut70[15] , \nScanOut46[10] , 
        \nOut1_8[29] , \nScanOut33[20] , \nScanOut10[11] , \nScanOut65[21] , 
        \nOut0_17[22] , \nOut0_34[13] , \nOut0_41[23] , \nOut0_47[5] , 
        \nScanOut51[9] , \nScanOut119[26] , \nOut1_19[12] , \nOut0_21[27] , 
        \nOut0_62[12] , \nScanOut30[0] , \nOut0_54[17] , \nScanOut58[31] , 
        \nOut1_3[25] , \nScanOut58[28] , \nOut1_19[6] , \nScanOut33[3] , 
        \nOut0_38[0] , \nScanOut80[18] , \nScanOut86[2] , \nOut1_1[4] , 
        \nScanOut1[6] , \nOut1_3[16] , \nOut1_2[7] , \nScanOut2[5] , 
        \nScanOut6[31] , \nOut1_24[31] , \nOut0_42[8] , \nScanOut54[4] , 
        \nScanOut57[7] , \nOut1_24[28] , \nScanOut85[1] , \nOut1_51[18] , 
        \nOut0_6[20] , \nScanOut6[28] , \nScanOut112[19] , \nScanOut93[5] , 
        \nOut0_6[13] , \nOut1_9[23] , \nOut0_16[31] , \nOut0_16[28] , 
        \nOut1_18[18] , \nOut0_40[30] , \nOut0_63[18] , \nOut0_35[19] , 
        \nScanOut41[3] , \nOut0_40[29] , \nScanOut42[0] , \nScanOut25[7] , 
        \nOut0_49[3] , \nScanOut90[6] , \nScanOut38[8] , \nScanOut7[22] , 
        \nOut0_9[3] , \nOut1_9[10] , \nScanOut11[28] , \nScanOut124[4] , 
        \nScanOut127[7] , \nScanOut47[30] , \nScanOut64[18] , \nScanOut11[31] , 
        \nOut1_13[27] , \nOut1_25[22] , \nScanOut26[4] , \nScanOut32[19] , 
        \nOut0_30[8] , \nScanOut47[29] , \nOut1_50[12] , \nScanOut106[27] , 
        \nScanOut94[15] , \nScanOut125[16] , \nScanOut81[21] , \nScanOut7[11] , 
        \nOut1_14[3] , \nScanOut23[9] , \nOut1_30[16] , \nScanOut39[15] , 
        \nOut1_45[26] , \nOut0_51[1] , \nScanOut88[4] , \nScanOut113[13] , 
        \nOut0_52[2] , \nScanOut59[1] , \nScanOut59[11] , \nScanOut96[8] , 
        \nOut0_35[5] , \nOut1_13[14] , \nOut1_17[0] , \nOut1_25[11] , 
        \nOut1_30[25] , \nOut1_45[15] , \nScanOut81[12] , \nScanOut113[20] , 
        \nOut1_50[21] , \nScanOut106[14] , \nScanOut39[26] , \nScanOut59[22] , 
        \nScanOut94[26] , \nScanOut125[25] , \nScanOut121[9] , 
        \nScanOut28[23] , \nOut0_36[6] , \nScanOut3[20] , \nOut0_11[3] , 
        \nOut0_12[0] , \nScanOut19[3] , \nScanOut48[27] , \nScanOut118[0] , 
        \nOut1_33[6] , \nOut1_17[25] , \nOut1_30[5] , \nOut1_62[15] , 
        \nScanOut85[23] , \nOut0_19[15] , \nOut1_21[20] , \nOut1_34[14] , 
        \nOut1_41[24] , \nScanOut117[11] , \nOut1_54[10] , \nScanOut102[25] , 
        \nScanOut90[17] , \nOut0_2[22] , \nScanOut3[13] , \nOut1_21[13] , 
        \nScanOut28[10] , \nScanOut48[14] , \nOut1_57[2] , \nScanOut60[8] , 
        \nScanOut121[14] , \nOut1_54[23] , \nScanOut102[16] , \nOut1_62[26] , 
        \nScanOut90[24] , \nScanOut121[27] , \nOut1_4[9] , \nOut1_17[16] , 
        \nOut0_19[26] , \nOut1_28[7] , \nOut1_34[27] , \nOut1_41[17] , 
        \nScanOut85[10] , \nScanOut117[22] , \nOut1_54[1] , \nScanOut103[1] , 
        \nScanOut15[19] , \nScanOut36[31] , \nScanOut60[29] , \nOut1_35[8] , 
        \nScanOut36[28] , \nScanOut43[18] , \nScanOut60[30] , \nScanOut100[2] , 
        \nOut0_2[18] , \nOut0_2[11] , \nScanOut66[6] , \nOut1_2[26] , 
        \nScanOut7[18] , \nOut0_12[19] , \nOut0_31[31] , \nScanOut23[0] , 
        \nOut0_31[28] , \nOut0_44[18] , \nScanOut65[5] , \nScanOut109[30] , 
        \nScanOut109[29] , \nOut1_25[18] , \nOut1_50[28] , \nScanOut122[3] , 
        \nOut1_50[31] , \nOut0_28[3] , \nScanOut113[30] , \nScanOut113[29] , 
        \nOut1_2[15] , \nOut1_17[9] , \nScanOut20[3] , \nScanOut121[0] , 
        \nScanOut44[7] , \nScanOut47[4] , \nScanOut81[31] , \nScanOut81[28] , 
        \nScanOut95[2] , \nOut0_51[8] , \nScanOut59[18] , \nOut0_6[30] , 
        \nOut1_9[19] , \nScanOut11[21] , \nOut1_12[4] , \nOut0_16[12] , 
        \nOut1_18[22] , \nScanOut59[8] , \nScanOut96[1] , \nOut0_63[22] , 
        \nOut0_20[17] , \nOut0_35[23] , \nOut0_40[13] , \nOut0_55[27] , 
        \nScanOut118[16] , \nScanOut27[24] , \nOut0_33[2] , \nScanOut38[1] , 
        \nScanOut52[14] , \nScanOut71[25] , \nOut1_11[7] , \nScanOut32[10] , 
        \nScanOut64[11] , \nScanOut47[20] , \nOut0_30[1] , \nOut0_6[29] , 
        \nScanOut9[7] , \nOut0_20[24] , \nOut0_55[14] , \nScanOut11[12] , 
        \nOut0_16[21] , \nOut1_18[11] , \nOut0_35[10] , \nOut0_63[11] , 
        \nOut0_40[20] , \nOut0_57[6] , \nScanOut118[25] , \nScanOut64[22] , 
        \nScanOut15[23] , \nScanOut27[17] , \nScanOut32[23] , \nScanOut47[13] , 
        \nScanOut42[9] , \nScanOut52[27] , \nOut0_54[5] , \nScanOut71[16] , 
        \nScanOut23[26] , \nScanOut36[12] , \nScanOut60[13] , \nScanOut43[22] , 
        \nOut1_51[5] , \nScanOut56[16] , \nScanOut75[27] , \nScanOut78[3] , 
        \nScanOut8[25] , \nOut0_24[15] , \nOut0_51[25] , \nOut1_52[6] , 
        \nScanOut109[20] , \nOut0_12[10] , \nOut0_31[21] , \nOut0_44[11] , 
        \nScanOut2[23] , \nOut0_3[21] , \nScanOut3[30] , \nScanOut3[29] , 
        \nOut1_4[0] , \nOut1_6[24] , \nOut1_7[3] , \nScanOut8[16] , 
        \nOut0_14[7] , \nScanOut56[25] , \nScanOut103[8] , \nScanOut15[10] , 
        \nScanOut23[15] , \nOut1_35[1] , \nScanOut60[20] , \nScanOut75[14] , 
        \nScanOut36[21] , \nScanOut43[11] , \nOut0_12[23] , \nOut0_17[4] , 
        \nOut0_31[12] , \nOut0_24[26] , \nOut1_36[2] , \nOut0_44[22] , 
        \nOut0_51[16] , \nScanOut109[13] , \nScanOut28[19] , \nScanOut60[1] , 
        \nOut1_6[17] , \nOut0_9[27] , \nOut1_49[7] , \nScanOut85[19] , 
        \nOut1_54[8] , \nScanOut63[2] , \nOut0_9[14] , \nOut0_12[9] , 
        \nScanOut105[6] , \nScanOut118[9] , \nOut1_21[30] , \nOut1_21[29] , 
        \nOut1_54[19] , \nScanOut106[5] , \nScanOut117[18] , \nOut0_3[12] , 
        \nOut1_9[5] , \nScanOut11[2] , \nScanOut110[1] , \nOut0_13[30] , 
        \nOut0_13[29] , \nOut1_26[8] , \nOut0_30[18] , \nOut0_45[28] , 
        \nOut0_45[31] , \nScanOut108[19] , \nScanOut12[1] , \nOut0_19[2] , 
        \nOut1_38[4] , \nScanOut75[6] , \nScanOut113[2] , \nScanOut14[30] , 
        \nScanOut68[9] , \nScanOut14[29] , \nScanOut37[18] , \nScanOut42[28] , 
        \nScanOut76[5] , \nOut0_60[9] , \nOut1_16[26] , \nOut1_20[23] , 
        \nScanOut42[31] , \nScanOut61[19] , \nScanOut91[14] , 
        \nScanOut120[17] , \nOut1_35[17] , \nOut1_55[13] , \nScanOut103[26] , 
        \nOut1_40[27] , \nScanOut116[12] , \nOut1_63[16] , \nScanOut84[20] , 
        \nOut0_18[16] , \nOut1_20[6] , \nOut1_23[5] , \nScanOut29[20] , 
        \nScanOut49[24] , \nScanOut108[3] , \nScanOut73[8] , \nOut0_1[2] , 
        \nOut0_2[1] , \nScanOut2[10] , \nOut1_35[24] , \nOut1_40[14] , 
        \nOut1_44[2] , \nScanOut116[21] , \nOut1_63[25] , \nScanOut6[21] , 
        \nOut1_12[24] , \nOut1_16[15] , \nOut0_18[25] , \nOut1_20[10] , 
        \nOut1_55[20] , \nScanOut84[13] , \nScanOut91[27] , \nScanOut120[24] , 
        \nScanOut103[15] , \nScanOut29[13] , \nOut1_31[15] , \nScanOut38[16] , 
        \nOut1_47[1] , \nScanOut49[17] , \nScanOut49[2] , \nScanOut58[12] , 
        \nOut0_41[2] , \nOut0_42[1] , \nOut1_63[7] , \nScanOut98[7] , 
        \nOut1_60[4] , \nOut1_44[25] , \nScanOut112[10] , \nScanOut80[22] , 
        \nOut1_24[21] , \nScanOut85[8] , \nScanOut95[16] , \nScanOut124[15] , 
        \nOut0_26[5] , \nScanOut30[9] , \nOut1_51[11] , \nScanOut107[24] , 
        \nScanOut38[25] , \nScanOut6[12] , \nOut1_24[12] , \nOut1_51[22] , 
        \nScanOut58[21] , \nScanOut95[25] , \nScanOut124[26] , 
        \nScanOut107[17] , \nOut1_31[26] , \nOut1_44[16] , \nScanOut112[23] , 
        \nOut0_38[9] , \nOut1_12[17] , \nOut1_1[0] , \nOut0_2[26] , 
        \nScanOut4[2] , \nOut0_7[23] , \nScanOut7[1] , \nOut0_25[6] , 
        \nScanOut80[11] , \nOut1_8[20] , \nScanOut33[29] , \nScanOut46[19] , 
        \nOut0_59[0] , \nScanOut80[5] , \nScanOut65[31] , \nScanOut65[28] , 
        \nScanOut10[18] , \nScanOut33[30] , \nScanOut51[0] , \nScanOut52[3] , 
        \nOut0_7[10] , \nOut1_8[13] , \nScanOut36[7] , \nScanOut83[6] , 
        \nOut0_17[18] , \nOut1_19[31] , \nOut1_19[28] , \nOut0_34[29] , 
        \nOut0_41[19] , \nOut0_62[31] , \nOut0_34[30] , \nOut0_62[28] , 
        \nOut0_23[8] , \nScanOut35[4] , \nOut0_2[15] , \nScanOut8[31] , 
        \nOut0_17[9] , \nScanOut100[6] , \nScanOut23[18] , \nScanOut56[31] , 
        \nScanOut56[28] , \nScanOut75[19] , \nOut0_24[18] , \nOut1_28[3] , 
        \nOut0_51[31] , \nScanOut103[5] , \nOut0_51[28] , \nScanOut65[1] , 
        \nScanOut8[28] , \nOut1_51[8] , \nScanOut66[2] , \nScanOut90[13] , 
        \nScanOut1[2] , \nOut1_2[18] , \nOut1_2[3] , \nScanOut3[24] , 
        \nOut1_17[21] , \nOut1_21[24] , \nScanOut121[10] , \nOut1_34[10] , 
        \nOut1_54[14] , \nScanOut102[21] , \nOut1_41[20] , \nScanOut106[8] , 
        \nScanOut117[15] , \nScanOut85[27] , \nOut0_9[19] , \nOut0_19[11] , 
        \nOut1_62[11] , \nOut0_11[7] , \nOut0_12[4] , \nOut1_30[1] , 
        \nScanOut19[7] , \nOut1_33[2] , \nScanOut118[4] , \nScanOut48[23] , 
        \nScanOut3[17] , \nScanOut28[27] , \nOut1_34[23] , \nOut1_41[13] , 
        \nOut1_54[5] , \nScanOut117[26] , \nOut1_6[30] , \nOut1_17[12] , 
        \nOut0_19[22] , \nOut1_62[22] , \nOut1_21[17] , \nOut1_54[27] , 
        \nScanOut85[14] , \nScanOut90[20] , \nScanOut121[23] , 
        \nScanOut102[12] , \nScanOut28[14] , \nOut1_6[29] , \nScanOut48[10] , 
        \nScanOut39[11] , \nOut1_57[6] , \nScanOut59[15] , \nScanOut59[5] , 
        \nScanOut2[1] , \nOut1_3[21] , \nOut0_6[24] , \nScanOut7[26] , 
        \nOut1_13[23] , \nOut1_30[12] , \nScanOut47[9] , \nOut0_52[6] , 
        \nScanOut88[0] , \nOut0_51[5] , \nOut1_45[22] , \nScanOut113[17] , 
        \nScanOut81[25] , \nScanOut7[15] , \nOut1_17[4] , \nOut1_25[26] , 
        \nScanOut94[11] , \nScanOut125[12] , \nOut1_50[16] , \nScanOut106[23] , 
        \nOut1_25[15] , \nOut0_36[2] , \nScanOut39[22] , \nOut1_50[25] , 
        \nScanOut59[26] , \nScanOut94[22] , \nScanOut125[21] , 
        \nScanOut106[10] , \nOut1_30[21] , \nOut1_45[11] , \nScanOut113[24] , 
        \nOut1_9[27] , \nOut1_13[10] , \nOut1_14[7] , \nScanOut81[16] , 
        \nOut0_35[1] , \nOut0_49[7] , \nScanOut90[2] , \nOut0_20[30] , 
        \nScanOut42[4] , \nOut0_54[8] , \nOut0_20[29] , \nScanOut41[7] , 
        \nOut0_55[19] , \nScanOut118[31] , \nScanOut118[28] , \nOut0_6[17] , 
        \nOut0_9[7] , \nOut1_9[14] , \nScanOut26[0] , \nScanOut27[30] , 
        \nScanOut93[1] , \nScanOut27[29] , \nScanOut71[28] , \nScanOut52[19] , 
        \nScanOut71[31] , \nScanOut124[0] , \nScanOut127[3] , \nOut1_12[9] , 
        \nScanOut25[3] , \nOut1_19[2] , \nScanOut33[7] , \nScanOut95[31] , 
        \nScanOut95[28] , \nOut0_38[4] , \nOut1_12[30] , \nOut1_12[29] , 
        \nOut0_26[8] , \nScanOut30[4] , \nScanOut38[31] , \nScanOut38[28] , 
        \nOut1_31[18] , \nOut1_44[31] , \nOut1_44[28] , \nScanOut54[0] , 
        \nScanOut57[3] , \nScanOut85[5] , \nScanOut107[30] , \nScanOut107[29] , 
        \nScanOut124[18] , \nOut1_60[9] , \nOut1_3[12] , \nOut0_4[2] , 
        \nOut0_7[1] , \nOut0_17[15] , \nOut1_19[25] , \nScanOut86[6] , 
        \nOut0_62[25] , \nOut0_21[10] , \nOut0_34[24] , \nOut0_41[14] , 
        \nScanOut35[9] , \nScanOut119[11] , \nOut0_54[20] , \nOut0_23[5] , 
        \nScanOut28[6] , \nOut1_7[23] , \nOut1_9[8] , \nScanOut9[22] , 
        \nScanOut10[26] , \nScanOut26[23] , \nScanOut53[13] , \nScanOut70[22] , 
        \nScanOut10[15] , \nOut0_17[26] , \nOut0_20[6] , \nScanOut33[17] , 
        \nScanOut65[16] , \nScanOut46[27] , \nOut0_21[23] , \nOut0_54[13] , 
        \nOut1_19[16] , \nOut0_34[17] , \nOut0_62[16] , \nOut0_41[27] , 
        \nOut0_47[1] , \nScanOut119[22] , \nScanOut65[25] , \nScanOut14[24] , 
        \nScanOut26[10] , \nScanOut33[24] , \nScanOut46[14] , \nOut0_44[2] , 
        \nScanOut53[20] , \nScanOut70[11] , \nScanOut80[8] , \nScanOut22[21] , 
        \nScanOut37[15] , \nScanOut61[14] , \nOut1_41[2] , \nScanOut42[25] , 
        \nScanOut76[8] , \nOut0_60[4] , \nOut0_25[12] , \nOut0_50[22] , 
        \nScanOut57[11] , \nScanOut68[4] , \nScanOut74[20] , \nOut1_42[1] , 
        \nScanOut108[27] , \nOut0_63[7] , \nOut0_13[17] , \nScanOut22[12] , 
        \nOut1_25[6] , \nOut0_30[26] , \nOut0_45[16] , \nOut1_38[9] , 
        \nScanOut57[22] , \nScanOut9[11] , \nScanOut14[17] , \nScanOut61[27] , 
        \nScanOut74[13] , \nScanOut37[26] , \nScanOut42[16] , \nOut0_13[24] , 
        \nOut0_25[21] , \nOut1_26[5] , \nOut0_30[15] , \nOut0_45[25] , 
        \nOut0_50[11] , \nScanOut108[14] , \nScanOut70[6] , \nOut1_7[10] , 
        \nOut0_8[20] , \nOut1_16[18] , \nOut0_18[28] , \nOut1_63[28] , 
        \nOut0_18[31] , \nOut1_35[30] , \nOut1_40[19] , \nOut1_63[31] , 
        \nOut1_35[29] , \nOut1_59[0] , \nScanOut73[5] , \nScanOut103[18] , 
        \nScanOut120[30] , \nScanOut120[29] , \nOut0_8[13] , \nScanOut14[2] , 
        \nScanOut49[30] , \nScanOut49[29] , \nScanOut115[1] , \nScanOut17[1] , 
        \nOut1_23[8] , \nOut0_1[6] , \nScanOut2[8] , \nScanOut4[6] , 
        \nScanOut83[2] , \nScanOut91[19] , \nScanOut116[2] , \nScanOut6[25] , 
        \nOut0_7[27] , \nOut0_7[14] , \nScanOut7[5] , \nOut1_8[24] , 
        \nScanOut26[19] , \nOut0_47[8] , \nScanOut51[4] , \nScanOut52[7] , 
        \nScanOut53[29] , \nScanOut53[30] , \nScanOut70[18] , \nOut0_59[4] , 
        \nScanOut80[1] , \nOut0_21[19] , \nScanOut35[0] , \nOut0_54[29] , 
        \nOut0_54[30] , \nScanOut119[18] , \nOut0_7[8] , \nOut1_8[17] , 
        \nOut1_12[20] , \nOut1_24[25] , \nScanOut36[3] , \nOut1_51[15] , 
        \nScanOut107[20] , \nScanOut95[12] , \nScanOut124[11] , 
        \nScanOut80[26] , \nOut1_31[11] , \nOut1_44[21] , \nScanOut6[16] , 
        \nOut0_25[2] , \nScanOut38[12] , \nOut0_41[6] , \nScanOut98[3] , 
        \nScanOut112[14] , \nOut0_42[5] , \nScanOut54[9] , \nOut1_60[0] , 
        \nScanOut49[6] , \nOut1_63[3] , \nScanOut58[16] , \nOut0_2[5] , 
        \nOut1_12[13] , \nOut1_24[16] , \nOut1_31[22] , \nOut1_44[12] , 
        \nScanOut80[15] , \nScanOut112[27] , \nOut1_51[26] , \nScanOut107[13] , 
        \nScanOut58[25] , \nScanOut95[21] , \nScanOut124[22] , \nOut1_3[31] , 
        \nOut1_3[28] , \nOut1_7[19] , \nOut0_26[1] , \nScanOut38[21] , 
        \nScanOut29[24] , \nScanOut115[8] , \nOut1_23[1] , \nScanOut49[20] , 
        \nScanOut108[7] , \nScanOut2[27] , \nOut1_16[22] , \nScanOut17[8] , 
        \nOut1_20[2] , \nScanOut84[24] , \nScanOut2[14] , \nOut0_18[12] , 
        \nOut1_63[12] , \nOut1_20[27] , \nOut1_35[13] , \nOut1_40[23] , 
        \nScanOut116[16] , \nOut1_20[14] , \nScanOut29[17] , \nOut1_47[5] , 
        \nOut1_55[17] , \nScanOut103[22] , \nScanOut91[10] , \nScanOut120[13] , 
        \nScanOut49[13] , \nOut1_55[24] , \nScanOut103[11] , \nScanOut91[23] , 
        \nScanOut120[20] , \nOut0_8[30] , \nOut1_16[11] , \nOut0_18[21] , 
        \nOut1_63[21] , \nOut1_35[20] , \nOut1_40[10] , \nScanOut84[17] , 
        \nScanOut116[25] , \nOut1_59[9] , \nOut0_8[29] , \nOut1_1[9] , 
        \nOut0_3[25] , \nOut1_9[1] , \nScanOut12[5] , \nOut0_19[6] , 
        \nOut1_44[6] , \nScanOut113[6] , \nOut1_38[0] , \nScanOut9[18] , 
        \nOut0_25[31] , \nOut0_25[28] , \nOut0_50[18] , \nScanOut11[6] , 
        \nScanOut110[5] , \nOut0_3[16] , \nScanOut22[31] , \nScanOut22[28] , 
        \nScanOut57[18] , \nScanOut74[30] , \nScanOut74[29] , \nScanOut76[1] , 
        \nOut1_6[20] , \nOut0_9[23] , \nOut1_42[8] , \nScanOut75[2] , 
        \nScanOut48[19] , \nOut1_49[3] , \nScanOut63[6] , \nScanOut90[30] , 
        \nScanOut90[29] , \nOut1_17[31] , \nOut1_34[19] , \nScanOut60[5] , 
        \nOut1_17[28] , \nOut1_41[29] , \nScanOut106[1] , \nOut0_19[18] , 
        \nOut1_41[30] , \nOut1_62[18] , \nOut1_4[4] , \nOut1_6[13] , 
        \nOut0_9[10] , \nScanOut102[31] , \nScanOut102[28] , \nScanOut121[19] , 
        \nOut1_30[8] , \nScanOut105[2] , \nOut1_7[7] , \nScanOut8[21] , 
        \nOut0_31[25] , \nOut0_44[15] , \nOut0_12[14] , \nScanOut15[27] , 
        \nScanOut23[22] , \nOut0_24[11] , \nOut0_51[21] , \nScanOut65[8] , 
        \nOut1_52[2] , \nScanOut109[24] , \nScanOut75[23] , \nScanOut78[7] , 
        \nScanOut36[16] , \nScanOut56[12] , \nScanOut43[26] , \nOut1_51[1] , 
        \nScanOut60[17] , \nScanOut8[12] , \nOut0_17[0] , \nOut0_24[22] , 
        \nOut0_31[16] , \nOut0_51[12] , \nScanOut109[17] , \nOut1_36[6] , 
        \nOut0_44[26] , \nOut0_12[27] , \nOut0_14[3] , \nScanOut15[14] , 
        \nScanOut36[25] , \nScanOut43[15] , \nScanOut60[24] , \nScanOut56[21] , 
        \nScanOut75[10] , \nScanOut23[11] , \nOut1_35[5] , \nOut1_2[22] , 
        \nScanOut9[3] , \nOut1_11[3] , \nScanOut26[9] , \nScanOut32[14] , 
        \nScanOut47[24] , \nScanOut11[25] , \nOut0_30[5] , \nScanOut11[16] , 
        \nOut1_12[0] , \nScanOut27[20] , \nScanOut64[15] , \nScanOut71[21] , 
        \nScanOut38[5] , \nScanOut52[10] , \nOut0_55[23] , \nScanOut124[9] , 
        \nOut0_16[16] , \nOut1_18[26] , \nOut0_20[13] , \nOut0_33[6] , 
        \nOut0_35[27] , \nOut0_40[17] , \nScanOut118[12] , \nOut0_63[26] , 
        \nScanOut27[13] , \nScanOut52[23] , \nScanOut71[12] , \nOut0_54[1] , 
        \nScanOut32[27] , \nScanOut47[17] , \nScanOut64[26] , \nOut0_16[25] , 
        \nOut0_35[14] , \nOut0_40[24] , \nOut0_57[2] , \nScanOut118[21] , 
        \nOut1_18[15] , \nOut0_20[20] , \nOut0_63[15] , \nOut0_55[10] , 
        \nScanOut20[7] , \nScanOut93[8] , \nScanOut121[4] , \nOut1_2[11] , 
        \nOut1_13[19] , \nOut0_28[7] , \nOut1_30[28] , \nOut1_45[18] , 
        \nScanOut23[4] , \nOut1_30[31] , \nScanOut106[19] , \nScanOut125[31] , 
        \nScanOut125[28] , \nScanOut122[7] , \nOut0_35[8] , \nScanOut39[18] , 
        \nScanOut96[5] , \nOut1_2[8] , \nOut1_6[22] , \nScanOut44[3] , 
        \nScanOut47[0] , \nScanOut88[9] , \nScanOut60[7] , \nScanOut94[18] , 
        \nScanOut95[6] , \nOut1_6[11] , \nOut0_9[21] , \nOut1_17[19] , 
        \nOut0_19[30] , \nOut1_34[28] , \nOut1_41[18] , \nOut1_49[1] , 
        \nOut1_62[30] , \nOut1_34[31] , \nOut0_19[29] , \nOut1_62[29] , 
        \nScanOut63[4] , \nScanOut102[19] , \nScanOut121[28] , 
        \nScanOut121[31] , \nScanOut48[31] , \nScanOut48[28] , \nOut1_4[6] , 
        \nScanOut8[23] , \nOut0_9[12] , \nOut1_33[9] , \nScanOut105[0] , 
        \nScanOut15[25] , \nScanOut36[14] , \nScanOut43[24] , \nScanOut90[18] , 
        \nScanOut106[3] , \nOut1_51[3] , \nScanOut60[15] , \nScanOut66[9] , 
        \nScanOut23[20] , \nScanOut56[10] , \nScanOut75[21] , \nOut0_24[13] , 
        \nOut1_52[0] , \nScanOut78[5] , \nScanOut109[26] , \nOut0_31[27] , 
        \nOut0_51[23] , \nOut0_44[17] , \nOut0_12[16] , \nOut1_28[8] , 
        \nOut0_1[4] , \nScanOut1[9] , \nOut1_2[20] , \nOut1_7[5] , 
        \nScanOut8[10] , \nOut0_14[1] , \nOut1_35[7] , \nScanOut75[12] , 
        \nScanOut15[16] , \nScanOut23[13] , \nScanOut36[27] , \nScanOut56[23] , 
        \nScanOut43[17] , \nOut0_17[2] , \nOut1_36[4] , \nOut0_44[24] , 
        \nScanOut60[26] , \nOut0_31[14] , \nOut0_12[25] , \nOut0_24[20] , 
        \nOut0_51[10] , \nScanOut109[15] , \nScanOut9[1] , \nOut1_11[1] , 
        \nOut1_12[2] , \nOut0_16[14] , \nOut0_35[25] , \nScanOut118[10] , 
        \nOut0_40[15] , \nOut1_18[24] , \nOut0_20[11] , \nOut0_33[4] , 
        \nOut0_63[24] , \nScanOut25[8] , \nOut0_55[21] , \nScanOut27[22] , 
        \nScanOut38[7] , \nScanOut52[12] , \nScanOut71[23] , \nScanOut127[8] , 
        \nOut0_30[7] , \nScanOut47[26] , \nScanOut11[27] , \nScanOut32[16] , 
        \nScanOut64[17] , \nOut0_55[12] , \nScanOut11[14] , \nOut0_16[27] , 
        \nOut1_18[17] , \nOut0_20[22] , \nOut0_35[16] , \nOut0_40[26] , 
        \nOut0_57[0] , \nScanOut118[23] , \nOut0_63[17] , \nScanOut32[25] , 
        \nScanOut47[15] , \nScanOut23[6] , \nScanOut27[11] , \nOut0_54[3] , 
        \nScanOut64[24] , \nScanOut71[10] , \nScanOut52[21] , \nScanOut90[9] , 
        \nOut0_28[5] , \nScanOut94[30] , \nScanOut94[29] , \nScanOut122[5] , 
        \nScanOut39[30] , \nScanOut39[29] , \nScanOut121[6] , \nOut1_2[13] , 
        \nOut1_13[31] , \nScanOut20[5] , \nOut0_36[9] , \nOut1_45[29] , 
        \nOut1_13[28] , \nOut1_30[19] , \nOut1_45[30] , \nScanOut44[1] , 
        \nScanOut47[2] , \nScanOut95[4] , \nScanOut106[31] , \nScanOut125[19] , 
        \nScanOut106[28] , \nScanOut96[7] , \nOut0_4[9] , \nScanOut4[4] , 
        \nScanOut7[7] , \nOut1_8[26] , \nOut0_59[6] , \nScanOut80[3] , 
        \nOut0_21[31] , \nOut0_21[28] , \nOut0_44[9] , \nScanOut52[5] , 
        \nOut0_54[18] , \nScanOut51[6] , \nScanOut119[30] , \nScanOut119[29] , 
        \nOut0_7[25] , \nOut1_8[15] , \nScanOut26[31] , \nScanOut26[28] , 
        \nScanOut53[18] , \nScanOut83[0] , \nScanOut70[30] , \nScanOut70[29] , 
        \nScanOut36[1] , \nOut0_7[16] , \nScanOut35[2] , \nOut0_2[7] , 
        \nOut1_3[19] , \nScanOut58[14] , \nScanOut6[27] , \nScanOut38[10] , 
        \nOut0_41[4] , \nOut0_42[7] , \nScanOut49[4] , \nOut1_63[1] , 
        \nOut1_60[2] , \nScanOut57[8] , \nScanOut98[1] , \nOut1_12[22] , 
        \nOut1_24[27] , \nOut1_31[13] , \nOut1_44[23] , \nScanOut80[24] , 
        \nScanOut112[16] , \nOut1_51[17] , \nScanOut107[22] , \nOut0_26[3] , 
        \nScanOut95[10] , \nScanOut124[13] , \nScanOut38[23] , 
        \nScanOut58[27] , \nOut1_12[11] , \nOut1_24[14] , \nOut1_51[24] , 
        \nScanOut107[11] , \nScanOut95[23] , \nScanOut124[20] , 
        \nScanOut2[25] , \nScanOut6[14] , \nScanOut80[17] , \nOut1_19[9] , 
        \nOut1_20[25] , \nOut0_25[0] , \nOut1_31[20] , \nOut1_44[10] , 
        \nScanOut112[25] , \nOut1_55[15] , \nScanOut103[20] , \nOut1_63[10] , 
        \nScanOut91[12] , \nScanOut120[11] , \nOut0_8[18] , \nOut1_16[20] , 
        \nOut0_18[10] , \nOut1_20[0] , \nOut1_35[11] , \nOut1_40[21] , 
        \nScanOut84[26] , \nScanOut116[14] , \nScanOut116[9] , \nScanOut14[9] , 
        \nOut1_23[3] , \nScanOut29[26] , \nScanOut49[22] , \nScanOut108[5] , 
        \nOut1_44[4] , \nScanOut1[0] , \nScanOut2[16] , \nOut1_16[13] , 
        \nOut1_63[23] , \nScanOut84[15] , \nOut0_3[27] , \nOut1_7[31] , 
        \nOut1_7[28] , \nOut0_18[23] , \nOut1_20[16] , \nOut1_35[22] , 
        \nOut1_40[12] , \nScanOut116[27] , \nScanOut29[15] , \nOut1_55[26] , 
        \nScanOut103[13] , \nScanOut91[21] , \nScanOut120[22] , 
        \nScanOut49[11] , \nOut1_47[7] , \nScanOut110[7] , \nOut0_3[14] , 
        \nOut1_9[3] , \nScanOut11[4] , \nScanOut12[7] , \nScanOut22[19] , 
        \nScanOut57[29] , \nScanOut9[30] , \nScanOut9[29] , \nOut0_19[4] , 
        \nOut1_38[2] , \nScanOut57[30] , \nScanOut74[18] , \nOut0_25[19] , 
        \nScanOut113[4] , \nOut0_50[30] , \nOut0_50[29] , \nScanOut75[0] , 
        \nOut1_3[23] , \nScanOut30[6] , \nOut1_41[9] , \nScanOut76[3] , 
        \nOut1_3[10] , \nOut1_12[18] , \nOut1_31[30] , \nOut1_19[0] , 
        \nOut1_31[29] , \nOut0_38[6] , \nOut0_25[9] , \nOut1_44[19] , 
        \nScanOut107[18] , \nScanOut124[30] , \nScanOut124[29] , 
        \nScanOut33[5] , \nScanOut38[19] , \nScanOut86[4] , \nScanOut2[3] , 
        \nScanOut54[2] , \nOut1_63[8] , \nScanOut57[1] , \nScanOut98[8] , 
        \nScanOut85[7] , \nScanOut95[19] , \nOut0_4[0] , \nScanOut10[24] , 
        \nScanOut65[14] , \nOut0_20[4] , \nScanOut46[25] , \nScanOut26[21] , 
        \nScanOut33[15] , \nScanOut36[8] , \nScanOut53[11] , \nScanOut70[20] , 
        \nOut0_7[3] , \nScanOut28[4] , \nOut0_8[22] , \nScanOut9[20] , 
        \nScanOut10[17] , \nOut0_17[17] , \nOut0_21[12] , \nOut0_23[7] , 
        \nOut0_54[22] , \nOut1_19[27] , \nScanOut26[12] , \nOut0_34[26] , 
        \nOut0_62[27] , \nScanOut119[13] , \nOut0_41[16] , \nOut0_44[0] , 
        \nScanOut53[22] , \nScanOut70[13] , \nOut0_17[24] , \nOut1_19[14] , 
        \nScanOut33[26] , \nScanOut65[27] , \nScanOut46[16] , \nOut0_62[14] , 
        \nOut0_21[21] , \nOut0_34[15] , \nOut0_41[25] , \nOut0_47[3] , 
        \nScanOut119[20] , \nOut0_54[11] , \nScanOut83[9] , \nScanOut9[13] , 
        \nOut0_13[15] , \nScanOut14[26] , \nScanOut22[23] , \nOut0_25[10] , 
        \nOut0_30[24] , \nOut1_42[3] , \nOut0_45[14] , \nOut0_63[5] , 
        \nScanOut108[25] , \nOut0_50[20] , \nScanOut57[13] , \nScanOut68[6] , 
        \nScanOut75[9] , \nScanOut61[16] , \nScanOut74[22] , \nOut0_25[23] , 
        \nScanOut37[17] , \nOut1_41[0] , \nScanOut42[27] , \nOut0_60[6] , 
        \nOut0_50[13] , \nScanOut108[16] , \nOut0_13[26] , \nScanOut14[15] , 
        \nOut1_26[7] , \nOut0_45[27] , \nOut0_30[17] , \nScanOut22[10] , 
        \nOut1_25[4] , \nScanOut37[24] , \nScanOut61[25] , \nScanOut42[14] , 
        \nScanOut57[20] , \nScanOut74[11] , \nScanOut73[7] , \nOut1_7[21] , 
        \nOut1_59[2] , \nScanOut91[31] , \nScanOut91[28] , \nOut1_7[12] , 
        \nOut0_8[11] , \nOut1_16[30] , \nOut1_16[29] , \nOut0_18[19] , 
        \nOut1_40[31] , \nScanOut49[18] , \nScanOut70[4] , \nOut1_63[19] , 
        \nOut1_40[28] , \nScanOut116[0] , \nScanOut17[3] , \nOut1_20[9] , 
        \nOut1_35[18] , \nScanOut103[30] , \nScanOut103[29] , 
        \nScanOut120[18] , \nScanOut14[0] , \nScanOut115[3] , \nOut1_28[1] , 
        \nScanOut103[7] , \nEnable[0] , \nOut1_1[2] , \nOut0_2[24] , 
        \nScanOut8[19] , \nOut0_14[8] , \nOut0_24[30] , \nOut0_24[29] , 
        \nOut0_51[19] , \nOut0_2[17] , \nScanOut23[30] , \nScanOut75[28] , 
        \nScanOut100[4] , \nScanOut23[29] , \nScanOut56[19] , \nScanOut75[31] , 
        \nScanOut66[0] , \nOut1_2[1] , \nOut1_6[18] , \nScanOut19[5] , 
        \nScanOut28[25] , \nOut1_52[9] , \nScanOut65[3] , \nScanOut105[9] , 
        \nScanOut48[21] , \nScanOut3[26] , \nOut0_11[5] , \nOut0_12[6] , 
        \nOut1_33[0] , \nScanOut118[6] , \nOut1_30[3] , \nOut1_34[12] , 
        \nOut1_41[22] , \nScanOut117[17] , \nOut1_62[13] , \nOut1_17[23] , 
        \nOut0_19[13] , \nScanOut85[25] , \nScanOut90[11] , \nScanOut121[12] , 
        \nScanOut3[15] , \nOut1_17[10] , \nOut1_21[26] , \nOut1_54[16] , 
        \nScanOut102[23] , \nOut1_21[15] , \nScanOut28[16] , \nScanOut48[12] , 
        \nOut1_57[4] , \nScanOut90[22] , \nScanOut121[21] , \nOut1_34[21] , 
        \nOut1_49[8] , \nOut1_54[25] , \nScanOut102[10] , \nOut1_41[11] , 
        \nScanOut117[24] , \nOut1_62[20] , \nScanOut85[16] , \nOut0_9[31] , 
        \nOut0_9[28] , \nOut0_19[20] , \nOut1_54[7] , \nScanOut94[13] , 
        \nScanOut125[10] , \nOut1_2[30] , \nScanOut7[24] , \nOut1_25[24] , 
        \nOut1_50[14] , \nScanOut106[21] , \nOut1_30[10] , \nOut1_45[20] , 
        \nScanOut113[15] , \nScanOut7[17] , \nOut1_13[21] , \nOut1_13[12] , 
        \nOut1_14[5] , \nOut0_35[3] , \nScanOut39[13] , \nScanOut44[8] , 
        \nOut0_51[7] , \nScanOut81[27] , \nOut0_52[4] , \nScanOut88[2] , 
        \nScanOut59[17] , \nScanOut59[7] , \nOut1_30[23] , \nOut1_45[13] , 
        \nScanOut113[26] , \nScanOut81[14] , \nOut1_25[17] , \nScanOut94[20] , 
        \nScanOut125[23] , \nScanOut39[20] , \nOut1_50[27] , \nScanOut106[12] , 
        \nScanOut59[24] , \nOut1_2[29] , \nOut0_3[23] , \nOut0_6[26] , 
        \nOut1_17[6] , \nOut0_36[0] , \nScanOut93[3] , \nOut0_6[15] , 
        \nOut1_9[25] , \nScanOut9[8] , \nScanOut41[5] , \nOut0_57[9] , 
        \nScanOut27[18] , \nScanOut52[31] , \nScanOut71[19] , \nScanOut42[6] , 
        \nScanOut52[28] , \nOut0_20[18] , \nOut0_49[5] , \nOut0_55[31] , 
        \nScanOut90[0] , \nScanOut25[1] , \nOut0_55[28] , \nScanOut118[19] , 
        \nOut0_9[5] , \nOut1_9[16] , \nOut1_11[8] , \nScanOut124[2] , 
        \nScanOut127[1] , \nScanOut26[2] , \nOut1_9[7] , \nScanOut14[18] , 
        \nOut0_19[0] , \nOut1_38[6] , \nScanOut113[0] , \nScanOut37[29] , 
        \nScanOut42[19] , \nScanOut61[31] , \nScanOut37[30] , \nScanOut61[28] , 
        \nScanOut11[0] , \nScanOut12[3] , \nOut1_25[9] , \nOut0_3[10] , 
        \nScanOut76[7] , \nScanOut110[3] , \nOut0_13[18] , \nOut0_30[29] , 
        \nOut0_45[19] , \nOut1_23[7] , \nScanOut29[22] , \nOut0_30[30] , 
        \nOut0_63[8] , \nScanOut108[31] , \nScanOut108[28] , \nScanOut75[4] , 
        \nScanOut49[26] , \nScanOut108[1] , \nScanOut2[21] , \nOut1_20[4] , 
        \nOut1_35[15] , \nOut1_40[25] , \nScanOut116[10] , \nScanOut2[12] , 
        \nOut1_16[24] , \nOut0_18[14] , \nOut1_63[14] , \nOut1_16[17] , 
        \nOut1_20[21] , \nOut1_55[11] , \nScanOut84[22] , \nScanOut91[16] , 
        \nScanOut120[15] , \nScanOut103[24] , \nOut1_20[12] , \nScanOut29[11] , 
        \nOut1_47[3] , \nScanOut49[15] , \nScanOut70[9] , \nScanOut91[25] , 
        \nScanOut120[26] , \nOut1_35[26] , \nOut1_55[22] , \nScanOut103[17] , 
        \nOut1_40[16] , \nScanOut116[23] , \nScanOut84[11] , \nOut0_18[27] , 
        \nOut1_63[27] , \nOut1_44[0] , \nOut0_1[0] , \nScanOut6[23] , 
        \nOut1_24[23] , \nOut1_51[13] , \nScanOut95[14] , \nScanOut124[17] , 
        \nScanOut107[26] , \nOut1_31[17] , \nOut1_44[27] , \nScanOut112[12] , 
        \nOut1_12[26] , \nOut0_25[4] , \nScanOut38[14] , \nOut0_41[0] , 
        \nOut1_60[6] , \nScanOut80[20] , \nOut0_42[3] , \nOut1_63[5] , 
        \nScanOut98[5] , \nScanOut49[0] , \nScanOut58[10] , \nScanOut86[9] , 
        \nOut1_31[24] , \nScanOut33[8] , \nOut1_44[14] , \nScanOut112[21] , 
        \nOut0_2[30] , \nOut0_2[3] , \nScanOut6[10] , \nOut1_12[15] , 
        \nScanOut80[13] , \nOut1_24[10] , \nScanOut95[27] , \nScanOut124[24] , 
        \nOut1_51[20] , \nScanOut107[15] , \nOut1_2[24] , \nScanOut4[0] , 
        \nOut0_7[21] , \nOut0_26[7] , \nScanOut38[27] , \nScanOut58[23] , 
        \nScanOut83[4] , \nOut0_7[12] , \nScanOut7[3] , \nOut1_8[22] , 
        \nOut0_17[30] , \nOut0_34[18] , \nOut0_41[28] , \nScanOut51[2] , 
        \nOut0_17[29] , \nOut1_19[19] , \nOut0_41[31] , \nOut0_62[19] , 
        \nScanOut52[1] , \nOut0_59[2] , \nScanOut80[7] , \nScanOut35[6] , 
        \nOut1_8[11] , \nScanOut10[30] , \nOut0_20[9] , \nScanOut28[9] , 
        \nScanOut46[28] , \nScanOut33[18] , \nScanOut36[5] , \nScanOut10[29] , 
        \nScanOut46[31] , \nScanOut65[19] , \nScanOut20[1] , \nScanOut59[30] , 
        \nScanOut59[29] , \nOut1_2[17] , \nOut1_14[8] , \nOut0_28[1] , 
        \nScanOut81[19] , \nScanOut121[2] , \nScanOut122[1] , \nScanOut23[2] , 
        \nOut0_6[18] , \nScanOut7[30] , \nScanOut7[29] , \nOut1_25[30] , 
        \nOut1_25[29] , \nScanOut44[5] , \nOut0_52[9] , \nScanOut96[3] , 
        \nScanOut47[6] , \nOut1_50[19] , \nScanOut95[0] , \nOut0_9[8] , 
        \nScanOut64[13] , \nScanOut113[18] , \nOut1_11[5] , \nScanOut11[23] , 
        \nOut0_30[3] , \nScanOut47[22] , \nScanOut27[26] , \nScanOut32[12] , 
        \nScanOut52[16] , \nScanOut38[3] , \nScanOut71[27] , \nScanOut8[27] , 
        \nOut1_9[31] , \nOut1_9[28] , \nScanOut11[10] , \nOut1_12[6] , 
        \nOut0_33[0] , \nOut0_16[10] , \nOut0_20[15] , \nOut0_55[25] , 
        \nOut1_18[20] , \nScanOut27[15] , \nOut0_35[21] , \nOut0_63[20] , 
        \nScanOut118[14] , \nOut0_40[11] , \nOut0_49[8] , \nOut0_54[7] , 
        \nScanOut52[25] , \nScanOut71[14] , \nScanOut64[20] , \nScanOut32[21] , 
        \nScanOut9[5] , \nOut0_16[23] , \nOut1_18[13] , \nScanOut47[11] , 
        \nOut0_63[13] , \nOut0_35[12] , \nOut0_40[22] , \nScanOut41[8] , 
        \nOut0_57[4] , \nScanOut118[27] , \nOut0_55[16] , \nOut0_20[26] , 
        \nOut0_12[12] , \nScanOut15[21] , \nScanOut23[24] , \nOut0_24[17] , 
        \nOut0_31[23] , \nOut0_44[13] , \nScanOut109[22] , \nOut0_51[27] , 
        \nOut1_52[4] , \nScanOut56[14] , \nScanOut78[1] , \nScanOut60[11] , 
        \nScanOut75[25] , \nScanOut36[10] , \nScanOut43[20] , \nOut1_51[7] , 
        \nScanOut100[9] , \nOut0_2[29] , \nOut1_7[1] , \nScanOut8[14] , 
        \nOut0_24[24] , \nOut0_51[14] , \nScanOut109[11] , \nOut0_12[21] , 
        \nOut0_14[5] , \nScanOut15[12] , \nOut0_17[6] , \nOut1_36[0] , 
        \nOut0_44[20] , \nOut0_31[10] , \nOut1_35[3] , \nScanOut36[23] , 
        \nScanOut60[22] , \nScanOut43[13] , \nScanOut23[17] , \nScanOut56[27] , 
        \nScanOut75[16] , \nOut0_1[9] , \nOut1_1[6] , \nScanOut3[18] , 
        \nOut1_4[2] , \nOut0_9[25] , \nOut1_21[18] , \nScanOut63[0] , 
        \nOut1_54[31] , \nOut1_54[28] , \nOut0_6[22] , \nOut1_6[26] , 
        \nOut1_49[5] , \nScanOut117[30] , \nScanOut117[29] , \nOut1_6[15] , 
        \nOut0_9[16] , \nOut0_11[8] , \nOut1_57[9] , \nScanOut60[3] , 
        \nScanOut85[31] , \nScanOut85[28] , \nScanOut106[7] , \nScanOut28[31] , 
        \nScanOut28[28] , \nScanOut105[4] , \nOut1_9[21] , \nScanOut11[19] , 
        \nScanOut19[8] , \nOut0_49[1] , \nScanOut90[4] , \nScanOut32[31] , 
        \nScanOut32[28] , \nScanOut64[29] , \nScanOut41[1] , \nScanOut42[2] , 
        \nScanOut47[18] , \nScanOut64[30] , \nOut0_6[11] , \nOut0_9[1] , 
        \nOut1_9[12] , \nScanOut93[7] , \nScanOut26[6] , \nScanOut124[6] , 
        \nScanOut127[5] , \nScanOut7[20] , \nOut0_16[19] , \nOut1_18[30] , 
        \nOut1_18[29] , \nOut0_35[31] , \nOut0_35[28] , \nOut0_63[29] , 
        \nScanOut25[5] , \nOut0_33[9] , \nOut0_40[18] , \nOut0_63[30] , 
        \nScanOut39[17] , \nScanOut59[13] , \nOut0_51[3] , \nOut0_52[0] , 
        \nScanOut59[3] , \nScanOut88[6] , \nScanOut7[13] , \nOut1_13[25] , 
        \nOut1_13[16] , \nOut1_17[2] , \nOut1_25[20] , \nOut1_30[14] , 
        \nOut1_45[24] , \nScanOut81[23] , \nScanOut113[11] , \nOut1_50[10] , 
        \nScanOut106[25] , \nScanOut95[9] , \nOut0_36[4] , \nScanOut94[17] , 
        \nScanOut125[14] , \nScanOut20[8] , \nOut1_25[13] , \nScanOut39[24] , 
        \nScanOut59[20] , \nScanOut122[8] , \nOut1_50[23] , \nScanOut106[16] , 
        \nScanOut94[24] , \nScanOut125[27] , \nScanOut81[10] , \nOut1_14[1] , 
        \nOut0_28[8] , \nOut1_30[27] , \nOut0_35[7] , \nOut1_45[17] , 
        \nScanOut113[22] , \nOut1_21[22] , \nOut1_54[12] , \nScanOut102[27] , 
        \nScanOut90[15] , \nScanOut121[16] , \nOut0_2[20] , \nOut1_2[5] , 
        \nScanOut3[22] , \nOut0_11[1] , \nOut1_17[27] , \nOut0_19[17] , 
        \nOut1_62[17] , \nOut1_30[7] , \nOut1_34[16] , \nOut1_41[26] , 
        \nScanOut85[21] , \nScanOut117[13] , \nOut0_12[2] , \nOut1_33[4] , 
        \nScanOut118[2] , \nScanOut3[11] , \nOut1_17[14] , \nScanOut19[1] , 
        \nScanOut48[25] , \nScanOut28[21] , \nOut1_54[3] , \nScanOut63[9] , 
        \nScanOut85[12] , \nOut1_7[8] , \nOut0_19[24] , \nOut1_62[24] , 
        \nOut1_21[11] , \nOut1_34[25] , \nOut1_41[15] , \nScanOut117[20] , 
        \nScanOut28[12] , \nOut1_54[21] , \nScanOut102[14] , \nScanOut90[26] , 
        \nScanOut121[25] , \nScanOut48[16] , \nOut1_57[0] , \nScanOut100[0] , 
        \nOut0_2[13] , \nOut0_12[31] , \nOut0_12[28] , \nOut0_44[30] , 
        \nOut0_31[19] , \nOut1_36[9] , \nOut0_44[29] , \nOut1_28[5] , 
        \nScanOut109[18] , \nScanOut65[7] , \nScanOut103[3] , \nScanOut78[8] , 
        \nScanOut2[31] , \nOut1_7[25] , \nScanOut15[31] , \nScanOut15[28] , 
        \nScanOut43[30] , \nScanOut60[18] , \nScanOut36[19] , \nScanOut43[29] , 
        \nScanOut29[18] , \nScanOut66[4] , \nScanOut70[0] , \nOut1_7[16] , 
        \nOut0_8[26] , \nOut1_44[9] , \nOut1_59[6] , \nScanOut84[18] , 
        \nScanOut73[3] , \nOut0_8[15] , \nScanOut14[4] , \nScanOut115[7] , 
        \nScanOut108[8] , \nScanOut17[7] , \nOut1_20[31] , \nOut1_20[28] , 
        \nOut1_55[18] , \nScanOut2[28] , \nScanOut116[19] , \nScanOut116[4] , 
        \nOut0_3[19] , \nScanOut14[22] , \nScanOut37[13] , \nOut1_41[4] , 
        \nScanOut42[23] , \nOut0_60[2] , \nScanOut61[12] , \nScanOut22[27] , 
        \nScanOut57[17] , \nScanOut74[26] , \nOut0_4[4] , \nOut0_7[7] , 
        \nScanOut9[24] , \nOut0_25[14] , \nOut0_63[1] , \nScanOut68[2] , 
        \nScanOut108[21] , \nOut0_30[20] , \nOut1_42[7] , \nOut0_50[24] , 
        \nOut0_45[10] , \nScanOut9[17] , \nScanOut11[9] , \nOut0_13[11] , 
        \nScanOut14[11] , \nOut0_19[9] , \nScanOut22[14] , \nOut1_25[0] , 
        \nScanOut74[15] , \nScanOut113[9] , \nScanOut37[20] , \nScanOut57[24] , 
        \nScanOut42[10] , \nOut1_26[3] , \nScanOut61[21] , \nOut0_45[23] , 
        \nOut0_30[13] , \nOut0_13[22] , \nOut0_17[13] , \nOut0_25[27] , 
        \nOut0_50[17] , \nScanOut108[12] , \nOut0_34[22] , \nScanOut119[17] , 
        \nOut0_41[12] , \nOut1_19[23] , \nOut0_21[16] , \nOut0_23[3] , 
        \nOut0_62[23] , \nOut0_54[26] , \nScanOut28[0] , \nScanOut4[9] , 
        \nOut0_7[28] , \nOut1_8[18] , \nOut0_20[0] , \nScanOut26[25] , 
        \nScanOut53[15] , \nScanOut70[24] , \nScanOut46[21] , \nScanOut33[11] , 
        \nScanOut65[10] , \nScanOut10[20] , \nOut0_7[31] , \nScanOut10[13] , 
        \nOut0_17[20] , \nOut1_19[10] , \nOut0_21[25] , \nOut0_54[15] , 
        \nOut0_34[11] , \nOut0_41[21] , \nOut0_47[7] , \nScanOut119[24] , 
        \nOut0_62[10] , \nScanOut33[22] , \nScanOut46[12] , \nOut1_19[4] , 
        \nOut1_24[19] , \nScanOut26[16] , \nOut0_44[4] , \nScanOut65[23] , 
        \nScanOut70[17] , \nScanOut33[1] , \nScanOut52[8] , \nScanOut53[26] , 
        \nOut1_51[30] , \nOut0_38[2] , \nOut1_51[29] , \nScanOut112[28] , 
        \nScanOut1[4] , \nScanOut2[7] , \nOut1_3[27] , \nScanOut6[19] , 
        \nScanOut112[31] , \nScanOut30[2] , \nOut0_41[9] , \nScanOut80[30] , 
        \nScanOut80[29] , \nScanOut85[3] , \nScanOut54[6] , \nScanOut57[5] , 
        \nOut1_3[14] , \nScanOut49[9] , \nScanOut58[19] , \nScanOut86[0] ;
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut4[31] , \nScanOut4[30] , \nScanOut4[29] , 
        \nScanOut4[28] , \nScanOut4[27] , \nScanOut4[26] , \nScanOut4[25] , 
        \nScanOut4[24] , \nScanOut4[23] , \nScanOut4[22] , \nScanOut4[21] , 
        \nScanOut4[20] , \nScanOut4[19] , \nScanOut4[18] , \nScanOut4[17] , 
        \nScanOut4[16] , \nScanOut4[15] , \nScanOut4[14] , \nScanOut4[13] , 
        \nScanOut4[12] , \nScanOut4[11] , \nScanOut4[10] , \nScanOut4[9] , 
        \nScanOut4[8] , \nScanOut4[7] , \nScanOut4[6] , \nScanOut4[5] , 
        \nScanOut4[4] , \nScanOut4[3] , \nScanOut4[2] , \nScanOut4[1] , 
        \nScanOut4[0] }), .ScanOut({\nScanOut3[31] , \nScanOut3[30] , 
        \nScanOut3[29] , \nScanOut3[28] , \nScanOut3[27] , \nScanOut3[26] , 
        \nScanOut3[25] , \nScanOut3[24] , \nScanOut3[23] , \nScanOut3[22] , 
        \nScanOut3[21] , \nScanOut3[20] , \nScanOut3[19] , \nScanOut3[18] , 
        \nScanOut3[17] , \nScanOut3[16] , \nScanOut3[15] , \nScanOut3[14] , 
        \nScanOut3[13] , \nScanOut3[12] , \nScanOut3[11] , \nScanOut3[10] , 
        \nScanOut3[9] , \nScanOut3[8] , \nScanOut3[7] , \nScanOut3[6] , 
        \nScanOut3[5] , \nScanOut3[4] , \nScanOut3[3] , \nScanOut3[2] , 
        \nScanOut3[1] , \nScanOut3[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_3[31] , 
        \nOut0_3[30] , \nOut0_3[29] , \nOut0_3[28] , \nOut0_3[27] , 
        \nOut0_3[26] , \nOut0_3[25] , \nOut0_3[24] , \nOut0_3[23] , 
        \nOut0_3[22] , \nOut0_3[21] , \nOut0_3[20] , \nOut0_3[19] , 
        \nOut0_3[18] , \nOut0_3[17] , \nOut0_3[16] , \nOut0_3[15] , 
        \nOut0_3[14] , \nOut0_3[13] , \nOut0_3[12] , \nOut0_3[11] , 
        \nOut0_3[10] , \nOut0_3[9] , \nOut0_3[8] , \nOut0_3[7] , \nOut0_3[6] , 
        \nOut0_3[5] , \nOut0_3[4] , \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , 
        \nOut0_3[0] }), .NORTH_EDGE({\nOut0_2[31] , \nOut0_2[30] , 
        \nOut0_2[29] , \nOut0_2[28] , \nOut0_2[27] , \nOut0_2[26] , 
        \nOut0_2[25] , \nOut0_2[24] , \nOut0_2[23] , \nOut0_2[22] , 
        \nOut0_2[21] , \nOut0_2[20] , \nOut0_2[19] , \nOut0_2[18] , 
        \nOut0_2[17] , \nOut0_2[16] , \nOut0_2[15] , \nOut0_2[14] , 
        \nOut0_2[13] , \nOut0_2[12] , \nOut0_2[11] , \nOut0_2[10] , 
        \nOut0_2[9] , \nOut0_2[8] , \nOut0_2[7] , \nOut0_2[6] , \nOut0_2[5] , 
        \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , \nOut0_2[0] }), 
        .SOUTH_EDGE({\nOut0_4[31] , \nOut0_4[30] , \nOut0_4[29] , 
        \nOut0_4[28] , \nOut0_4[27] , \nOut0_4[26] , \nOut0_4[25] , 
        \nOut0_4[24] , \nOut0_4[23] , \nOut0_4[22] , \nOut0_4[21] , 
        \nOut0_4[20] , \nOut0_4[19] , \nOut0_4[18] , \nOut0_4[17] , 
        \nOut0_4[16] , \nOut0_4[15] , \nOut0_4[14] , \nOut0_4[13] , 
        \nOut0_4[12] , \nOut0_4[11] , \nOut0_4[10] , \nOut0_4[9] , 
        \nOut0_4[8] , \nOut0_4[7] , \nOut0_4[6] , \nOut0_4[5] , \nOut0_4[4] , 
        \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , \nOut0_4[0] }), .EAST_EDGE(
        \nOut1_3[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_2[31] ), .SE_EDGE(\nOut1_4[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_54 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut55[31] , \nScanOut55[30] , \nScanOut55[29] , 
        \nScanOut55[28] , \nScanOut55[27] , \nScanOut55[26] , \nScanOut55[25] , 
        \nScanOut55[24] , \nScanOut55[23] , \nScanOut55[22] , \nScanOut55[21] , 
        \nScanOut55[20] , \nScanOut55[19] , \nScanOut55[18] , \nScanOut55[17] , 
        \nScanOut55[16] , \nScanOut55[15] , \nScanOut55[14] , \nScanOut55[13] , 
        \nScanOut55[12] , \nScanOut55[11] , \nScanOut55[10] , \nScanOut55[9] , 
        \nScanOut55[8] , \nScanOut55[7] , \nScanOut55[6] , \nScanOut55[5] , 
        \nScanOut55[4] , \nScanOut55[3] , \nScanOut55[2] , \nScanOut55[1] , 
        \nScanOut55[0] }), .ScanOut({\nScanOut54[31] , \nScanOut54[30] , 
        \nScanOut54[29] , \nScanOut54[28] , \nScanOut54[27] , \nScanOut54[26] , 
        \nScanOut54[25] , \nScanOut54[24] , \nScanOut54[23] , \nScanOut54[22] , 
        \nScanOut54[21] , \nScanOut54[20] , \nScanOut54[19] , \nScanOut54[18] , 
        \nScanOut54[17] , \nScanOut54[16] , \nScanOut54[15] , \nScanOut54[14] , 
        \nScanOut54[13] , \nScanOut54[12] , \nScanOut54[11] , \nScanOut54[10] , 
        \nScanOut54[9] , \nScanOut54[8] , \nScanOut54[7] , \nScanOut54[6] , 
        \nScanOut54[5] , \nScanOut54[4] , \nScanOut54[3] , \nScanOut54[2] , 
        \nScanOut54[1] , \nScanOut54[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_54[31] , 
        \nOut0_54[30] , \nOut0_54[29] , \nOut0_54[28] , \nOut0_54[27] , 
        \nOut0_54[26] , \nOut0_54[25] , \nOut0_54[24] , \nOut0_54[23] , 
        \nOut0_54[22] , \nOut0_54[21] , \nOut0_54[20] , \nOut0_54[19] , 
        \nOut0_54[18] , \nOut0_54[17] , \nOut0_54[16] , \nOut0_54[15] , 
        \nOut0_54[14] , \nOut0_54[13] , \nOut0_54[12] , \nOut0_54[11] , 
        \nOut0_54[10] , \nOut0_54[9] , \nOut0_54[8] , \nOut0_54[7] , 
        \nOut0_54[6] , \nOut0_54[5] , \nOut0_54[4] , \nOut0_54[3] , 
        \nOut0_54[2] , \nOut0_54[1] , \nOut0_54[0] }), .NORTH_EDGE({
        \nOut0_53[31] , \nOut0_53[30] , \nOut0_53[29] , \nOut0_53[28] , 
        \nOut0_53[27] , \nOut0_53[26] , \nOut0_53[25] , \nOut0_53[24] , 
        \nOut0_53[23] , \nOut0_53[22] , \nOut0_53[21] , \nOut0_53[20] , 
        \nOut0_53[19] , \nOut0_53[18] , \nOut0_53[17] , \nOut0_53[16] , 
        \nOut0_53[15] , \nOut0_53[14] , \nOut0_53[13] , \nOut0_53[12] , 
        \nOut0_53[11] , \nOut0_53[10] , \nOut0_53[9] , \nOut0_53[8] , 
        \nOut0_53[7] , \nOut0_53[6] , \nOut0_53[5] , \nOut0_53[4] , 
        \nOut0_53[3] , \nOut0_53[2] , \nOut0_53[1] , \nOut0_53[0] }), 
        .SOUTH_EDGE({\nOut0_55[31] , \nOut0_55[30] , \nOut0_55[29] , 
        \nOut0_55[28] , \nOut0_55[27] , \nOut0_55[26] , \nOut0_55[25] , 
        \nOut0_55[24] , \nOut0_55[23] , \nOut0_55[22] , \nOut0_55[21] , 
        \nOut0_55[20] , \nOut0_55[19] , \nOut0_55[18] , \nOut0_55[17] , 
        \nOut0_55[16] , \nOut0_55[15] , \nOut0_55[14] , \nOut0_55[13] , 
        \nOut0_55[12] , \nOut0_55[11] , \nOut0_55[10] , \nOut0_55[9] , 
        \nOut0_55[8] , \nOut0_55[7] , \nOut0_55[6] , \nOut0_55[5] , 
        \nOut0_55[4] , \nOut0_55[3] , \nOut0_55[2] , \nOut0_55[1] , 
        \nOut0_55[0] }), .EAST_EDGE(\nOut1_54[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_53[31] ), .SE_EDGE(
        \nOut1_55[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_96 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut97[31] , \nScanOut97[30] , \nScanOut97[29] , 
        \nScanOut97[28] , \nScanOut97[27] , \nScanOut97[26] , \nScanOut97[25] , 
        \nScanOut97[24] , \nScanOut97[23] , \nScanOut97[22] , \nScanOut97[21] , 
        \nScanOut97[20] , \nScanOut97[19] , \nScanOut97[18] , \nScanOut97[17] , 
        \nScanOut97[16] , \nScanOut97[15] , \nScanOut97[14] , \nScanOut97[13] , 
        \nScanOut97[12] , \nScanOut97[11] , \nScanOut97[10] , \nScanOut97[9] , 
        \nScanOut97[8] , \nScanOut97[7] , \nScanOut97[6] , \nScanOut97[5] , 
        \nScanOut97[4] , \nScanOut97[3] , \nScanOut97[2] , \nScanOut97[1] , 
        \nScanOut97[0] }), .ScanOut({\nScanOut96[31] , \nScanOut96[30] , 
        \nScanOut96[29] , \nScanOut96[28] , \nScanOut96[27] , \nScanOut96[26] , 
        \nScanOut96[25] , \nScanOut96[24] , \nScanOut96[23] , \nScanOut96[22] , 
        \nScanOut96[21] , \nScanOut96[20] , \nScanOut96[19] , \nScanOut96[18] , 
        \nScanOut96[17] , \nScanOut96[16] , \nScanOut96[15] , \nScanOut96[14] , 
        \nScanOut96[13] , \nScanOut96[12] , \nScanOut96[11] , \nScanOut96[10] , 
        \nScanOut96[9] , \nScanOut96[8] , \nScanOut96[7] , \nScanOut96[6] , 
        \nScanOut96[5] , \nScanOut96[4] , \nScanOut96[3] , \nScanOut96[2] , 
        \nScanOut96[1] , \nScanOut96[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_32[31] , 
        \nOut1_32[30] , \nOut1_32[29] , \nOut1_32[28] , \nOut1_32[27] , 
        \nOut1_32[26] , \nOut1_32[25] , \nOut1_32[24] , \nOut1_32[23] , 
        \nOut1_32[22] , \nOut1_32[21] , \nOut1_32[20] , \nOut1_32[19] , 
        \nOut1_32[18] , \nOut1_32[17] , \nOut1_32[16] , \nOut1_32[15] , 
        \nOut1_32[14] , \nOut1_32[13] , \nOut1_32[12] , \nOut1_32[11] , 
        \nOut1_32[10] , \nOut1_32[9] , \nOut1_32[8] , \nOut1_32[7] , 
        \nOut1_32[6] , \nOut1_32[5] , \nOut1_32[4] , \nOut1_32[3] , 
        \nOut1_32[2] , \nOut1_32[1] , \nOut1_32[0] }), .NORTH_EDGE({
        \nOut1_31[31] , \nOut1_31[30] , \nOut1_31[29] , \nOut1_31[28] , 
        \nOut1_31[27] , \nOut1_31[26] , \nOut1_31[25] , \nOut1_31[24] , 
        \nOut1_31[23] , \nOut1_31[22] , \nOut1_31[21] , \nOut1_31[20] , 
        \nOut1_31[19] , \nOut1_31[18] , \nOut1_31[17] , \nOut1_31[16] , 
        \nOut1_31[15] , \nOut1_31[14] , \nOut1_31[13] , \nOut1_31[12] , 
        \nOut1_31[11] , \nOut1_31[10] , \nOut1_31[9] , \nOut1_31[8] , 
        \nOut1_31[7] , \nOut1_31[6] , \nOut1_31[5] , \nOut1_31[4] , 
        \nOut1_31[3] , \nOut1_31[2] , \nOut1_31[1] , \nOut1_31[0] }), 
        .SOUTH_EDGE({\nOut1_33[31] , \nOut1_33[30] , \nOut1_33[29] , 
        \nOut1_33[28] , \nOut1_33[27] , \nOut1_33[26] , \nOut1_33[25] , 
        \nOut1_33[24] , \nOut1_33[23] , \nOut1_33[22] , \nOut1_33[21] , 
        \nOut1_33[20] , \nOut1_33[19] , \nOut1_33[18] , \nOut1_33[17] , 
        \nOut1_33[16] , \nOut1_33[15] , \nOut1_33[14] , \nOut1_33[13] , 
        \nOut1_33[12] , \nOut1_33[11] , \nOut1_33[10] , \nOut1_33[9] , 
        \nOut1_33[8] , \nOut1_33[7] , \nOut1_33[6] , \nOut1_33[5] , 
        \nOut1_33[4] , \nOut1_33[3] , \nOut1_33[2] , \nOut1_33[1] , 
        \nOut1_33[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_32[0] ), 
        .NW_EDGE(\nOut0_31[0] ), .SW_EDGE(\nOut0_33[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_73 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut74[31] , \nScanOut74[30] , \nScanOut74[29] , 
        \nScanOut74[28] , \nScanOut74[27] , \nScanOut74[26] , \nScanOut74[25] , 
        \nScanOut74[24] , \nScanOut74[23] , \nScanOut74[22] , \nScanOut74[21] , 
        \nScanOut74[20] , \nScanOut74[19] , \nScanOut74[18] , \nScanOut74[17] , 
        \nScanOut74[16] , \nScanOut74[15] , \nScanOut74[14] , \nScanOut74[13] , 
        \nScanOut74[12] , \nScanOut74[11] , \nScanOut74[10] , \nScanOut74[9] , 
        \nScanOut74[8] , \nScanOut74[7] , \nScanOut74[6] , \nScanOut74[5] , 
        \nScanOut74[4] , \nScanOut74[3] , \nScanOut74[2] , \nScanOut74[1] , 
        \nScanOut74[0] }), .ScanOut({\nScanOut73[31] , \nScanOut73[30] , 
        \nScanOut73[29] , \nScanOut73[28] , \nScanOut73[27] , \nScanOut73[26] , 
        \nScanOut73[25] , \nScanOut73[24] , \nScanOut73[23] , \nScanOut73[22] , 
        \nScanOut73[21] , \nScanOut73[20] , \nScanOut73[19] , \nScanOut73[18] , 
        \nScanOut73[17] , \nScanOut73[16] , \nScanOut73[15] , \nScanOut73[14] , 
        \nScanOut73[13] , \nScanOut73[12] , \nScanOut73[11] , \nScanOut73[10] , 
        \nScanOut73[9] , \nScanOut73[8] , \nScanOut73[7] , \nScanOut73[6] , 
        \nScanOut73[5] , \nScanOut73[4] , \nScanOut73[3] , \nScanOut73[2] , 
        \nScanOut73[1] , \nScanOut73[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_9[31] , 
        \nOut1_9[30] , \nOut1_9[29] , \nOut1_9[28] , \nOut1_9[27] , 
        \nOut1_9[26] , \nOut1_9[25] , \nOut1_9[24] , \nOut1_9[23] , 
        \nOut1_9[22] , \nOut1_9[21] , \nOut1_9[20] , \nOut1_9[19] , 
        \nOut1_9[18] , \nOut1_9[17] , \nOut1_9[16] , \nOut1_9[15] , 
        \nOut1_9[14] , \nOut1_9[13] , \nOut1_9[12] , \nOut1_9[11] , 
        \nOut1_9[10] , \nOut1_9[9] , \nOut1_9[8] , \nOut1_9[7] , \nOut1_9[6] , 
        \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , \nOut1_9[1] , 
        \nOut1_9[0] }), .NORTH_EDGE({\nOut1_8[31] , \nOut1_8[30] , 
        \nOut1_8[29] , \nOut1_8[28] , \nOut1_8[27] , \nOut1_8[26] , 
        \nOut1_8[25] , \nOut1_8[24] , \nOut1_8[23] , \nOut1_8[22] , 
        \nOut1_8[21] , \nOut1_8[20] , \nOut1_8[19] , \nOut1_8[18] , 
        \nOut1_8[17] , \nOut1_8[16] , \nOut1_8[15] , \nOut1_8[14] , 
        \nOut1_8[13] , \nOut1_8[12] , \nOut1_8[11] , \nOut1_8[10] , 
        \nOut1_8[9] , \nOut1_8[8] , \nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , 
        \nOut1_8[4] , \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }), 
        .SOUTH_EDGE({\nOut1_10[31] , \nOut1_10[30] , \nOut1_10[29] , 
        \nOut1_10[28] , \nOut1_10[27] , \nOut1_10[26] , \nOut1_10[25] , 
        \nOut1_10[24] , \nOut1_10[23] , \nOut1_10[22] , \nOut1_10[21] , 
        \nOut1_10[20] , \nOut1_10[19] , \nOut1_10[18] , \nOut1_10[17] , 
        \nOut1_10[16] , \nOut1_10[15] , \nOut1_10[14] , \nOut1_10[13] , 
        \nOut1_10[12] , \nOut1_10[11] , \nOut1_10[10] , \nOut1_10[9] , 
        \nOut1_10[8] , \nOut1_10[7] , \nOut1_10[6] , \nOut1_10[5] , 
        \nOut1_10[4] , \nOut1_10[3] , \nOut1_10[2] , \nOut1_10[1] , 
        \nOut1_10[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_9[0] ), .NW_EDGE(
        \nOut0_8[0] ), .SW_EDGE(\nOut0_10[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0)
         );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_102 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut103[31] , \nScanOut103[30] , \nScanOut103[29] , 
        \nScanOut103[28] , \nScanOut103[27] , \nScanOut103[26] , 
        \nScanOut103[25] , \nScanOut103[24] , \nScanOut103[23] , 
        \nScanOut103[22] , \nScanOut103[21] , \nScanOut103[20] , 
        \nScanOut103[19] , \nScanOut103[18] , \nScanOut103[17] , 
        \nScanOut103[16] , \nScanOut103[15] , \nScanOut103[14] , 
        \nScanOut103[13] , \nScanOut103[12] , \nScanOut103[11] , 
        \nScanOut103[10] , \nScanOut103[9] , \nScanOut103[8] , 
        \nScanOut103[7] , \nScanOut103[6] , \nScanOut103[5] , \nScanOut103[4] , 
        \nScanOut103[3] , \nScanOut103[2] , \nScanOut103[1] , \nScanOut103[0] 
        }), .ScanOut({\nScanOut102[31] , \nScanOut102[30] , \nScanOut102[29] , 
        \nScanOut102[28] , \nScanOut102[27] , \nScanOut102[26] , 
        \nScanOut102[25] , \nScanOut102[24] , \nScanOut102[23] , 
        \nScanOut102[22] , \nScanOut102[21] , \nScanOut102[20] , 
        \nScanOut102[19] , \nScanOut102[18] , \nScanOut102[17] , 
        \nScanOut102[16] , \nScanOut102[15] , \nScanOut102[14] , 
        \nScanOut102[13] , \nScanOut102[12] , \nScanOut102[11] , 
        \nScanOut102[10] , \nScanOut102[9] , \nScanOut102[8] , 
        \nScanOut102[7] , \nScanOut102[6] , \nScanOut102[5] , \nScanOut102[4] , 
        \nScanOut102[3] , \nScanOut102[2] , \nScanOut102[1] , \nScanOut102[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_38[31] , \nOut1_38[30] , \nOut1_38[29] , 
        \nOut1_38[28] , \nOut1_38[27] , \nOut1_38[26] , \nOut1_38[25] , 
        \nOut1_38[24] , \nOut1_38[23] , \nOut1_38[22] , \nOut1_38[21] , 
        \nOut1_38[20] , \nOut1_38[19] , \nOut1_38[18] , \nOut1_38[17] , 
        \nOut1_38[16] , \nOut1_38[15] , \nOut1_38[14] , \nOut1_38[13] , 
        \nOut1_38[12] , \nOut1_38[11] , \nOut1_38[10] , \nOut1_38[9] , 
        \nOut1_38[8] , \nOut1_38[7] , \nOut1_38[6] , \nOut1_38[5] , 
        \nOut1_38[4] , \nOut1_38[3] , \nOut1_38[2] , \nOut1_38[1] , 
        \nOut1_38[0] }), .NORTH_EDGE({\nOut1_37[31] , \nOut1_37[30] , 
        \nOut1_37[29] , \nOut1_37[28] , \nOut1_37[27] , \nOut1_37[26] , 
        \nOut1_37[25] , \nOut1_37[24] , \nOut1_37[23] , \nOut1_37[22] , 
        \nOut1_37[21] , \nOut1_37[20] , \nOut1_37[19] , \nOut1_37[18] , 
        \nOut1_37[17] , \nOut1_37[16] , \nOut1_37[15] , \nOut1_37[14] , 
        \nOut1_37[13] , \nOut1_37[12] , \nOut1_37[11] , \nOut1_37[10] , 
        \nOut1_37[9] , \nOut1_37[8] , \nOut1_37[7] , \nOut1_37[6] , 
        \nOut1_37[5] , \nOut1_37[4] , \nOut1_37[3] , \nOut1_37[2] , 
        \nOut1_37[1] , \nOut1_37[0] }), .SOUTH_EDGE({\nOut1_39[31] , 
        \nOut1_39[30] , \nOut1_39[29] , \nOut1_39[28] , \nOut1_39[27] , 
        \nOut1_39[26] , \nOut1_39[25] , \nOut1_39[24] , \nOut1_39[23] , 
        \nOut1_39[22] , \nOut1_39[21] , \nOut1_39[20] , \nOut1_39[19] , 
        \nOut1_39[18] , \nOut1_39[17] , \nOut1_39[16] , \nOut1_39[15] , 
        \nOut1_39[14] , \nOut1_39[13] , \nOut1_39[12] , \nOut1_39[11] , 
        \nOut1_39[10] , \nOut1_39[9] , \nOut1_39[8] , \nOut1_39[7] , 
        \nOut1_39[6] , \nOut1_39[5] , \nOut1_39[4] , \nOut1_39[3] , 
        \nOut1_39[2] , \nOut1_39[1] , \nOut1_39[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_38[0] ), .NW_EDGE(\nOut0_37[0] ), .SW_EDGE(
        \nOut0_39[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_125 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut126[31] , \nScanOut126[30] , \nScanOut126[29] , 
        \nScanOut126[28] , \nScanOut126[27] , \nScanOut126[26] , 
        \nScanOut126[25] , \nScanOut126[24] , \nScanOut126[23] , 
        \nScanOut126[22] , \nScanOut126[21] , \nScanOut126[20] , 
        \nScanOut126[19] , \nScanOut126[18] , \nScanOut126[17] , 
        \nScanOut126[16] , \nScanOut126[15] , \nScanOut126[14] , 
        \nScanOut126[13] , \nScanOut126[12] , \nScanOut126[11] , 
        \nScanOut126[10] , \nScanOut126[9] , \nScanOut126[8] , 
        \nScanOut126[7] , \nScanOut126[6] , \nScanOut126[5] , \nScanOut126[4] , 
        \nScanOut126[3] , \nScanOut126[2] , \nScanOut126[1] , \nScanOut126[0] 
        }), .ScanOut({\nScanOut125[31] , \nScanOut125[30] , \nScanOut125[29] , 
        \nScanOut125[28] , \nScanOut125[27] , \nScanOut125[26] , 
        \nScanOut125[25] , \nScanOut125[24] , \nScanOut125[23] , 
        \nScanOut125[22] , \nScanOut125[21] , \nScanOut125[20] , 
        \nScanOut125[19] , \nScanOut125[18] , \nScanOut125[17] , 
        \nScanOut125[16] , \nScanOut125[15] , \nScanOut125[14] , 
        \nScanOut125[13] , \nScanOut125[12] , \nScanOut125[11] , 
        \nScanOut125[10] , \nScanOut125[9] , \nScanOut125[8] , 
        \nScanOut125[7] , \nScanOut125[6] , \nScanOut125[5] , \nScanOut125[4] , 
        \nScanOut125[3] , \nScanOut125[2] , \nScanOut125[1] , \nScanOut125[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_61[31] , \nOut1_61[30] , \nOut1_61[29] , 
        \nOut1_61[28] , \nOut1_61[27] , \nOut1_61[26] , \nOut1_61[25] , 
        \nOut1_61[24] , \nOut1_61[23] , \nOut1_61[22] , \nOut1_61[21] , 
        \nOut1_61[20] , \nOut1_61[19] , \nOut1_61[18] , \nOut1_61[17] , 
        \nOut1_61[16] , \nOut1_61[15] , \nOut1_61[14] , \nOut1_61[13] , 
        \nOut1_61[12] , \nOut1_61[11] , \nOut1_61[10] , \nOut1_61[9] , 
        \nOut1_61[8] , \nOut1_61[7] , \nOut1_61[6] , \nOut1_61[5] , 
        \nOut1_61[4] , \nOut1_61[3] , \nOut1_61[2] , \nOut1_61[1] , 
        \nOut1_61[0] }), .NORTH_EDGE({\nOut1_60[31] , \nOut1_60[30] , 
        \nOut1_60[29] , \nOut1_60[28] , \nOut1_60[27] , \nOut1_60[26] , 
        \nOut1_60[25] , \nOut1_60[24] , \nOut1_60[23] , \nOut1_60[22] , 
        \nOut1_60[21] , \nOut1_60[20] , \nOut1_60[19] , \nOut1_60[18] , 
        \nOut1_60[17] , \nOut1_60[16] , \nOut1_60[15] , \nOut1_60[14] , 
        \nOut1_60[13] , \nOut1_60[12] , \nOut1_60[11] , \nOut1_60[10] , 
        \nOut1_60[9] , \nOut1_60[8] , \nOut1_60[7] , \nOut1_60[6] , 
        \nOut1_60[5] , \nOut1_60[4] , \nOut1_60[3] , \nOut1_60[2] , 
        \nOut1_60[1] , \nOut1_60[0] }), .SOUTH_EDGE({\nOut1_62[31] , 
        \nOut1_62[30] , \nOut1_62[29] , \nOut1_62[28] , \nOut1_62[27] , 
        \nOut1_62[26] , \nOut1_62[25] , \nOut1_62[24] , \nOut1_62[23] , 
        \nOut1_62[22] , \nOut1_62[21] , \nOut1_62[20] , \nOut1_62[19] , 
        \nOut1_62[18] , \nOut1_62[17] , \nOut1_62[16] , \nOut1_62[15] , 
        \nOut1_62[14] , \nOut1_62[13] , \nOut1_62[12] , \nOut1_62[11] , 
        \nOut1_62[10] , \nOut1_62[9] , \nOut1_62[8] , \nOut1_62[7] , 
        \nOut1_62[6] , \nOut1_62[5] , \nOut1_62[4] , \nOut1_62[3] , 
        \nOut1_62[2] , \nOut1_62[1] , \nOut1_62[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_61[0] ), .NW_EDGE(\nOut0_60[0] ), .SW_EDGE(
        \nOut0_62[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_21 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut22[31] , \nScanOut22[30] , \nScanOut22[29] , 
        \nScanOut22[28] , \nScanOut22[27] , \nScanOut22[26] , \nScanOut22[25] , 
        \nScanOut22[24] , \nScanOut22[23] , \nScanOut22[22] , \nScanOut22[21] , 
        \nScanOut22[20] , \nScanOut22[19] , \nScanOut22[18] , \nScanOut22[17] , 
        \nScanOut22[16] , \nScanOut22[15] , \nScanOut22[14] , \nScanOut22[13] , 
        \nScanOut22[12] , \nScanOut22[11] , \nScanOut22[10] , \nScanOut22[9] , 
        \nScanOut22[8] , \nScanOut22[7] , \nScanOut22[6] , \nScanOut22[5] , 
        \nScanOut22[4] , \nScanOut22[3] , \nScanOut22[2] , \nScanOut22[1] , 
        \nScanOut22[0] }), .ScanOut({\nScanOut21[31] , \nScanOut21[30] , 
        \nScanOut21[29] , \nScanOut21[28] , \nScanOut21[27] , \nScanOut21[26] , 
        \nScanOut21[25] , \nScanOut21[24] , \nScanOut21[23] , \nScanOut21[22] , 
        \nScanOut21[21] , \nScanOut21[20] , \nScanOut21[19] , \nScanOut21[18] , 
        \nScanOut21[17] , \nScanOut21[16] , \nScanOut21[15] , \nScanOut21[14] , 
        \nScanOut21[13] , \nScanOut21[12] , \nScanOut21[11] , \nScanOut21[10] , 
        \nScanOut21[9] , \nScanOut21[8] , \nScanOut21[7] , \nScanOut21[6] , 
        \nScanOut21[5] , \nScanOut21[4] , \nScanOut21[3] , \nScanOut21[2] , 
        \nScanOut21[1] , \nScanOut21[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_21[31] , 
        \nOut0_21[30] , \nOut0_21[29] , \nOut0_21[28] , \nOut0_21[27] , 
        \nOut0_21[26] , \nOut0_21[25] , \nOut0_21[24] , \nOut0_21[23] , 
        \nOut0_21[22] , \nOut0_21[21] , \nOut0_21[20] , \nOut0_21[19] , 
        \nOut0_21[18] , \nOut0_21[17] , \nOut0_21[16] , \nOut0_21[15] , 
        \nOut0_21[14] , \nOut0_21[13] , \nOut0_21[12] , \nOut0_21[11] , 
        \nOut0_21[10] , \nOut0_21[9] , \nOut0_21[8] , \nOut0_21[7] , 
        \nOut0_21[6] , \nOut0_21[5] , \nOut0_21[4] , \nOut0_21[3] , 
        \nOut0_21[2] , \nOut0_21[1] , \nOut0_21[0] }), .NORTH_EDGE({
        \nOut0_20[31] , \nOut0_20[30] , \nOut0_20[29] , \nOut0_20[28] , 
        \nOut0_20[27] , \nOut0_20[26] , \nOut0_20[25] , \nOut0_20[24] , 
        \nOut0_20[23] , \nOut0_20[22] , \nOut0_20[21] , \nOut0_20[20] , 
        \nOut0_20[19] , \nOut0_20[18] , \nOut0_20[17] , \nOut0_20[16] , 
        \nOut0_20[15] , \nOut0_20[14] , \nOut0_20[13] , \nOut0_20[12] , 
        \nOut0_20[11] , \nOut0_20[10] , \nOut0_20[9] , \nOut0_20[8] , 
        \nOut0_20[7] , \nOut0_20[6] , \nOut0_20[5] , \nOut0_20[4] , 
        \nOut0_20[3] , \nOut0_20[2] , \nOut0_20[1] , \nOut0_20[0] }), 
        .SOUTH_EDGE({\nOut0_22[31] , \nOut0_22[30] , \nOut0_22[29] , 
        \nOut0_22[28] , \nOut0_22[27] , \nOut0_22[26] , \nOut0_22[25] , 
        \nOut0_22[24] , \nOut0_22[23] , \nOut0_22[22] , \nOut0_22[21] , 
        \nOut0_22[20] , \nOut0_22[19] , \nOut0_22[18] , \nOut0_22[17] , 
        \nOut0_22[16] , \nOut0_22[15] , \nOut0_22[14] , \nOut0_22[13] , 
        \nOut0_22[12] , \nOut0_22[11] , \nOut0_22[10] , \nOut0_22[9] , 
        \nOut0_22[8] , \nOut0_22[7] , \nOut0_22[6] , \nOut0_22[5] , 
        \nOut0_22[4] , \nOut0_22[3] , \nOut0_22[2] , \nOut0_22[1] , 
        \nOut0_22[0] }), .EAST_EDGE(\nOut1_21[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_20[31] ), .SE_EDGE(
        \nOut1_22[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_68 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut69[31] , \nScanOut69[30] , \nScanOut69[29] , 
        \nScanOut69[28] , \nScanOut69[27] , \nScanOut69[26] , \nScanOut69[25] , 
        \nScanOut69[24] , \nScanOut69[23] , \nScanOut69[22] , \nScanOut69[21] , 
        \nScanOut69[20] , \nScanOut69[19] , \nScanOut69[18] , \nScanOut69[17] , 
        \nScanOut69[16] , \nScanOut69[15] , \nScanOut69[14] , \nScanOut69[13] , 
        \nScanOut69[12] , \nScanOut69[11] , \nScanOut69[10] , \nScanOut69[9] , 
        \nScanOut69[8] , \nScanOut69[7] , \nScanOut69[6] , \nScanOut69[5] , 
        \nScanOut69[4] , \nScanOut69[3] , \nScanOut69[2] , \nScanOut69[1] , 
        \nScanOut69[0] }), .ScanOut({\nScanOut68[31] , \nScanOut68[30] , 
        \nScanOut68[29] , \nScanOut68[28] , \nScanOut68[27] , \nScanOut68[26] , 
        \nScanOut68[25] , \nScanOut68[24] , \nScanOut68[23] , \nScanOut68[22] , 
        \nScanOut68[21] , \nScanOut68[20] , \nScanOut68[19] , \nScanOut68[18] , 
        \nScanOut68[17] , \nScanOut68[16] , \nScanOut68[15] , \nScanOut68[14] , 
        \nScanOut68[13] , \nScanOut68[12] , \nScanOut68[11] , \nScanOut68[10] , 
        \nScanOut68[9] , \nScanOut68[8] , \nScanOut68[7] , \nScanOut68[6] , 
        \nScanOut68[5] , \nScanOut68[4] , \nScanOut68[3] , \nScanOut68[2] , 
        \nScanOut68[1] , \nScanOut68[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_4[31] , 
        \nOut1_4[30] , \nOut1_4[29] , \nOut1_4[28] , \nOut1_4[27] , 
        \nOut1_4[26] , \nOut1_4[25] , \nOut1_4[24] , \nOut1_4[23] , 
        \nOut1_4[22] , \nOut1_4[21] , \nOut1_4[20] , \nOut1_4[19] , 
        \nOut1_4[18] , \nOut1_4[17] , \nOut1_4[16] , \nOut1_4[15] , 
        \nOut1_4[14] , \nOut1_4[13] , \nOut1_4[12] , \nOut1_4[11] , 
        \nOut1_4[10] , \nOut1_4[9] , \nOut1_4[8] , \nOut1_4[7] , \nOut1_4[6] , 
        \nOut1_4[5] , \nOut1_4[4] , \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , 
        \nOut1_4[0] }), .NORTH_EDGE({\nOut1_3[31] , \nOut1_3[30] , 
        \nOut1_3[29] , \nOut1_3[28] , \nOut1_3[27] , \nOut1_3[26] , 
        \nOut1_3[25] , \nOut1_3[24] , \nOut1_3[23] , \nOut1_3[22] , 
        \nOut1_3[21] , \nOut1_3[20] , \nOut1_3[19] , \nOut1_3[18] , 
        \nOut1_3[17] , \nOut1_3[16] , \nOut1_3[15] , \nOut1_3[14] , 
        \nOut1_3[13] , \nOut1_3[12] , \nOut1_3[11] , \nOut1_3[10] , 
        \nOut1_3[9] , \nOut1_3[8] , \nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , 
        \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }), 
        .SOUTH_EDGE({\nOut1_5[31] , \nOut1_5[30] , \nOut1_5[29] , 
        \nOut1_5[28] , \nOut1_5[27] , \nOut1_5[26] , \nOut1_5[25] , 
        \nOut1_5[24] , \nOut1_5[23] , \nOut1_5[22] , \nOut1_5[21] , 
        \nOut1_5[20] , \nOut1_5[19] , \nOut1_5[18] , \nOut1_5[17] , 
        \nOut1_5[16] , \nOut1_5[15] , \nOut1_5[14] , \nOut1_5[13] , 
        \nOut1_5[12] , \nOut1_5[11] , \nOut1_5[10] , \nOut1_5[9] , 
        \nOut1_5[8] , \nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , \nOut1_5[4] , 
        \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_4[0] ), .NW_EDGE(\nOut0_3[0] ), .SW_EDGE(
        \nOut0_5[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_119 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut120[31] , \nScanOut120[30] , \nScanOut120[29] , 
        \nScanOut120[28] , \nScanOut120[27] , \nScanOut120[26] , 
        \nScanOut120[25] , \nScanOut120[24] , \nScanOut120[23] , 
        \nScanOut120[22] , \nScanOut120[21] , \nScanOut120[20] , 
        \nScanOut120[19] , \nScanOut120[18] , \nScanOut120[17] , 
        \nScanOut120[16] , \nScanOut120[15] , \nScanOut120[14] , 
        \nScanOut120[13] , \nScanOut120[12] , \nScanOut120[11] , 
        \nScanOut120[10] , \nScanOut120[9] , \nScanOut120[8] , 
        \nScanOut120[7] , \nScanOut120[6] , \nScanOut120[5] , \nScanOut120[4] , 
        \nScanOut120[3] , \nScanOut120[2] , \nScanOut120[1] , \nScanOut120[0] 
        }), .ScanOut({\nScanOut119[31] , \nScanOut119[30] , \nScanOut119[29] , 
        \nScanOut119[28] , \nScanOut119[27] , \nScanOut119[26] , 
        \nScanOut119[25] , \nScanOut119[24] , \nScanOut119[23] , 
        \nScanOut119[22] , \nScanOut119[21] , \nScanOut119[20] , 
        \nScanOut119[19] , \nScanOut119[18] , \nScanOut119[17] , 
        \nScanOut119[16] , \nScanOut119[15] , \nScanOut119[14] , 
        \nScanOut119[13] , \nScanOut119[12] , \nScanOut119[11] , 
        \nScanOut119[10] , \nScanOut119[9] , \nScanOut119[8] , 
        \nScanOut119[7] , \nScanOut119[6] , \nScanOut119[5] , \nScanOut119[4] , 
        \nScanOut119[3] , \nScanOut119[2] , \nScanOut119[1] , \nScanOut119[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_55[31] , \nOut1_55[30] , \nOut1_55[29] , 
        \nOut1_55[28] , \nOut1_55[27] , \nOut1_55[26] , \nOut1_55[25] , 
        \nOut1_55[24] , \nOut1_55[23] , \nOut1_55[22] , \nOut1_55[21] , 
        \nOut1_55[20] , \nOut1_55[19] , \nOut1_55[18] , \nOut1_55[17] , 
        \nOut1_55[16] , \nOut1_55[15] , \nOut1_55[14] , \nOut1_55[13] , 
        \nOut1_55[12] , \nOut1_55[11] , \nOut1_55[10] , \nOut1_55[9] , 
        \nOut1_55[8] , \nOut1_55[7] , \nOut1_55[6] , \nOut1_55[5] , 
        \nOut1_55[4] , \nOut1_55[3] , \nOut1_55[2] , \nOut1_55[1] , 
        \nOut1_55[0] }), .NORTH_EDGE({\nOut1_54[31] , \nOut1_54[30] , 
        \nOut1_54[29] , \nOut1_54[28] , \nOut1_54[27] , \nOut1_54[26] , 
        \nOut1_54[25] , \nOut1_54[24] , \nOut1_54[23] , \nOut1_54[22] , 
        \nOut1_54[21] , \nOut1_54[20] , \nOut1_54[19] , \nOut1_54[18] , 
        \nOut1_54[17] , \nOut1_54[16] , \nOut1_54[15] , \nOut1_54[14] , 
        \nOut1_54[13] , \nOut1_54[12] , \nOut1_54[11] , \nOut1_54[10] , 
        \nOut1_54[9] , \nOut1_54[8] , \nOut1_54[7] , \nOut1_54[6] , 
        \nOut1_54[5] , \nOut1_54[4] , \nOut1_54[3] , \nOut1_54[2] , 
        \nOut1_54[1] , \nOut1_54[0] }), .SOUTH_EDGE({\nOut1_56[31] , 
        \nOut1_56[30] , \nOut1_56[29] , \nOut1_56[28] , \nOut1_56[27] , 
        \nOut1_56[26] , \nOut1_56[25] , \nOut1_56[24] , \nOut1_56[23] , 
        \nOut1_56[22] , \nOut1_56[21] , \nOut1_56[20] , \nOut1_56[19] , 
        \nOut1_56[18] , \nOut1_56[17] , \nOut1_56[16] , \nOut1_56[15] , 
        \nOut1_56[14] , \nOut1_56[13] , \nOut1_56[12] , \nOut1_56[11] , 
        \nOut1_56[10] , \nOut1_56[9] , \nOut1_56[8] , \nOut1_56[7] , 
        \nOut1_56[6] , \nOut1_56[5] , \nOut1_56[4] , \nOut1_56[3] , 
        \nOut1_56[2] , \nOut1_56[1] , \nOut1_56[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_55[0] ), .NW_EDGE(\nOut0_54[0] ), .SW_EDGE(
        \nOut0_56[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut1[31] , \nScanOut1[30] , \nScanOut1[29] , 
        \nScanOut1[28] , \nScanOut1[27] , \nScanOut1[26] , \nScanOut1[25] , 
        \nScanOut1[24] , \nScanOut1[23] , \nScanOut1[22] , \nScanOut1[21] , 
        \nScanOut1[20] , \nScanOut1[19] , \nScanOut1[18] , \nScanOut1[17] , 
        \nScanOut1[16] , \nScanOut1[15] , \nScanOut1[14] , \nScanOut1[13] , 
        \nScanOut1[12] , \nScanOut1[11] , \nScanOut1[10] , \nScanOut1[9] , 
        \nScanOut1[8] , \nScanOut1[7] , \nScanOut1[6] , \nScanOut1[5] , 
        \nScanOut1[4] , \nScanOut1[3] , \nScanOut1[2] , \nScanOut1[1] , 
        \nScanOut1[0] }), .ScanOut({\nScanOut0[31] , \nScanOut0[30] , 
        \nScanOut0[29] , \nScanOut0[28] , \nScanOut0[27] , \nScanOut0[26] , 
        \nScanOut0[25] , \nScanOut0[24] , \nScanOut0[23] , \nScanOut0[22] , 
        \nScanOut0[21] , \nScanOut0[20] , \nScanOut0[19] , \nScanOut0[18] , 
        \nScanOut0[17] , \nScanOut0[16] , \nScanOut0[15] , \nScanOut0[14] , 
        \nScanOut0[13] , \nScanOut0[12] , \nScanOut0[11] , \nScanOut0[10] , 
        \nScanOut0[9] , \nScanOut0[8] , \nScanOut0[7] , \nScanOut0[6] , 
        \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , \nScanOut0[2] , 
        \nScanOut0[1] , \nScanOut0[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_0[31] , 
        \nOut0_0[30] , \nOut0_0[29] , \nOut0_0[28] , \nOut0_0[27] , 
        \nOut0_0[26] , \nOut0_0[25] , \nOut0_0[24] , \nOut0_0[23] , 
        \nOut0_0[22] , \nOut0_0[21] , \nOut0_0[20] , \nOut0_0[19] , 
        \nOut0_0[18] , \nOut0_0[17] , \nOut0_0[16] , \nOut0_0[15] , 
        \nOut0_0[14] , \nOut0_0[13] , \nOut0_0[12] , \nOut0_0[11] , 
        \nOut0_0[10] , \nOut0_0[9] , \nOut0_0[8] , \nOut0_0[7] , \nOut0_0[6] , 
        \nOut0_0[5] , \nOut0_0[4] , \nOut0_0[3] , \nOut0_0[2] , \nOut0_0[1] , 
        \nOut0_0[0] }), .NORTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .SOUTH_EDGE({\nOut0_1[31] , \nOut0_1[30] , \nOut0_1[29] , 
        \nOut0_1[28] , \nOut0_1[27] , \nOut0_1[26] , \nOut0_1[25] , 
        \nOut0_1[24] , \nOut0_1[23] , \nOut0_1[22] , \nOut0_1[21] , 
        \nOut0_1[20] , \nOut0_1[19] , \nOut0_1[18] , \nOut0_1[17] , 
        \nOut0_1[16] , \nOut0_1[15] , \nOut0_1[14] , \nOut0_1[13] , 
        \nOut0_1[12] , \nOut0_1[11] , \nOut0_1[10] , \nOut0_1[9] , 
        \nOut0_1[8] , \nOut0_1[7] , \nOut0_1[6] , \nOut0_1[5] , \nOut0_1[4] , 
        \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , \nOut0_1[0] }), .EAST_EDGE(
        \nOut1_0[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(1'b0), .SE_EDGE(\nOut1_1[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut3[31] , \nScanOut3[30] , \nScanOut3[29] , 
        \nScanOut3[28] , \nScanOut3[27] , \nScanOut3[26] , \nScanOut3[25] , 
        \nScanOut3[24] , \nScanOut3[23] , \nScanOut3[22] , \nScanOut3[21] , 
        \nScanOut3[20] , \nScanOut3[19] , \nScanOut3[18] , \nScanOut3[17] , 
        \nScanOut3[16] , \nScanOut3[15] , \nScanOut3[14] , \nScanOut3[13] , 
        \nScanOut3[12] , \nScanOut3[11] , \nScanOut3[10] , \nScanOut3[9] , 
        \nScanOut3[8] , \nScanOut3[7] , \nScanOut3[6] , \nScanOut3[5] , 
        \nScanOut3[4] , \nScanOut3[3] , \nScanOut3[2] , \nScanOut3[1] , 
        \nScanOut3[0] }), .ScanOut({\nScanOut2[31] , \nScanOut2[30] , 
        \nScanOut2[29] , \nScanOut2[28] , \nScanOut2[27] , \nScanOut2[26] , 
        \nScanOut2[25] , \nScanOut2[24] , \nScanOut2[23] , \nScanOut2[22] , 
        \nScanOut2[21] , \nScanOut2[20] , \nScanOut2[19] , \nScanOut2[18] , 
        \nScanOut2[17] , \nScanOut2[16] , \nScanOut2[15] , \nScanOut2[14] , 
        \nScanOut2[13] , \nScanOut2[12] , \nScanOut2[11] , \nScanOut2[10] , 
        \nScanOut2[9] , \nScanOut2[8] , \nScanOut2[7] , \nScanOut2[6] , 
        \nScanOut2[5] , \nScanOut2[4] , \nScanOut2[3] , \nScanOut2[2] , 
        \nScanOut2[1] , \nScanOut2[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_2[31] , 
        \nOut0_2[30] , \nOut0_2[29] , \nOut0_2[28] , \nOut0_2[27] , 
        \nOut0_2[26] , \nOut0_2[25] , \nOut0_2[24] , \nOut0_2[23] , 
        \nOut0_2[22] , \nOut0_2[21] , \nOut0_2[20] , \nOut0_2[19] , 
        \nOut0_2[18] , \nOut0_2[17] , \nOut0_2[16] , \nOut0_2[15] , 
        \nOut0_2[14] , \nOut0_2[13] , \nOut0_2[12] , \nOut0_2[11] , 
        \nOut0_2[10] , \nOut0_2[9] , \nOut0_2[8] , \nOut0_2[7] , \nOut0_2[6] , 
        \nOut0_2[5] , \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , 
        \nOut0_2[0] }), .NORTH_EDGE({\nOut0_1[31] , \nOut0_1[30] , 
        \nOut0_1[29] , \nOut0_1[28] , \nOut0_1[27] , \nOut0_1[26] , 
        \nOut0_1[25] , \nOut0_1[24] , \nOut0_1[23] , \nOut0_1[22] , 
        \nOut0_1[21] , \nOut0_1[20] , \nOut0_1[19] , \nOut0_1[18] , 
        \nOut0_1[17] , \nOut0_1[16] , \nOut0_1[15] , \nOut0_1[14] , 
        \nOut0_1[13] , \nOut0_1[12] , \nOut0_1[11] , \nOut0_1[10] , 
        \nOut0_1[9] , \nOut0_1[8] , \nOut0_1[7] , \nOut0_1[6] , \nOut0_1[5] , 
        \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , \nOut0_1[0] }), 
        .SOUTH_EDGE({\nOut0_3[31] , \nOut0_3[30] , \nOut0_3[29] , 
        \nOut0_3[28] , \nOut0_3[27] , \nOut0_3[26] , \nOut0_3[25] , 
        \nOut0_3[24] , \nOut0_3[23] , \nOut0_3[22] , \nOut0_3[21] , 
        \nOut0_3[20] , \nOut0_3[19] , \nOut0_3[18] , \nOut0_3[17] , 
        \nOut0_3[16] , \nOut0_3[15] , \nOut0_3[14] , \nOut0_3[13] , 
        \nOut0_3[12] , \nOut0_3[11] , \nOut0_3[10] , \nOut0_3[9] , 
        \nOut0_3[8] , \nOut0_3[7] , \nOut0_3[6] , \nOut0_3[5] , \nOut0_3[4] , 
        \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , \nOut0_3[0] }), .EAST_EDGE(
        \nOut1_2[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_1[31] ), .SE_EDGE(\nOut1_3[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut5[31] , \nScanOut5[30] , \nScanOut5[29] , 
        \nScanOut5[28] , \nScanOut5[27] , \nScanOut5[26] , \nScanOut5[25] , 
        \nScanOut5[24] , \nScanOut5[23] , \nScanOut5[22] , \nScanOut5[21] , 
        \nScanOut5[20] , \nScanOut5[19] , \nScanOut5[18] , \nScanOut5[17] , 
        \nScanOut5[16] , \nScanOut5[15] , \nScanOut5[14] , \nScanOut5[13] , 
        \nScanOut5[12] , \nScanOut5[11] , \nScanOut5[10] , \nScanOut5[9] , 
        \nScanOut5[8] , \nScanOut5[7] , \nScanOut5[6] , \nScanOut5[5] , 
        \nScanOut5[4] , \nScanOut5[3] , \nScanOut5[2] , \nScanOut5[1] , 
        \nScanOut5[0] }), .ScanOut({\nScanOut4[31] , \nScanOut4[30] , 
        \nScanOut4[29] , \nScanOut4[28] , \nScanOut4[27] , \nScanOut4[26] , 
        \nScanOut4[25] , \nScanOut4[24] , \nScanOut4[23] , \nScanOut4[22] , 
        \nScanOut4[21] , \nScanOut4[20] , \nScanOut4[19] , \nScanOut4[18] , 
        \nScanOut4[17] , \nScanOut4[16] , \nScanOut4[15] , \nScanOut4[14] , 
        \nScanOut4[13] , \nScanOut4[12] , \nScanOut4[11] , \nScanOut4[10] , 
        \nScanOut4[9] , \nScanOut4[8] , \nScanOut4[7] , \nScanOut4[6] , 
        \nScanOut4[5] , \nScanOut4[4] , \nScanOut4[3] , \nScanOut4[2] , 
        \nScanOut4[1] , \nScanOut4[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_4[31] , 
        \nOut0_4[30] , \nOut0_4[29] , \nOut0_4[28] , \nOut0_4[27] , 
        \nOut0_4[26] , \nOut0_4[25] , \nOut0_4[24] , \nOut0_4[23] , 
        \nOut0_4[22] , \nOut0_4[21] , \nOut0_4[20] , \nOut0_4[19] , 
        \nOut0_4[18] , \nOut0_4[17] , \nOut0_4[16] , \nOut0_4[15] , 
        \nOut0_4[14] , \nOut0_4[13] , \nOut0_4[12] , \nOut0_4[11] , 
        \nOut0_4[10] , \nOut0_4[9] , \nOut0_4[8] , \nOut0_4[7] , \nOut0_4[6] , 
        \nOut0_4[5] , \nOut0_4[4] , \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , 
        \nOut0_4[0] }), .NORTH_EDGE({\nOut0_3[31] , \nOut0_3[30] , 
        \nOut0_3[29] , \nOut0_3[28] , \nOut0_3[27] , \nOut0_3[26] , 
        \nOut0_3[25] , \nOut0_3[24] , \nOut0_3[23] , \nOut0_3[22] , 
        \nOut0_3[21] , \nOut0_3[20] , \nOut0_3[19] , \nOut0_3[18] , 
        \nOut0_3[17] , \nOut0_3[16] , \nOut0_3[15] , \nOut0_3[14] , 
        \nOut0_3[13] , \nOut0_3[12] , \nOut0_3[11] , \nOut0_3[10] , 
        \nOut0_3[9] , \nOut0_3[8] , \nOut0_3[7] , \nOut0_3[6] , \nOut0_3[5] , 
        \nOut0_3[4] , \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , \nOut0_3[0] }), 
        .SOUTH_EDGE({\nOut0_5[31] , \nOut0_5[30] , \nOut0_5[29] , 
        \nOut0_5[28] , \nOut0_5[27] , \nOut0_5[26] , \nOut0_5[25] , 
        \nOut0_5[24] , \nOut0_5[23] , \nOut0_5[22] , \nOut0_5[21] , 
        \nOut0_5[20] , \nOut0_5[19] , \nOut0_5[18] , \nOut0_5[17] , 
        \nOut0_5[16] , \nOut0_5[15] , \nOut0_5[14] , \nOut0_5[13] , 
        \nOut0_5[12] , \nOut0_5[11] , \nOut0_5[10] , \nOut0_5[9] , 
        \nOut0_5[8] , \nOut0_5[7] , \nOut0_5[6] , \nOut0_5[5] , \nOut0_5[4] , 
        \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , \nOut0_5[0] }), .EAST_EDGE(
        \nOut1_4[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_3[31] ), .SE_EDGE(\nOut1_5[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut14[31] , \nScanOut14[30] , \nScanOut14[29] , 
        \nScanOut14[28] , \nScanOut14[27] , \nScanOut14[26] , \nScanOut14[25] , 
        \nScanOut14[24] , \nScanOut14[23] , \nScanOut14[22] , \nScanOut14[21] , 
        \nScanOut14[20] , \nScanOut14[19] , \nScanOut14[18] , \nScanOut14[17] , 
        \nScanOut14[16] , \nScanOut14[15] , \nScanOut14[14] , \nScanOut14[13] , 
        \nScanOut14[12] , \nScanOut14[11] , \nScanOut14[10] , \nScanOut14[9] , 
        \nScanOut14[8] , \nScanOut14[7] , \nScanOut14[6] , \nScanOut14[5] , 
        \nScanOut14[4] , \nScanOut14[3] , \nScanOut14[2] , \nScanOut14[1] , 
        \nScanOut14[0] }), .ScanOut({\nScanOut13[31] , \nScanOut13[30] , 
        \nScanOut13[29] , \nScanOut13[28] , \nScanOut13[27] , \nScanOut13[26] , 
        \nScanOut13[25] , \nScanOut13[24] , \nScanOut13[23] , \nScanOut13[22] , 
        \nScanOut13[21] , \nScanOut13[20] , \nScanOut13[19] , \nScanOut13[18] , 
        \nScanOut13[17] , \nScanOut13[16] , \nScanOut13[15] , \nScanOut13[14] , 
        \nScanOut13[13] , \nScanOut13[12] , \nScanOut13[11] , \nScanOut13[10] , 
        \nScanOut13[9] , \nScanOut13[8] , \nScanOut13[7] , \nScanOut13[6] , 
        \nScanOut13[5] , \nScanOut13[4] , \nScanOut13[3] , \nScanOut13[2] , 
        \nScanOut13[1] , \nScanOut13[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_13[31] , 
        \nOut0_13[30] , \nOut0_13[29] , \nOut0_13[28] , \nOut0_13[27] , 
        \nOut0_13[26] , \nOut0_13[25] , \nOut0_13[24] , \nOut0_13[23] , 
        \nOut0_13[22] , \nOut0_13[21] , \nOut0_13[20] , \nOut0_13[19] , 
        \nOut0_13[18] , \nOut0_13[17] , \nOut0_13[16] , \nOut0_13[15] , 
        \nOut0_13[14] , \nOut0_13[13] , \nOut0_13[12] , \nOut0_13[11] , 
        \nOut0_13[10] , \nOut0_13[9] , \nOut0_13[8] , \nOut0_13[7] , 
        \nOut0_13[6] , \nOut0_13[5] , \nOut0_13[4] , \nOut0_13[3] , 
        \nOut0_13[2] , \nOut0_13[1] , \nOut0_13[0] }), .NORTH_EDGE({
        \nOut0_12[31] , \nOut0_12[30] , \nOut0_12[29] , \nOut0_12[28] , 
        \nOut0_12[27] , \nOut0_12[26] , \nOut0_12[25] , \nOut0_12[24] , 
        \nOut0_12[23] , \nOut0_12[22] , \nOut0_12[21] , \nOut0_12[20] , 
        \nOut0_12[19] , \nOut0_12[18] , \nOut0_12[17] , \nOut0_12[16] , 
        \nOut0_12[15] , \nOut0_12[14] , \nOut0_12[13] , \nOut0_12[12] , 
        \nOut0_12[11] , \nOut0_12[10] , \nOut0_12[9] , \nOut0_12[8] , 
        \nOut0_12[7] , \nOut0_12[6] , \nOut0_12[5] , \nOut0_12[4] , 
        \nOut0_12[3] , \nOut0_12[2] , \nOut0_12[1] , \nOut0_12[0] }), 
        .SOUTH_EDGE({\nOut0_14[31] , \nOut0_14[30] , \nOut0_14[29] , 
        \nOut0_14[28] , \nOut0_14[27] , \nOut0_14[26] , \nOut0_14[25] , 
        \nOut0_14[24] , \nOut0_14[23] , \nOut0_14[22] , \nOut0_14[21] , 
        \nOut0_14[20] , \nOut0_14[19] , \nOut0_14[18] , \nOut0_14[17] , 
        \nOut0_14[16] , \nOut0_14[15] , \nOut0_14[14] , \nOut0_14[13] , 
        \nOut0_14[12] , \nOut0_14[11] , \nOut0_14[10] , \nOut0_14[9] , 
        \nOut0_14[8] , \nOut0_14[7] , \nOut0_14[6] , \nOut0_14[5] , 
        \nOut0_14[4] , \nOut0_14[3] , \nOut0_14[2] , \nOut0_14[1] , 
        \nOut0_14[0] }), .EAST_EDGE(\nOut1_13[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_12[31] ), .SE_EDGE(
        \nOut1_14[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut15[31] , \nScanOut15[30] , \nScanOut15[29] , 
        \nScanOut15[28] , \nScanOut15[27] , \nScanOut15[26] , \nScanOut15[25] , 
        \nScanOut15[24] , \nScanOut15[23] , \nScanOut15[22] , \nScanOut15[21] , 
        \nScanOut15[20] , \nScanOut15[19] , \nScanOut15[18] , \nScanOut15[17] , 
        \nScanOut15[16] , \nScanOut15[15] , \nScanOut15[14] , \nScanOut15[13] , 
        \nScanOut15[12] , \nScanOut15[11] , \nScanOut15[10] , \nScanOut15[9] , 
        \nScanOut15[8] , \nScanOut15[7] , \nScanOut15[6] , \nScanOut15[5] , 
        \nScanOut15[4] , \nScanOut15[3] , \nScanOut15[2] , \nScanOut15[1] , 
        \nScanOut15[0] }), .ScanOut({\nScanOut14[31] , \nScanOut14[30] , 
        \nScanOut14[29] , \nScanOut14[28] , \nScanOut14[27] , \nScanOut14[26] , 
        \nScanOut14[25] , \nScanOut14[24] , \nScanOut14[23] , \nScanOut14[22] , 
        \nScanOut14[21] , \nScanOut14[20] , \nScanOut14[19] , \nScanOut14[18] , 
        \nScanOut14[17] , \nScanOut14[16] , \nScanOut14[15] , \nScanOut14[14] , 
        \nScanOut14[13] , \nScanOut14[12] , \nScanOut14[11] , \nScanOut14[10] , 
        \nScanOut14[9] , \nScanOut14[8] , \nScanOut14[7] , \nScanOut14[6] , 
        \nScanOut14[5] , \nScanOut14[4] , \nScanOut14[3] , \nScanOut14[2] , 
        \nScanOut14[1] , \nScanOut14[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_14[31] , 
        \nOut0_14[30] , \nOut0_14[29] , \nOut0_14[28] , \nOut0_14[27] , 
        \nOut0_14[26] , \nOut0_14[25] , \nOut0_14[24] , \nOut0_14[23] , 
        \nOut0_14[22] , \nOut0_14[21] , \nOut0_14[20] , \nOut0_14[19] , 
        \nOut0_14[18] , \nOut0_14[17] , \nOut0_14[16] , \nOut0_14[15] , 
        \nOut0_14[14] , \nOut0_14[13] , \nOut0_14[12] , \nOut0_14[11] , 
        \nOut0_14[10] , \nOut0_14[9] , \nOut0_14[8] , \nOut0_14[7] , 
        \nOut0_14[6] , \nOut0_14[5] , \nOut0_14[4] , \nOut0_14[3] , 
        \nOut0_14[2] , \nOut0_14[1] , \nOut0_14[0] }), .NORTH_EDGE({
        \nOut0_13[31] , \nOut0_13[30] , \nOut0_13[29] , \nOut0_13[28] , 
        \nOut0_13[27] , \nOut0_13[26] , \nOut0_13[25] , \nOut0_13[24] , 
        \nOut0_13[23] , \nOut0_13[22] , \nOut0_13[21] , \nOut0_13[20] , 
        \nOut0_13[19] , \nOut0_13[18] , \nOut0_13[17] , \nOut0_13[16] , 
        \nOut0_13[15] , \nOut0_13[14] , \nOut0_13[13] , \nOut0_13[12] , 
        \nOut0_13[11] , \nOut0_13[10] , \nOut0_13[9] , \nOut0_13[8] , 
        \nOut0_13[7] , \nOut0_13[6] , \nOut0_13[5] , \nOut0_13[4] , 
        \nOut0_13[3] , \nOut0_13[2] , \nOut0_13[1] , \nOut0_13[0] }), 
        .SOUTH_EDGE({\nOut0_15[31] , \nOut0_15[30] , \nOut0_15[29] , 
        \nOut0_15[28] , \nOut0_15[27] , \nOut0_15[26] , \nOut0_15[25] , 
        \nOut0_15[24] , \nOut0_15[23] , \nOut0_15[22] , \nOut0_15[21] , 
        \nOut0_15[20] , \nOut0_15[19] , \nOut0_15[18] , \nOut0_15[17] , 
        \nOut0_15[16] , \nOut0_15[15] , \nOut0_15[14] , \nOut0_15[13] , 
        \nOut0_15[12] , \nOut0_15[11] , \nOut0_15[10] , \nOut0_15[9] , 
        \nOut0_15[8] , \nOut0_15[7] , \nOut0_15[6] , \nOut0_15[5] , 
        \nOut0_15[4] , \nOut0_15[3] , \nOut0_15[2] , \nOut0_15[1] , 
        \nOut0_15[0] }), .EAST_EDGE(\nOut1_14[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_13[31] ), .SE_EDGE(
        \nOut1_15[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_33 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut34[31] , \nScanOut34[30] , \nScanOut34[29] , 
        \nScanOut34[28] , \nScanOut34[27] , \nScanOut34[26] , \nScanOut34[25] , 
        \nScanOut34[24] , \nScanOut34[23] , \nScanOut34[22] , \nScanOut34[21] , 
        \nScanOut34[20] , \nScanOut34[19] , \nScanOut34[18] , \nScanOut34[17] , 
        \nScanOut34[16] , \nScanOut34[15] , \nScanOut34[14] , \nScanOut34[13] , 
        \nScanOut34[12] , \nScanOut34[11] , \nScanOut34[10] , \nScanOut34[9] , 
        \nScanOut34[8] , \nScanOut34[7] , \nScanOut34[6] , \nScanOut34[5] , 
        \nScanOut34[4] , \nScanOut34[3] , \nScanOut34[2] , \nScanOut34[1] , 
        \nScanOut34[0] }), .ScanOut({\nScanOut33[31] , \nScanOut33[30] , 
        \nScanOut33[29] , \nScanOut33[28] , \nScanOut33[27] , \nScanOut33[26] , 
        \nScanOut33[25] , \nScanOut33[24] , \nScanOut33[23] , \nScanOut33[22] , 
        \nScanOut33[21] , \nScanOut33[20] , \nScanOut33[19] , \nScanOut33[18] , 
        \nScanOut33[17] , \nScanOut33[16] , \nScanOut33[15] , \nScanOut33[14] , 
        \nScanOut33[13] , \nScanOut33[12] , \nScanOut33[11] , \nScanOut33[10] , 
        \nScanOut33[9] , \nScanOut33[8] , \nScanOut33[7] , \nScanOut33[6] , 
        \nScanOut33[5] , \nScanOut33[4] , \nScanOut33[3] , \nScanOut33[2] , 
        \nScanOut33[1] , \nScanOut33[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_33[31] , 
        \nOut0_33[30] , \nOut0_33[29] , \nOut0_33[28] , \nOut0_33[27] , 
        \nOut0_33[26] , \nOut0_33[25] , \nOut0_33[24] , \nOut0_33[23] , 
        \nOut0_33[22] , \nOut0_33[21] , \nOut0_33[20] , \nOut0_33[19] , 
        \nOut0_33[18] , \nOut0_33[17] , \nOut0_33[16] , \nOut0_33[15] , 
        \nOut0_33[14] , \nOut0_33[13] , \nOut0_33[12] , \nOut0_33[11] , 
        \nOut0_33[10] , \nOut0_33[9] , \nOut0_33[8] , \nOut0_33[7] , 
        \nOut0_33[6] , \nOut0_33[5] , \nOut0_33[4] , \nOut0_33[3] , 
        \nOut0_33[2] , \nOut0_33[1] , \nOut0_33[0] }), .NORTH_EDGE({
        \nOut0_32[31] , \nOut0_32[30] , \nOut0_32[29] , \nOut0_32[28] , 
        \nOut0_32[27] , \nOut0_32[26] , \nOut0_32[25] , \nOut0_32[24] , 
        \nOut0_32[23] , \nOut0_32[22] , \nOut0_32[21] , \nOut0_32[20] , 
        \nOut0_32[19] , \nOut0_32[18] , \nOut0_32[17] , \nOut0_32[16] , 
        \nOut0_32[15] , \nOut0_32[14] , \nOut0_32[13] , \nOut0_32[12] , 
        \nOut0_32[11] , \nOut0_32[10] , \nOut0_32[9] , \nOut0_32[8] , 
        \nOut0_32[7] , \nOut0_32[6] , \nOut0_32[5] , \nOut0_32[4] , 
        \nOut0_32[3] , \nOut0_32[2] , \nOut0_32[1] , \nOut0_32[0] }), 
        .SOUTH_EDGE({\nOut0_34[31] , \nOut0_34[30] , \nOut0_34[29] , 
        \nOut0_34[28] , \nOut0_34[27] , \nOut0_34[26] , \nOut0_34[25] , 
        \nOut0_34[24] , \nOut0_34[23] , \nOut0_34[22] , \nOut0_34[21] , 
        \nOut0_34[20] , \nOut0_34[19] , \nOut0_34[18] , \nOut0_34[17] , 
        \nOut0_34[16] , \nOut0_34[15] , \nOut0_34[14] , \nOut0_34[13] , 
        \nOut0_34[12] , \nOut0_34[11] , \nOut0_34[10] , \nOut0_34[9] , 
        \nOut0_34[8] , \nOut0_34[7] , \nOut0_34[6] , \nOut0_34[5] , 
        \nOut0_34[4] , \nOut0_34[3] , \nOut0_34[2] , \nOut0_34[1] , 
        \nOut0_34[0] }), .EAST_EDGE(\nOut1_33[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_32[31] ), .SE_EDGE(
        \nOut1_34[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_28 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut29[31] , \nScanOut29[30] , \nScanOut29[29] , 
        \nScanOut29[28] , \nScanOut29[27] , \nScanOut29[26] , \nScanOut29[25] , 
        \nScanOut29[24] , \nScanOut29[23] , \nScanOut29[22] , \nScanOut29[21] , 
        \nScanOut29[20] , \nScanOut29[19] , \nScanOut29[18] , \nScanOut29[17] , 
        \nScanOut29[16] , \nScanOut29[15] , \nScanOut29[14] , \nScanOut29[13] , 
        \nScanOut29[12] , \nScanOut29[11] , \nScanOut29[10] , \nScanOut29[9] , 
        \nScanOut29[8] , \nScanOut29[7] , \nScanOut29[6] , \nScanOut29[5] , 
        \nScanOut29[4] , \nScanOut29[3] , \nScanOut29[2] , \nScanOut29[1] , 
        \nScanOut29[0] }), .ScanOut({\nScanOut28[31] , \nScanOut28[30] , 
        \nScanOut28[29] , \nScanOut28[28] , \nScanOut28[27] , \nScanOut28[26] , 
        \nScanOut28[25] , \nScanOut28[24] , \nScanOut28[23] , \nScanOut28[22] , 
        \nScanOut28[21] , \nScanOut28[20] , \nScanOut28[19] , \nScanOut28[18] , 
        \nScanOut28[17] , \nScanOut28[16] , \nScanOut28[15] , \nScanOut28[14] , 
        \nScanOut28[13] , \nScanOut28[12] , \nScanOut28[11] , \nScanOut28[10] , 
        \nScanOut28[9] , \nScanOut28[8] , \nScanOut28[7] , \nScanOut28[6] , 
        \nScanOut28[5] , \nScanOut28[4] , \nScanOut28[3] , \nScanOut28[2] , 
        \nScanOut28[1] , \nScanOut28[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_28[31] , 
        \nOut0_28[30] , \nOut0_28[29] , \nOut0_28[28] , \nOut0_28[27] , 
        \nOut0_28[26] , \nOut0_28[25] , \nOut0_28[24] , \nOut0_28[23] , 
        \nOut0_28[22] , \nOut0_28[21] , \nOut0_28[20] , \nOut0_28[19] , 
        \nOut0_28[18] , \nOut0_28[17] , \nOut0_28[16] , \nOut0_28[15] , 
        \nOut0_28[14] , \nOut0_28[13] , \nOut0_28[12] , \nOut0_28[11] , 
        \nOut0_28[10] , \nOut0_28[9] , \nOut0_28[8] , \nOut0_28[7] , 
        \nOut0_28[6] , \nOut0_28[5] , \nOut0_28[4] , \nOut0_28[3] , 
        \nOut0_28[2] , \nOut0_28[1] , \nOut0_28[0] }), .NORTH_EDGE({
        \nOut0_27[31] , \nOut0_27[30] , \nOut0_27[29] , \nOut0_27[28] , 
        \nOut0_27[27] , \nOut0_27[26] , \nOut0_27[25] , \nOut0_27[24] , 
        \nOut0_27[23] , \nOut0_27[22] , \nOut0_27[21] , \nOut0_27[20] , 
        \nOut0_27[19] , \nOut0_27[18] , \nOut0_27[17] , \nOut0_27[16] , 
        \nOut0_27[15] , \nOut0_27[14] , \nOut0_27[13] , \nOut0_27[12] , 
        \nOut0_27[11] , \nOut0_27[10] , \nOut0_27[9] , \nOut0_27[8] , 
        \nOut0_27[7] , \nOut0_27[6] , \nOut0_27[5] , \nOut0_27[4] , 
        \nOut0_27[3] , \nOut0_27[2] , \nOut0_27[1] , \nOut0_27[0] }), 
        .SOUTH_EDGE({\nOut0_29[31] , \nOut0_29[30] , \nOut0_29[29] , 
        \nOut0_29[28] , \nOut0_29[27] , \nOut0_29[26] , \nOut0_29[25] , 
        \nOut0_29[24] , \nOut0_29[23] , \nOut0_29[22] , \nOut0_29[21] , 
        \nOut0_29[20] , \nOut0_29[19] , \nOut0_29[18] , \nOut0_29[17] , 
        \nOut0_29[16] , \nOut0_29[15] , \nOut0_29[14] , \nOut0_29[13] , 
        \nOut0_29[12] , \nOut0_29[11] , \nOut0_29[10] , \nOut0_29[9] , 
        \nOut0_29[8] , \nOut0_29[7] , \nOut0_29[6] , \nOut0_29[5] , 
        \nOut0_29[4] , \nOut0_29[3] , \nOut0_29[2] , \nOut0_29[1] , 
        \nOut0_29[0] }), .EAST_EDGE(\nOut1_28[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_27[31] ), .SE_EDGE(
        \nOut1_29[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_46 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut47[31] , \nScanOut47[30] , \nScanOut47[29] , 
        \nScanOut47[28] , \nScanOut47[27] , \nScanOut47[26] , \nScanOut47[25] , 
        \nScanOut47[24] , \nScanOut47[23] , \nScanOut47[22] , \nScanOut47[21] , 
        \nScanOut47[20] , \nScanOut47[19] , \nScanOut47[18] , \nScanOut47[17] , 
        \nScanOut47[16] , \nScanOut47[15] , \nScanOut47[14] , \nScanOut47[13] , 
        \nScanOut47[12] , \nScanOut47[11] , \nScanOut47[10] , \nScanOut47[9] , 
        \nScanOut47[8] , \nScanOut47[7] , \nScanOut47[6] , \nScanOut47[5] , 
        \nScanOut47[4] , \nScanOut47[3] , \nScanOut47[2] , \nScanOut47[1] , 
        \nScanOut47[0] }), .ScanOut({\nScanOut46[31] , \nScanOut46[30] , 
        \nScanOut46[29] , \nScanOut46[28] , \nScanOut46[27] , \nScanOut46[26] , 
        \nScanOut46[25] , \nScanOut46[24] , \nScanOut46[23] , \nScanOut46[22] , 
        \nScanOut46[21] , \nScanOut46[20] , \nScanOut46[19] , \nScanOut46[18] , 
        \nScanOut46[17] , \nScanOut46[16] , \nScanOut46[15] , \nScanOut46[14] , 
        \nScanOut46[13] , \nScanOut46[12] , \nScanOut46[11] , \nScanOut46[10] , 
        \nScanOut46[9] , \nScanOut46[8] , \nScanOut46[7] , \nScanOut46[6] , 
        \nScanOut46[5] , \nScanOut46[4] , \nScanOut46[3] , \nScanOut46[2] , 
        \nScanOut46[1] , \nScanOut46[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_46[31] , 
        \nOut0_46[30] , \nOut0_46[29] , \nOut0_46[28] , \nOut0_46[27] , 
        \nOut0_46[26] , \nOut0_46[25] , \nOut0_46[24] , \nOut0_46[23] , 
        \nOut0_46[22] , \nOut0_46[21] , \nOut0_46[20] , \nOut0_46[19] , 
        \nOut0_46[18] , \nOut0_46[17] , \nOut0_46[16] , \nOut0_46[15] , 
        \nOut0_46[14] , \nOut0_46[13] , \nOut0_46[12] , \nOut0_46[11] , 
        \nOut0_46[10] , \nOut0_46[9] , \nOut0_46[8] , \nOut0_46[7] , 
        \nOut0_46[6] , \nOut0_46[5] , \nOut0_46[4] , \nOut0_46[3] , 
        \nOut0_46[2] , \nOut0_46[1] , \nOut0_46[0] }), .NORTH_EDGE({
        \nOut0_45[31] , \nOut0_45[30] , \nOut0_45[29] , \nOut0_45[28] , 
        \nOut0_45[27] , \nOut0_45[26] , \nOut0_45[25] , \nOut0_45[24] , 
        \nOut0_45[23] , \nOut0_45[22] , \nOut0_45[21] , \nOut0_45[20] , 
        \nOut0_45[19] , \nOut0_45[18] , \nOut0_45[17] , \nOut0_45[16] , 
        \nOut0_45[15] , \nOut0_45[14] , \nOut0_45[13] , \nOut0_45[12] , 
        \nOut0_45[11] , \nOut0_45[10] , \nOut0_45[9] , \nOut0_45[8] , 
        \nOut0_45[7] , \nOut0_45[6] , \nOut0_45[5] , \nOut0_45[4] , 
        \nOut0_45[3] , \nOut0_45[2] , \nOut0_45[1] , \nOut0_45[0] }), 
        .SOUTH_EDGE({\nOut0_47[31] , \nOut0_47[30] , \nOut0_47[29] , 
        \nOut0_47[28] , \nOut0_47[27] , \nOut0_47[26] , \nOut0_47[25] , 
        \nOut0_47[24] , \nOut0_47[23] , \nOut0_47[22] , \nOut0_47[21] , 
        \nOut0_47[20] , \nOut0_47[19] , \nOut0_47[18] , \nOut0_47[17] , 
        \nOut0_47[16] , \nOut0_47[15] , \nOut0_47[14] , \nOut0_47[13] , 
        \nOut0_47[12] , \nOut0_47[11] , \nOut0_47[10] , \nOut0_47[9] , 
        \nOut0_47[8] , \nOut0_47[7] , \nOut0_47[6] , \nOut0_47[5] , 
        \nOut0_47[4] , \nOut0_47[3] , \nOut0_47[2] , \nOut0_47[1] , 
        \nOut0_47[0] }), .EAST_EDGE(\nOut1_46[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_45[31] ), .SE_EDGE(
        \nOut1_47[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_61 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut62[31] , \nScanOut62[30] , \nScanOut62[29] , 
        \nScanOut62[28] , \nScanOut62[27] , \nScanOut62[26] , \nScanOut62[25] , 
        \nScanOut62[24] , \nScanOut62[23] , \nScanOut62[22] , \nScanOut62[21] , 
        \nScanOut62[20] , \nScanOut62[19] , \nScanOut62[18] , \nScanOut62[17] , 
        \nScanOut62[16] , \nScanOut62[15] , \nScanOut62[14] , \nScanOut62[13] , 
        \nScanOut62[12] , \nScanOut62[11] , \nScanOut62[10] , \nScanOut62[9] , 
        \nScanOut62[8] , \nScanOut62[7] , \nScanOut62[6] , \nScanOut62[5] , 
        \nScanOut62[4] , \nScanOut62[3] , \nScanOut62[2] , \nScanOut62[1] , 
        \nScanOut62[0] }), .ScanOut({\nScanOut61[31] , \nScanOut61[30] , 
        \nScanOut61[29] , \nScanOut61[28] , \nScanOut61[27] , \nScanOut61[26] , 
        \nScanOut61[25] , \nScanOut61[24] , \nScanOut61[23] , \nScanOut61[22] , 
        \nScanOut61[21] , \nScanOut61[20] , \nScanOut61[19] , \nScanOut61[18] , 
        \nScanOut61[17] , \nScanOut61[16] , \nScanOut61[15] , \nScanOut61[14] , 
        \nScanOut61[13] , \nScanOut61[12] , \nScanOut61[11] , \nScanOut61[10] , 
        \nScanOut61[9] , \nScanOut61[8] , \nScanOut61[7] , \nScanOut61[6] , 
        \nScanOut61[5] , \nScanOut61[4] , \nScanOut61[3] , \nScanOut61[2] , 
        \nScanOut61[1] , \nScanOut61[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_61[31] , 
        \nOut0_61[30] , \nOut0_61[29] , \nOut0_61[28] , \nOut0_61[27] , 
        \nOut0_61[26] , \nOut0_61[25] , \nOut0_61[24] , \nOut0_61[23] , 
        \nOut0_61[22] , \nOut0_61[21] , \nOut0_61[20] , \nOut0_61[19] , 
        \nOut0_61[18] , \nOut0_61[17] , \nOut0_61[16] , \nOut0_61[15] , 
        \nOut0_61[14] , \nOut0_61[13] , \nOut0_61[12] , \nOut0_61[11] , 
        \nOut0_61[10] , \nOut0_61[9] , \nOut0_61[8] , \nOut0_61[7] , 
        \nOut0_61[6] , \nOut0_61[5] , \nOut0_61[4] , \nOut0_61[3] , 
        \nOut0_61[2] , \nOut0_61[1] , \nOut0_61[0] }), .NORTH_EDGE({
        \nOut0_60[31] , \nOut0_60[30] , \nOut0_60[29] , \nOut0_60[28] , 
        \nOut0_60[27] , \nOut0_60[26] , \nOut0_60[25] , \nOut0_60[24] , 
        \nOut0_60[23] , \nOut0_60[22] , \nOut0_60[21] , \nOut0_60[20] , 
        \nOut0_60[19] , \nOut0_60[18] , \nOut0_60[17] , \nOut0_60[16] , 
        \nOut0_60[15] , \nOut0_60[14] , \nOut0_60[13] , \nOut0_60[12] , 
        \nOut0_60[11] , \nOut0_60[10] , \nOut0_60[9] , \nOut0_60[8] , 
        \nOut0_60[7] , \nOut0_60[6] , \nOut0_60[5] , \nOut0_60[4] , 
        \nOut0_60[3] , \nOut0_60[2] , \nOut0_60[1] , \nOut0_60[0] }), 
        .SOUTH_EDGE({\nOut0_62[31] , \nOut0_62[30] , \nOut0_62[29] , 
        \nOut0_62[28] , \nOut0_62[27] , \nOut0_62[26] , \nOut0_62[25] , 
        \nOut0_62[24] , \nOut0_62[23] , \nOut0_62[22] , \nOut0_62[21] , 
        \nOut0_62[20] , \nOut0_62[19] , \nOut0_62[18] , \nOut0_62[17] , 
        \nOut0_62[16] , \nOut0_62[15] , \nOut0_62[14] , \nOut0_62[13] , 
        \nOut0_62[12] , \nOut0_62[11] , \nOut0_62[10] , \nOut0_62[9] , 
        \nOut0_62[8] , \nOut0_62[7] , \nOut0_62[6] , \nOut0_62[5] , 
        \nOut0_62[4] , \nOut0_62[3] , \nOut0_62[2] , \nOut0_62[1] , 
        \nOut0_62[0] }), .EAST_EDGE(\nOut1_61[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_60[31] ), .SE_EDGE(
        \nOut1_62[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_110 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut111[31] , \nScanOut111[30] , \nScanOut111[29] , 
        \nScanOut111[28] , \nScanOut111[27] , \nScanOut111[26] , 
        \nScanOut111[25] , \nScanOut111[24] , \nScanOut111[23] , 
        \nScanOut111[22] , \nScanOut111[21] , \nScanOut111[20] , 
        \nScanOut111[19] , \nScanOut111[18] , \nScanOut111[17] , 
        \nScanOut111[16] , \nScanOut111[15] , \nScanOut111[14] , 
        \nScanOut111[13] , \nScanOut111[12] , \nScanOut111[11] , 
        \nScanOut111[10] , \nScanOut111[9] , \nScanOut111[8] , 
        \nScanOut111[7] , \nScanOut111[6] , \nScanOut111[5] , \nScanOut111[4] , 
        \nScanOut111[3] , \nScanOut111[2] , \nScanOut111[1] , \nScanOut111[0] 
        }), .ScanOut({\nScanOut110[31] , \nScanOut110[30] , \nScanOut110[29] , 
        \nScanOut110[28] , \nScanOut110[27] , \nScanOut110[26] , 
        \nScanOut110[25] , \nScanOut110[24] , \nScanOut110[23] , 
        \nScanOut110[22] , \nScanOut110[21] , \nScanOut110[20] , 
        \nScanOut110[19] , \nScanOut110[18] , \nScanOut110[17] , 
        \nScanOut110[16] , \nScanOut110[15] , \nScanOut110[14] , 
        \nScanOut110[13] , \nScanOut110[12] , \nScanOut110[11] , 
        \nScanOut110[10] , \nScanOut110[9] , \nScanOut110[8] , 
        \nScanOut110[7] , \nScanOut110[6] , \nScanOut110[5] , \nScanOut110[4] , 
        \nScanOut110[3] , \nScanOut110[2] , \nScanOut110[1] , \nScanOut110[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_46[31] , \nOut1_46[30] , \nOut1_46[29] , 
        \nOut1_46[28] , \nOut1_46[27] , \nOut1_46[26] , \nOut1_46[25] , 
        \nOut1_46[24] , \nOut1_46[23] , \nOut1_46[22] , \nOut1_46[21] , 
        \nOut1_46[20] , \nOut1_46[19] , \nOut1_46[18] , \nOut1_46[17] , 
        \nOut1_46[16] , \nOut1_46[15] , \nOut1_46[14] , \nOut1_46[13] , 
        \nOut1_46[12] , \nOut1_46[11] , \nOut1_46[10] , \nOut1_46[9] , 
        \nOut1_46[8] , \nOut1_46[7] , \nOut1_46[6] , \nOut1_46[5] , 
        \nOut1_46[4] , \nOut1_46[3] , \nOut1_46[2] , \nOut1_46[1] , 
        \nOut1_46[0] }), .NORTH_EDGE({\nOut1_45[31] , \nOut1_45[30] , 
        \nOut1_45[29] , \nOut1_45[28] , \nOut1_45[27] , \nOut1_45[26] , 
        \nOut1_45[25] , \nOut1_45[24] , \nOut1_45[23] , \nOut1_45[22] , 
        \nOut1_45[21] , \nOut1_45[20] , \nOut1_45[19] , \nOut1_45[18] , 
        \nOut1_45[17] , \nOut1_45[16] , \nOut1_45[15] , \nOut1_45[14] , 
        \nOut1_45[13] , \nOut1_45[12] , \nOut1_45[11] , \nOut1_45[10] , 
        \nOut1_45[9] , \nOut1_45[8] , \nOut1_45[7] , \nOut1_45[6] , 
        \nOut1_45[5] , \nOut1_45[4] , \nOut1_45[3] , \nOut1_45[2] , 
        \nOut1_45[1] , \nOut1_45[0] }), .SOUTH_EDGE({\nOut1_47[31] , 
        \nOut1_47[30] , \nOut1_47[29] , \nOut1_47[28] , \nOut1_47[27] , 
        \nOut1_47[26] , \nOut1_47[25] , \nOut1_47[24] , \nOut1_47[23] , 
        \nOut1_47[22] , \nOut1_47[21] , \nOut1_47[20] , \nOut1_47[19] , 
        \nOut1_47[18] , \nOut1_47[17] , \nOut1_47[16] , \nOut1_47[15] , 
        \nOut1_47[14] , \nOut1_47[13] , \nOut1_47[12] , \nOut1_47[11] , 
        \nOut1_47[10] , \nOut1_47[9] , \nOut1_47[8] , \nOut1_47[7] , 
        \nOut1_47[6] , \nOut1_47[5] , \nOut1_47[4] , \nOut1_47[3] , 
        \nOut1_47[2] , \nOut1_47[1] , \nOut1_47[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_46[0] ), .NW_EDGE(\nOut0_45[0] ), .SW_EDGE(
        \nOut0_47[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_41 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut42[31] , \nScanOut42[30] , \nScanOut42[29] , 
        \nScanOut42[28] , \nScanOut42[27] , \nScanOut42[26] , \nScanOut42[25] , 
        \nScanOut42[24] , \nScanOut42[23] , \nScanOut42[22] , \nScanOut42[21] , 
        \nScanOut42[20] , \nScanOut42[19] , \nScanOut42[18] , \nScanOut42[17] , 
        \nScanOut42[16] , \nScanOut42[15] , \nScanOut42[14] , \nScanOut42[13] , 
        \nScanOut42[12] , \nScanOut42[11] , \nScanOut42[10] , \nScanOut42[9] , 
        \nScanOut42[8] , \nScanOut42[7] , \nScanOut42[6] , \nScanOut42[5] , 
        \nScanOut42[4] , \nScanOut42[3] , \nScanOut42[2] , \nScanOut42[1] , 
        \nScanOut42[0] }), .ScanOut({\nScanOut41[31] , \nScanOut41[30] , 
        \nScanOut41[29] , \nScanOut41[28] , \nScanOut41[27] , \nScanOut41[26] , 
        \nScanOut41[25] , \nScanOut41[24] , \nScanOut41[23] , \nScanOut41[22] , 
        \nScanOut41[21] , \nScanOut41[20] , \nScanOut41[19] , \nScanOut41[18] , 
        \nScanOut41[17] , \nScanOut41[16] , \nScanOut41[15] , \nScanOut41[14] , 
        \nScanOut41[13] , \nScanOut41[12] , \nScanOut41[11] , \nScanOut41[10] , 
        \nScanOut41[9] , \nScanOut41[8] , \nScanOut41[7] , \nScanOut41[6] , 
        \nScanOut41[5] , \nScanOut41[4] , \nScanOut41[3] , \nScanOut41[2] , 
        \nScanOut41[1] , \nScanOut41[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_41[31] , 
        \nOut0_41[30] , \nOut0_41[29] , \nOut0_41[28] , \nOut0_41[27] , 
        \nOut0_41[26] , \nOut0_41[25] , \nOut0_41[24] , \nOut0_41[23] , 
        \nOut0_41[22] , \nOut0_41[21] , \nOut0_41[20] , \nOut0_41[19] , 
        \nOut0_41[18] , \nOut0_41[17] , \nOut0_41[16] , \nOut0_41[15] , 
        \nOut0_41[14] , \nOut0_41[13] , \nOut0_41[12] , \nOut0_41[11] , 
        \nOut0_41[10] , \nOut0_41[9] , \nOut0_41[8] , \nOut0_41[7] , 
        \nOut0_41[6] , \nOut0_41[5] , \nOut0_41[4] , \nOut0_41[3] , 
        \nOut0_41[2] , \nOut0_41[1] , \nOut0_41[0] }), .NORTH_EDGE({
        \nOut0_40[31] , \nOut0_40[30] , \nOut0_40[29] , \nOut0_40[28] , 
        \nOut0_40[27] , \nOut0_40[26] , \nOut0_40[25] , \nOut0_40[24] , 
        \nOut0_40[23] , \nOut0_40[22] , \nOut0_40[21] , \nOut0_40[20] , 
        \nOut0_40[19] , \nOut0_40[18] , \nOut0_40[17] , \nOut0_40[16] , 
        \nOut0_40[15] , \nOut0_40[14] , \nOut0_40[13] , \nOut0_40[12] , 
        \nOut0_40[11] , \nOut0_40[10] , \nOut0_40[9] , \nOut0_40[8] , 
        \nOut0_40[7] , \nOut0_40[6] , \nOut0_40[5] , \nOut0_40[4] , 
        \nOut0_40[3] , \nOut0_40[2] , \nOut0_40[1] , \nOut0_40[0] }), 
        .SOUTH_EDGE({\nOut0_42[31] , \nOut0_42[30] , \nOut0_42[29] , 
        \nOut0_42[28] , \nOut0_42[27] , \nOut0_42[26] , \nOut0_42[25] , 
        \nOut0_42[24] , \nOut0_42[23] , \nOut0_42[22] , \nOut0_42[21] , 
        \nOut0_42[20] , \nOut0_42[19] , \nOut0_42[18] , \nOut0_42[17] , 
        \nOut0_42[16] , \nOut0_42[15] , \nOut0_42[14] , \nOut0_42[13] , 
        \nOut0_42[12] , \nOut0_42[11] , \nOut0_42[10] , \nOut0_42[9] , 
        \nOut0_42[8] , \nOut0_42[7] , \nOut0_42[6] , \nOut0_42[5] , 
        \nOut0_42[4] , \nOut0_42[3] , \nOut0_42[2] , \nOut0_42[1] , 
        \nOut0_42[0] }), .EAST_EDGE(\nOut1_41[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_40[31] ), .SE_EDGE(
        \nOut1_42[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_66 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut67[31] , \nScanOut67[30] , \nScanOut67[29] , 
        \nScanOut67[28] , \nScanOut67[27] , \nScanOut67[26] , \nScanOut67[25] , 
        \nScanOut67[24] , \nScanOut67[23] , \nScanOut67[22] , \nScanOut67[21] , 
        \nScanOut67[20] , \nScanOut67[19] , \nScanOut67[18] , \nScanOut67[17] , 
        \nScanOut67[16] , \nScanOut67[15] , \nScanOut67[14] , \nScanOut67[13] , 
        \nScanOut67[12] , \nScanOut67[11] , \nScanOut67[10] , \nScanOut67[9] , 
        \nScanOut67[8] , \nScanOut67[7] , \nScanOut67[6] , \nScanOut67[5] , 
        \nScanOut67[4] , \nScanOut67[3] , \nScanOut67[2] , \nScanOut67[1] , 
        \nScanOut67[0] }), .ScanOut({\nScanOut66[31] , \nScanOut66[30] , 
        \nScanOut66[29] , \nScanOut66[28] , \nScanOut66[27] , \nScanOut66[26] , 
        \nScanOut66[25] , \nScanOut66[24] , \nScanOut66[23] , \nScanOut66[22] , 
        \nScanOut66[21] , \nScanOut66[20] , \nScanOut66[19] , \nScanOut66[18] , 
        \nScanOut66[17] , \nScanOut66[16] , \nScanOut66[15] , \nScanOut66[14] , 
        \nScanOut66[13] , \nScanOut66[12] , \nScanOut66[11] , \nScanOut66[10] , 
        \nScanOut66[9] , \nScanOut66[8] , \nScanOut66[7] , \nScanOut66[6] , 
        \nScanOut66[5] , \nScanOut66[4] , \nScanOut66[3] , \nScanOut66[2] , 
        \nScanOut66[1] , \nScanOut66[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_2[31] , 
        \nOut1_2[30] , \nOut1_2[29] , \nOut1_2[28] , \nOut1_2[27] , 
        \nOut1_2[26] , \nOut1_2[25] , \nOut1_2[24] , \nOut1_2[23] , 
        \nOut1_2[22] , \nOut1_2[21] , \nOut1_2[20] , \nOut1_2[19] , 
        \nOut1_2[18] , \nOut1_2[17] , \nOut1_2[16] , \nOut1_2[15] , 
        \nOut1_2[14] , \nOut1_2[13] , \nOut1_2[12] , \nOut1_2[11] , 
        \nOut1_2[10] , \nOut1_2[9] , \nOut1_2[8] , \nOut1_2[7] , \nOut1_2[6] , 
        \nOut1_2[5] , \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , 
        \nOut1_2[0] }), .NORTH_EDGE({\nOut1_1[31] , \nOut1_1[30] , 
        \nOut1_1[29] , \nOut1_1[28] , \nOut1_1[27] , \nOut1_1[26] , 
        \nOut1_1[25] , \nOut1_1[24] , \nOut1_1[23] , \nOut1_1[22] , 
        \nOut1_1[21] , \nOut1_1[20] , \nOut1_1[19] , \nOut1_1[18] , 
        \nOut1_1[17] , \nOut1_1[16] , \nOut1_1[15] , \nOut1_1[14] , 
        \nOut1_1[13] , \nOut1_1[12] , \nOut1_1[11] , \nOut1_1[10] , 
        \nOut1_1[9] , \nOut1_1[8] , \nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , 
        \nOut1_1[4] , \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), 
        .SOUTH_EDGE({\nOut1_3[31] , \nOut1_3[30] , \nOut1_3[29] , 
        \nOut1_3[28] , \nOut1_3[27] , \nOut1_3[26] , \nOut1_3[25] , 
        \nOut1_3[24] , \nOut1_3[23] , \nOut1_3[22] , \nOut1_3[21] , 
        \nOut1_3[20] , \nOut1_3[19] , \nOut1_3[18] , \nOut1_3[17] , 
        \nOut1_3[16] , \nOut1_3[15] , \nOut1_3[14] , \nOut1_3[13] , 
        \nOut1_3[12] , \nOut1_3[11] , \nOut1_3[10] , \nOut1_3[9] , 
        \nOut1_3[8] , \nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , 
        \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_2[0] ), .NW_EDGE(\nOut0_1[0] ), .SW_EDGE(
        \nOut0_3[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_83 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut84[31] , \nScanOut84[30] , \nScanOut84[29] , 
        \nScanOut84[28] , \nScanOut84[27] , \nScanOut84[26] , \nScanOut84[25] , 
        \nScanOut84[24] , \nScanOut84[23] , \nScanOut84[22] , \nScanOut84[21] , 
        \nScanOut84[20] , \nScanOut84[19] , \nScanOut84[18] , \nScanOut84[17] , 
        \nScanOut84[16] , \nScanOut84[15] , \nScanOut84[14] , \nScanOut84[13] , 
        \nScanOut84[12] , \nScanOut84[11] , \nScanOut84[10] , \nScanOut84[9] , 
        \nScanOut84[8] , \nScanOut84[7] , \nScanOut84[6] , \nScanOut84[5] , 
        \nScanOut84[4] , \nScanOut84[3] , \nScanOut84[2] , \nScanOut84[1] , 
        \nScanOut84[0] }), .ScanOut({\nScanOut83[31] , \nScanOut83[30] , 
        \nScanOut83[29] , \nScanOut83[28] , \nScanOut83[27] , \nScanOut83[26] , 
        \nScanOut83[25] , \nScanOut83[24] , \nScanOut83[23] , \nScanOut83[22] , 
        \nScanOut83[21] , \nScanOut83[20] , \nScanOut83[19] , \nScanOut83[18] , 
        \nScanOut83[17] , \nScanOut83[16] , \nScanOut83[15] , \nScanOut83[14] , 
        \nScanOut83[13] , \nScanOut83[12] , \nScanOut83[11] , \nScanOut83[10] , 
        \nScanOut83[9] , \nScanOut83[8] , \nScanOut83[7] , \nScanOut83[6] , 
        \nScanOut83[5] , \nScanOut83[4] , \nScanOut83[3] , \nScanOut83[2] , 
        \nScanOut83[1] , \nScanOut83[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_19[31] , 
        \nOut1_19[30] , \nOut1_19[29] , \nOut1_19[28] , \nOut1_19[27] , 
        \nOut1_19[26] , \nOut1_19[25] , \nOut1_19[24] , \nOut1_19[23] , 
        \nOut1_19[22] , \nOut1_19[21] , \nOut1_19[20] , \nOut1_19[19] , 
        \nOut1_19[18] , \nOut1_19[17] , \nOut1_19[16] , \nOut1_19[15] , 
        \nOut1_19[14] , \nOut1_19[13] , \nOut1_19[12] , \nOut1_19[11] , 
        \nOut1_19[10] , \nOut1_19[9] , \nOut1_19[8] , \nOut1_19[7] , 
        \nOut1_19[6] , \nOut1_19[5] , \nOut1_19[4] , \nOut1_19[3] , 
        \nOut1_19[2] , \nOut1_19[1] , \nOut1_19[0] }), .NORTH_EDGE({
        \nOut1_18[31] , \nOut1_18[30] , \nOut1_18[29] , \nOut1_18[28] , 
        \nOut1_18[27] , \nOut1_18[26] , \nOut1_18[25] , \nOut1_18[24] , 
        \nOut1_18[23] , \nOut1_18[22] , \nOut1_18[21] , \nOut1_18[20] , 
        \nOut1_18[19] , \nOut1_18[18] , \nOut1_18[17] , \nOut1_18[16] , 
        \nOut1_18[15] , \nOut1_18[14] , \nOut1_18[13] , \nOut1_18[12] , 
        \nOut1_18[11] , \nOut1_18[10] , \nOut1_18[9] , \nOut1_18[8] , 
        \nOut1_18[7] , \nOut1_18[6] , \nOut1_18[5] , \nOut1_18[4] , 
        \nOut1_18[3] , \nOut1_18[2] , \nOut1_18[1] , \nOut1_18[0] }), 
        .SOUTH_EDGE({\nOut1_20[31] , \nOut1_20[30] , \nOut1_20[29] , 
        \nOut1_20[28] , \nOut1_20[27] , \nOut1_20[26] , \nOut1_20[25] , 
        \nOut1_20[24] , \nOut1_20[23] , \nOut1_20[22] , \nOut1_20[21] , 
        \nOut1_20[20] , \nOut1_20[19] , \nOut1_20[18] , \nOut1_20[17] , 
        \nOut1_20[16] , \nOut1_20[15] , \nOut1_20[14] , \nOut1_20[13] , 
        \nOut1_20[12] , \nOut1_20[11] , \nOut1_20[10] , \nOut1_20[9] , 
        \nOut1_20[8] , \nOut1_20[7] , \nOut1_20[6] , \nOut1_20[5] , 
        \nOut1_20[4] , \nOut1_20[3] , \nOut1_20[2] , \nOut1_20[1] , 
        \nOut1_20[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_19[0] ), 
        .NW_EDGE(\nOut0_18[0] ), .SW_EDGE(\nOut0_20[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_84 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut85[31] , \nScanOut85[30] , \nScanOut85[29] , 
        \nScanOut85[28] , \nScanOut85[27] , \nScanOut85[26] , \nScanOut85[25] , 
        \nScanOut85[24] , \nScanOut85[23] , \nScanOut85[22] , \nScanOut85[21] , 
        \nScanOut85[20] , \nScanOut85[19] , \nScanOut85[18] , \nScanOut85[17] , 
        \nScanOut85[16] , \nScanOut85[15] , \nScanOut85[14] , \nScanOut85[13] , 
        \nScanOut85[12] , \nScanOut85[11] , \nScanOut85[10] , \nScanOut85[9] , 
        \nScanOut85[8] , \nScanOut85[7] , \nScanOut85[6] , \nScanOut85[5] , 
        \nScanOut85[4] , \nScanOut85[3] , \nScanOut85[2] , \nScanOut85[1] , 
        \nScanOut85[0] }), .ScanOut({\nScanOut84[31] , \nScanOut84[30] , 
        \nScanOut84[29] , \nScanOut84[28] , \nScanOut84[27] , \nScanOut84[26] , 
        \nScanOut84[25] , \nScanOut84[24] , \nScanOut84[23] , \nScanOut84[22] , 
        \nScanOut84[21] , \nScanOut84[20] , \nScanOut84[19] , \nScanOut84[18] , 
        \nScanOut84[17] , \nScanOut84[16] , \nScanOut84[15] , \nScanOut84[14] , 
        \nScanOut84[13] , \nScanOut84[12] , \nScanOut84[11] , \nScanOut84[10] , 
        \nScanOut84[9] , \nScanOut84[8] , \nScanOut84[7] , \nScanOut84[6] , 
        \nScanOut84[5] , \nScanOut84[4] , \nScanOut84[3] , \nScanOut84[2] , 
        \nScanOut84[1] , \nScanOut84[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_20[31] , 
        \nOut1_20[30] , \nOut1_20[29] , \nOut1_20[28] , \nOut1_20[27] , 
        \nOut1_20[26] , \nOut1_20[25] , \nOut1_20[24] , \nOut1_20[23] , 
        \nOut1_20[22] , \nOut1_20[21] , \nOut1_20[20] , \nOut1_20[19] , 
        \nOut1_20[18] , \nOut1_20[17] , \nOut1_20[16] , \nOut1_20[15] , 
        \nOut1_20[14] , \nOut1_20[13] , \nOut1_20[12] , \nOut1_20[11] , 
        \nOut1_20[10] , \nOut1_20[9] , \nOut1_20[8] , \nOut1_20[7] , 
        \nOut1_20[6] , \nOut1_20[5] , \nOut1_20[4] , \nOut1_20[3] , 
        \nOut1_20[2] , \nOut1_20[1] , \nOut1_20[0] }), .NORTH_EDGE({
        \nOut1_19[31] , \nOut1_19[30] , \nOut1_19[29] , \nOut1_19[28] , 
        \nOut1_19[27] , \nOut1_19[26] , \nOut1_19[25] , \nOut1_19[24] , 
        \nOut1_19[23] , \nOut1_19[22] , \nOut1_19[21] , \nOut1_19[20] , 
        \nOut1_19[19] , \nOut1_19[18] , \nOut1_19[17] , \nOut1_19[16] , 
        \nOut1_19[15] , \nOut1_19[14] , \nOut1_19[13] , \nOut1_19[12] , 
        \nOut1_19[11] , \nOut1_19[10] , \nOut1_19[9] , \nOut1_19[8] , 
        \nOut1_19[7] , \nOut1_19[6] , \nOut1_19[5] , \nOut1_19[4] , 
        \nOut1_19[3] , \nOut1_19[2] , \nOut1_19[1] , \nOut1_19[0] }), 
        .SOUTH_EDGE({\nOut1_21[31] , \nOut1_21[30] , \nOut1_21[29] , 
        \nOut1_21[28] , \nOut1_21[27] , \nOut1_21[26] , \nOut1_21[25] , 
        \nOut1_21[24] , \nOut1_21[23] , \nOut1_21[22] , \nOut1_21[21] , 
        \nOut1_21[20] , \nOut1_21[19] , \nOut1_21[18] , \nOut1_21[17] , 
        \nOut1_21[16] , \nOut1_21[15] , \nOut1_21[14] , \nOut1_21[13] , 
        \nOut1_21[12] , \nOut1_21[11] , \nOut1_21[10] , \nOut1_21[9] , 
        \nOut1_21[8] , \nOut1_21[7] , \nOut1_21[6] , \nOut1_21[5] , 
        \nOut1_21[4] , \nOut1_21[3] , \nOut1_21[2] , \nOut1_21[1] , 
        \nOut1_21[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_20[0] ), 
        .NW_EDGE(\nOut0_19[0] ), .SW_EDGE(\nOut0_21[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_117 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut118[31] , \nScanOut118[30] , \nScanOut118[29] , 
        \nScanOut118[28] , \nScanOut118[27] , \nScanOut118[26] , 
        \nScanOut118[25] , \nScanOut118[24] , \nScanOut118[23] , 
        \nScanOut118[22] , \nScanOut118[21] , \nScanOut118[20] , 
        \nScanOut118[19] , \nScanOut118[18] , \nScanOut118[17] , 
        \nScanOut118[16] , \nScanOut118[15] , \nScanOut118[14] , 
        \nScanOut118[13] , \nScanOut118[12] , \nScanOut118[11] , 
        \nScanOut118[10] , \nScanOut118[9] , \nScanOut118[8] , 
        \nScanOut118[7] , \nScanOut118[6] , \nScanOut118[5] , \nScanOut118[4] , 
        \nScanOut118[3] , \nScanOut118[2] , \nScanOut118[1] , \nScanOut118[0] 
        }), .ScanOut({\nScanOut117[31] , \nScanOut117[30] , \nScanOut117[29] , 
        \nScanOut117[28] , \nScanOut117[27] , \nScanOut117[26] , 
        \nScanOut117[25] , \nScanOut117[24] , \nScanOut117[23] , 
        \nScanOut117[22] , \nScanOut117[21] , \nScanOut117[20] , 
        \nScanOut117[19] , \nScanOut117[18] , \nScanOut117[17] , 
        \nScanOut117[16] , \nScanOut117[15] , \nScanOut117[14] , 
        \nScanOut117[13] , \nScanOut117[12] , \nScanOut117[11] , 
        \nScanOut117[10] , \nScanOut117[9] , \nScanOut117[8] , 
        \nScanOut117[7] , \nScanOut117[6] , \nScanOut117[5] , \nScanOut117[4] , 
        \nScanOut117[3] , \nScanOut117[2] , \nScanOut117[1] , \nScanOut117[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_53[31] , \nOut1_53[30] , \nOut1_53[29] , 
        \nOut1_53[28] , \nOut1_53[27] , \nOut1_53[26] , \nOut1_53[25] , 
        \nOut1_53[24] , \nOut1_53[23] , \nOut1_53[22] , \nOut1_53[21] , 
        \nOut1_53[20] , \nOut1_53[19] , \nOut1_53[18] , \nOut1_53[17] , 
        \nOut1_53[16] , \nOut1_53[15] , \nOut1_53[14] , \nOut1_53[13] , 
        \nOut1_53[12] , \nOut1_53[11] , \nOut1_53[10] , \nOut1_53[9] , 
        \nOut1_53[8] , \nOut1_53[7] , \nOut1_53[6] , \nOut1_53[5] , 
        \nOut1_53[4] , \nOut1_53[3] , \nOut1_53[2] , \nOut1_53[1] , 
        \nOut1_53[0] }), .NORTH_EDGE({\nOut1_52[31] , \nOut1_52[30] , 
        \nOut1_52[29] , \nOut1_52[28] , \nOut1_52[27] , \nOut1_52[26] , 
        \nOut1_52[25] , \nOut1_52[24] , \nOut1_52[23] , \nOut1_52[22] , 
        \nOut1_52[21] , \nOut1_52[20] , \nOut1_52[19] , \nOut1_52[18] , 
        \nOut1_52[17] , \nOut1_52[16] , \nOut1_52[15] , \nOut1_52[14] , 
        \nOut1_52[13] , \nOut1_52[12] , \nOut1_52[11] , \nOut1_52[10] , 
        \nOut1_52[9] , \nOut1_52[8] , \nOut1_52[7] , \nOut1_52[6] , 
        \nOut1_52[5] , \nOut1_52[4] , \nOut1_52[3] , \nOut1_52[2] , 
        \nOut1_52[1] , \nOut1_52[0] }), .SOUTH_EDGE({\nOut1_54[31] , 
        \nOut1_54[30] , \nOut1_54[29] , \nOut1_54[28] , \nOut1_54[27] , 
        \nOut1_54[26] , \nOut1_54[25] , \nOut1_54[24] , \nOut1_54[23] , 
        \nOut1_54[22] , \nOut1_54[21] , \nOut1_54[20] , \nOut1_54[19] , 
        \nOut1_54[18] , \nOut1_54[17] , \nOut1_54[16] , \nOut1_54[15] , 
        \nOut1_54[14] , \nOut1_54[13] , \nOut1_54[12] , \nOut1_54[11] , 
        \nOut1_54[10] , \nOut1_54[9] , \nOut1_54[8] , \nOut1_54[7] , 
        \nOut1_54[6] , \nOut1_54[5] , \nOut1_54[4] , \nOut1_54[3] , 
        \nOut1_54[2] , \nOut1_54[1] , \nOut1_54[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_53[0] ), .NW_EDGE(\nOut0_52[0] ), .SW_EDGE(
        \nOut0_54[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_98 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut99[31] , \nScanOut99[30] , \nScanOut99[29] , 
        \nScanOut99[28] , \nScanOut99[27] , \nScanOut99[26] , \nScanOut99[25] , 
        \nScanOut99[24] , \nScanOut99[23] , \nScanOut99[22] , \nScanOut99[21] , 
        \nScanOut99[20] , \nScanOut99[19] , \nScanOut99[18] , \nScanOut99[17] , 
        \nScanOut99[16] , \nScanOut99[15] , \nScanOut99[14] , \nScanOut99[13] , 
        \nScanOut99[12] , \nScanOut99[11] , \nScanOut99[10] , \nScanOut99[9] , 
        \nScanOut99[8] , \nScanOut99[7] , \nScanOut99[6] , \nScanOut99[5] , 
        \nScanOut99[4] , \nScanOut99[3] , \nScanOut99[2] , \nScanOut99[1] , 
        \nScanOut99[0] }), .ScanOut({\nScanOut98[31] , \nScanOut98[30] , 
        \nScanOut98[29] , \nScanOut98[28] , \nScanOut98[27] , \nScanOut98[26] , 
        \nScanOut98[25] , \nScanOut98[24] , \nScanOut98[23] , \nScanOut98[22] , 
        \nScanOut98[21] , \nScanOut98[20] , \nScanOut98[19] , \nScanOut98[18] , 
        \nScanOut98[17] , \nScanOut98[16] , \nScanOut98[15] , \nScanOut98[14] , 
        \nScanOut98[13] , \nScanOut98[12] , \nScanOut98[11] , \nScanOut98[10] , 
        \nScanOut98[9] , \nScanOut98[8] , \nScanOut98[7] , \nScanOut98[6] , 
        \nScanOut98[5] , \nScanOut98[4] , \nScanOut98[3] , \nScanOut98[2] , 
        \nScanOut98[1] , \nScanOut98[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_34[31] , 
        \nOut1_34[30] , \nOut1_34[29] , \nOut1_34[28] , \nOut1_34[27] , 
        \nOut1_34[26] , \nOut1_34[25] , \nOut1_34[24] , \nOut1_34[23] , 
        \nOut1_34[22] , \nOut1_34[21] , \nOut1_34[20] , \nOut1_34[19] , 
        \nOut1_34[18] , \nOut1_34[17] , \nOut1_34[16] , \nOut1_34[15] , 
        \nOut1_34[14] , \nOut1_34[13] , \nOut1_34[12] , \nOut1_34[11] , 
        \nOut1_34[10] , \nOut1_34[9] , \nOut1_34[8] , \nOut1_34[7] , 
        \nOut1_34[6] , \nOut1_34[5] , \nOut1_34[4] , \nOut1_34[3] , 
        \nOut1_34[2] , \nOut1_34[1] , \nOut1_34[0] }), .NORTH_EDGE({
        \nOut1_33[31] , \nOut1_33[30] , \nOut1_33[29] , \nOut1_33[28] , 
        \nOut1_33[27] , \nOut1_33[26] , \nOut1_33[25] , \nOut1_33[24] , 
        \nOut1_33[23] , \nOut1_33[22] , \nOut1_33[21] , \nOut1_33[20] , 
        \nOut1_33[19] , \nOut1_33[18] , \nOut1_33[17] , \nOut1_33[16] , 
        \nOut1_33[15] , \nOut1_33[14] , \nOut1_33[13] , \nOut1_33[12] , 
        \nOut1_33[11] , \nOut1_33[10] , \nOut1_33[9] , \nOut1_33[8] , 
        \nOut1_33[7] , \nOut1_33[6] , \nOut1_33[5] , \nOut1_33[4] , 
        \nOut1_33[3] , \nOut1_33[2] , \nOut1_33[1] , \nOut1_33[0] }), 
        .SOUTH_EDGE({\nOut1_35[31] , \nOut1_35[30] , \nOut1_35[29] , 
        \nOut1_35[28] , \nOut1_35[27] , \nOut1_35[26] , \nOut1_35[25] , 
        \nOut1_35[24] , \nOut1_35[23] , \nOut1_35[22] , \nOut1_35[21] , 
        \nOut1_35[20] , \nOut1_35[19] , \nOut1_35[18] , \nOut1_35[17] , 
        \nOut1_35[16] , \nOut1_35[15] , \nOut1_35[14] , \nOut1_35[13] , 
        \nOut1_35[12] , \nOut1_35[11] , \nOut1_35[10] , \nOut1_35[9] , 
        \nOut1_35[8] , \nOut1_35[7] , \nOut1_35[6] , \nOut1_35[5] , 
        \nOut1_35[4] , \nOut1_35[3] , \nOut1_35[2] , \nOut1_35[1] , 
        \nOut1_35[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_34[0] ), 
        .NW_EDGE(\nOut0_33[0] ), .SW_EDGE(\nOut0_35[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_26 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut27[31] , \nScanOut27[30] , \nScanOut27[29] , 
        \nScanOut27[28] , \nScanOut27[27] , \nScanOut27[26] , \nScanOut27[25] , 
        \nScanOut27[24] , \nScanOut27[23] , \nScanOut27[22] , \nScanOut27[21] , 
        \nScanOut27[20] , \nScanOut27[19] , \nScanOut27[18] , \nScanOut27[17] , 
        \nScanOut27[16] , \nScanOut27[15] , \nScanOut27[14] , \nScanOut27[13] , 
        \nScanOut27[12] , \nScanOut27[11] , \nScanOut27[10] , \nScanOut27[9] , 
        \nScanOut27[8] , \nScanOut27[7] , \nScanOut27[6] , \nScanOut27[5] , 
        \nScanOut27[4] , \nScanOut27[3] , \nScanOut27[2] , \nScanOut27[1] , 
        \nScanOut27[0] }), .ScanOut({\nScanOut26[31] , \nScanOut26[30] , 
        \nScanOut26[29] , \nScanOut26[28] , \nScanOut26[27] , \nScanOut26[26] , 
        \nScanOut26[25] , \nScanOut26[24] , \nScanOut26[23] , \nScanOut26[22] , 
        \nScanOut26[21] , \nScanOut26[20] , \nScanOut26[19] , \nScanOut26[18] , 
        \nScanOut26[17] , \nScanOut26[16] , \nScanOut26[15] , \nScanOut26[14] , 
        \nScanOut26[13] , \nScanOut26[12] , \nScanOut26[11] , \nScanOut26[10] , 
        \nScanOut26[9] , \nScanOut26[8] , \nScanOut26[7] , \nScanOut26[6] , 
        \nScanOut26[5] , \nScanOut26[4] , \nScanOut26[3] , \nScanOut26[2] , 
        \nScanOut26[1] , \nScanOut26[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_26[31] , 
        \nOut0_26[30] , \nOut0_26[29] , \nOut0_26[28] , \nOut0_26[27] , 
        \nOut0_26[26] , \nOut0_26[25] , \nOut0_26[24] , \nOut0_26[23] , 
        \nOut0_26[22] , \nOut0_26[21] , \nOut0_26[20] , \nOut0_26[19] , 
        \nOut0_26[18] , \nOut0_26[17] , \nOut0_26[16] , \nOut0_26[15] , 
        \nOut0_26[14] , \nOut0_26[13] , \nOut0_26[12] , \nOut0_26[11] , 
        \nOut0_26[10] , \nOut0_26[9] , \nOut0_26[8] , \nOut0_26[7] , 
        \nOut0_26[6] , \nOut0_26[5] , \nOut0_26[4] , \nOut0_26[3] , 
        \nOut0_26[2] , \nOut0_26[1] , \nOut0_26[0] }), .NORTH_EDGE({
        \nOut0_25[31] , \nOut0_25[30] , \nOut0_25[29] , \nOut0_25[28] , 
        \nOut0_25[27] , \nOut0_25[26] , \nOut0_25[25] , \nOut0_25[24] , 
        \nOut0_25[23] , \nOut0_25[22] , \nOut0_25[21] , \nOut0_25[20] , 
        \nOut0_25[19] , \nOut0_25[18] , \nOut0_25[17] , \nOut0_25[16] , 
        \nOut0_25[15] , \nOut0_25[14] , \nOut0_25[13] , \nOut0_25[12] , 
        \nOut0_25[11] , \nOut0_25[10] , \nOut0_25[9] , \nOut0_25[8] , 
        \nOut0_25[7] , \nOut0_25[6] , \nOut0_25[5] , \nOut0_25[4] , 
        \nOut0_25[3] , \nOut0_25[2] , \nOut0_25[1] , \nOut0_25[0] }), 
        .SOUTH_EDGE({\nOut0_27[31] , \nOut0_27[30] , \nOut0_27[29] , 
        \nOut0_27[28] , \nOut0_27[27] , \nOut0_27[26] , \nOut0_27[25] , 
        \nOut0_27[24] , \nOut0_27[23] , \nOut0_27[22] , \nOut0_27[21] , 
        \nOut0_27[20] , \nOut0_27[19] , \nOut0_27[18] , \nOut0_27[17] , 
        \nOut0_27[16] , \nOut0_27[15] , \nOut0_27[14] , \nOut0_27[13] , 
        \nOut0_27[12] , \nOut0_27[11] , \nOut0_27[10] , \nOut0_27[9] , 
        \nOut0_27[8] , \nOut0_27[7] , \nOut0_27[6] , \nOut0_27[5] , 
        \nOut0_27[4] , \nOut0_27[3] , \nOut0_27[2] , \nOut0_27[1] , 
        \nOut0_27[0] }), .EAST_EDGE(\nOut1_26[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_25[31] ), .SE_EDGE(
        \nOut1_27[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_34 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut35[31] , \nScanOut35[30] , \nScanOut35[29] , 
        \nScanOut35[28] , \nScanOut35[27] , \nScanOut35[26] , \nScanOut35[25] , 
        \nScanOut35[24] , \nScanOut35[23] , \nScanOut35[22] , \nScanOut35[21] , 
        \nScanOut35[20] , \nScanOut35[19] , \nScanOut35[18] , \nScanOut35[17] , 
        \nScanOut35[16] , \nScanOut35[15] , \nScanOut35[14] , \nScanOut35[13] , 
        \nScanOut35[12] , \nScanOut35[11] , \nScanOut35[10] , \nScanOut35[9] , 
        \nScanOut35[8] , \nScanOut35[7] , \nScanOut35[6] , \nScanOut35[5] , 
        \nScanOut35[4] , \nScanOut35[3] , \nScanOut35[2] , \nScanOut35[1] , 
        \nScanOut35[0] }), .ScanOut({\nScanOut34[31] , \nScanOut34[30] , 
        \nScanOut34[29] , \nScanOut34[28] , \nScanOut34[27] , \nScanOut34[26] , 
        \nScanOut34[25] , \nScanOut34[24] , \nScanOut34[23] , \nScanOut34[22] , 
        \nScanOut34[21] , \nScanOut34[20] , \nScanOut34[19] , \nScanOut34[18] , 
        \nScanOut34[17] , \nScanOut34[16] , \nScanOut34[15] , \nScanOut34[14] , 
        \nScanOut34[13] , \nScanOut34[12] , \nScanOut34[11] , \nScanOut34[10] , 
        \nScanOut34[9] , \nScanOut34[8] , \nScanOut34[7] , \nScanOut34[6] , 
        \nScanOut34[5] , \nScanOut34[4] , \nScanOut34[3] , \nScanOut34[2] , 
        \nScanOut34[1] , \nScanOut34[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_34[31] , 
        \nOut0_34[30] , \nOut0_34[29] , \nOut0_34[28] , \nOut0_34[27] , 
        \nOut0_34[26] , \nOut0_34[25] , \nOut0_34[24] , \nOut0_34[23] , 
        \nOut0_34[22] , \nOut0_34[21] , \nOut0_34[20] , \nOut0_34[19] , 
        \nOut0_34[18] , \nOut0_34[17] , \nOut0_34[16] , \nOut0_34[15] , 
        \nOut0_34[14] , \nOut0_34[13] , \nOut0_34[12] , \nOut0_34[11] , 
        \nOut0_34[10] , \nOut0_34[9] , \nOut0_34[8] , \nOut0_34[7] , 
        \nOut0_34[6] , \nOut0_34[5] , \nOut0_34[4] , \nOut0_34[3] , 
        \nOut0_34[2] , \nOut0_34[1] , \nOut0_34[0] }), .NORTH_EDGE({
        \nOut0_33[31] , \nOut0_33[30] , \nOut0_33[29] , \nOut0_33[28] , 
        \nOut0_33[27] , \nOut0_33[26] , \nOut0_33[25] , \nOut0_33[24] , 
        \nOut0_33[23] , \nOut0_33[22] , \nOut0_33[21] , \nOut0_33[20] , 
        \nOut0_33[19] , \nOut0_33[18] , \nOut0_33[17] , \nOut0_33[16] , 
        \nOut0_33[15] , \nOut0_33[14] , \nOut0_33[13] , \nOut0_33[12] , 
        \nOut0_33[11] , \nOut0_33[10] , \nOut0_33[9] , \nOut0_33[8] , 
        \nOut0_33[7] , \nOut0_33[6] , \nOut0_33[5] , \nOut0_33[4] , 
        \nOut0_33[3] , \nOut0_33[2] , \nOut0_33[1] , \nOut0_33[0] }), 
        .SOUTH_EDGE({\nOut0_35[31] , \nOut0_35[30] , \nOut0_35[29] , 
        \nOut0_35[28] , \nOut0_35[27] , \nOut0_35[26] , \nOut0_35[25] , 
        \nOut0_35[24] , \nOut0_35[23] , \nOut0_35[22] , \nOut0_35[21] , 
        \nOut0_35[20] , \nOut0_35[19] , \nOut0_35[18] , \nOut0_35[17] , 
        \nOut0_35[16] , \nOut0_35[15] , \nOut0_35[14] , \nOut0_35[13] , 
        \nOut0_35[12] , \nOut0_35[11] , \nOut0_35[10] , \nOut0_35[9] , 
        \nOut0_35[8] , \nOut0_35[7] , \nOut0_35[6] , \nOut0_35[5] , 
        \nOut0_35[4] , \nOut0_35[3] , \nOut0_35[2] , \nOut0_35[1] , 
        \nOut0_35[0] }), .EAST_EDGE(\nOut1_34[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_33[31] ), .SE_EDGE(
        \nOut1_35[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_48 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut49[31] , \nScanOut49[30] , \nScanOut49[29] , 
        \nScanOut49[28] , \nScanOut49[27] , \nScanOut49[26] , \nScanOut49[25] , 
        \nScanOut49[24] , \nScanOut49[23] , \nScanOut49[22] , \nScanOut49[21] , 
        \nScanOut49[20] , \nScanOut49[19] , \nScanOut49[18] , \nScanOut49[17] , 
        \nScanOut49[16] , \nScanOut49[15] , \nScanOut49[14] , \nScanOut49[13] , 
        \nScanOut49[12] , \nScanOut49[11] , \nScanOut49[10] , \nScanOut49[9] , 
        \nScanOut49[8] , \nScanOut49[7] , \nScanOut49[6] , \nScanOut49[5] , 
        \nScanOut49[4] , \nScanOut49[3] , \nScanOut49[2] , \nScanOut49[1] , 
        \nScanOut49[0] }), .ScanOut({\nScanOut48[31] , \nScanOut48[30] , 
        \nScanOut48[29] , \nScanOut48[28] , \nScanOut48[27] , \nScanOut48[26] , 
        \nScanOut48[25] , \nScanOut48[24] , \nScanOut48[23] , \nScanOut48[22] , 
        \nScanOut48[21] , \nScanOut48[20] , \nScanOut48[19] , \nScanOut48[18] , 
        \nScanOut48[17] , \nScanOut48[16] , \nScanOut48[15] , \nScanOut48[14] , 
        \nScanOut48[13] , \nScanOut48[12] , \nScanOut48[11] , \nScanOut48[10] , 
        \nScanOut48[9] , \nScanOut48[8] , \nScanOut48[7] , \nScanOut48[6] , 
        \nScanOut48[5] , \nScanOut48[4] , \nScanOut48[3] , \nScanOut48[2] , 
        \nScanOut48[1] , \nScanOut48[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_48[31] , 
        \nOut0_48[30] , \nOut0_48[29] , \nOut0_48[28] , \nOut0_48[27] , 
        \nOut0_48[26] , \nOut0_48[25] , \nOut0_48[24] , \nOut0_48[23] , 
        \nOut0_48[22] , \nOut0_48[21] , \nOut0_48[20] , \nOut0_48[19] , 
        \nOut0_48[18] , \nOut0_48[17] , \nOut0_48[16] , \nOut0_48[15] , 
        \nOut0_48[14] , \nOut0_48[13] , \nOut0_48[12] , \nOut0_48[11] , 
        \nOut0_48[10] , \nOut0_48[9] , \nOut0_48[8] , \nOut0_48[7] , 
        \nOut0_48[6] , \nOut0_48[5] , \nOut0_48[4] , \nOut0_48[3] , 
        \nOut0_48[2] , \nOut0_48[1] , \nOut0_48[0] }), .NORTH_EDGE({
        \nOut0_47[31] , \nOut0_47[30] , \nOut0_47[29] , \nOut0_47[28] , 
        \nOut0_47[27] , \nOut0_47[26] , \nOut0_47[25] , \nOut0_47[24] , 
        \nOut0_47[23] , \nOut0_47[22] , \nOut0_47[21] , \nOut0_47[20] , 
        \nOut0_47[19] , \nOut0_47[18] , \nOut0_47[17] , \nOut0_47[16] , 
        \nOut0_47[15] , \nOut0_47[14] , \nOut0_47[13] , \nOut0_47[12] , 
        \nOut0_47[11] , \nOut0_47[10] , \nOut0_47[9] , \nOut0_47[8] , 
        \nOut0_47[7] , \nOut0_47[6] , \nOut0_47[5] , \nOut0_47[4] , 
        \nOut0_47[3] , \nOut0_47[2] , \nOut0_47[1] , \nOut0_47[0] }), 
        .SOUTH_EDGE({\nOut0_49[31] , \nOut0_49[30] , \nOut0_49[29] , 
        \nOut0_49[28] , \nOut0_49[27] , \nOut0_49[26] , \nOut0_49[25] , 
        \nOut0_49[24] , \nOut0_49[23] , \nOut0_49[22] , \nOut0_49[21] , 
        \nOut0_49[20] , \nOut0_49[19] , \nOut0_49[18] , \nOut0_49[17] , 
        \nOut0_49[16] , \nOut0_49[15] , \nOut0_49[14] , \nOut0_49[13] , 
        \nOut0_49[12] , \nOut0_49[11] , \nOut0_49[10] , \nOut0_49[9] , 
        \nOut0_49[8] , \nOut0_49[7] , \nOut0_49[6] , \nOut0_49[5] , 
        \nOut0_49[4] , \nOut0_49[3] , \nOut0_49[2] , \nOut0_49[1] , 
        \nOut0_49[0] }), .EAST_EDGE(\nOut1_48[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_47[31] ), .SE_EDGE(
        \nOut1_49[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_53 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut54[31] , \nScanOut54[30] , \nScanOut54[29] , 
        \nScanOut54[28] , \nScanOut54[27] , \nScanOut54[26] , \nScanOut54[25] , 
        \nScanOut54[24] , \nScanOut54[23] , \nScanOut54[22] , \nScanOut54[21] , 
        \nScanOut54[20] , \nScanOut54[19] , \nScanOut54[18] , \nScanOut54[17] , 
        \nScanOut54[16] , \nScanOut54[15] , \nScanOut54[14] , \nScanOut54[13] , 
        \nScanOut54[12] , \nScanOut54[11] , \nScanOut54[10] , \nScanOut54[9] , 
        \nScanOut54[8] , \nScanOut54[7] , \nScanOut54[6] , \nScanOut54[5] , 
        \nScanOut54[4] , \nScanOut54[3] , \nScanOut54[2] , \nScanOut54[1] , 
        \nScanOut54[0] }), .ScanOut({\nScanOut53[31] , \nScanOut53[30] , 
        \nScanOut53[29] , \nScanOut53[28] , \nScanOut53[27] , \nScanOut53[26] , 
        \nScanOut53[25] , \nScanOut53[24] , \nScanOut53[23] , \nScanOut53[22] , 
        \nScanOut53[21] , \nScanOut53[20] , \nScanOut53[19] , \nScanOut53[18] , 
        \nScanOut53[17] , \nScanOut53[16] , \nScanOut53[15] , \nScanOut53[14] , 
        \nScanOut53[13] , \nScanOut53[12] , \nScanOut53[11] , \nScanOut53[10] , 
        \nScanOut53[9] , \nScanOut53[8] , \nScanOut53[7] , \nScanOut53[6] , 
        \nScanOut53[5] , \nScanOut53[4] , \nScanOut53[3] , \nScanOut53[2] , 
        \nScanOut53[1] , \nScanOut53[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_53[31] , 
        \nOut0_53[30] , \nOut0_53[29] , \nOut0_53[28] , \nOut0_53[27] , 
        \nOut0_53[26] , \nOut0_53[25] , \nOut0_53[24] , \nOut0_53[23] , 
        \nOut0_53[22] , \nOut0_53[21] , \nOut0_53[20] , \nOut0_53[19] , 
        \nOut0_53[18] , \nOut0_53[17] , \nOut0_53[16] , \nOut0_53[15] , 
        \nOut0_53[14] , \nOut0_53[13] , \nOut0_53[12] , \nOut0_53[11] , 
        \nOut0_53[10] , \nOut0_53[9] , \nOut0_53[8] , \nOut0_53[7] , 
        \nOut0_53[6] , \nOut0_53[5] , \nOut0_53[4] , \nOut0_53[3] , 
        \nOut0_53[2] , \nOut0_53[1] , \nOut0_53[0] }), .NORTH_EDGE({
        \nOut0_52[31] , \nOut0_52[30] , \nOut0_52[29] , \nOut0_52[28] , 
        \nOut0_52[27] , \nOut0_52[26] , \nOut0_52[25] , \nOut0_52[24] , 
        \nOut0_52[23] , \nOut0_52[22] , \nOut0_52[21] , \nOut0_52[20] , 
        \nOut0_52[19] , \nOut0_52[18] , \nOut0_52[17] , \nOut0_52[16] , 
        \nOut0_52[15] , \nOut0_52[14] , \nOut0_52[13] , \nOut0_52[12] , 
        \nOut0_52[11] , \nOut0_52[10] , \nOut0_52[9] , \nOut0_52[8] , 
        \nOut0_52[7] , \nOut0_52[6] , \nOut0_52[5] , \nOut0_52[4] , 
        \nOut0_52[3] , \nOut0_52[2] , \nOut0_52[1] , \nOut0_52[0] }), 
        .SOUTH_EDGE({\nOut0_54[31] , \nOut0_54[30] , \nOut0_54[29] , 
        \nOut0_54[28] , \nOut0_54[27] , \nOut0_54[26] , \nOut0_54[25] , 
        \nOut0_54[24] , \nOut0_54[23] , \nOut0_54[22] , \nOut0_54[21] , 
        \nOut0_54[20] , \nOut0_54[19] , \nOut0_54[18] , \nOut0_54[17] , 
        \nOut0_54[16] , \nOut0_54[15] , \nOut0_54[14] , \nOut0_54[13] , 
        \nOut0_54[12] , \nOut0_54[11] , \nOut0_54[10] , \nOut0_54[9] , 
        \nOut0_54[8] , \nOut0_54[7] , \nOut0_54[6] , \nOut0_54[5] , 
        \nOut0_54[4] , \nOut0_54[3] , \nOut0_54[2] , \nOut0_54[1] , 
        \nOut0_54[0] }), .EAST_EDGE(\nOut1_53[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_52[31] ), .SE_EDGE(
        \nOut1_54[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_74 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut75[31] , \nScanOut75[30] , \nScanOut75[29] , 
        \nScanOut75[28] , \nScanOut75[27] , \nScanOut75[26] , \nScanOut75[25] , 
        \nScanOut75[24] , \nScanOut75[23] , \nScanOut75[22] , \nScanOut75[21] , 
        \nScanOut75[20] , \nScanOut75[19] , \nScanOut75[18] , \nScanOut75[17] , 
        \nScanOut75[16] , \nScanOut75[15] , \nScanOut75[14] , \nScanOut75[13] , 
        \nScanOut75[12] , \nScanOut75[11] , \nScanOut75[10] , \nScanOut75[9] , 
        \nScanOut75[8] , \nScanOut75[7] , \nScanOut75[6] , \nScanOut75[5] , 
        \nScanOut75[4] , \nScanOut75[3] , \nScanOut75[2] , \nScanOut75[1] , 
        \nScanOut75[0] }), .ScanOut({\nScanOut74[31] , \nScanOut74[30] , 
        \nScanOut74[29] , \nScanOut74[28] , \nScanOut74[27] , \nScanOut74[26] , 
        \nScanOut74[25] , \nScanOut74[24] , \nScanOut74[23] , \nScanOut74[22] , 
        \nScanOut74[21] , \nScanOut74[20] , \nScanOut74[19] , \nScanOut74[18] , 
        \nScanOut74[17] , \nScanOut74[16] , \nScanOut74[15] , \nScanOut74[14] , 
        \nScanOut74[13] , \nScanOut74[12] , \nScanOut74[11] , \nScanOut74[10] , 
        \nScanOut74[9] , \nScanOut74[8] , \nScanOut74[7] , \nScanOut74[6] , 
        \nScanOut74[5] , \nScanOut74[4] , \nScanOut74[3] , \nScanOut74[2] , 
        \nScanOut74[1] , \nScanOut74[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_10[31] , 
        \nOut1_10[30] , \nOut1_10[29] , \nOut1_10[28] , \nOut1_10[27] , 
        \nOut1_10[26] , \nOut1_10[25] , \nOut1_10[24] , \nOut1_10[23] , 
        \nOut1_10[22] , \nOut1_10[21] , \nOut1_10[20] , \nOut1_10[19] , 
        \nOut1_10[18] , \nOut1_10[17] , \nOut1_10[16] , \nOut1_10[15] , 
        \nOut1_10[14] , \nOut1_10[13] , \nOut1_10[12] , \nOut1_10[11] , 
        \nOut1_10[10] , \nOut1_10[9] , \nOut1_10[8] , \nOut1_10[7] , 
        \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , \nOut1_10[3] , 
        \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), .NORTH_EDGE({
        \nOut1_9[31] , \nOut1_9[30] , \nOut1_9[29] , \nOut1_9[28] , 
        \nOut1_9[27] , \nOut1_9[26] , \nOut1_9[25] , \nOut1_9[24] , 
        \nOut1_9[23] , \nOut1_9[22] , \nOut1_9[21] , \nOut1_9[20] , 
        \nOut1_9[19] , \nOut1_9[18] , \nOut1_9[17] , \nOut1_9[16] , 
        \nOut1_9[15] , \nOut1_9[14] , \nOut1_9[13] , \nOut1_9[12] , 
        \nOut1_9[11] , \nOut1_9[10] , \nOut1_9[9] , \nOut1_9[8] , \nOut1_9[7] , 
        \nOut1_9[6] , \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , 
        \nOut1_9[1] , \nOut1_9[0] }), .SOUTH_EDGE({\nOut1_11[31] , 
        \nOut1_11[30] , \nOut1_11[29] , \nOut1_11[28] , \nOut1_11[27] , 
        \nOut1_11[26] , \nOut1_11[25] , \nOut1_11[24] , \nOut1_11[23] , 
        \nOut1_11[22] , \nOut1_11[21] , \nOut1_11[20] , \nOut1_11[19] , 
        \nOut1_11[18] , \nOut1_11[17] , \nOut1_11[16] , \nOut1_11[15] , 
        \nOut1_11[14] , \nOut1_11[13] , \nOut1_11[12] , \nOut1_11[11] , 
        \nOut1_11[10] , \nOut1_11[9] , \nOut1_11[8] , \nOut1_11[7] , 
        \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , \nOut1_11[3] , 
        \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_10[0] ), .NW_EDGE(\nOut0_9[0] ), .SW_EDGE(
        \nOut0_11[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_105 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut106[31] , \nScanOut106[30] , \nScanOut106[29] , 
        \nScanOut106[28] , \nScanOut106[27] , \nScanOut106[26] , 
        \nScanOut106[25] , \nScanOut106[24] , \nScanOut106[23] , 
        \nScanOut106[22] , \nScanOut106[21] , \nScanOut106[20] , 
        \nScanOut106[19] , \nScanOut106[18] , \nScanOut106[17] , 
        \nScanOut106[16] , \nScanOut106[15] , \nScanOut106[14] , 
        \nScanOut106[13] , \nScanOut106[12] , \nScanOut106[11] , 
        \nScanOut106[10] , \nScanOut106[9] , \nScanOut106[8] , 
        \nScanOut106[7] , \nScanOut106[6] , \nScanOut106[5] , \nScanOut106[4] , 
        \nScanOut106[3] , \nScanOut106[2] , \nScanOut106[1] , \nScanOut106[0] 
        }), .ScanOut({\nScanOut105[31] , \nScanOut105[30] , \nScanOut105[29] , 
        \nScanOut105[28] , \nScanOut105[27] , \nScanOut105[26] , 
        \nScanOut105[25] , \nScanOut105[24] , \nScanOut105[23] , 
        \nScanOut105[22] , \nScanOut105[21] , \nScanOut105[20] , 
        \nScanOut105[19] , \nScanOut105[18] , \nScanOut105[17] , 
        \nScanOut105[16] , \nScanOut105[15] , \nScanOut105[14] , 
        \nScanOut105[13] , \nScanOut105[12] , \nScanOut105[11] , 
        \nScanOut105[10] , \nScanOut105[9] , \nScanOut105[8] , 
        \nScanOut105[7] , \nScanOut105[6] , \nScanOut105[5] , \nScanOut105[4] , 
        \nScanOut105[3] , \nScanOut105[2] , \nScanOut105[1] , \nScanOut105[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_41[31] , \nOut1_41[30] , \nOut1_41[29] , 
        \nOut1_41[28] , \nOut1_41[27] , \nOut1_41[26] , \nOut1_41[25] , 
        \nOut1_41[24] , \nOut1_41[23] , \nOut1_41[22] , \nOut1_41[21] , 
        \nOut1_41[20] , \nOut1_41[19] , \nOut1_41[18] , \nOut1_41[17] , 
        \nOut1_41[16] , \nOut1_41[15] , \nOut1_41[14] , \nOut1_41[13] , 
        \nOut1_41[12] , \nOut1_41[11] , \nOut1_41[10] , \nOut1_41[9] , 
        \nOut1_41[8] , \nOut1_41[7] , \nOut1_41[6] , \nOut1_41[5] , 
        \nOut1_41[4] , \nOut1_41[3] , \nOut1_41[2] , \nOut1_41[1] , 
        \nOut1_41[0] }), .NORTH_EDGE({\nOut1_40[31] , \nOut1_40[30] , 
        \nOut1_40[29] , \nOut1_40[28] , \nOut1_40[27] , \nOut1_40[26] , 
        \nOut1_40[25] , \nOut1_40[24] , \nOut1_40[23] , \nOut1_40[22] , 
        \nOut1_40[21] , \nOut1_40[20] , \nOut1_40[19] , \nOut1_40[18] , 
        \nOut1_40[17] , \nOut1_40[16] , \nOut1_40[15] , \nOut1_40[14] , 
        \nOut1_40[13] , \nOut1_40[12] , \nOut1_40[11] , \nOut1_40[10] , 
        \nOut1_40[9] , \nOut1_40[8] , \nOut1_40[7] , \nOut1_40[6] , 
        \nOut1_40[5] , \nOut1_40[4] , \nOut1_40[3] , \nOut1_40[2] , 
        \nOut1_40[1] , \nOut1_40[0] }), .SOUTH_EDGE({\nOut1_42[31] , 
        \nOut1_42[30] , \nOut1_42[29] , \nOut1_42[28] , \nOut1_42[27] , 
        \nOut1_42[26] , \nOut1_42[25] , \nOut1_42[24] , \nOut1_42[23] , 
        \nOut1_42[22] , \nOut1_42[21] , \nOut1_42[20] , \nOut1_42[19] , 
        \nOut1_42[18] , \nOut1_42[17] , \nOut1_42[16] , \nOut1_42[15] , 
        \nOut1_42[14] , \nOut1_42[13] , \nOut1_42[12] , \nOut1_42[11] , 
        \nOut1_42[10] , \nOut1_42[9] , \nOut1_42[8] , \nOut1_42[7] , 
        \nOut1_42[6] , \nOut1_42[5] , \nOut1_42[4] , \nOut1_42[3] , 
        \nOut1_42[2] , \nOut1_42[1] , \nOut1_42[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_41[0] ), .NW_EDGE(\nOut0_40[0] ), .SW_EDGE(
        \nOut0_42[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_122 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut123[31] , \nScanOut123[30] , \nScanOut123[29] , 
        \nScanOut123[28] , \nScanOut123[27] , \nScanOut123[26] , 
        \nScanOut123[25] , \nScanOut123[24] , \nScanOut123[23] , 
        \nScanOut123[22] , \nScanOut123[21] , \nScanOut123[20] , 
        \nScanOut123[19] , \nScanOut123[18] , \nScanOut123[17] , 
        \nScanOut123[16] , \nScanOut123[15] , \nScanOut123[14] , 
        \nScanOut123[13] , \nScanOut123[12] , \nScanOut123[11] , 
        \nScanOut123[10] , \nScanOut123[9] , \nScanOut123[8] , 
        \nScanOut123[7] , \nScanOut123[6] , \nScanOut123[5] , \nScanOut123[4] , 
        \nScanOut123[3] , \nScanOut123[2] , \nScanOut123[1] , \nScanOut123[0] 
        }), .ScanOut({\nScanOut122[31] , \nScanOut122[30] , \nScanOut122[29] , 
        \nScanOut122[28] , \nScanOut122[27] , \nScanOut122[26] , 
        \nScanOut122[25] , \nScanOut122[24] , \nScanOut122[23] , 
        \nScanOut122[22] , \nScanOut122[21] , \nScanOut122[20] , 
        \nScanOut122[19] , \nScanOut122[18] , \nScanOut122[17] , 
        \nScanOut122[16] , \nScanOut122[15] , \nScanOut122[14] , 
        \nScanOut122[13] , \nScanOut122[12] , \nScanOut122[11] , 
        \nScanOut122[10] , \nScanOut122[9] , \nScanOut122[8] , 
        \nScanOut122[7] , \nScanOut122[6] , \nScanOut122[5] , \nScanOut122[4] , 
        \nScanOut122[3] , \nScanOut122[2] , \nScanOut122[1] , \nScanOut122[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_58[31] , \nOut1_58[30] , \nOut1_58[29] , 
        \nOut1_58[28] , \nOut1_58[27] , \nOut1_58[26] , \nOut1_58[25] , 
        \nOut1_58[24] , \nOut1_58[23] , \nOut1_58[22] , \nOut1_58[21] , 
        \nOut1_58[20] , \nOut1_58[19] , \nOut1_58[18] , \nOut1_58[17] , 
        \nOut1_58[16] , \nOut1_58[15] , \nOut1_58[14] , \nOut1_58[13] , 
        \nOut1_58[12] , \nOut1_58[11] , \nOut1_58[10] , \nOut1_58[9] , 
        \nOut1_58[8] , \nOut1_58[7] , \nOut1_58[6] , \nOut1_58[5] , 
        \nOut1_58[4] , \nOut1_58[3] , \nOut1_58[2] , \nOut1_58[1] , 
        \nOut1_58[0] }), .NORTH_EDGE({\nOut1_57[31] , \nOut1_57[30] , 
        \nOut1_57[29] , \nOut1_57[28] , \nOut1_57[27] , \nOut1_57[26] , 
        \nOut1_57[25] , \nOut1_57[24] , \nOut1_57[23] , \nOut1_57[22] , 
        \nOut1_57[21] , \nOut1_57[20] , \nOut1_57[19] , \nOut1_57[18] , 
        \nOut1_57[17] , \nOut1_57[16] , \nOut1_57[15] , \nOut1_57[14] , 
        \nOut1_57[13] , \nOut1_57[12] , \nOut1_57[11] , \nOut1_57[10] , 
        \nOut1_57[9] , \nOut1_57[8] , \nOut1_57[7] , \nOut1_57[6] , 
        \nOut1_57[5] , \nOut1_57[4] , \nOut1_57[3] , \nOut1_57[2] , 
        \nOut1_57[1] , \nOut1_57[0] }), .SOUTH_EDGE({\nOut1_59[31] , 
        \nOut1_59[30] , \nOut1_59[29] , \nOut1_59[28] , \nOut1_59[27] , 
        \nOut1_59[26] , \nOut1_59[25] , \nOut1_59[24] , \nOut1_59[23] , 
        \nOut1_59[22] , \nOut1_59[21] , \nOut1_59[20] , \nOut1_59[19] , 
        \nOut1_59[18] , \nOut1_59[17] , \nOut1_59[16] , \nOut1_59[15] , 
        \nOut1_59[14] , \nOut1_59[13] , \nOut1_59[12] , \nOut1_59[11] , 
        \nOut1_59[10] , \nOut1_59[9] , \nOut1_59[8] , \nOut1_59[7] , 
        \nOut1_59[6] , \nOut1_59[5] , \nOut1_59[4] , \nOut1_59[3] , 
        \nOut1_59[2] , \nOut1_59[1] , \nOut1_59[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_58[0] ), .NW_EDGE(\nOut0_57[0] ), .SW_EDGE(
        \nOut0_59[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut6[31] , \nScanOut6[30] , \nScanOut6[29] , 
        \nScanOut6[28] , \nScanOut6[27] , \nScanOut6[26] , \nScanOut6[25] , 
        \nScanOut6[24] , \nScanOut6[23] , \nScanOut6[22] , \nScanOut6[21] , 
        \nScanOut6[20] , \nScanOut6[19] , \nScanOut6[18] , \nScanOut6[17] , 
        \nScanOut6[16] , \nScanOut6[15] , \nScanOut6[14] , \nScanOut6[13] , 
        \nScanOut6[12] , \nScanOut6[11] , \nScanOut6[10] , \nScanOut6[9] , 
        \nScanOut6[8] , \nScanOut6[7] , \nScanOut6[6] , \nScanOut6[5] , 
        \nScanOut6[4] , \nScanOut6[3] , \nScanOut6[2] , \nScanOut6[1] , 
        \nScanOut6[0] }), .ScanOut({\nScanOut5[31] , \nScanOut5[30] , 
        \nScanOut5[29] , \nScanOut5[28] , \nScanOut5[27] , \nScanOut5[26] , 
        \nScanOut5[25] , \nScanOut5[24] , \nScanOut5[23] , \nScanOut5[22] , 
        \nScanOut5[21] , \nScanOut5[20] , \nScanOut5[19] , \nScanOut5[18] , 
        \nScanOut5[17] , \nScanOut5[16] , \nScanOut5[15] , \nScanOut5[14] , 
        \nScanOut5[13] , \nScanOut5[12] , \nScanOut5[11] , \nScanOut5[10] , 
        \nScanOut5[9] , \nScanOut5[8] , \nScanOut5[7] , \nScanOut5[6] , 
        \nScanOut5[5] , \nScanOut5[4] , \nScanOut5[3] , \nScanOut5[2] , 
        \nScanOut5[1] , \nScanOut5[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_5[31] , 
        \nOut0_5[30] , \nOut0_5[29] , \nOut0_5[28] , \nOut0_5[27] , 
        \nOut0_5[26] , \nOut0_5[25] , \nOut0_5[24] , \nOut0_5[23] , 
        \nOut0_5[22] , \nOut0_5[21] , \nOut0_5[20] , \nOut0_5[19] , 
        \nOut0_5[18] , \nOut0_5[17] , \nOut0_5[16] , \nOut0_5[15] , 
        \nOut0_5[14] , \nOut0_5[13] , \nOut0_5[12] , \nOut0_5[11] , 
        \nOut0_5[10] , \nOut0_5[9] , \nOut0_5[8] , \nOut0_5[7] , \nOut0_5[6] , 
        \nOut0_5[5] , \nOut0_5[4] , \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , 
        \nOut0_5[0] }), .NORTH_EDGE({\nOut0_4[31] , \nOut0_4[30] , 
        \nOut0_4[29] , \nOut0_4[28] , \nOut0_4[27] , \nOut0_4[26] , 
        \nOut0_4[25] , \nOut0_4[24] , \nOut0_4[23] , \nOut0_4[22] , 
        \nOut0_4[21] , \nOut0_4[20] , \nOut0_4[19] , \nOut0_4[18] , 
        \nOut0_4[17] , \nOut0_4[16] , \nOut0_4[15] , \nOut0_4[14] , 
        \nOut0_4[13] , \nOut0_4[12] , \nOut0_4[11] , \nOut0_4[10] , 
        \nOut0_4[9] , \nOut0_4[8] , \nOut0_4[7] , \nOut0_4[6] , \nOut0_4[5] , 
        \nOut0_4[4] , \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , \nOut0_4[0] }), 
        .SOUTH_EDGE({\nOut0_6[31] , \nOut0_6[30] , \nOut0_6[29] , 
        \nOut0_6[28] , \nOut0_6[27] , \nOut0_6[26] , \nOut0_6[25] , 
        \nOut0_6[24] , \nOut0_6[23] , \nOut0_6[22] , \nOut0_6[21] , 
        \nOut0_6[20] , \nOut0_6[19] , \nOut0_6[18] , \nOut0_6[17] , 
        \nOut0_6[16] , \nOut0_6[15] , \nOut0_6[14] , \nOut0_6[13] , 
        \nOut0_6[12] , \nOut0_6[11] , \nOut0_6[10] , \nOut0_6[9] , 
        \nOut0_6[8] , \nOut0_6[7] , \nOut0_6[6] , \nOut0_6[5] , \nOut0_6[4] , 
        \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , \nOut0_6[0] }), .EAST_EDGE(
        \nOut1_5[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_4[31] ), .SE_EDGE(\nOut1_6[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut13[31] , \nScanOut13[30] , \nScanOut13[29] , 
        \nScanOut13[28] , \nScanOut13[27] , \nScanOut13[26] , \nScanOut13[25] , 
        \nScanOut13[24] , \nScanOut13[23] , \nScanOut13[22] , \nScanOut13[21] , 
        \nScanOut13[20] , \nScanOut13[19] , \nScanOut13[18] , \nScanOut13[17] , 
        \nScanOut13[16] , \nScanOut13[15] , \nScanOut13[14] , \nScanOut13[13] , 
        \nScanOut13[12] , \nScanOut13[11] , \nScanOut13[10] , \nScanOut13[9] , 
        \nScanOut13[8] , \nScanOut13[7] , \nScanOut13[6] , \nScanOut13[5] , 
        \nScanOut13[4] , \nScanOut13[3] , \nScanOut13[2] , \nScanOut13[1] , 
        \nScanOut13[0] }), .ScanOut({\nScanOut12[31] , \nScanOut12[30] , 
        \nScanOut12[29] , \nScanOut12[28] , \nScanOut12[27] , \nScanOut12[26] , 
        \nScanOut12[25] , \nScanOut12[24] , \nScanOut12[23] , \nScanOut12[22] , 
        \nScanOut12[21] , \nScanOut12[20] , \nScanOut12[19] , \nScanOut12[18] , 
        \nScanOut12[17] , \nScanOut12[16] , \nScanOut12[15] , \nScanOut12[14] , 
        \nScanOut12[13] , \nScanOut12[12] , \nScanOut12[11] , \nScanOut12[10] , 
        \nScanOut12[9] , \nScanOut12[8] , \nScanOut12[7] , \nScanOut12[6] , 
        \nScanOut12[5] , \nScanOut12[4] , \nScanOut12[3] , \nScanOut12[2] , 
        \nScanOut12[1] , \nScanOut12[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_12[31] , 
        \nOut0_12[30] , \nOut0_12[29] , \nOut0_12[28] , \nOut0_12[27] , 
        \nOut0_12[26] , \nOut0_12[25] , \nOut0_12[24] , \nOut0_12[23] , 
        \nOut0_12[22] , \nOut0_12[21] , \nOut0_12[20] , \nOut0_12[19] , 
        \nOut0_12[18] , \nOut0_12[17] , \nOut0_12[16] , \nOut0_12[15] , 
        \nOut0_12[14] , \nOut0_12[13] , \nOut0_12[12] , \nOut0_12[11] , 
        \nOut0_12[10] , \nOut0_12[9] , \nOut0_12[8] , \nOut0_12[7] , 
        \nOut0_12[6] , \nOut0_12[5] , \nOut0_12[4] , \nOut0_12[3] , 
        \nOut0_12[2] , \nOut0_12[1] , \nOut0_12[0] }), .NORTH_EDGE({
        \nOut0_11[31] , \nOut0_11[30] , \nOut0_11[29] , \nOut0_11[28] , 
        \nOut0_11[27] , \nOut0_11[26] , \nOut0_11[25] , \nOut0_11[24] , 
        \nOut0_11[23] , \nOut0_11[22] , \nOut0_11[21] , \nOut0_11[20] , 
        \nOut0_11[19] , \nOut0_11[18] , \nOut0_11[17] , \nOut0_11[16] , 
        \nOut0_11[15] , \nOut0_11[14] , \nOut0_11[13] , \nOut0_11[12] , 
        \nOut0_11[11] , \nOut0_11[10] , \nOut0_11[9] , \nOut0_11[8] , 
        \nOut0_11[7] , \nOut0_11[6] , \nOut0_11[5] , \nOut0_11[4] , 
        \nOut0_11[3] , \nOut0_11[2] , \nOut0_11[1] , \nOut0_11[0] }), 
        .SOUTH_EDGE({\nOut0_13[31] , \nOut0_13[30] , \nOut0_13[29] , 
        \nOut0_13[28] , \nOut0_13[27] , \nOut0_13[26] , \nOut0_13[25] , 
        \nOut0_13[24] , \nOut0_13[23] , \nOut0_13[22] , \nOut0_13[21] , 
        \nOut0_13[20] , \nOut0_13[19] , \nOut0_13[18] , \nOut0_13[17] , 
        \nOut0_13[16] , \nOut0_13[15] , \nOut0_13[14] , \nOut0_13[13] , 
        \nOut0_13[12] , \nOut0_13[11] , \nOut0_13[10] , \nOut0_13[9] , 
        \nOut0_13[8] , \nOut0_13[7] , \nOut0_13[6] , \nOut0_13[5] , 
        \nOut0_13[4] , \nOut0_13[3] , \nOut0_13[2] , \nOut0_13[1] , 
        \nOut0_13[0] }), .EAST_EDGE(\nOut1_12[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_11[31] ), .SE_EDGE(
        \nOut1_13[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_91 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut92[31] , \nScanOut92[30] , \nScanOut92[29] , 
        \nScanOut92[28] , \nScanOut92[27] , \nScanOut92[26] , \nScanOut92[25] , 
        \nScanOut92[24] , \nScanOut92[23] , \nScanOut92[22] , \nScanOut92[21] , 
        \nScanOut92[20] , \nScanOut92[19] , \nScanOut92[18] , \nScanOut92[17] , 
        \nScanOut92[16] , \nScanOut92[15] , \nScanOut92[14] , \nScanOut92[13] , 
        \nScanOut92[12] , \nScanOut92[11] , \nScanOut92[10] , \nScanOut92[9] , 
        \nScanOut92[8] , \nScanOut92[7] , \nScanOut92[6] , \nScanOut92[5] , 
        \nScanOut92[4] , \nScanOut92[3] , \nScanOut92[2] , \nScanOut92[1] , 
        \nScanOut92[0] }), .ScanOut({\nScanOut91[31] , \nScanOut91[30] , 
        \nScanOut91[29] , \nScanOut91[28] , \nScanOut91[27] , \nScanOut91[26] , 
        \nScanOut91[25] , \nScanOut91[24] , \nScanOut91[23] , \nScanOut91[22] , 
        \nScanOut91[21] , \nScanOut91[20] , \nScanOut91[19] , \nScanOut91[18] , 
        \nScanOut91[17] , \nScanOut91[16] , \nScanOut91[15] , \nScanOut91[14] , 
        \nScanOut91[13] , \nScanOut91[12] , \nScanOut91[11] , \nScanOut91[10] , 
        \nScanOut91[9] , \nScanOut91[8] , \nScanOut91[7] , \nScanOut91[6] , 
        \nScanOut91[5] , \nScanOut91[4] , \nScanOut91[3] , \nScanOut91[2] , 
        \nScanOut91[1] , \nScanOut91[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_27[31] , 
        \nOut1_27[30] , \nOut1_27[29] , \nOut1_27[28] , \nOut1_27[27] , 
        \nOut1_27[26] , \nOut1_27[25] , \nOut1_27[24] , \nOut1_27[23] , 
        \nOut1_27[22] , \nOut1_27[21] , \nOut1_27[20] , \nOut1_27[19] , 
        \nOut1_27[18] , \nOut1_27[17] , \nOut1_27[16] , \nOut1_27[15] , 
        \nOut1_27[14] , \nOut1_27[13] , \nOut1_27[12] , \nOut1_27[11] , 
        \nOut1_27[10] , \nOut1_27[9] , \nOut1_27[8] , \nOut1_27[7] , 
        \nOut1_27[6] , \nOut1_27[5] , \nOut1_27[4] , \nOut1_27[3] , 
        \nOut1_27[2] , \nOut1_27[1] , \nOut1_27[0] }), .NORTH_EDGE({
        \nOut1_26[31] , \nOut1_26[30] , \nOut1_26[29] , \nOut1_26[28] , 
        \nOut1_26[27] , \nOut1_26[26] , \nOut1_26[25] , \nOut1_26[24] , 
        \nOut1_26[23] , \nOut1_26[22] , \nOut1_26[21] , \nOut1_26[20] , 
        \nOut1_26[19] , \nOut1_26[18] , \nOut1_26[17] , \nOut1_26[16] , 
        \nOut1_26[15] , \nOut1_26[14] , \nOut1_26[13] , \nOut1_26[12] , 
        \nOut1_26[11] , \nOut1_26[10] , \nOut1_26[9] , \nOut1_26[8] , 
        \nOut1_26[7] , \nOut1_26[6] , \nOut1_26[5] , \nOut1_26[4] , 
        \nOut1_26[3] , \nOut1_26[2] , \nOut1_26[1] , \nOut1_26[0] }), 
        .SOUTH_EDGE({\nOut1_28[31] , \nOut1_28[30] , \nOut1_28[29] , 
        \nOut1_28[28] , \nOut1_28[27] , \nOut1_28[26] , \nOut1_28[25] , 
        \nOut1_28[24] , \nOut1_28[23] , \nOut1_28[22] , \nOut1_28[21] , 
        \nOut1_28[20] , \nOut1_28[19] , \nOut1_28[18] , \nOut1_28[17] , 
        \nOut1_28[16] , \nOut1_28[15] , \nOut1_28[14] , \nOut1_28[13] , 
        \nOut1_28[12] , \nOut1_28[11] , \nOut1_28[10] , \nOut1_28[9] , 
        \nOut1_28[8] , \nOut1_28[7] , \nOut1_28[6] , \nOut1_28[5] , 
        \nOut1_28[4] , \nOut1_28[3] , \nOut1_28[2] , \nOut1_28[1] , 
        \nOut1_28[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_27[0] ), 
        .NW_EDGE(\nOut0_26[0] ), .SW_EDGE(\nOut0_28[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_99 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut100[31] , \nScanOut100[30] , \nScanOut100[29] , 
        \nScanOut100[28] , \nScanOut100[27] , \nScanOut100[26] , 
        \nScanOut100[25] , \nScanOut100[24] , \nScanOut100[23] , 
        \nScanOut100[22] , \nScanOut100[21] , \nScanOut100[20] , 
        \nScanOut100[19] , \nScanOut100[18] , \nScanOut100[17] , 
        \nScanOut100[16] , \nScanOut100[15] , \nScanOut100[14] , 
        \nScanOut100[13] , \nScanOut100[12] , \nScanOut100[11] , 
        \nScanOut100[10] , \nScanOut100[9] , \nScanOut100[8] , 
        \nScanOut100[7] , \nScanOut100[6] , \nScanOut100[5] , \nScanOut100[4] , 
        \nScanOut100[3] , \nScanOut100[2] , \nScanOut100[1] , \nScanOut100[0] 
        }), .ScanOut({\nScanOut99[31] , \nScanOut99[30] , \nScanOut99[29] , 
        \nScanOut99[28] , \nScanOut99[27] , \nScanOut99[26] , \nScanOut99[25] , 
        \nScanOut99[24] , \nScanOut99[23] , \nScanOut99[22] , \nScanOut99[21] , 
        \nScanOut99[20] , \nScanOut99[19] , \nScanOut99[18] , \nScanOut99[17] , 
        \nScanOut99[16] , \nScanOut99[15] , \nScanOut99[14] , \nScanOut99[13] , 
        \nScanOut99[12] , \nScanOut99[11] , \nScanOut99[10] , \nScanOut99[9] , 
        \nScanOut99[8] , \nScanOut99[7] , \nScanOut99[6] , \nScanOut99[5] , 
        \nScanOut99[4] , \nScanOut99[3] , \nScanOut99[2] , \nScanOut99[1] , 
        \nScanOut99[0] }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(
        \nEnable[0] ), .BLOCK_VALUE({\nOut1_35[31] , \nOut1_35[30] , 
        \nOut1_35[29] , \nOut1_35[28] , \nOut1_35[27] , \nOut1_35[26] , 
        \nOut1_35[25] , \nOut1_35[24] , \nOut1_35[23] , \nOut1_35[22] , 
        \nOut1_35[21] , \nOut1_35[20] , \nOut1_35[19] , \nOut1_35[18] , 
        \nOut1_35[17] , \nOut1_35[16] , \nOut1_35[15] , \nOut1_35[14] , 
        \nOut1_35[13] , \nOut1_35[12] , \nOut1_35[11] , \nOut1_35[10] , 
        \nOut1_35[9] , \nOut1_35[8] , \nOut1_35[7] , \nOut1_35[6] , 
        \nOut1_35[5] , \nOut1_35[4] , \nOut1_35[3] , \nOut1_35[2] , 
        \nOut1_35[1] , \nOut1_35[0] }), .NORTH_EDGE({\nOut1_34[31] , 
        \nOut1_34[30] , \nOut1_34[29] , \nOut1_34[28] , \nOut1_34[27] , 
        \nOut1_34[26] , \nOut1_34[25] , \nOut1_34[24] , \nOut1_34[23] , 
        \nOut1_34[22] , \nOut1_34[21] , \nOut1_34[20] , \nOut1_34[19] , 
        \nOut1_34[18] , \nOut1_34[17] , \nOut1_34[16] , \nOut1_34[15] , 
        \nOut1_34[14] , \nOut1_34[13] , \nOut1_34[12] , \nOut1_34[11] , 
        \nOut1_34[10] , \nOut1_34[9] , \nOut1_34[8] , \nOut1_34[7] , 
        \nOut1_34[6] , \nOut1_34[5] , \nOut1_34[4] , \nOut1_34[3] , 
        \nOut1_34[2] , \nOut1_34[1] , \nOut1_34[0] }), .SOUTH_EDGE({
        \nOut1_36[31] , \nOut1_36[30] , \nOut1_36[29] , \nOut1_36[28] , 
        \nOut1_36[27] , \nOut1_36[26] , \nOut1_36[25] , \nOut1_36[24] , 
        \nOut1_36[23] , \nOut1_36[22] , \nOut1_36[21] , \nOut1_36[20] , 
        \nOut1_36[19] , \nOut1_36[18] , \nOut1_36[17] , \nOut1_36[16] , 
        \nOut1_36[15] , \nOut1_36[14] , \nOut1_36[13] , \nOut1_36[12] , 
        \nOut1_36[11] , \nOut1_36[10] , \nOut1_36[9] , \nOut1_36[8] , 
        \nOut1_36[7] , \nOut1_36[6] , \nOut1_36[5] , \nOut1_36[4] , 
        \nOut1_36[3] , \nOut1_36[2] , \nOut1_36[1] , \nOut1_36[0] }), 
        .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_35[0] ), .NW_EDGE(\nOut0_34[0] ), 
        .SW_EDGE(\nOut0_36[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_35 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut36[31] , \nScanOut36[30] , \nScanOut36[29] , 
        \nScanOut36[28] , \nScanOut36[27] , \nScanOut36[26] , \nScanOut36[25] , 
        \nScanOut36[24] , \nScanOut36[23] , \nScanOut36[22] , \nScanOut36[21] , 
        \nScanOut36[20] , \nScanOut36[19] , \nScanOut36[18] , \nScanOut36[17] , 
        \nScanOut36[16] , \nScanOut36[15] , \nScanOut36[14] , \nScanOut36[13] , 
        \nScanOut36[12] , \nScanOut36[11] , \nScanOut36[10] , \nScanOut36[9] , 
        \nScanOut36[8] , \nScanOut36[7] , \nScanOut36[6] , \nScanOut36[5] , 
        \nScanOut36[4] , \nScanOut36[3] , \nScanOut36[2] , \nScanOut36[1] , 
        \nScanOut36[0] }), .ScanOut({\nScanOut35[31] , \nScanOut35[30] , 
        \nScanOut35[29] , \nScanOut35[28] , \nScanOut35[27] , \nScanOut35[26] , 
        \nScanOut35[25] , \nScanOut35[24] , \nScanOut35[23] , \nScanOut35[22] , 
        \nScanOut35[21] , \nScanOut35[20] , \nScanOut35[19] , \nScanOut35[18] , 
        \nScanOut35[17] , \nScanOut35[16] , \nScanOut35[15] , \nScanOut35[14] , 
        \nScanOut35[13] , \nScanOut35[12] , \nScanOut35[11] , \nScanOut35[10] , 
        \nScanOut35[9] , \nScanOut35[8] , \nScanOut35[7] , \nScanOut35[6] , 
        \nScanOut35[5] , \nScanOut35[4] , \nScanOut35[3] , \nScanOut35[2] , 
        \nScanOut35[1] , \nScanOut35[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_35[31] , 
        \nOut0_35[30] , \nOut0_35[29] , \nOut0_35[28] , \nOut0_35[27] , 
        \nOut0_35[26] , \nOut0_35[25] , \nOut0_35[24] , \nOut0_35[23] , 
        \nOut0_35[22] , \nOut0_35[21] , \nOut0_35[20] , \nOut0_35[19] , 
        \nOut0_35[18] , \nOut0_35[17] , \nOut0_35[16] , \nOut0_35[15] , 
        \nOut0_35[14] , \nOut0_35[13] , \nOut0_35[12] , \nOut0_35[11] , 
        \nOut0_35[10] , \nOut0_35[9] , \nOut0_35[8] , \nOut0_35[7] , 
        \nOut0_35[6] , \nOut0_35[5] , \nOut0_35[4] , \nOut0_35[3] , 
        \nOut0_35[2] , \nOut0_35[1] , \nOut0_35[0] }), .NORTH_EDGE({
        \nOut0_34[31] , \nOut0_34[30] , \nOut0_34[29] , \nOut0_34[28] , 
        \nOut0_34[27] , \nOut0_34[26] , \nOut0_34[25] , \nOut0_34[24] , 
        \nOut0_34[23] , \nOut0_34[22] , \nOut0_34[21] , \nOut0_34[20] , 
        \nOut0_34[19] , \nOut0_34[18] , \nOut0_34[17] , \nOut0_34[16] , 
        \nOut0_34[15] , \nOut0_34[14] , \nOut0_34[13] , \nOut0_34[12] , 
        \nOut0_34[11] , \nOut0_34[10] , \nOut0_34[9] , \nOut0_34[8] , 
        \nOut0_34[7] , \nOut0_34[6] , \nOut0_34[5] , \nOut0_34[4] , 
        \nOut0_34[3] , \nOut0_34[2] , \nOut0_34[1] , \nOut0_34[0] }), 
        .SOUTH_EDGE({\nOut0_36[31] , \nOut0_36[30] , \nOut0_36[29] , 
        \nOut0_36[28] , \nOut0_36[27] , \nOut0_36[26] , \nOut0_36[25] , 
        \nOut0_36[24] , \nOut0_36[23] , \nOut0_36[22] , \nOut0_36[21] , 
        \nOut0_36[20] , \nOut0_36[19] , \nOut0_36[18] , \nOut0_36[17] , 
        \nOut0_36[16] , \nOut0_36[15] , \nOut0_36[14] , \nOut0_36[13] , 
        \nOut0_36[12] , \nOut0_36[11] , \nOut0_36[10] , \nOut0_36[9] , 
        \nOut0_36[8] , \nOut0_36[7] , \nOut0_36[6] , \nOut0_36[5] , 
        \nOut0_36[4] , \nOut0_36[3] , \nOut0_36[2] , \nOut0_36[1] , 
        \nOut0_36[0] }), .EAST_EDGE(\nOut1_35[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_34[31] ), .SE_EDGE(
        \nOut1_36[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_40 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut41[31] , \nScanOut41[30] , \nScanOut41[29] , 
        \nScanOut41[28] , \nScanOut41[27] , \nScanOut41[26] , \nScanOut41[25] , 
        \nScanOut41[24] , \nScanOut41[23] , \nScanOut41[22] , \nScanOut41[21] , 
        \nScanOut41[20] , \nScanOut41[19] , \nScanOut41[18] , \nScanOut41[17] , 
        \nScanOut41[16] , \nScanOut41[15] , \nScanOut41[14] , \nScanOut41[13] , 
        \nScanOut41[12] , \nScanOut41[11] , \nScanOut41[10] , \nScanOut41[9] , 
        \nScanOut41[8] , \nScanOut41[7] , \nScanOut41[6] , \nScanOut41[5] , 
        \nScanOut41[4] , \nScanOut41[3] , \nScanOut41[2] , \nScanOut41[1] , 
        \nScanOut41[0] }), .ScanOut({\nScanOut40[31] , \nScanOut40[30] , 
        \nScanOut40[29] , \nScanOut40[28] , \nScanOut40[27] , \nScanOut40[26] , 
        \nScanOut40[25] , \nScanOut40[24] , \nScanOut40[23] , \nScanOut40[22] , 
        \nScanOut40[21] , \nScanOut40[20] , \nScanOut40[19] , \nScanOut40[18] , 
        \nScanOut40[17] , \nScanOut40[16] , \nScanOut40[15] , \nScanOut40[14] , 
        \nScanOut40[13] , \nScanOut40[12] , \nScanOut40[11] , \nScanOut40[10] , 
        \nScanOut40[9] , \nScanOut40[8] , \nScanOut40[7] , \nScanOut40[6] , 
        \nScanOut40[5] , \nScanOut40[4] , \nScanOut40[3] , \nScanOut40[2] , 
        \nScanOut40[1] , \nScanOut40[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_40[31] , 
        \nOut0_40[30] , \nOut0_40[29] , \nOut0_40[28] , \nOut0_40[27] , 
        \nOut0_40[26] , \nOut0_40[25] , \nOut0_40[24] , \nOut0_40[23] , 
        \nOut0_40[22] , \nOut0_40[21] , \nOut0_40[20] , \nOut0_40[19] , 
        \nOut0_40[18] , \nOut0_40[17] , \nOut0_40[16] , \nOut0_40[15] , 
        \nOut0_40[14] , \nOut0_40[13] , \nOut0_40[12] , \nOut0_40[11] , 
        \nOut0_40[10] , \nOut0_40[9] , \nOut0_40[8] , \nOut0_40[7] , 
        \nOut0_40[6] , \nOut0_40[5] , \nOut0_40[4] , \nOut0_40[3] , 
        \nOut0_40[2] , \nOut0_40[1] , \nOut0_40[0] }), .NORTH_EDGE({
        \nOut0_39[31] , \nOut0_39[30] , \nOut0_39[29] , \nOut0_39[28] , 
        \nOut0_39[27] , \nOut0_39[26] , \nOut0_39[25] , \nOut0_39[24] , 
        \nOut0_39[23] , \nOut0_39[22] , \nOut0_39[21] , \nOut0_39[20] , 
        \nOut0_39[19] , \nOut0_39[18] , \nOut0_39[17] , \nOut0_39[16] , 
        \nOut0_39[15] , \nOut0_39[14] , \nOut0_39[13] , \nOut0_39[12] , 
        \nOut0_39[11] , \nOut0_39[10] , \nOut0_39[9] , \nOut0_39[8] , 
        \nOut0_39[7] , \nOut0_39[6] , \nOut0_39[5] , \nOut0_39[4] , 
        \nOut0_39[3] , \nOut0_39[2] , \nOut0_39[1] , \nOut0_39[0] }), 
        .SOUTH_EDGE({\nOut0_41[31] , \nOut0_41[30] , \nOut0_41[29] , 
        \nOut0_41[28] , \nOut0_41[27] , \nOut0_41[26] , \nOut0_41[25] , 
        \nOut0_41[24] , \nOut0_41[23] , \nOut0_41[22] , \nOut0_41[21] , 
        \nOut0_41[20] , \nOut0_41[19] , \nOut0_41[18] , \nOut0_41[17] , 
        \nOut0_41[16] , \nOut0_41[15] , \nOut0_41[14] , \nOut0_41[13] , 
        \nOut0_41[12] , \nOut0_41[11] , \nOut0_41[10] , \nOut0_41[9] , 
        \nOut0_41[8] , \nOut0_41[7] , \nOut0_41[6] , \nOut0_41[5] , 
        \nOut0_41[4] , \nOut0_41[3] , \nOut0_41[2] , \nOut0_41[1] , 
        \nOut0_41[0] }), .EAST_EDGE(\nOut1_40[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_39[31] ), .SE_EDGE(
        \nOut1_41[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_67 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut68[31] , \nScanOut68[30] , \nScanOut68[29] , 
        \nScanOut68[28] , \nScanOut68[27] , \nScanOut68[26] , \nScanOut68[25] , 
        \nScanOut68[24] , \nScanOut68[23] , \nScanOut68[22] , \nScanOut68[21] , 
        \nScanOut68[20] , \nScanOut68[19] , \nScanOut68[18] , \nScanOut68[17] , 
        \nScanOut68[16] , \nScanOut68[15] , \nScanOut68[14] , \nScanOut68[13] , 
        \nScanOut68[12] , \nScanOut68[11] , \nScanOut68[10] , \nScanOut68[9] , 
        \nScanOut68[8] , \nScanOut68[7] , \nScanOut68[6] , \nScanOut68[5] , 
        \nScanOut68[4] , \nScanOut68[3] , \nScanOut68[2] , \nScanOut68[1] , 
        \nScanOut68[0] }), .ScanOut({\nScanOut67[31] , \nScanOut67[30] , 
        \nScanOut67[29] , \nScanOut67[28] , \nScanOut67[27] , \nScanOut67[26] , 
        \nScanOut67[25] , \nScanOut67[24] , \nScanOut67[23] , \nScanOut67[22] , 
        \nScanOut67[21] , \nScanOut67[20] , \nScanOut67[19] , \nScanOut67[18] , 
        \nScanOut67[17] , \nScanOut67[16] , \nScanOut67[15] , \nScanOut67[14] , 
        \nScanOut67[13] , \nScanOut67[12] , \nScanOut67[11] , \nScanOut67[10] , 
        \nScanOut67[9] , \nScanOut67[8] , \nScanOut67[7] , \nScanOut67[6] , 
        \nScanOut67[5] , \nScanOut67[4] , \nScanOut67[3] , \nScanOut67[2] , 
        \nScanOut67[1] , \nScanOut67[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_3[31] , 
        \nOut1_3[30] , \nOut1_3[29] , \nOut1_3[28] , \nOut1_3[27] , 
        \nOut1_3[26] , \nOut1_3[25] , \nOut1_3[24] , \nOut1_3[23] , 
        \nOut1_3[22] , \nOut1_3[21] , \nOut1_3[20] , \nOut1_3[19] , 
        \nOut1_3[18] , \nOut1_3[17] , \nOut1_3[16] , \nOut1_3[15] , 
        \nOut1_3[14] , \nOut1_3[13] , \nOut1_3[12] , \nOut1_3[11] , 
        \nOut1_3[10] , \nOut1_3[9] , \nOut1_3[8] , \nOut1_3[7] , \nOut1_3[6] , 
        \nOut1_3[5] , \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , 
        \nOut1_3[0] }), .NORTH_EDGE({\nOut1_2[31] , \nOut1_2[30] , 
        \nOut1_2[29] , \nOut1_2[28] , \nOut1_2[27] , \nOut1_2[26] , 
        \nOut1_2[25] , \nOut1_2[24] , \nOut1_2[23] , \nOut1_2[22] , 
        \nOut1_2[21] , \nOut1_2[20] , \nOut1_2[19] , \nOut1_2[18] , 
        \nOut1_2[17] , \nOut1_2[16] , \nOut1_2[15] , \nOut1_2[14] , 
        \nOut1_2[13] , \nOut1_2[12] , \nOut1_2[11] , \nOut1_2[10] , 
        \nOut1_2[9] , \nOut1_2[8] , \nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , 
        \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), 
        .SOUTH_EDGE({\nOut1_4[31] , \nOut1_4[30] , \nOut1_4[29] , 
        \nOut1_4[28] , \nOut1_4[27] , \nOut1_4[26] , \nOut1_4[25] , 
        \nOut1_4[24] , \nOut1_4[23] , \nOut1_4[22] , \nOut1_4[21] , 
        \nOut1_4[20] , \nOut1_4[19] , \nOut1_4[18] , \nOut1_4[17] , 
        \nOut1_4[16] , \nOut1_4[15] , \nOut1_4[14] , \nOut1_4[13] , 
        \nOut1_4[12] , \nOut1_4[11] , \nOut1_4[10] , \nOut1_4[9] , 
        \nOut1_4[8] , \nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , \nOut1_4[4] , 
        \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_3[0] ), .NW_EDGE(\nOut0_2[0] ), .SW_EDGE(
        \nOut0_4[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_116 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut117[31] , \nScanOut117[30] , \nScanOut117[29] , 
        \nScanOut117[28] , \nScanOut117[27] , \nScanOut117[26] , 
        \nScanOut117[25] , \nScanOut117[24] , \nScanOut117[23] , 
        \nScanOut117[22] , \nScanOut117[21] , \nScanOut117[20] , 
        \nScanOut117[19] , \nScanOut117[18] , \nScanOut117[17] , 
        \nScanOut117[16] , \nScanOut117[15] , \nScanOut117[14] , 
        \nScanOut117[13] , \nScanOut117[12] , \nScanOut117[11] , 
        \nScanOut117[10] , \nScanOut117[9] , \nScanOut117[8] , 
        \nScanOut117[7] , \nScanOut117[6] , \nScanOut117[5] , \nScanOut117[4] , 
        \nScanOut117[3] , \nScanOut117[2] , \nScanOut117[1] , \nScanOut117[0] 
        }), .ScanOut({\nScanOut116[31] , \nScanOut116[30] , \nScanOut116[29] , 
        \nScanOut116[28] , \nScanOut116[27] , \nScanOut116[26] , 
        \nScanOut116[25] , \nScanOut116[24] , \nScanOut116[23] , 
        \nScanOut116[22] , \nScanOut116[21] , \nScanOut116[20] , 
        \nScanOut116[19] , \nScanOut116[18] , \nScanOut116[17] , 
        \nScanOut116[16] , \nScanOut116[15] , \nScanOut116[14] , 
        \nScanOut116[13] , \nScanOut116[12] , \nScanOut116[11] , 
        \nScanOut116[10] , \nScanOut116[9] , \nScanOut116[8] , 
        \nScanOut116[7] , \nScanOut116[6] , \nScanOut116[5] , \nScanOut116[4] , 
        \nScanOut116[3] , \nScanOut116[2] , \nScanOut116[1] , \nScanOut116[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_52[31] , \nOut1_52[30] , \nOut1_52[29] , 
        \nOut1_52[28] , \nOut1_52[27] , \nOut1_52[26] , \nOut1_52[25] , 
        \nOut1_52[24] , \nOut1_52[23] , \nOut1_52[22] , \nOut1_52[21] , 
        \nOut1_52[20] , \nOut1_52[19] , \nOut1_52[18] , \nOut1_52[17] , 
        \nOut1_52[16] , \nOut1_52[15] , \nOut1_52[14] , \nOut1_52[13] , 
        \nOut1_52[12] , \nOut1_52[11] , \nOut1_52[10] , \nOut1_52[9] , 
        \nOut1_52[8] , \nOut1_52[7] , \nOut1_52[6] , \nOut1_52[5] , 
        \nOut1_52[4] , \nOut1_52[3] , \nOut1_52[2] , \nOut1_52[1] , 
        \nOut1_52[0] }), .NORTH_EDGE({\nOut1_51[31] , \nOut1_51[30] , 
        \nOut1_51[29] , \nOut1_51[28] , \nOut1_51[27] , \nOut1_51[26] , 
        \nOut1_51[25] , \nOut1_51[24] , \nOut1_51[23] , \nOut1_51[22] , 
        \nOut1_51[21] , \nOut1_51[20] , \nOut1_51[19] , \nOut1_51[18] , 
        \nOut1_51[17] , \nOut1_51[16] , \nOut1_51[15] , \nOut1_51[14] , 
        \nOut1_51[13] , \nOut1_51[12] , \nOut1_51[11] , \nOut1_51[10] , 
        \nOut1_51[9] , \nOut1_51[8] , \nOut1_51[7] , \nOut1_51[6] , 
        \nOut1_51[5] , \nOut1_51[4] , \nOut1_51[3] , \nOut1_51[2] , 
        \nOut1_51[1] , \nOut1_51[0] }), .SOUTH_EDGE({\nOut1_53[31] , 
        \nOut1_53[30] , \nOut1_53[29] , \nOut1_53[28] , \nOut1_53[27] , 
        \nOut1_53[26] , \nOut1_53[25] , \nOut1_53[24] , \nOut1_53[23] , 
        \nOut1_53[22] , \nOut1_53[21] , \nOut1_53[20] , \nOut1_53[19] , 
        \nOut1_53[18] , \nOut1_53[17] , \nOut1_53[16] , \nOut1_53[15] , 
        \nOut1_53[14] , \nOut1_53[13] , \nOut1_53[12] , \nOut1_53[11] , 
        \nOut1_53[10] , \nOut1_53[9] , \nOut1_53[8] , \nOut1_53[7] , 
        \nOut1_53[6] , \nOut1_53[5] , \nOut1_53[4] , \nOut1_53[3] , 
        \nOut1_53[2] , \nOut1_53[1] , \nOut1_53[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_52[0] ), .NW_EDGE(\nOut0_51[0] ), .SW_EDGE(
        \nOut0_53[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_52 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut53[31] , \nScanOut53[30] , \nScanOut53[29] , 
        \nScanOut53[28] , \nScanOut53[27] , \nScanOut53[26] , \nScanOut53[25] , 
        \nScanOut53[24] , \nScanOut53[23] , \nScanOut53[22] , \nScanOut53[21] , 
        \nScanOut53[20] , \nScanOut53[19] , \nScanOut53[18] , \nScanOut53[17] , 
        \nScanOut53[16] , \nScanOut53[15] , \nScanOut53[14] , \nScanOut53[13] , 
        \nScanOut53[12] , \nScanOut53[11] , \nScanOut53[10] , \nScanOut53[9] , 
        \nScanOut53[8] , \nScanOut53[7] , \nScanOut53[6] , \nScanOut53[5] , 
        \nScanOut53[4] , \nScanOut53[3] , \nScanOut53[2] , \nScanOut53[1] , 
        \nScanOut53[0] }), .ScanOut({\nScanOut52[31] , \nScanOut52[30] , 
        \nScanOut52[29] , \nScanOut52[28] , \nScanOut52[27] , \nScanOut52[26] , 
        \nScanOut52[25] , \nScanOut52[24] , \nScanOut52[23] , \nScanOut52[22] , 
        \nScanOut52[21] , \nScanOut52[20] , \nScanOut52[19] , \nScanOut52[18] , 
        \nScanOut52[17] , \nScanOut52[16] , \nScanOut52[15] , \nScanOut52[14] , 
        \nScanOut52[13] , \nScanOut52[12] , \nScanOut52[11] , \nScanOut52[10] , 
        \nScanOut52[9] , \nScanOut52[8] , \nScanOut52[7] , \nScanOut52[6] , 
        \nScanOut52[5] , \nScanOut52[4] , \nScanOut52[3] , \nScanOut52[2] , 
        \nScanOut52[1] , \nScanOut52[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_52[31] , 
        \nOut0_52[30] , \nOut0_52[29] , \nOut0_52[28] , \nOut0_52[27] , 
        \nOut0_52[26] , \nOut0_52[25] , \nOut0_52[24] , \nOut0_52[23] , 
        \nOut0_52[22] , \nOut0_52[21] , \nOut0_52[20] , \nOut0_52[19] , 
        \nOut0_52[18] , \nOut0_52[17] , \nOut0_52[16] , \nOut0_52[15] , 
        \nOut0_52[14] , \nOut0_52[13] , \nOut0_52[12] , \nOut0_52[11] , 
        \nOut0_52[10] , \nOut0_52[9] , \nOut0_52[8] , \nOut0_52[7] , 
        \nOut0_52[6] , \nOut0_52[5] , \nOut0_52[4] , \nOut0_52[3] , 
        \nOut0_52[2] , \nOut0_52[1] , \nOut0_52[0] }), .NORTH_EDGE({
        \nOut0_51[31] , \nOut0_51[30] , \nOut0_51[29] , \nOut0_51[28] , 
        \nOut0_51[27] , \nOut0_51[26] , \nOut0_51[25] , \nOut0_51[24] , 
        \nOut0_51[23] , \nOut0_51[22] , \nOut0_51[21] , \nOut0_51[20] , 
        \nOut0_51[19] , \nOut0_51[18] , \nOut0_51[17] , \nOut0_51[16] , 
        \nOut0_51[15] , \nOut0_51[14] , \nOut0_51[13] , \nOut0_51[12] , 
        \nOut0_51[11] , \nOut0_51[10] , \nOut0_51[9] , \nOut0_51[8] , 
        \nOut0_51[7] , \nOut0_51[6] , \nOut0_51[5] , \nOut0_51[4] , 
        \nOut0_51[3] , \nOut0_51[2] , \nOut0_51[1] , \nOut0_51[0] }), 
        .SOUTH_EDGE({\nOut0_53[31] , \nOut0_53[30] , \nOut0_53[29] , 
        \nOut0_53[28] , \nOut0_53[27] , \nOut0_53[26] , \nOut0_53[25] , 
        \nOut0_53[24] , \nOut0_53[23] , \nOut0_53[22] , \nOut0_53[21] , 
        \nOut0_53[20] , \nOut0_53[19] , \nOut0_53[18] , \nOut0_53[17] , 
        \nOut0_53[16] , \nOut0_53[15] , \nOut0_53[14] , \nOut0_53[13] , 
        \nOut0_53[12] , \nOut0_53[11] , \nOut0_53[10] , \nOut0_53[9] , 
        \nOut0_53[8] , \nOut0_53[7] , \nOut0_53[6] , \nOut0_53[5] , 
        \nOut0_53[4] , \nOut0_53[3] , \nOut0_53[2] , \nOut0_53[1] , 
        \nOut0_53[0] }), .EAST_EDGE(\nOut1_52[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_51[31] ), .SE_EDGE(
        \nOut1_53[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_75 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut76[31] , \nScanOut76[30] , \nScanOut76[29] , 
        \nScanOut76[28] , \nScanOut76[27] , \nScanOut76[26] , \nScanOut76[25] , 
        \nScanOut76[24] , \nScanOut76[23] , \nScanOut76[22] , \nScanOut76[21] , 
        \nScanOut76[20] , \nScanOut76[19] , \nScanOut76[18] , \nScanOut76[17] , 
        \nScanOut76[16] , \nScanOut76[15] , \nScanOut76[14] , \nScanOut76[13] , 
        \nScanOut76[12] , \nScanOut76[11] , \nScanOut76[10] , \nScanOut76[9] , 
        \nScanOut76[8] , \nScanOut76[7] , \nScanOut76[6] , \nScanOut76[5] , 
        \nScanOut76[4] , \nScanOut76[3] , \nScanOut76[2] , \nScanOut76[1] , 
        \nScanOut76[0] }), .ScanOut({\nScanOut75[31] , \nScanOut75[30] , 
        \nScanOut75[29] , \nScanOut75[28] , \nScanOut75[27] , \nScanOut75[26] , 
        \nScanOut75[25] , \nScanOut75[24] , \nScanOut75[23] , \nScanOut75[22] , 
        \nScanOut75[21] , \nScanOut75[20] , \nScanOut75[19] , \nScanOut75[18] , 
        \nScanOut75[17] , \nScanOut75[16] , \nScanOut75[15] , \nScanOut75[14] , 
        \nScanOut75[13] , \nScanOut75[12] , \nScanOut75[11] , \nScanOut75[10] , 
        \nScanOut75[9] , \nScanOut75[8] , \nScanOut75[7] , \nScanOut75[6] , 
        \nScanOut75[5] , \nScanOut75[4] , \nScanOut75[3] , \nScanOut75[2] , 
        \nScanOut75[1] , \nScanOut75[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_11[31] , 
        \nOut1_11[30] , \nOut1_11[29] , \nOut1_11[28] , \nOut1_11[27] , 
        \nOut1_11[26] , \nOut1_11[25] , \nOut1_11[24] , \nOut1_11[23] , 
        \nOut1_11[22] , \nOut1_11[21] , \nOut1_11[20] , \nOut1_11[19] , 
        \nOut1_11[18] , \nOut1_11[17] , \nOut1_11[16] , \nOut1_11[15] , 
        \nOut1_11[14] , \nOut1_11[13] , \nOut1_11[12] , \nOut1_11[11] , 
        \nOut1_11[10] , \nOut1_11[9] , \nOut1_11[8] , \nOut1_11[7] , 
        \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , \nOut1_11[3] , 
        \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), .NORTH_EDGE({
        \nOut1_10[31] , \nOut1_10[30] , \nOut1_10[29] , \nOut1_10[28] , 
        \nOut1_10[27] , \nOut1_10[26] , \nOut1_10[25] , \nOut1_10[24] , 
        \nOut1_10[23] , \nOut1_10[22] , \nOut1_10[21] , \nOut1_10[20] , 
        \nOut1_10[19] , \nOut1_10[18] , \nOut1_10[17] , \nOut1_10[16] , 
        \nOut1_10[15] , \nOut1_10[14] , \nOut1_10[13] , \nOut1_10[12] , 
        \nOut1_10[11] , \nOut1_10[10] , \nOut1_10[9] , \nOut1_10[8] , 
        \nOut1_10[7] , \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , 
        \nOut1_10[3] , \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), 
        .SOUTH_EDGE({\nOut1_12[31] , \nOut1_12[30] , \nOut1_12[29] , 
        \nOut1_12[28] , \nOut1_12[27] , \nOut1_12[26] , \nOut1_12[25] , 
        \nOut1_12[24] , \nOut1_12[23] , \nOut1_12[22] , \nOut1_12[21] , 
        \nOut1_12[20] , \nOut1_12[19] , \nOut1_12[18] , \nOut1_12[17] , 
        \nOut1_12[16] , \nOut1_12[15] , \nOut1_12[14] , \nOut1_12[13] , 
        \nOut1_12[12] , \nOut1_12[11] , \nOut1_12[10] , \nOut1_12[9] , 
        \nOut1_12[8] , \nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , 
        \nOut1_12[4] , \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , 
        \nOut1_12[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_11[0] ), 
        .NW_EDGE(\nOut0_10[0] ), .SW_EDGE(\nOut0_12[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_82 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut83[31] , \nScanOut83[30] , \nScanOut83[29] , 
        \nScanOut83[28] , \nScanOut83[27] , \nScanOut83[26] , \nScanOut83[25] , 
        \nScanOut83[24] , \nScanOut83[23] , \nScanOut83[22] , \nScanOut83[21] , 
        \nScanOut83[20] , \nScanOut83[19] , \nScanOut83[18] , \nScanOut83[17] , 
        \nScanOut83[16] , \nScanOut83[15] , \nScanOut83[14] , \nScanOut83[13] , 
        \nScanOut83[12] , \nScanOut83[11] , \nScanOut83[10] , \nScanOut83[9] , 
        \nScanOut83[8] , \nScanOut83[7] , \nScanOut83[6] , \nScanOut83[5] , 
        \nScanOut83[4] , \nScanOut83[3] , \nScanOut83[2] , \nScanOut83[1] , 
        \nScanOut83[0] }), .ScanOut({\nScanOut82[31] , \nScanOut82[30] , 
        \nScanOut82[29] , \nScanOut82[28] , \nScanOut82[27] , \nScanOut82[26] , 
        \nScanOut82[25] , \nScanOut82[24] , \nScanOut82[23] , \nScanOut82[22] , 
        \nScanOut82[21] , \nScanOut82[20] , \nScanOut82[19] , \nScanOut82[18] , 
        \nScanOut82[17] , \nScanOut82[16] , \nScanOut82[15] , \nScanOut82[14] , 
        \nScanOut82[13] , \nScanOut82[12] , \nScanOut82[11] , \nScanOut82[10] , 
        \nScanOut82[9] , \nScanOut82[8] , \nScanOut82[7] , \nScanOut82[6] , 
        \nScanOut82[5] , \nScanOut82[4] , \nScanOut82[3] , \nScanOut82[2] , 
        \nScanOut82[1] , \nScanOut82[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_18[31] , 
        \nOut1_18[30] , \nOut1_18[29] , \nOut1_18[28] , \nOut1_18[27] , 
        \nOut1_18[26] , \nOut1_18[25] , \nOut1_18[24] , \nOut1_18[23] , 
        \nOut1_18[22] , \nOut1_18[21] , \nOut1_18[20] , \nOut1_18[19] , 
        \nOut1_18[18] , \nOut1_18[17] , \nOut1_18[16] , \nOut1_18[15] , 
        \nOut1_18[14] , \nOut1_18[13] , \nOut1_18[12] , \nOut1_18[11] , 
        \nOut1_18[10] , \nOut1_18[9] , \nOut1_18[8] , \nOut1_18[7] , 
        \nOut1_18[6] , \nOut1_18[5] , \nOut1_18[4] , \nOut1_18[3] , 
        \nOut1_18[2] , \nOut1_18[1] , \nOut1_18[0] }), .NORTH_EDGE({
        \nOut1_17[31] , \nOut1_17[30] , \nOut1_17[29] , \nOut1_17[28] , 
        \nOut1_17[27] , \nOut1_17[26] , \nOut1_17[25] , \nOut1_17[24] , 
        \nOut1_17[23] , \nOut1_17[22] , \nOut1_17[21] , \nOut1_17[20] , 
        \nOut1_17[19] , \nOut1_17[18] , \nOut1_17[17] , \nOut1_17[16] , 
        \nOut1_17[15] , \nOut1_17[14] , \nOut1_17[13] , \nOut1_17[12] , 
        \nOut1_17[11] , \nOut1_17[10] , \nOut1_17[9] , \nOut1_17[8] , 
        \nOut1_17[7] , \nOut1_17[6] , \nOut1_17[5] , \nOut1_17[4] , 
        \nOut1_17[3] , \nOut1_17[2] , \nOut1_17[1] , \nOut1_17[0] }), 
        .SOUTH_EDGE({\nOut1_19[31] , \nOut1_19[30] , \nOut1_19[29] , 
        \nOut1_19[28] , \nOut1_19[27] , \nOut1_19[26] , \nOut1_19[25] , 
        \nOut1_19[24] , \nOut1_19[23] , \nOut1_19[22] , \nOut1_19[21] , 
        \nOut1_19[20] , \nOut1_19[19] , \nOut1_19[18] , \nOut1_19[17] , 
        \nOut1_19[16] , \nOut1_19[15] , \nOut1_19[14] , \nOut1_19[13] , 
        \nOut1_19[12] , \nOut1_19[11] , \nOut1_19[10] , \nOut1_19[9] , 
        \nOut1_19[8] , \nOut1_19[7] , \nOut1_19[6] , \nOut1_19[5] , 
        \nOut1_19[4] , \nOut1_19[3] , \nOut1_19[2] , \nOut1_19[1] , 
        \nOut1_19[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_18[0] ), 
        .NW_EDGE(\nOut0_17[0] ), .SW_EDGE(\nOut0_19[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_90 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut91[31] , \nScanOut91[30] , \nScanOut91[29] , 
        \nScanOut91[28] , \nScanOut91[27] , \nScanOut91[26] , \nScanOut91[25] , 
        \nScanOut91[24] , \nScanOut91[23] , \nScanOut91[22] , \nScanOut91[21] , 
        \nScanOut91[20] , \nScanOut91[19] , \nScanOut91[18] , \nScanOut91[17] , 
        \nScanOut91[16] , \nScanOut91[15] , \nScanOut91[14] , \nScanOut91[13] , 
        \nScanOut91[12] , \nScanOut91[11] , \nScanOut91[10] , \nScanOut91[9] , 
        \nScanOut91[8] , \nScanOut91[7] , \nScanOut91[6] , \nScanOut91[5] , 
        \nScanOut91[4] , \nScanOut91[3] , \nScanOut91[2] , \nScanOut91[1] , 
        \nScanOut91[0] }), .ScanOut({\nScanOut90[31] , \nScanOut90[30] , 
        \nScanOut90[29] , \nScanOut90[28] , \nScanOut90[27] , \nScanOut90[26] , 
        \nScanOut90[25] , \nScanOut90[24] , \nScanOut90[23] , \nScanOut90[22] , 
        \nScanOut90[21] , \nScanOut90[20] , \nScanOut90[19] , \nScanOut90[18] , 
        \nScanOut90[17] , \nScanOut90[16] , \nScanOut90[15] , \nScanOut90[14] , 
        \nScanOut90[13] , \nScanOut90[12] , \nScanOut90[11] , \nScanOut90[10] , 
        \nScanOut90[9] , \nScanOut90[8] , \nScanOut90[7] , \nScanOut90[6] , 
        \nScanOut90[5] , \nScanOut90[4] , \nScanOut90[3] , \nScanOut90[2] , 
        \nScanOut90[1] , \nScanOut90[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_26[31] , 
        \nOut1_26[30] , \nOut1_26[29] , \nOut1_26[28] , \nOut1_26[27] , 
        \nOut1_26[26] , \nOut1_26[25] , \nOut1_26[24] , \nOut1_26[23] , 
        \nOut1_26[22] , \nOut1_26[21] , \nOut1_26[20] , \nOut1_26[19] , 
        \nOut1_26[18] , \nOut1_26[17] , \nOut1_26[16] , \nOut1_26[15] , 
        \nOut1_26[14] , \nOut1_26[13] , \nOut1_26[12] , \nOut1_26[11] , 
        \nOut1_26[10] , \nOut1_26[9] , \nOut1_26[8] , \nOut1_26[7] , 
        \nOut1_26[6] , \nOut1_26[5] , \nOut1_26[4] , \nOut1_26[3] , 
        \nOut1_26[2] , \nOut1_26[1] , \nOut1_26[0] }), .NORTH_EDGE({
        \nOut1_25[31] , \nOut1_25[30] , \nOut1_25[29] , \nOut1_25[28] , 
        \nOut1_25[27] , \nOut1_25[26] , \nOut1_25[25] , \nOut1_25[24] , 
        \nOut1_25[23] , \nOut1_25[22] , \nOut1_25[21] , \nOut1_25[20] , 
        \nOut1_25[19] , \nOut1_25[18] , \nOut1_25[17] , \nOut1_25[16] , 
        \nOut1_25[15] , \nOut1_25[14] , \nOut1_25[13] , \nOut1_25[12] , 
        \nOut1_25[11] , \nOut1_25[10] , \nOut1_25[9] , \nOut1_25[8] , 
        \nOut1_25[7] , \nOut1_25[6] , \nOut1_25[5] , \nOut1_25[4] , 
        \nOut1_25[3] , \nOut1_25[2] , \nOut1_25[1] , \nOut1_25[0] }), 
        .SOUTH_EDGE({\nOut1_27[31] , \nOut1_27[30] , \nOut1_27[29] , 
        \nOut1_27[28] , \nOut1_27[27] , \nOut1_27[26] , \nOut1_27[25] , 
        \nOut1_27[24] , \nOut1_27[23] , \nOut1_27[22] , \nOut1_27[21] , 
        \nOut1_27[20] , \nOut1_27[19] , \nOut1_27[18] , \nOut1_27[17] , 
        \nOut1_27[16] , \nOut1_27[15] , \nOut1_27[14] , \nOut1_27[13] , 
        \nOut1_27[12] , \nOut1_27[11] , \nOut1_27[10] , \nOut1_27[9] , 
        \nOut1_27[8] , \nOut1_27[7] , \nOut1_27[6] , \nOut1_27[5] , 
        \nOut1_27[4] , \nOut1_27[3] , \nOut1_27[2] , \nOut1_27[1] , 
        \nOut1_27[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_26[0] ), 
        .NW_EDGE(\nOut0_25[0] ), .SW_EDGE(\nOut0_27[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_104 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut105[31] , \nScanOut105[30] , \nScanOut105[29] , 
        \nScanOut105[28] , \nScanOut105[27] , \nScanOut105[26] , 
        \nScanOut105[25] , \nScanOut105[24] , \nScanOut105[23] , 
        \nScanOut105[22] , \nScanOut105[21] , \nScanOut105[20] , 
        \nScanOut105[19] , \nScanOut105[18] , \nScanOut105[17] , 
        \nScanOut105[16] , \nScanOut105[15] , \nScanOut105[14] , 
        \nScanOut105[13] , \nScanOut105[12] , \nScanOut105[11] , 
        \nScanOut105[10] , \nScanOut105[9] , \nScanOut105[8] , 
        \nScanOut105[7] , \nScanOut105[6] , \nScanOut105[5] , \nScanOut105[4] , 
        \nScanOut105[3] , \nScanOut105[2] , \nScanOut105[1] , \nScanOut105[0] 
        }), .ScanOut({\nScanOut104[31] , \nScanOut104[30] , \nScanOut104[29] , 
        \nScanOut104[28] , \nScanOut104[27] , \nScanOut104[26] , 
        \nScanOut104[25] , \nScanOut104[24] , \nScanOut104[23] , 
        \nScanOut104[22] , \nScanOut104[21] , \nScanOut104[20] , 
        \nScanOut104[19] , \nScanOut104[18] , \nScanOut104[17] , 
        \nScanOut104[16] , \nScanOut104[15] , \nScanOut104[14] , 
        \nScanOut104[13] , \nScanOut104[12] , \nScanOut104[11] , 
        \nScanOut104[10] , \nScanOut104[9] , \nScanOut104[8] , 
        \nScanOut104[7] , \nScanOut104[6] , \nScanOut104[5] , \nScanOut104[4] , 
        \nScanOut104[3] , \nScanOut104[2] , \nScanOut104[1] , \nScanOut104[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_40[31] , \nOut1_40[30] , \nOut1_40[29] , 
        \nOut1_40[28] , \nOut1_40[27] , \nOut1_40[26] , \nOut1_40[25] , 
        \nOut1_40[24] , \nOut1_40[23] , \nOut1_40[22] , \nOut1_40[21] , 
        \nOut1_40[20] , \nOut1_40[19] , \nOut1_40[18] , \nOut1_40[17] , 
        \nOut1_40[16] , \nOut1_40[15] , \nOut1_40[14] , \nOut1_40[13] , 
        \nOut1_40[12] , \nOut1_40[11] , \nOut1_40[10] , \nOut1_40[9] , 
        \nOut1_40[8] , \nOut1_40[7] , \nOut1_40[6] , \nOut1_40[5] , 
        \nOut1_40[4] , \nOut1_40[3] , \nOut1_40[2] , \nOut1_40[1] , 
        \nOut1_40[0] }), .NORTH_EDGE({\nOut1_39[31] , \nOut1_39[30] , 
        \nOut1_39[29] , \nOut1_39[28] , \nOut1_39[27] , \nOut1_39[26] , 
        \nOut1_39[25] , \nOut1_39[24] , \nOut1_39[23] , \nOut1_39[22] , 
        \nOut1_39[21] , \nOut1_39[20] , \nOut1_39[19] , \nOut1_39[18] , 
        \nOut1_39[17] , \nOut1_39[16] , \nOut1_39[15] , \nOut1_39[14] , 
        \nOut1_39[13] , \nOut1_39[12] , \nOut1_39[11] , \nOut1_39[10] , 
        \nOut1_39[9] , \nOut1_39[8] , \nOut1_39[7] , \nOut1_39[6] , 
        \nOut1_39[5] , \nOut1_39[4] , \nOut1_39[3] , \nOut1_39[2] , 
        \nOut1_39[1] , \nOut1_39[0] }), .SOUTH_EDGE({\nOut1_41[31] , 
        \nOut1_41[30] , \nOut1_41[29] , \nOut1_41[28] , \nOut1_41[27] , 
        \nOut1_41[26] , \nOut1_41[25] , \nOut1_41[24] , \nOut1_41[23] , 
        \nOut1_41[22] , \nOut1_41[21] , \nOut1_41[20] , \nOut1_41[19] , 
        \nOut1_41[18] , \nOut1_41[17] , \nOut1_41[16] , \nOut1_41[15] , 
        \nOut1_41[14] , \nOut1_41[13] , \nOut1_41[12] , \nOut1_41[11] , 
        \nOut1_41[10] , \nOut1_41[9] , \nOut1_41[8] , \nOut1_41[7] , 
        \nOut1_41[6] , \nOut1_41[5] , \nOut1_41[4] , \nOut1_41[3] , 
        \nOut1_41[2] , \nOut1_41[1] , \nOut1_41[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_40[0] ), .NW_EDGE(\nOut0_39[0] ), .SW_EDGE(
        \nOut0_41[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_123 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut124[31] , \nScanOut124[30] , \nScanOut124[29] , 
        \nScanOut124[28] , \nScanOut124[27] , \nScanOut124[26] , 
        \nScanOut124[25] , \nScanOut124[24] , \nScanOut124[23] , 
        \nScanOut124[22] , \nScanOut124[21] , \nScanOut124[20] , 
        \nScanOut124[19] , \nScanOut124[18] , \nScanOut124[17] , 
        \nScanOut124[16] , \nScanOut124[15] , \nScanOut124[14] , 
        \nScanOut124[13] , \nScanOut124[12] , \nScanOut124[11] , 
        \nScanOut124[10] , \nScanOut124[9] , \nScanOut124[8] , 
        \nScanOut124[7] , \nScanOut124[6] , \nScanOut124[5] , \nScanOut124[4] , 
        \nScanOut124[3] , \nScanOut124[2] , \nScanOut124[1] , \nScanOut124[0] 
        }), .ScanOut({\nScanOut123[31] , \nScanOut123[30] , \nScanOut123[29] , 
        \nScanOut123[28] , \nScanOut123[27] , \nScanOut123[26] , 
        \nScanOut123[25] , \nScanOut123[24] , \nScanOut123[23] , 
        \nScanOut123[22] , \nScanOut123[21] , \nScanOut123[20] , 
        \nScanOut123[19] , \nScanOut123[18] , \nScanOut123[17] , 
        \nScanOut123[16] , \nScanOut123[15] , \nScanOut123[14] , 
        \nScanOut123[13] , \nScanOut123[12] , \nScanOut123[11] , 
        \nScanOut123[10] , \nScanOut123[9] , \nScanOut123[8] , 
        \nScanOut123[7] , \nScanOut123[6] , \nScanOut123[5] , \nScanOut123[4] , 
        \nScanOut123[3] , \nScanOut123[2] , \nScanOut123[1] , \nScanOut123[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_59[31] , \nOut1_59[30] , \nOut1_59[29] , 
        \nOut1_59[28] , \nOut1_59[27] , \nOut1_59[26] , \nOut1_59[25] , 
        \nOut1_59[24] , \nOut1_59[23] , \nOut1_59[22] , \nOut1_59[21] , 
        \nOut1_59[20] , \nOut1_59[19] , \nOut1_59[18] , \nOut1_59[17] , 
        \nOut1_59[16] , \nOut1_59[15] , \nOut1_59[14] , \nOut1_59[13] , 
        \nOut1_59[12] , \nOut1_59[11] , \nOut1_59[10] , \nOut1_59[9] , 
        \nOut1_59[8] , \nOut1_59[7] , \nOut1_59[6] , \nOut1_59[5] , 
        \nOut1_59[4] , \nOut1_59[3] , \nOut1_59[2] , \nOut1_59[1] , 
        \nOut1_59[0] }), .NORTH_EDGE({\nOut1_58[31] , \nOut1_58[30] , 
        \nOut1_58[29] , \nOut1_58[28] , \nOut1_58[27] , \nOut1_58[26] , 
        \nOut1_58[25] , \nOut1_58[24] , \nOut1_58[23] , \nOut1_58[22] , 
        \nOut1_58[21] , \nOut1_58[20] , \nOut1_58[19] , \nOut1_58[18] , 
        \nOut1_58[17] , \nOut1_58[16] , \nOut1_58[15] , \nOut1_58[14] , 
        \nOut1_58[13] , \nOut1_58[12] , \nOut1_58[11] , \nOut1_58[10] , 
        \nOut1_58[9] , \nOut1_58[8] , \nOut1_58[7] , \nOut1_58[6] , 
        \nOut1_58[5] , \nOut1_58[4] , \nOut1_58[3] , \nOut1_58[2] , 
        \nOut1_58[1] , \nOut1_58[0] }), .SOUTH_EDGE({\nOut1_60[31] , 
        \nOut1_60[30] , \nOut1_60[29] , \nOut1_60[28] , \nOut1_60[27] , 
        \nOut1_60[26] , \nOut1_60[25] , \nOut1_60[24] , \nOut1_60[23] , 
        \nOut1_60[22] , \nOut1_60[21] , \nOut1_60[20] , \nOut1_60[19] , 
        \nOut1_60[18] , \nOut1_60[17] , \nOut1_60[16] , \nOut1_60[15] , 
        \nOut1_60[14] , \nOut1_60[13] , \nOut1_60[12] , \nOut1_60[11] , 
        \nOut1_60[10] , \nOut1_60[9] , \nOut1_60[8] , \nOut1_60[7] , 
        \nOut1_60[6] , \nOut1_60[5] , \nOut1_60[4] , \nOut1_60[3] , 
        \nOut1_60[2] , \nOut1_60[1] , \nOut1_60[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_59[0] ), .NW_EDGE(\nOut0_58[0] ), .SW_EDGE(
        \nOut0_60[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_20 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut21[31] , \nScanOut21[30] , \nScanOut21[29] , 
        \nScanOut21[28] , \nScanOut21[27] , \nScanOut21[26] , \nScanOut21[25] , 
        \nScanOut21[24] , \nScanOut21[23] , \nScanOut21[22] , \nScanOut21[21] , 
        \nScanOut21[20] , \nScanOut21[19] , \nScanOut21[18] , \nScanOut21[17] , 
        \nScanOut21[16] , \nScanOut21[15] , \nScanOut21[14] , \nScanOut21[13] , 
        \nScanOut21[12] , \nScanOut21[11] , \nScanOut21[10] , \nScanOut21[9] , 
        \nScanOut21[8] , \nScanOut21[7] , \nScanOut21[6] , \nScanOut21[5] , 
        \nScanOut21[4] , \nScanOut21[3] , \nScanOut21[2] , \nScanOut21[1] , 
        \nScanOut21[0] }), .ScanOut({\nScanOut20[31] , \nScanOut20[30] , 
        \nScanOut20[29] , \nScanOut20[28] , \nScanOut20[27] , \nScanOut20[26] , 
        \nScanOut20[25] , \nScanOut20[24] , \nScanOut20[23] , \nScanOut20[22] , 
        \nScanOut20[21] , \nScanOut20[20] , \nScanOut20[19] , \nScanOut20[18] , 
        \nScanOut20[17] , \nScanOut20[16] , \nScanOut20[15] , \nScanOut20[14] , 
        \nScanOut20[13] , \nScanOut20[12] , \nScanOut20[11] , \nScanOut20[10] , 
        \nScanOut20[9] , \nScanOut20[8] , \nScanOut20[7] , \nScanOut20[6] , 
        \nScanOut20[5] , \nScanOut20[4] , \nScanOut20[3] , \nScanOut20[2] , 
        \nScanOut20[1] , \nScanOut20[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_20[31] , 
        \nOut0_20[30] , \nOut0_20[29] , \nOut0_20[28] , \nOut0_20[27] , 
        \nOut0_20[26] , \nOut0_20[25] , \nOut0_20[24] , \nOut0_20[23] , 
        \nOut0_20[22] , \nOut0_20[21] , \nOut0_20[20] , \nOut0_20[19] , 
        \nOut0_20[18] , \nOut0_20[17] , \nOut0_20[16] , \nOut0_20[15] , 
        \nOut0_20[14] , \nOut0_20[13] , \nOut0_20[12] , \nOut0_20[11] , 
        \nOut0_20[10] , \nOut0_20[9] , \nOut0_20[8] , \nOut0_20[7] , 
        \nOut0_20[6] , \nOut0_20[5] , \nOut0_20[4] , \nOut0_20[3] , 
        \nOut0_20[2] , \nOut0_20[1] , \nOut0_20[0] }), .NORTH_EDGE({
        \nOut0_19[31] , \nOut0_19[30] , \nOut0_19[29] , \nOut0_19[28] , 
        \nOut0_19[27] , \nOut0_19[26] , \nOut0_19[25] , \nOut0_19[24] , 
        \nOut0_19[23] , \nOut0_19[22] , \nOut0_19[21] , \nOut0_19[20] , 
        \nOut0_19[19] , \nOut0_19[18] , \nOut0_19[17] , \nOut0_19[16] , 
        \nOut0_19[15] , \nOut0_19[14] , \nOut0_19[13] , \nOut0_19[12] , 
        \nOut0_19[11] , \nOut0_19[10] , \nOut0_19[9] , \nOut0_19[8] , 
        \nOut0_19[7] , \nOut0_19[6] , \nOut0_19[5] , \nOut0_19[4] , 
        \nOut0_19[3] , \nOut0_19[2] , \nOut0_19[1] , \nOut0_19[0] }), 
        .SOUTH_EDGE({\nOut0_21[31] , \nOut0_21[30] , \nOut0_21[29] , 
        \nOut0_21[28] , \nOut0_21[27] , \nOut0_21[26] , \nOut0_21[25] , 
        \nOut0_21[24] , \nOut0_21[23] , \nOut0_21[22] , \nOut0_21[21] , 
        \nOut0_21[20] , \nOut0_21[19] , \nOut0_21[18] , \nOut0_21[17] , 
        \nOut0_21[16] , \nOut0_21[15] , \nOut0_21[14] , \nOut0_21[13] , 
        \nOut0_21[12] , \nOut0_21[11] , \nOut0_21[10] , \nOut0_21[9] , 
        \nOut0_21[8] , \nOut0_21[7] , \nOut0_21[6] , \nOut0_21[5] , 
        \nOut0_21[4] , \nOut0_21[3] , \nOut0_21[2] , \nOut0_21[1] , 
        \nOut0_21[0] }), .EAST_EDGE(\nOut1_20[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_19[31] ), .SE_EDGE(
        \nOut1_21[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_27 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut28[31] , \nScanOut28[30] , \nScanOut28[29] , 
        \nScanOut28[28] , \nScanOut28[27] , \nScanOut28[26] , \nScanOut28[25] , 
        \nScanOut28[24] , \nScanOut28[23] , \nScanOut28[22] , \nScanOut28[21] , 
        \nScanOut28[20] , \nScanOut28[19] , \nScanOut28[18] , \nScanOut28[17] , 
        \nScanOut28[16] , \nScanOut28[15] , \nScanOut28[14] , \nScanOut28[13] , 
        \nScanOut28[12] , \nScanOut28[11] , \nScanOut28[10] , \nScanOut28[9] , 
        \nScanOut28[8] , \nScanOut28[7] , \nScanOut28[6] , \nScanOut28[5] , 
        \nScanOut28[4] , \nScanOut28[3] , \nScanOut28[2] , \nScanOut28[1] , 
        \nScanOut28[0] }), .ScanOut({\nScanOut27[31] , \nScanOut27[30] , 
        \nScanOut27[29] , \nScanOut27[28] , \nScanOut27[27] , \nScanOut27[26] , 
        \nScanOut27[25] , \nScanOut27[24] , \nScanOut27[23] , \nScanOut27[22] , 
        \nScanOut27[21] , \nScanOut27[20] , \nScanOut27[19] , \nScanOut27[18] , 
        \nScanOut27[17] , \nScanOut27[16] , \nScanOut27[15] , \nScanOut27[14] , 
        \nScanOut27[13] , \nScanOut27[12] , \nScanOut27[11] , \nScanOut27[10] , 
        \nScanOut27[9] , \nScanOut27[8] , \nScanOut27[7] , \nScanOut27[6] , 
        \nScanOut27[5] , \nScanOut27[4] , \nScanOut27[3] , \nScanOut27[2] , 
        \nScanOut27[1] , \nScanOut27[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_27[31] , 
        \nOut0_27[30] , \nOut0_27[29] , \nOut0_27[28] , \nOut0_27[27] , 
        \nOut0_27[26] , \nOut0_27[25] , \nOut0_27[24] , \nOut0_27[23] , 
        \nOut0_27[22] , \nOut0_27[21] , \nOut0_27[20] , \nOut0_27[19] , 
        \nOut0_27[18] , \nOut0_27[17] , \nOut0_27[16] , \nOut0_27[15] , 
        \nOut0_27[14] , \nOut0_27[13] , \nOut0_27[12] , \nOut0_27[11] , 
        \nOut0_27[10] , \nOut0_27[9] , \nOut0_27[8] , \nOut0_27[7] , 
        \nOut0_27[6] , \nOut0_27[5] , \nOut0_27[4] , \nOut0_27[3] , 
        \nOut0_27[2] , \nOut0_27[1] , \nOut0_27[0] }), .NORTH_EDGE({
        \nOut0_26[31] , \nOut0_26[30] , \nOut0_26[29] , \nOut0_26[28] , 
        \nOut0_26[27] , \nOut0_26[26] , \nOut0_26[25] , \nOut0_26[24] , 
        \nOut0_26[23] , \nOut0_26[22] , \nOut0_26[21] , \nOut0_26[20] , 
        \nOut0_26[19] , \nOut0_26[18] , \nOut0_26[17] , \nOut0_26[16] , 
        \nOut0_26[15] , \nOut0_26[14] , \nOut0_26[13] , \nOut0_26[12] , 
        \nOut0_26[11] , \nOut0_26[10] , \nOut0_26[9] , \nOut0_26[8] , 
        \nOut0_26[7] , \nOut0_26[6] , \nOut0_26[5] , \nOut0_26[4] , 
        \nOut0_26[3] , \nOut0_26[2] , \nOut0_26[1] , \nOut0_26[0] }), 
        .SOUTH_EDGE({\nOut0_28[31] , \nOut0_28[30] , \nOut0_28[29] , 
        \nOut0_28[28] , \nOut0_28[27] , \nOut0_28[26] , \nOut0_28[25] , 
        \nOut0_28[24] , \nOut0_28[23] , \nOut0_28[22] , \nOut0_28[21] , 
        \nOut0_28[20] , \nOut0_28[19] , \nOut0_28[18] , \nOut0_28[17] , 
        \nOut0_28[16] , \nOut0_28[15] , \nOut0_28[14] , \nOut0_28[13] , 
        \nOut0_28[12] , \nOut0_28[11] , \nOut0_28[10] , \nOut0_28[9] , 
        \nOut0_28[8] , \nOut0_28[7] , \nOut0_28[6] , \nOut0_28[5] , 
        \nOut0_28[4] , \nOut0_28[3] , \nOut0_28[2] , \nOut0_28[1] , 
        \nOut0_28[0] }), .EAST_EDGE(\nOut1_27[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_26[31] ), .SE_EDGE(
        \nOut1_28[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_49 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut50[31] , \nScanOut50[30] , \nScanOut50[29] , 
        \nScanOut50[28] , \nScanOut50[27] , \nScanOut50[26] , \nScanOut50[25] , 
        \nScanOut50[24] , \nScanOut50[23] , \nScanOut50[22] , \nScanOut50[21] , 
        \nScanOut50[20] , \nScanOut50[19] , \nScanOut50[18] , \nScanOut50[17] , 
        \nScanOut50[16] , \nScanOut50[15] , \nScanOut50[14] , \nScanOut50[13] , 
        \nScanOut50[12] , \nScanOut50[11] , \nScanOut50[10] , \nScanOut50[9] , 
        \nScanOut50[8] , \nScanOut50[7] , \nScanOut50[6] , \nScanOut50[5] , 
        \nScanOut50[4] , \nScanOut50[3] , \nScanOut50[2] , \nScanOut50[1] , 
        \nScanOut50[0] }), .ScanOut({\nScanOut49[31] , \nScanOut49[30] , 
        \nScanOut49[29] , \nScanOut49[28] , \nScanOut49[27] , \nScanOut49[26] , 
        \nScanOut49[25] , \nScanOut49[24] , \nScanOut49[23] , \nScanOut49[22] , 
        \nScanOut49[21] , \nScanOut49[20] , \nScanOut49[19] , \nScanOut49[18] , 
        \nScanOut49[17] , \nScanOut49[16] , \nScanOut49[15] , \nScanOut49[14] , 
        \nScanOut49[13] , \nScanOut49[12] , \nScanOut49[11] , \nScanOut49[10] , 
        \nScanOut49[9] , \nScanOut49[8] , \nScanOut49[7] , \nScanOut49[6] , 
        \nScanOut49[5] , \nScanOut49[4] , \nScanOut49[3] , \nScanOut49[2] , 
        \nScanOut49[1] , \nScanOut49[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_49[31] , 
        \nOut0_49[30] , \nOut0_49[29] , \nOut0_49[28] , \nOut0_49[27] , 
        \nOut0_49[26] , \nOut0_49[25] , \nOut0_49[24] , \nOut0_49[23] , 
        \nOut0_49[22] , \nOut0_49[21] , \nOut0_49[20] , \nOut0_49[19] , 
        \nOut0_49[18] , \nOut0_49[17] , \nOut0_49[16] , \nOut0_49[15] , 
        \nOut0_49[14] , \nOut0_49[13] , \nOut0_49[12] , \nOut0_49[11] , 
        \nOut0_49[10] , \nOut0_49[9] , \nOut0_49[8] , \nOut0_49[7] , 
        \nOut0_49[6] , \nOut0_49[5] , \nOut0_49[4] , \nOut0_49[3] , 
        \nOut0_49[2] , \nOut0_49[1] , \nOut0_49[0] }), .NORTH_EDGE({
        \nOut0_48[31] , \nOut0_48[30] , \nOut0_48[29] , \nOut0_48[28] , 
        \nOut0_48[27] , \nOut0_48[26] , \nOut0_48[25] , \nOut0_48[24] , 
        \nOut0_48[23] , \nOut0_48[22] , \nOut0_48[21] , \nOut0_48[20] , 
        \nOut0_48[19] , \nOut0_48[18] , \nOut0_48[17] , \nOut0_48[16] , 
        \nOut0_48[15] , \nOut0_48[14] , \nOut0_48[13] , \nOut0_48[12] , 
        \nOut0_48[11] , \nOut0_48[10] , \nOut0_48[9] , \nOut0_48[8] , 
        \nOut0_48[7] , \nOut0_48[6] , \nOut0_48[5] , \nOut0_48[4] , 
        \nOut0_48[3] , \nOut0_48[2] , \nOut0_48[1] , \nOut0_48[0] }), 
        .SOUTH_EDGE({\nOut0_50[31] , \nOut0_50[30] , \nOut0_50[29] , 
        \nOut0_50[28] , \nOut0_50[27] , \nOut0_50[26] , \nOut0_50[25] , 
        \nOut0_50[24] , \nOut0_50[23] , \nOut0_50[22] , \nOut0_50[21] , 
        \nOut0_50[20] , \nOut0_50[19] , \nOut0_50[18] , \nOut0_50[17] , 
        \nOut0_50[16] , \nOut0_50[15] , \nOut0_50[14] , \nOut0_50[13] , 
        \nOut0_50[12] , \nOut0_50[11] , \nOut0_50[10] , \nOut0_50[9] , 
        \nOut0_50[8] , \nOut0_50[7] , \nOut0_50[6] , \nOut0_50[5] , 
        \nOut0_50[4] , \nOut0_50[3] , \nOut0_50[2] , \nOut0_50[1] , 
        \nOut0_50[0] }), .EAST_EDGE(\nOut1_49[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_48[31] ), .SE_EDGE(
        \nOut1_50[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_55 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut56[31] , \nScanOut56[30] , \nScanOut56[29] , 
        \nScanOut56[28] , \nScanOut56[27] , \nScanOut56[26] , \nScanOut56[25] , 
        \nScanOut56[24] , \nScanOut56[23] , \nScanOut56[22] , \nScanOut56[21] , 
        \nScanOut56[20] , \nScanOut56[19] , \nScanOut56[18] , \nScanOut56[17] , 
        \nScanOut56[16] , \nScanOut56[15] , \nScanOut56[14] , \nScanOut56[13] , 
        \nScanOut56[12] , \nScanOut56[11] , \nScanOut56[10] , \nScanOut56[9] , 
        \nScanOut56[8] , \nScanOut56[7] , \nScanOut56[6] , \nScanOut56[5] , 
        \nScanOut56[4] , \nScanOut56[3] , \nScanOut56[2] , \nScanOut56[1] , 
        \nScanOut56[0] }), .ScanOut({\nScanOut55[31] , \nScanOut55[30] , 
        \nScanOut55[29] , \nScanOut55[28] , \nScanOut55[27] , \nScanOut55[26] , 
        \nScanOut55[25] , \nScanOut55[24] , \nScanOut55[23] , \nScanOut55[22] , 
        \nScanOut55[21] , \nScanOut55[20] , \nScanOut55[19] , \nScanOut55[18] , 
        \nScanOut55[17] , \nScanOut55[16] , \nScanOut55[15] , \nScanOut55[14] , 
        \nScanOut55[13] , \nScanOut55[12] , \nScanOut55[11] , \nScanOut55[10] , 
        \nScanOut55[9] , \nScanOut55[8] , \nScanOut55[7] , \nScanOut55[6] , 
        \nScanOut55[5] , \nScanOut55[4] , \nScanOut55[3] , \nScanOut55[2] , 
        \nScanOut55[1] , \nScanOut55[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_55[31] , 
        \nOut0_55[30] , \nOut0_55[29] , \nOut0_55[28] , \nOut0_55[27] , 
        \nOut0_55[26] , \nOut0_55[25] , \nOut0_55[24] , \nOut0_55[23] , 
        \nOut0_55[22] , \nOut0_55[21] , \nOut0_55[20] , \nOut0_55[19] , 
        \nOut0_55[18] , \nOut0_55[17] , \nOut0_55[16] , \nOut0_55[15] , 
        \nOut0_55[14] , \nOut0_55[13] , \nOut0_55[12] , \nOut0_55[11] , 
        \nOut0_55[10] , \nOut0_55[9] , \nOut0_55[8] , \nOut0_55[7] , 
        \nOut0_55[6] , \nOut0_55[5] , \nOut0_55[4] , \nOut0_55[3] , 
        \nOut0_55[2] , \nOut0_55[1] , \nOut0_55[0] }), .NORTH_EDGE({
        \nOut0_54[31] , \nOut0_54[30] , \nOut0_54[29] , \nOut0_54[28] , 
        \nOut0_54[27] , \nOut0_54[26] , \nOut0_54[25] , \nOut0_54[24] , 
        \nOut0_54[23] , \nOut0_54[22] , \nOut0_54[21] , \nOut0_54[20] , 
        \nOut0_54[19] , \nOut0_54[18] , \nOut0_54[17] , \nOut0_54[16] , 
        \nOut0_54[15] , \nOut0_54[14] , \nOut0_54[13] , \nOut0_54[12] , 
        \nOut0_54[11] , \nOut0_54[10] , \nOut0_54[9] , \nOut0_54[8] , 
        \nOut0_54[7] , \nOut0_54[6] , \nOut0_54[5] , \nOut0_54[4] , 
        \nOut0_54[3] , \nOut0_54[2] , \nOut0_54[1] , \nOut0_54[0] }), 
        .SOUTH_EDGE({\nOut0_56[31] , \nOut0_56[30] , \nOut0_56[29] , 
        \nOut0_56[28] , \nOut0_56[27] , \nOut0_56[26] , \nOut0_56[25] , 
        \nOut0_56[24] , \nOut0_56[23] , \nOut0_56[22] , \nOut0_56[21] , 
        \nOut0_56[20] , \nOut0_56[19] , \nOut0_56[18] , \nOut0_56[17] , 
        \nOut0_56[16] , \nOut0_56[15] , \nOut0_56[14] , \nOut0_56[13] , 
        \nOut0_56[12] , \nOut0_56[11] , \nOut0_56[10] , \nOut0_56[9] , 
        \nOut0_56[8] , \nOut0_56[7] , \nOut0_56[6] , \nOut0_56[5] , 
        \nOut0_56[4] , \nOut0_56[3] , \nOut0_56[2] , \nOut0_56[1] , 
        \nOut0_56[0] }), .EAST_EDGE(\nOut1_55[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_54[31] ), .SE_EDGE(
        \nOut1_56[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_69 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut70[31] , \nScanOut70[30] , \nScanOut70[29] , 
        \nScanOut70[28] , \nScanOut70[27] , \nScanOut70[26] , \nScanOut70[25] , 
        \nScanOut70[24] , \nScanOut70[23] , \nScanOut70[22] , \nScanOut70[21] , 
        \nScanOut70[20] , \nScanOut70[19] , \nScanOut70[18] , \nScanOut70[17] , 
        \nScanOut70[16] , \nScanOut70[15] , \nScanOut70[14] , \nScanOut70[13] , 
        \nScanOut70[12] , \nScanOut70[11] , \nScanOut70[10] , \nScanOut70[9] , 
        \nScanOut70[8] , \nScanOut70[7] , \nScanOut70[6] , \nScanOut70[5] , 
        \nScanOut70[4] , \nScanOut70[3] , \nScanOut70[2] , \nScanOut70[1] , 
        \nScanOut70[0] }), .ScanOut({\nScanOut69[31] , \nScanOut69[30] , 
        \nScanOut69[29] , \nScanOut69[28] , \nScanOut69[27] , \nScanOut69[26] , 
        \nScanOut69[25] , \nScanOut69[24] , \nScanOut69[23] , \nScanOut69[22] , 
        \nScanOut69[21] , \nScanOut69[20] , \nScanOut69[19] , \nScanOut69[18] , 
        \nScanOut69[17] , \nScanOut69[16] , \nScanOut69[15] , \nScanOut69[14] , 
        \nScanOut69[13] , \nScanOut69[12] , \nScanOut69[11] , \nScanOut69[10] , 
        \nScanOut69[9] , \nScanOut69[8] , \nScanOut69[7] , \nScanOut69[6] , 
        \nScanOut69[5] , \nScanOut69[4] , \nScanOut69[3] , \nScanOut69[2] , 
        \nScanOut69[1] , \nScanOut69[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_5[31] , 
        \nOut1_5[30] , \nOut1_5[29] , \nOut1_5[28] , \nOut1_5[27] , 
        \nOut1_5[26] , \nOut1_5[25] , \nOut1_5[24] , \nOut1_5[23] , 
        \nOut1_5[22] , \nOut1_5[21] , \nOut1_5[20] , \nOut1_5[19] , 
        \nOut1_5[18] , \nOut1_5[17] , \nOut1_5[16] , \nOut1_5[15] , 
        \nOut1_5[14] , \nOut1_5[13] , \nOut1_5[12] , \nOut1_5[11] , 
        \nOut1_5[10] , \nOut1_5[9] , \nOut1_5[8] , \nOut1_5[7] , \nOut1_5[6] , 
        \nOut1_5[5] , \nOut1_5[4] , \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , 
        \nOut1_5[0] }), .NORTH_EDGE({\nOut1_4[31] , \nOut1_4[30] , 
        \nOut1_4[29] , \nOut1_4[28] , \nOut1_4[27] , \nOut1_4[26] , 
        \nOut1_4[25] , \nOut1_4[24] , \nOut1_4[23] , \nOut1_4[22] , 
        \nOut1_4[21] , \nOut1_4[20] , \nOut1_4[19] , \nOut1_4[18] , 
        \nOut1_4[17] , \nOut1_4[16] , \nOut1_4[15] , \nOut1_4[14] , 
        \nOut1_4[13] , \nOut1_4[12] , \nOut1_4[11] , \nOut1_4[10] , 
        \nOut1_4[9] , \nOut1_4[8] , \nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , 
        \nOut1_4[4] , \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }), 
        .SOUTH_EDGE({\nOut1_6[31] , \nOut1_6[30] , \nOut1_6[29] , 
        \nOut1_6[28] , \nOut1_6[27] , \nOut1_6[26] , \nOut1_6[25] , 
        \nOut1_6[24] , \nOut1_6[23] , \nOut1_6[22] , \nOut1_6[21] , 
        \nOut1_6[20] , \nOut1_6[19] , \nOut1_6[18] , \nOut1_6[17] , 
        \nOut1_6[16] , \nOut1_6[15] , \nOut1_6[14] , \nOut1_6[13] , 
        \nOut1_6[12] , \nOut1_6[11] , \nOut1_6[10] , \nOut1_6[9] , 
        \nOut1_6[8] , \nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , \nOut1_6[4] , 
        \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_5[0] ), .NW_EDGE(\nOut0_4[0] ), .SW_EDGE(
        \nOut0_6[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_118 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut119[31] , \nScanOut119[30] , \nScanOut119[29] , 
        \nScanOut119[28] , \nScanOut119[27] , \nScanOut119[26] , 
        \nScanOut119[25] , \nScanOut119[24] , \nScanOut119[23] , 
        \nScanOut119[22] , \nScanOut119[21] , \nScanOut119[20] , 
        \nScanOut119[19] , \nScanOut119[18] , \nScanOut119[17] , 
        \nScanOut119[16] , \nScanOut119[15] , \nScanOut119[14] , 
        \nScanOut119[13] , \nScanOut119[12] , \nScanOut119[11] , 
        \nScanOut119[10] , \nScanOut119[9] , \nScanOut119[8] , 
        \nScanOut119[7] , \nScanOut119[6] , \nScanOut119[5] , \nScanOut119[4] , 
        \nScanOut119[3] , \nScanOut119[2] , \nScanOut119[1] , \nScanOut119[0] 
        }), .ScanOut({\nScanOut118[31] , \nScanOut118[30] , \nScanOut118[29] , 
        \nScanOut118[28] , \nScanOut118[27] , \nScanOut118[26] , 
        \nScanOut118[25] , \nScanOut118[24] , \nScanOut118[23] , 
        \nScanOut118[22] , \nScanOut118[21] , \nScanOut118[20] , 
        \nScanOut118[19] , \nScanOut118[18] , \nScanOut118[17] , 
        \nScanOut118[16] , \nScanOut118[15] , \nScanOut118[14] , 
        \nScanOut118[13] , \nScanOut118[12] , \nScanOut118[11] , 
        \nScanOut118[10] , \nScanOut118[9] , \nScanOut118[8] , 
        \nScanOut118[7] , \nScanOut118[6] , \nScanOut118[5] , \nScanOut118[4] , 
        \nScanOut118[3] , \nScanOut118[2] , \nScanOut118[1] , \nScanOut118[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_54[31] , \nOut1_54[30] , \nOut1_54[29] , 
        \nOut1_54[28] , \nOut1_54[27] , \nOut1_54[26] , \nOut1_54[25] , 
        \nOut1_54[24] , \nOut1_54[23] , \nOut1_54[22] , \nOut1_54[21] , 
        \nOut1_54[20] , \nOut1_54[19] , \nOut1_54[18] , \nOut1_54[17] , 
        \nOut1_54[16] , \nOut1_54[15] , \nOut1_54[14] , \nOut1_54[13] , 
        \nOut1_54[12] , \nOut1_54[11] , \nOut1_54[10] , \nOut1_54[9] , 
        \nOut1_54[8] , \nOut1_54[7] , \nOut1_54[6] , \nOut1_54[5] , 
        \nOut1_54[4] , \nOut1_54[3] , \nOut1_54[2] , \nOut1_54[1] , 
        \nOut1_54[0] }), .NORTH_EDGE({\nOut1_53[31] , \nOut1_53[30] , 
        \nOut1_53[29] , \nOut1_53[28] , \nOut1_53[27] , \nOut1_53[26] , 
        \nOut1_53[25] , \nOut1_53[24] , \nOut1_53[23] , \nOut1_53[22] , 
        \nOut1_53[21] , \nOut1_53[20] , \nOut1_53[19] , \nOut1_53[18] , 
        \nOut1_53[17] , \nOut1_53[16] , \nOut1_53[15] , \nOut1_53[14] , 
        \nOut1_53[13] , \nOut1_53[12] , \nOut1_53[11] , \nOut1_53[10] , 
        \nOut1_53[9] , \nOut1_53[8] , \nOut1_53[7] , \nOut1_53[6] , 
        \nOut1_53[5] , \nOut1_53[4] , \nOut1_53[3] , \nOut1_53[2] , 
        \nOut1_53[1] , \nOut1_53[0] }), .SOUTH_EDGE({\nOut1_55[31] , 
        \nOut1_55[30] , \nOut1_55[29] , \nOut1_55[28] , \nOut1_55[27] , 
        \nOut1_55[26] , \nOut1_55[25] , \nOut1_55[24] , \nOut1_55[23] , 
        \nOut1_55[22] , \nOut1_55[21] , \nOut1_55[20] , \nOut1_55[19] , 
        \nOut1_55[18] , \nOut1_55[17] , \nOut1_55[16] , \nOut1_55[15] , 
        \nOut1_55[14] , \nOut1_55[13] , \nOut1_55[12] , \nOut1_55[11] , 
        \nOut1_55[10] , \nOut1_55[9] , \nOut1_55[8] , \nOut1_55[7] , 
        \nOut1_55[6] , \nOut1_55[5] , \nOut1_55[4] , \nOut1_55[3] , 
        \nOut1_55[2] , \nOut1_55[1] , \nOut1_55[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_54[0] ), .NW_EDGE(\nOut0_53[0] ), .SW_EDGE(
        \nOut0_55[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_72 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut73[31] , \nScanOut73[30] , \nScanOut73[29] , 
        \nScanOut73[28] , \nScanOut73[27] , \nScanOut73[26] , \nScanOut73[25] , 
        \nScanOut73[24] , \nScanOut73[23] , \nScanOut73[22] , \nScanOut73[21] , 
        \nScanOut73[20] , \nScanOut73[19] , \nScanOut73[18] , \nScanOut73[17] , 
        \nScanOut73[16] , \nScanOut73[15] , \nScanOut73[14] , \nScanOut73[13] , 
        \nScanOut73[12] , \nScanOut73[11] , \nScanOut73[10] , \nScanOut73[9] , 
        \nScanOut73[8] , \nScanOut73[7] , \nScanOut73[6] , \nScanOut73[5] , 
        \nScanOut73[4] , \nScanOut73[3] , \nScanOut73[2] , \nScanOut73[1] , 
        \nScanOut73[0] }), .ScanOut({\nScanOut72[31] , \nScanOut72[30] , 
        \nScanOut72[29] , \nScanOut72[28] , \nScanOut72[27] , \nScanOut72[26] , 
        \nScanOut72[25] , \nScanOut72[24] , \nScanOut72[23] , \nScanOut72[22] , 
        \nScanOut72[21] , \nScanOut72[20] , \nScanOut72[19] , \nScanOut72[18] , 
        \nScanOut72[17] , \nScanOut72[16] , \nScanOut72[15] , \nScanOut72[14] , 
        \nScanOut72[13] , \nScanOut72[12] , \nScanOut72[11] , \nScanOut72[10] , 
        \nScanOut72[9] , \nScanOut72[8] , \nScanOut72[7] , \nScanOut72[6] , 
        \nScanOut72[5] , \nScanOut72[4] , \nScanOut72[3] , \nScanOut72[2] , 
        \nScanOut72[1] , \nScanOut72[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_8[31] , 
        \nOut1_8[30] , \nOut1_8[29] , \nOut1_8[28] , \nOut1_8[27] , 
        \nOut1_8[26] , \nOut1_8[25] , \nOut1_8[24] , \nOut1_8[23] , 
        \nOut1_8[22] , \nOut1_8[21] , \nOut1_8[20] , \nOut1_8[19] , 
        \nOut1_8[18] , \nOut1_8[17] , \nOut1_8[16] , \nOut1_8[15] , 
        \nOut1_8[14] , \nOut1_8[13] , \nOut1_8[12] , \nOut1_8[11] , 
        \nOut1_8[10] , \nOut1_8[9] , \nOut1_8[8] , \nOut1_8[7] , \nOut1_8[6] , 
        \nOut1_8[5] , \nOut1_8[4] , \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , 
        \nOut1_8[0] }), .NORTH_EDGE({\nOut1_7[31] , \nOut1_7[30] , 
        \nOut1_7[29] , \nOut1_7[28] , \nOut1_7[27] , \nOut1_7[26] , 
        \nOut1_7[25] , \nOut1_7[24] , \nOut1_7[23] , \nOut1_7[22] , 
        \nOut1_7[21] , \nOut1_7[20] , \nOut1_7[19] , \nOut1_7[18] , 
        \nOut1_7[17] , \nOut1_7[16] , \nOut1_7[15] , \nOut1_7[14] , 
        \nOut1_7[13] , \nOut1_7[12] , \nOut1_7[11] , \nOut1_7[10] , 
        \nOut1_7[9] , \nOut1_7[8] , \nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , 
        \nOut1_7[4] , \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }), 
        .SOUTH_EDGE({\nOut1_9[31] , \nOut1_9[30] , \nOut1_9[29] , 
        \nOut1_9[28] , \nOut1_9[27] , \nOut1_9[26] , \nOut1_9[25] , 
        \nOut1_9[24] , \nOut1_9[23] , \nOut1_9[22] , \nOut1_9[21] , 
        \nOut1_9[20] , \nOut1_9[19] , \nOut1_9[18] , \nOut1_9[17] , 
        \nOut1_9[16] , \nOut1_9[15] , \nOut1_9[14] , \nOut1_9[13] , 
        \nOut1_9[12] , \nOut1_9[11] , \nOut1_9[10] , \nOut1_9[9] , 
        \nOut1_9[8] , \nOut1_9[7] , \nOut1_9[6] , \nOut1_9[5] , \nOut1_9[4] , 
        \nOut1_9[3] , \nOut1_9[2] , \nOut1_9[1] , \nOut1_9[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_8[0] ), .NW_EDGE(\nOut0_7[0] ), .SW_EDGE(
        \nOut0_9[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_103 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut104[31] , \nScanOut104[30] , \nScanOut104[29] , 
        \nScanOut104[28] , \nScanOut104[27] , \nScanOut104[26] , 
        \nScanOut104[25] , \nScanOut104[24] , \nScanOut104[23] , 
        \nScanOut104[22] , \nScanOut104[21] , \nScanOut104[20] , 
        \nScanOut104[19] , \nScanOut104[18] , \nScanOut104[17] , 
        \nScanOut104[16] , \nScanOut104[15] , \nScanOut104[14] , 
        \nScanOut104[13] , \nScanOut104[12] , \nScanOut104[11] , 
        \nScanOut104[10] , \nScanOut104[9] , \nScanOut104[8] , 
        \nScanOut104[7] , \nScanOut104[6] , \nScanOut104[5] , \nScanOut104[4] , 
        \nScanOut104[3] , \nScanOut104[2] , \nScanOut104[1] , \nScanOut104[0] 
        }), .ScanOut({\nScanOut103[31] , \nScanOut103[30] , \nScanOut103[29] , 
        \nScanOut103[28] , \nScanOut103[27] , \nScanOut103[26] , 
        \nScanOut103[25] , \nScanOut103[24] , \nScanOut103[23] , 
        \nScanOut103[22] , \nScanOut103[21] , \nScanOut103[20] , 
        \nScanOut103[19] , \nScanOut103[18] , \nScanOut103[17] , 
        \nScanOut103[16] , \nScanOut103[15] , \nScanOut103[14] , 
        \nScanOut103[13] , \nScanOut103[12] , \nScanOut103[11] , 
        \nScanOut103[10] , \nScanOut103[9] , \nScanOut103[8] , 
        \nScanOut103[7] , \nScanOut103[6] , \nScanOut103[5] , \nScanOut103[4] , 
        \nScanOut103[3] , \nScanOut103[2] , \nScanOut103[1] , \nScanOut103[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_39[31] , \nOut1_39[30] , \nOut1_39[29] , 
        \nOut1_39[28] , \nOut1_39[27] , \nOut1_39[26] , \nOut1_39[25] , 
        \nOut1_39[24] , \nOut1_39[23] , \nOut1_39[22] , \nOut1_39[21] , 
        \nOut1_39[20] , \nOut1_39[19] , \nOut1_39[18] , \nOut1_39[17] , 
        \nOut1_39[16] , \nOut1_39[15] , \nOut1_39[14] , \nOut1_39[13] , 
        \nOut1_39[12] , \nOut1_39[11] , \nOut1_39[10] , \nOut1_39[9] , 
        \nOut1_39[8] , \nOut1_39[7] , \nOut1_39[6] , \nOut1_39[5] , 
        \nOut1_39[4] , \nOut1_39[3] , \nOut1_39[2] , \nOut1_39[1] , 
        \nOut1_39[0] }), .NORTH_EDGE({\nOut1_38[31] , \nOut1_38[30] , 
        \nOut1_38[29] , \nOut1_38[28] , \nOut1_38[27] , \nOut1_38[26] , 
        \nOut1_38[25] , \nOut1_38[24] , \nOut1_38[23] , \nOut1_38[22] , 
        \nOut1_38[21] , \nOut1_38[20] , \nOut1_38[19] , \nOut1_38[18] , 
        \nOut1_38[17] , \nOut1_38[16] , \nOut1_38[15] , \nOut1_38[14] , 
        \nOut1_38[13] , \nOut1_38[12] , \nOut1_38[11] , \nOut1_38[10] , 
        \nOut1_38[9] , \nOut1_38[8] , \nOut1_38[7] , \nOut1_38[6] , 
        \nOut1_38[5] , \nOut1_38[4] , \nOut1_38[3] , \nOut1_38[2] , 
        \nOut1_38[1] , \nOut1_38[0] }), .SOUTH_EDGE({\nOut1_40[31] , 
        \nOut1_40[30] , \nOut1_40[29] , \nOut1_40[28] , \nOut1_40[27] , 
        \nOut1_40[26] , \nOut1_40[25] , \nOut1_40[24] , \nOut1_40[23] , 
        \nOut1_40[22] , \nOut1_40[21] , \nOut1_40[20] , \nOut1_40[19] , 
        \nOut1_40[18] , \nOut1_40[17] , \nOut1_40[16] , \nOut1_40[15] , 
        \nOut1_40[14] , \nOut1_40[13] , \nOut1_40[12] , \nOut1_40[11] , 
        \nOut1_40[10] , \nOut1_40[9] , \nOut1_40[8] , \nOut1_40[7] , 
        \nOut1_40[6] , \nOut1_40[5] , \nOut1_40[4] , \nOut1_40[3] , 
        \nOut1_40[2] , \nOut1_40[1] , \nOut1_40[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_39[0] ), .NW_EDGE(\nOut0_38[0] ), .SW_EDGE(
        \nOut0_40[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_124 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut125[31] , \nScanOut125[30] , \nScanOut125[29] , 
        \nScanOut125[28] , \nScanOut125[27] , \nScanOut125[26] , 
        \nScanOut125[25] , \nScanOut125[24] , \nScanOut125[23] , 
        \nScanOut125[22] , \nScanOut125[21] , \nScanOut125[20] , 
        \nScanOut125[19] , \nScanOut125[18] , \nScanOut125[17] , 
        \nScanOut125[16] , \nScanOut125[15] , \nScanOut125[14] , 
        \nScanOut125[13] , \nScanOut125[12] , \nScanOut125[11] , 
        \nScanOut125[10] , \nScanOut125[9] , \nScanOut125[8] , 
        \nScanOut125[7] , \nScanOut125[6] , \nScanOut125[5] , \nScanOut125[4] , 
        \nScanOut125[3] , \nScanOut125[2] , \nScanOut125[1] , \nScanOut125[0] 
        }), .ScanOut({\nScanOut124[31] , \nScanOut124[30] , \nScanOut124[29] , 
        \nScanOut124[28] , \nScanOut124[27] , \nScanOut124[26] , 
        \nScanOut124[25] , \nScanOut124[24] , \nScanOut124[23] , 
        \nScanOut124[22] , \nScanOut124[21] , \nScanOut124[20] , 
        \nScanOut124[19] , \nScanOut124[18] , \nScanOut124[17] , 
        \nScanOut124[16] , \nScanOut124[15] , \nScanOut124[14] , 
        \nScanOut124[13] , \nScanOut124[12] , \nScanOut124[11] , 
        \nScanOut124[10] , \nScanOut124[9] , \nScanOut124[8] , 
        \nScanOut124[7] , \nScanOut124[6] , \nScanOut124[5] , \nScanOut124[4] , 
        \nScanOut124[3] , \nScanOut124[2] , \nScanOut124[1] , \nScanOut124[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_60[31] , \nOut1_60[30] , \nOut1_60[29] , 
        \nOut1_60[28] , \nOut1_60[27] , \nOut1_60[26] , \nOut1_60[25] , 
        \nOut1_60[24] , \nOut1_60[23] , \nOut1_60[22] , \nOut1_60[21] , 
        \nOut1_60[20] , \nOut1_60[19] , \nOut1_60[18] , \nOut1_60[17] , 
        \nOut1_60[16] , \nOut1_60[15] , \nOut1_60[14] , \nOut1_60[13] , 
        \nOut1_60[12] , \nOut1_60[11] , \nOut1_60[10] , \nOut1_60[9] , 
        \nOut1_60[8] , \nOut1_60[7] , \nOut1_60[6] , \nOut1_60[5] , 
        \nOut1_60[4] , \nOut1_60[3] , \nOut1_60[2] , \nOut1_60[1] , 
        \nOut1_60[0] }), .NORTH_EDGE({\nOut1_59[31] , \nOut1_59[30] , 
        \nOut1_59[29] , \nOut1_59[28] , \nOut1_59[27] , \nOut1_59[26] , 
        \nOut1_59[25] , \nOut1_59[24] , \nOut1_59[23] , \nOut1_59[22] , 
        \nOut1_59[21] , \nOut1_59[20] , \nOut1_59[19] , \nOut1_59[18] , 
        \nOut1_59[17] , \nOut1_59[16] , \nOut1_59[15] , \nOut1_59[14] , 
        \nOut1_59[13] , \nOut1_59[12] , \nOut1_59[11] , \nOut1_59[10] , 
        \nOut1_59[9] , \nOut1_59[8] , \nOut1_59[7] , \nOut1_59[6] , 
        \nOut1_59[5] , \nOut1_59[4] , \nOut1_59[3] , \nOut1_59[2] , 
        \nOut1_59[1] , \nOut1_59[0] }), .SOUTH_EDGE({\nOut1_61[31] , 
        \nOut1_61[30] , \nOut1_61[29] , \nOut1_61[28] , \nOut1_61[27] , 
        \nOut1_61[26] , \nOut1_61[25] , \nOut1_61[24] , \nOut1_61[23] , 
        \nOut1_61[22] , \nOut1_61[21] , \nOut1_61[20] , \nOut1_61[19] , 
        \nOut1_61[18] , \nOut1_61[17] , \nOut1_61[16] , \nOut1_61[15] , 
        \nOut1_61[14] , \nOut1_61[13] , \nOut1_61[12] , \nOut1_61[11] , 
        \nOut1_61[10] , \nOut1_61[9] , \nOut1_61[8] , \nOut1_61[7] , 
        \nOut1_61[6] , \nOut1_61[5] , \nOut1_61[4] , \nOut1_61[3] , 
        \nOut1_61[2] , \nOut1_61[1] , \nOut1_61[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_60[0] ), .NW_EDGE(\nOut0_59[0] ), .SW_EDGE(
        \nOut0_61[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut16[31] , \nScanOut16[30] , \nScanOut16[29] , 
        \nScanOut16[28] , \nScanOut16[27] , \nScanOut16[26] , \nScanOut16[25] , 
        \nScanOut16[24] , \nScanOut16[23] , \nScanOut16[22] , \nScanOut16[21] , 
        \nScanOut16[20] , \nScanOut16[19] , \nScanOut16[18] , \nScanOut16[17] , 
        \nScanOut16[16] , \nScanOut16[15] , \nScanOut16[14] , \nScanOut16[13] , 
        \nScanOut16[12] , \nScanOut16[11] , \nScanOut16[10] , \nScanOut16[9] , 
        \nScanOut16[8] , \nScanOut16[7] , \nScanOut16[6] , \nScanOut16[5] , 
        \nScanOut16[4] , \nScanOut16[3] , \nScanOut16[2] , \nScanOut16[1] , 
        \nScanOut16[0] }), .ScanOut({\nScanOut15[31] , \nScanOut15[30] , 
        \nScanOut15[29] , \nScanOut15[28] , \nScanOut15[27] , \nScanOut15[26] , 
        \nScanOut15[25] , \nScanOut15[24] , \nScanOut15[23] , \nScanOut15[22] , 
        \nScanOut15[21] , \nScanOut15[20] , \nScanOut15[19] , \nScanOut15[18] , 
        \nScanOut15[17] , \nScanOut15[16] , \nScanOut15[15] , \nScanOut15[14] , 
        \nScanOut15[13] , \nScanOut15[12] , \nScanOut15[11] , \nScanOut15[10] , 
        \nScanOut15[9] , \nScanOut15[8] , \nScanOut15[7] , \nScanOut15[6] , 
        \nScanOut15[5] , \nScanOut15[4] , \nScanOut15[3] , \nScanOut15[2] , 
        \nScanOut15[1] , \nScanOut15[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_15[31] , 
        \nOut0_15[30] , \nOut0_15[29] , \nOut0_15[28] , \nOut0_15[27] , 
        \nOut0_15[26] , \nOut0_15[25] , \nOut0_15[24] , \nOut0_15[23] , 
        \nOut0_15[22] , \nOut0_15[21] , \nOut0_15[20] , \nOut0_15[19] , 
        \nOut0_15[18] , \nOut0_15[17] , \nOut0_15[16] , \nOut0_15[15] , 
        \nOut0_15[14] , \nOut0_15[13] , \nOut0_15[12] , \nOut0_15[11] , 
        \nOut0_15[10] , \nOut0_15[9] , \nOut0_15[8] , \nOut0_15[7] , 
        \nOut0_15[6] , \nOut0_15[5] , \nOut0_15[4] , \nOut0_15[3] , 
        \nOut0_15[2] , \nOut0_15[1] , \nOut0_15[0] }), .NORTH_EDGE({
        \nOut0_14[31] , \nOut0_14[30] , \nOut0_14[29] , \nOut0_14[28] , 
        \nOut0_14[27] , \nOut0_14[26] , \nOut0_14[25] , \nOut0_14[24] , 
        \nOut0_14[23] , \nOut0_14[22] , \nOut0_14[21] , \nOut0_14[20] , 
        \nOut0_14[19] , \nOut0_14[18] , \nOut0_14[17] , \nOut0_14[16] , 
        \nOut0_14[15] , \nOut0_14[14] , \nOut0_14[13] , \nOut0_14[12] , 
        \nOut0_14[11] , \nOut0_14[10] , \nOut0_14[9] , \nOut0_14[8] , 
        \nOut0_14[7] , \nOut0_14[6] , \nOut0_14[5] , \nOut0_14[4] , 
        \nOut0_14[3] , \nOut0_14[2] , \nOut0_14[1] , \nOut0_14[0] }), 
        .SOUTH_EDGE({\nOut0_16[31] , \nOut0_16[30] , \nOut0_16[29] , 
        \nOut0_16[28] , \nOut0_16[27] , \nOut0_16[26] , \nOut0_16[25] , 
        \nOut0_16[24] , \nOut0_16[23] , \nOut0_16[22] , \nOut0_16[21] , 
        \nOut0_16[20] , \nOut0_16[19] , \nOut0_16[18] , \nOut0_16[17] , 
        \nOut0_16[16] , \nOut0_16[15] , \nOut0_16[14] , \nOut0_16[13] , 
        \nOut0_16[12] , \nOut0_16[11] , \nOut0_16[10] , \nOut0_16[9] , 
        \nOut0_16[8] , \nOut0_16[7] , \nOut0_16[6] , \nOut0_16[5] , 
        \nOut0_16[4] , \nOut0_16[3] , \nOut0_16[2] , \nOut0_16[1] , 
        \nOut0_16[0] }), .EAST_EDGE(\nOut1_15[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_14[31] ), .SE_EDGE(
        \nOut1_16[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_29 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut30[31] , \nScanOut30[30] , \nScanOut30[29] , 
        \nScanOut30[28] , \nScanOut30[27] , \nScanOut30[26] , \nScanOut30[25] , 
        \nScanOut30[24] , \nScanOut30[23] , \nScanOut30[22] , \nScanOut30[21] , 
        \nScanOut30[20] , \nScanOut30[19] , \nScanOut30[18] , \nScanOut30[17] , 
        \nScanOut30[16] , \nScanOut30[15] , \nScanOut30[14] , \nScanOut30[13] , 
        \nScanOut30[12] , \nScanOut30[11] , \nScanOut30[10] , \nScanOut30[9] , 
        \nScanOut30[8] , \nScanOut30[7] , \nScanOut30[6] , \nScanOut30[5] , 
        \nScanOut30[4] , \nScanOut30[3] , \nScanOut30[2] , \nScanOut30[1] , 
        \nScanOut30[0] }), .ScanOut({\nScanOut29[31] , \nScanOut29[30] , 
        \nScanOut29[29] , \nScanOut29[28] , \nScanOut29[27] , \nScanOut29[26] , 
        \nScanOut29[25] , \nScanOut29[24] , \nScanOut29[23] , \nScanOut29[22] , 
        \nScanOut29[21] , \nScanOut29[20] , \nScanOut29[19] , \nScanOut29[18] , 
        \nScanOut29[17] , \nScanOut29[16] , \nScanOut29[15] , \nScanOut29[14] , 
        \nScanOut29[13] , \nScanOut29[12] , \nScanOut29[11] , \nScanOut29[10] , 
        \nScanOut29[9] , \nScanOut29[8] , \nScanOut29[7] , \nScanOut29[6] , 
        \nScanOut29[5] , \nScanOut29[4] , \nScanOut29[3] , \nScanOut29[2] , 
        \nScanOut29[1] , \nScanOut29[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_29[31] , 
        \nOut0_29[30] , \nOut0_29[29] , \nOut0_29[28] , \nOut0_29[27] , 
        \nOut0_29[26] , \nOut0_29[25] , \nOut0_29[24] , \nOut0_29[23] , 
        \nOut0_29[22] , \nOut0_29[21] , \nOut0_29[20] , \nOut0_29[19] , 
        \nOut0_29[18] , \nOut0_29[17] , \nOut0_29[16] , \nOut0_29[15] , 
        \nOut0_29[14] , \nOut0_29[13] , \nOut0_29[12] , \nOut0_29[11] , 
        \nOut0_29[10] , \nOut0_29[9] , \nOut0_29[8] , \nOut0_29[7] , 
        \nOut0_29[6] , \nOut0_29[5] , \nOut0_29[4] , \nOut0_29[3] , 
        \nOut0_29[2] , \nOut0_29[1] , \nOut0_29[0] }), .NORTH_EDGE({
        \nOut0_28[31] , \nOut0_28[30] , \nOut0_28[29] , \nOut0_28[28] , 
        \nOut0_28[27] , \nOut0_28[26] , \nOut0_28[25] , \nOut0_28[24] , 
        \nOut0_28[23] , \nOut0_28[22] , \nOut0_28[21] , \nOut0_28[20] , 
        \nOut0_28[19] , \nOut0_28[18] , \nOut0_28[17] , \nOut0_28[16] , 
        \nOut0_28[15] , \nOut0_28[14] , \nOut0_28[13] , \nOut0_28[12] , 
        \nOut0_28[11] , \nOut0_28[10] , \nOut0_28[9] , \nOut0_28[8] , 
        \nOut0_28[7] , \nOut0_28[6] , \nOut0_28[5] , \nOut0_28[4] , 
        \nOut0_28[3] , \nOut0_28[2] , \nOut0_28[1] , \nOut0_28[0] }), 
        .SOUTH_EDGE({\nOut0_30[31] , \nOut0_30[30] , \nOut0_30[29] , 
        \nOut0_30[28] , \nOut0_30[27] , \nOut0_30[26] , \nOut0_30[25] , 
        \nOut0_30[24] , \nOut0_30[23] , \nOut0_30[22] , \nOut0_30[21] , 
        \nOut0_30[20] , \nOut0_30[19] , \nOut0_30[18] , \nOut0_30[17] , 
        \nOut0_30[16] , \nOut0_30[15] , \nOut0_30[14] , \nOut0_30[13] , 
        \nOut0_30[12] , \nOut0_30[11] , \nOut0_30[10] , \nOut0_30[9] , 
        \nOut0_30[8] , \nOut0_30[7] , \nOut0_30[6] , \nOut0_30[5] , 
        \nOut0_30[4] , \nOut0_30[3] , \nOut0_30[2] , \nOut0_30[1] , 
        \nOut0_30[0] }), .EAST_EDGE(\nOut1_29[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_28[31] ), .SE_EDGE(
        \nOut1_30[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_97 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut98[31] , \nScanOut98[30] , \nScanOut98[29] , 
        \nScanOut98[28] , \nScanOut98[27] , \nScanOut98[26] , \nScanOut98[25] , 
        \nScanOut98[24] , \nScanOut98[23] , \nScanOut98[22] , \nScanOut98[21] , 
        \nScanOut98[20] , \nScanOut98[19] , \nScanOut98[18] , \nScanOut98[17] , 
        \nScanOut98[16] , \nScanOut98[15] , \nScanOut98[14] , \nScanOut98[13] , 
        \nScanOut98[12] , \nScanOut98[11] , \nScanOut98[10] , \nScanOut98[9] , 
        \nScanOut98[8] , \nScanOut98[7] , \nScanOut98[6] , \nScanOut98[5] , 
        \nScanOut98[4] , \nScanOut98[3] , \nScanOut98[2] , \nScanOut98[1] , 
        \nScanOut98[0] }), .ScanOut({\nScanOut97[31] , \nScanOut97[30] , 
        \nScanOut97[29] , \nScanOut97[28] , \nScanOut97[27] , \nScanOut97[26] , 
        \nScanOut97[25] , \nScanOut97[24] , \nScanOut97[23] , \nScanOut97[22] , 
        \nScanOut97[21] , \nScanOut97[20] , \nScanOut97[19] , \nScanOut97[18] , 
        \nScanOut97[17] , \nScanOut97[16] , \nScanOut97[15] , \nScanOut97[14] , 
        \nScanOut97[13] , \nScanOut97[12] , \nScanOut97[11] , \nScanOut97[10] , 
        \nScanOut97[9] , \nScanOut97[8] , \nScanOut97[7] , \nScanOut97[6] , 
        \nScanOut97[5] , \nScanOut97[4] , \nScanOut97[3] , \nScanOut97[2] , 
        \nScanOut97[1] , \nScanOut97[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_33[31] , 
        \nOut1_33[30] , \nOut1_33[29] , \nOut1_33[28] , \nOut1_33[27] , 
        \nOut1_33[26] , \nOut1_33[25] , \nOut1_33[24] , \nOut1_33[23] , 
        \nOut1_33[22] , \nOut1_33[21] , \nOut1_33[20] , \nOut1_33[19] , 
        \nOut1_33[18] , \nOut1_33[17] , \nOut1_33[16] , \nOut1_33[15] , 
        \nOut1_33[14] , \nOut1_33[13] , \nOut1_33[12] , \nOut1_33[11] , 
        \nOut1_33[10] , \nOut1_33[9] , \nOut1_33[8] , \nOut1_33[7] , 
        \nOut1_33[6] , \nOut1_33[5] , \nOut1_33[4] , \nOut1_33[3] , 
        \nOut1_33[2] , \nOut1_33[1] , \nOut1_33[0] }), .NORTH_EDGE({
        \nOut1_32[31] , \nOut1_32[30] , \nOut1_32[29] , \nOut1_32[28] , 
        \nOut1_32[27] , \nOut1_32[26] , \nOut1_32[25] , \nOut1_32[24] , 
        \nOut1_32[23] , \nOut1_32[22] , \nOut1_32[21] , \nOut1_32[20] , 
        \nOut1_32[19] , \nOut1_32[18] , \nOut1_32[17] , \nOut1_32[16] , 
        \nOut1_32[15] , \nOut1_32[14] , \nOut1_32[13] , \nOut1_32[12] , 
        \nOut1_32[11] , \nOut1_32[10] , \nOut1_32[9] , \nOut1_32[8] , 
        \nOut1_32[7] , \nOut1_32[6] , \nOut1_32[5] , \nOut1_32[4] , 
        \nOut1_32[3] , \nOut1_32[2] , \nOut1_32[1] , \nOut1_32[0] }), 
        .SOUTH_EDGE({\nOut1_34[31] , \nOut1_34[30] , \nOut1_34[29] , 
        \nOut1_34[28] , \nOut1_34[27] , \nOut1_34[26] , \nOut1_34[25] , 
        \nOut1_34[24] , \nOut1_34[23] , \nOut1_34[22] , \nOut1_34[21] , 
        \nOut1_34[20] , \nOut1_34[19] , \nOut1_34[18] , \nOut1_34[17] , 
        \nOut1_34[16] , \nOut1_34[15] , \nOut1_34[14] , \nOut1_34[13] , 
        \nOut1_34[12] , \nOut1_34[11] , \nOut1_34[10] , \nOut1_34[9] , 
        \nOut1_34[8] , \nOut1_34[7] , \nOut1_34[6] , \nOut1_34[5] , 
        \nOut1_34[4] , \nOut1_34[3] , \nOut1_34[2] , \nOut1_34[1] , 
        \nOut1_34[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_33[0] ), 
        .NW_EDGE(\nOut0_32[0] ), .SW_EDGE(\nOut0_34[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_32 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut33[31] , \nScanOut33[30] , \nScanOut33[29] , 
        \nScanOut33[28] , \nScanOut33[27] , \nScanOut33[26] , \nScanOut33[25] , 
        \nScanOut33[24] , \nScanOut33[23] , \nScanOut33[22] , \nScanOut33[21] , 
        \nScanOut33[20] , \nScanOut33[19] , \nScanOut33[18] , \nScanOut33[17] , 
        \nScanOut33[16] , \nScanOut33[15] , \nScanOut33[14] , \nScanOut33[13] , 
        \nScanOut33[12] , \nScanOut33[11] , \nScanOut33[10] , \nScanOut33[9] , 
        \nScanOut33[8] , \nScanOut33[7] , \nScanOut33[6] , \nScanOut33[5] , 
        \nScanOut33[4] , \nScanOut33[3] , \nScanOut33[2] , \nScanOut33[1] , 
        \nScanOut33[0] }), .ScanOut({\nScanOut32[31] , \nScanOut32[30] , 
        \nScanOut32[29] , \nScanOut32[28] , \nScanOut32[27] , \nScanOut32[26] , 
        \nScanOut32[25] , \nScanOut32[24] , \nScanOut32[23] , \nScanOut32[22] , 
        \nScanOut32[21] , \nScanOut32[20] , \nScanOut32[19] , \nScanOut32[18] , 
        \nScanOut32[17] , \nScanOut32[16] , \nScanOut32[15] , \nScanOut32[14] , 
        \nScanOut32[13] , \nScanOut32[12] , \nScanOut32[11] , \nScanOut32[10] , 
        \nScanOut32[9] , \nScanOut32[8] , \nScanOut32[7] , \nScanOut32[6] , 
        \nScanOut32[5] , \nScanOut32[4] , \nScanOut32[3] , \nScanOut32[2] , 
        \nScanOut32[1] , \nScanOut32[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_32[31] , 
        \nOut0_32[30] , \nOut0_32[29] , \nOut0_32[28] , \nOut0_32[27] , 
        \nOut0_32[26] , \nOut0_32[25] , \nOut0_32[24] , \nOut0_32[23] , 
        \nOut0_32[22] , \nOut0_32[21] , \nOut0_32[20] , \nOut0_32[19] , 
        \nOut0_32[18] , \nOut0_32[17] , \nOut0_32[16] , \nOut0_32[15] , 
        \nOut0_32[14] , \nOut0_32[13] , \nOut0_32[12] , \nOut0_32[11] , 
        \nOut0_32[10] , \nOut0_32[9] , \nOut0_32[8] , \nOut0_32[7] , 
        \nOut0_32[6] , \nOut0_32[5] , \nOut0_32[4] , \nOut0_32[3] , 
        \nOut0_32[2] , \nOut0_32[1] , \nOut0_32[0] }), .NORTH_EDGE({
        \nOut0_31[31] , \nOut0_31[30] , \nOut0_31[29] , \nOut0_31[28] , 
        \nOut0_31[27] , \nOut0_31[26] , \nOut0_31[25] , \nOut0_31[24] , 
        \nOut0_31[23] , \nOut0_31[22] , \nOut0_31[21] , \nOut0_31[20] , 
        \nOut0_31[19] , \nOut0_31[18] , \nOut0_31[17] , \nOut0_31[16] , 
        \nOut0_31[15] , \nOut0_31[14] , \nOut0_31[13] , \nOut0_31[12] , 
        \nOut0_31[11] , \nOut0_31[10] , \nOut0_31[9] , \nOut0_31[8] , 
        \nOut0_31[7] , \nOut0_31[6] , \nOut0_31[5] , \nOut0_31[4] , 
        \nOut0_31[3] , \nOut0_31[2] , \nOut0_31[1] , \nOut0_31[0] }), 
        .SOUTH_EDGE({\nOut0_33[31] , \nOut0_33[30] , \nOut0_33[29] , 
        \nOut0_33[28] , \nOut0_33[27] , \nOut0_33[26] , \nOut0_33[25] , 
        \nOut0_33[24] , \nOut0_33[23] , \nOut0_33[22] , \nOut0_33[21] , 
        \nOut0_33[20] , \nOut0_33[19] , \nOut0_33[18] , \nOut0_33[17] , 
        \nOut0_33[16] , \nOut0_33[15] , \nOut0_33[14] , \nOut0_33[13] , 
        \nOut0_33[12] , \nOut0_33[11] , \nOut0_33[10] , \nOut0_33[9] , 
        \nOut0_33[8] , \nOut0_33[7] , \nOut0_33[6] , \nOut0_33[5] , 
        \nOut0_33[4] , \nOut0_33[3] , \nOut0_33[2] , \nOut0_33[1] , 
        \nOut0_33[0] }), .EAST_EDGE(\nOut1_32[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_31[31] ), .SE_EDGE(
        \nOut1_33[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_47 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut48[31] , \nScanOut48[30] , \nScanOut48[29] , 
        \nScanOut48[28] , \nScanOut48[27] , \nScanOut48[26] , \nScanOut48[25] , 
        \nScanOut48[24] , \nScanOut48[23] , \nScanOut48[22] , \nScanOut48[21] , 
        \nScanOut48[20] , \nScanOut48[19] , \nScanOut48[18] , \nScanOut48[17] , 
        \nScanOut48[16] , \nScanOut48[15] , \nScanOut48[14] , \nScanOut48[13] , 
        \nScanOut48[12] , \nScanOut48[11] , \nScanOut48[10] , \nScanOut48[9] , 
        \nScanOut48[8] , \nScanOut48[7] , \nScanOut48[6] , \nScanOut48[5] , 
        \nScanOut48[4] , \nScanOut48[3] , \nScanOut48[2] , \nScanOut48[1] , 
        \nScanOut48[0] }), .ScanOut({\nScanOut47[31] , \nScanOut47[30] , 
        \nScanOut47[29] , \nScanOut47[28] , \nScanOut47[27] , \nScanOut47[26] , 
        \nScanOut47[25] , \nScanOut47[24] , \nScanOut47[23] , \nScanOut47[22] , 
        \nScanOut47[21] , \nScanOut47[20] , \nScanOut47[19] , \nScanOut47[18] , 
        \nScanOut47[17] , \nScanOut47[16] , \nScanOut47[15] , \nScanOut47[14] , 
        \nScanOut47[13] , \nScanOut47[12] , \nScanOut47[11] , \nScanOut47[10] , 
        \nScanOut47[9] , \nScanOut47[8] , \nScanOut47[7] , \nScanOut47[6] , 
        \nScanOut47[5] , \nScanOut47[4] , \nScanOut47[3] , \nScanOut47[2] , 
        \nScanOut47[1] , \nScanOut47[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_47[31] , 
        \nOut0_47[30] , \nOut0_47[29] , \nOut0_47[28] , \nOut0_47[27] , 
        \nOut0_47[26] , \nOut0_47[25] , \nOut0_47[24] , \nOut0_47[23] , 
        \nOut0_47[22] , \nOut0_47[21] , \nOut0_47[20] , \nOut0_47[19] , 
        \nOut0_47[18] , \nOut0_47[17] , \nOut0_47[16] , \nOut0_47[15] , 
        \nOut0_47[14] , \nOut0_47[13] , \nOut0_47[12] , \nOut0_47[11] , 
        \nOut0_47[10] , \nOut0_47[9] , \nOut0_47[8] , \nOut0_47[7] , 
        \nOut0_47[6] , \nOut0_47[5] , \nOut0_47[4] , \nOut0_47[3] , 
        \nOut0_47[2] , \nOut0_47[1] , \nOut0_47[0] }), .NORTH_EDGE({
        \nOut0_46[31] , \nOut0_46[30] , \nOut0_46[29] , \nOut0_46[28] , 
        \nOut0_46[27] , \nOut0_46[26] , \nOut0_46[25] , \nOut0_46[24] , 
        \nOut0_46[23] , \nOut0_46[22] , \nOut0_46[21] , \nOut0_46[20] , 
        \nOut0_46[19] , \nOut0_46[18] , \nOut0_46[17] , \nOut0_46[16] , 
        \nOut0_46[15] , \nOut0_46[14] , \nOut0_46[13] , \nOut0_46[12] , 
        \nOut0_46[11] , \nOut0_46[10] , \nOut0_46[9] , \nOut0_46[8] , 
        \nOut0_46[7] , \nOut0_46[6] , \nOut0_46[5] , \nOut0_46[4] , 
        \nOut0_46[3] , \nOut0_46[2] , \nOut0_46[1] , \nOut0_46[0] }), 
        .SOUTH_EDGE({\nOut0_48[31] , \nOut0_48[30] , \nOut0_48[29] , 
        \nOut0_48[28] , \nOut0_48[27] , \nOut0_48[26] , \nOut0_48[25] , 
        \nOut0_48[24] , \nOut0_48[23] , \nOut0_48[22] , \nOut0_48[21] , 
        \nOut0_48[20] , \nOut0_48[19] , \nOut0_48[18] , \nOut0_48[17] , 
        \nOut0_48[16] , \nOut0_48[15] , \nOut0_48[14] , \nOut0_48[13] , 
        \nOut0_48[12] , \nOut0_48[11] , \nOut0_48[10] , \nOut0_48[9] , 
        \nOut0_48[8] , \nOut0_48[7] , \nOut0_48[6] , \nOut0_48[5] , 
        \nOut0_48[4] , \nOut0_48[3] , \nOut0_48[2] , \nOut0_48[1] , 
        \nOut0_48[0] }), .EAST_EDGE(\nOut1_47[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_46[31] ), .SE_EDGE(
        \nOut1_48[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_85 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut86[31] , \nScanOut86[30] , \nScanOut86[29] , 
        \nScanOut86[28] , \nScanOut86[27] , \nScanOut86[26] , \nScanOut86[25] , 
        \nScanOut86[24] , \nScanOut86[23] , \nScanOut86[22] , \nScanOut86[21] , 
        \nScanOut86[20] , \nScanOut86[19] , \nScanOut86[18] , \nScanOut86[17] , 
        \nScanOut86[16] , \nScanOut86[15] , \nScanOut86[14] , \nScanOut86[13] , 
        \nScanOut86[12] , \nScanOut86[11] , \nScanOut86[10] , \nScanOut86[9] , 
        \nScanOut86[8] , \nScanOut86[7] , \nScanOut86[6] , \nScanOut86[5] , 
        \nScanOut86[4] , \nScanOut86[3] , \nScanOut86[2] , \nScanOut86[1] , 
        \nScanOut86[0] }), .ScanOut({\nScanOut85[31] , \nScanOut85[30] , 
        \nScanOut85[29] , \nScanOut85[28] , \nScanOut85[27] , \nScanOut85[26] , 
        \nScanOut85[25] , \nScanOut85[24] , \nScanOut85[23] , \nScanOut85[22] , 
        \nScanOut85[21] , \nScanOut85[20] , \nScanOut85[19] , \nScanOut85[18] , 
        \nScanOut85[17] , \nScanOut85[16] , \nScanOut85[15] , \nScanOut85[14] , 
        \nScanOut85[13] , \nScanOut85[12] , \nScanOut85[11] , \nScanOut85[10] , 
        \nScanOut85[9] , \nScanOut85[8] , \nScanOut85[7] , \nScanOut85[6] , 
        \nScanOut85[5] , \nScanOut85[4] , \nScanOut85[3] , \nScanOut85[2] , 
        \nScanOut85[1] , \nScanOut85[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_21[31] , 
        \nOut1_21[30] , \nOut1_21[29] , \nOut1_21[28] , \nOut1_21[27] , 
        \nOut1_21[26] , \nOut1_21[25] , \nOut1_21[24] , \nOut1_21[23] , 
        \nOut1_21[22] , \nOut1_21[21] , \nOut1_21[20] , \nOut1_21[19] , 
        \nOut1_21[18] , \nOut1_21[17] , \nOut1_21[16] , \nOut1_21[15] , 
        \nOut1_21[14] , \nOut1_21[13] , \nOut1_21[12] , \nOut1_21[11] , 
        \nOut1_21[10] , \nOut1_21[9] , \nOut1_21[8] , \nOut1_21[7] , 
        \nOut1_21[6] , \nOut1_21[5] , \nOut1_21[4] , \nOut1_21[3] , 
        \nOut1_21[2] , \nOut1_21[1] , \nOut1_21[0] }), .NORTH_EDGE({
        \nOut1_20[31] , \nOut1_20[30] , \nOut1_20[29] , \nOut1_20[28] , 
        \nOut1_20[27] , \nOut1_20[26] , \nOut1_20[25] , \nOut1_20[24] , 
        \nOut1_20[23] , \nOut1_20[22] , \nOut1_20[21] , \nOut1_20[20] , 
        \nOut1_20[19] , \nOut1_20[18] , \nOut1_20[17] , \nOut1_20[16] , 
        \nOut1_20[15] , \nOut1_20[14] , \nOut1_20[13] , \nOut1_20[12] , 
        \nOut1_20[11] , \nOut1_20[10] , \nOut1_20[9] , \nOut1_20[8] , 
        \nOut1_20[7] , \nOut1_20[6] , \nOut1_20[5] , \nOut1_20[4] , 
        \nOut1_20[3] , \nOut1_20[2] , \nOut1_20[1] , \nOut1_20[0] }), 
        .SOUTH_EDGE({\nOut1_22[31] , \nOut1_22[30] , \nOut1_22[29] , 
        \nOut1_22[28] , \nOut1_22[27] , \nOut1_22[26] , \nOut1_22[25] , 
        \nOut1_22[24] , \nOut1_22[23] , \nOut1_22[22] , \nOut1_22[21] , 
        \nOut1_22[20] , \nOut1_22[19] , \nOut1_22[18] , \nOut1_22[17] , 
        \nOut1_22[16] , \nOut1_22[15] , \nOut1_22[14] , \nOut1_22[13] , 
        \nOut1_22[12] , \nOut1_22[11] , \nOut1_22[10] , \nOut1_22[9] , 
        \nOut1_22[8] , \nOut1_22[7] , \nOut1_22[6] , \nOut1_22[5] , 
        \nOut1_22[4] , \nOut1_22[3] , \nOut1_22[2] , \nOut1_22[1] , 
        \nOut1_22[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_21[0] ), 
        .NW_EDGE(\nOut0_20[0] ), .SW_EDGE(\nOut0_22[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_60 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut61[31] , \nScanOut61[30] , \nScanOut61[29] , 
        \nScanOut61[28] , \nScanOut61[27] , \nScanOut61[26] , \nScanOut61[25] , 
        \nScanOut61[24] , \nScanOut61[23] , \nScanOut61[22] , \nScanOut61[21] , 
        \nScanOut61[20] , \nScanOut61[19] , \nScanOut61[18] , \nScanOut61[17] , 
        \nScanOut61[16] , \nScanOut61[15] , \nScanOut61[14] , \nScanOut61[13] , 
        \nScanOut61[12] , \nScanOut61[11] , \nScanOut61[10] , \nScanOut61[9] , 
        \nScanOut61[8] , \nScanOut61[7] , \nScanOut61[6] , \nScanOut61[5] , 
        \nScanOut61[4] , \nScanOut61[3] , \nScanOut61[2] , \nScanOut61[1] , 
        \nScanOut61[0] }), .ScanOut({\nScanOut60[31] , \nScanOut60[30] , 
        \nScanOut60[29] , \nScanOut60[28] , \nScanOut60[27] , \nScanOut60[26] , 
        \nScanOut60[25] , \nScanOut60[24] , \nScanOut60[23] , \nScanOut60[22] , 
        \nScanOut60[21] , \nScanOut60[20] , \nScanOut60[19] , \nScanOut60[18] , 
        \nScanOut60[17] , \nScanOut60[16] , \nScanOut60[15] , \nScanOut60[14] , 
        \nScanOut60[13] , \nScanOut60[12] , \nScanOut60[11] , \nScanOut60[10] , 
        \nScanOut60[9] , \nScanOut60[8] , \nScanOut60[7] , \nScanOut60[6] , 
        \nScanOut60[5] , \nScanOut60[4] , \nScanOut60[3] , \nScanOut60[2] , 
        \nScanOut60[1] , \nScanOut60[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_60[31] , 
        \nOut0_60[30] , \nOut0_60[29] , \nOut0_60[28] , \nOut0_60[27] , 
        \nOut0_60[26] , \nOut0_60[25] , \nOut0_60[24] , \nOut0_60[23] , 
        \nOut0_60[22] , \nOut0_60[21] , \nOut0_60[20] , \nOut0_60[19] , 
        \nOut0_60[18] , \nOut0_60[17] , \nOut0_60[16] , \nOut0_60[15] , 
        \nOut0_60[14] , \nOut0_60[13] , \nOut0_60[12] , \nOut0_60[11] , 
        \nOut0_60[10] , \nOut0_60[9] , \nOut0_60[8] , \nOut0_60[7] , 
        \nOut0_60[6] , \nOut0_60[5] , \nOut0_60[4] , \nOut0_60[3] , 
        \nOut0_60[2] , \nOut0_60[1] , \nOut0_60[0] }), .NORTH_EDGE({
        \nOut0_59[31] , \nOut0_59[30] , \nOut0_59[29] , \nOut0_59[28] , 
        \nOut0_59[27] , \nOut0_59[26] , \nOut0_59[25] , \nOut0_59[24] , 
        \nOut0_59[23] , \nOut0_59[22] , \nOut0_59[21] , \nOut0_59[20] , 
        \nOut0_59[19] , \nOut0_59[18] , \nOut0_59[17] , \nOut0_59[16] , 
        \nOut0_59[15] , \nOut0_59[14] , \nOut0_59[13] , \nOut0_59[12] , 
        \nOut0_59[11] , \nOut0_59[10] , \nOut0_59[9] , \nOut0_59[8] , 
        \nOut0_59[7] , \nOut0_59[6] , \nOut0_59[5] , \nOut0_59[4] , 
        \nOut0_59[3] , \nOut0_59[2] , \nOut0_59[1] , \nOut0_59[0] }), 
        .SOUTH_EDGE({\nOut0_61[31] , \nOut0_61[30] , \nOut0_61[29] , 
        \nOut0_61[28] , \nOut0_61[27] , \nOut0_61[26] , \nOut0_61[25] , 
        \nOut0_61[24] , \nOut0_61[23] , \nOut0_61[22] , \nOut0_61[21] , 
        \nOut0_61[20] , \nOut0_61[19] , \nOut0_61[18] , \nOut0_61[17] , 
        \nOut0_61[16] , \nOut0_61[15] , \nOut0_61[14] , \nOut0_61[13] , 
        \nOut0_61[12] , \nOut0_61[11] , \nOut0_61[10] , \nOut0_61[9] , 
        \nOut0_61[8] , \nOut0_61[7] , \nOut0_61[6] , \nOut0_61[5] , 
        \nOut0_61[4] , \nOut0_61[3] , \nOut0_61[2] , \nOut0_61[1] , 
        \nOut0_61[0] }), .EAST_EDGE(\nOut1_60[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_59[31] ), .SE_EDGE(
        \nOut1_61[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_111 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut112[31] , \nScanOut112[30] , \nScanOut112[29] , 
        \nScanOut112[28] , \nScanOut112[27] , \nScanOut112[26] , 
        \nScanOut112[25] , \nScanOut112[24] , \nScanOut112[23] , 
        \nScanOut112[22] , \nScanOut112[21] , \nScanOut112[20] , 
        \nScanOut112[19] , \nScanOut112[18] , \nScanOut112[17] , 
        \nScanOut112[16] , \nScanOut112[15] , \nScanOut112[14] , 
        \nScanOut112[13] , \nScanOut112[12] , \nScanOut112[11] , 
        \nScanOut112[10] , \nScanOut112[9] , \nScanOut112[8] , 
        \nScanOut112[7] , \nScanOut112[6] , \nScanOut112[5] , \nScanOut112[4] , 
        \nScanOut112[3] , \nScanOut112[2] , \nScanOut112[1] , \nScanOut112[0] 
        }), .ScanOut({\nScanOut111[31] , \nScanOut111[30] , \nScanOut111[29] , 
        \nScanOut111[28] , \nScanOut111[27] , \nScanOut111[26] , 
        \nScanOut111[25] , \nScanOut111[24] , \nScanOut111[23] , 
        \nScanOut111[22] , \nScanOut111[21] , \nScanOut111[20] , 
        \nScanOut111[19] , \nScanOut111[18] , \nScanOut111[17] , 
        \nScanOut111[16] , \nScanOut111[15] , \nScanOut111[14] , 
        \nScanOut111[13] , \nScanOut111[12] , \nScanOut111[11] , 
        \nScanOut111[10] , \nScanOut111[9] , \nScanOut111[8] , 
        \nScanOut111[7] , \nScanOut111[6] , \nScanOut111[5] , \nScanOut111[4] , 
        \nScanOut111[3] , \nScanOut111[2] , \nScanOut111[1] , \nScanOut111[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_47[31] , \nOut1_47[30] , \nOut1_47[29] , 
        \nOut1_47[28] , \nOut1_47[27] , \nOut1_47[26] , \nOut1_47[25] , 
        \nOut1_47[24] , \nOut1_47[23] , \nOut1_47[22] , \nOut1_47[21] , 
        \nOut1_47[20] , \nOut1_47[19] , \nOut1_47[18] , \nOut1_47[17] , 
        \nOut1_47[16] , \nOut1_47[15] , \nOut1_47[14] , \nOut1_47[13] , 
        \nOut1_47[12] , \nOut1_47[11] , \nOut1_47[10] , \nOut1_47[9] , 
        \nOut1_47[8] , \nOut1_47[7] , \nOut1_47[6] , \nOut1_47[5] , 
        \nOut1_47[4] , \nOut1_47[3] , \nOut1_47[2] , \nOut1_47[1] , 
        \nOut1_47[0] }), .NORTH_EDGE({\nOut1_46[31] , \nOut1_46[30] , 
        \nOut1_46[29] , \nOut1_46[28] , \nOut1_46[27] , \nOut1_46[26] , 
        \nOut1_46[25] , \nOut1_46[24] , \nOut1_46[23] , \nOut1_46[22] , 
        \nOut1_46[21] , \nOut1_46[20] , \nOut1_46[19] , \nOut1_46[18] , 
        \nOut1_46[17] , \nOut1_46[16] , \nOut1_46[15] , \nOut1_46[14] , 
        \nOut1_46[13] , \nOut1_46[12] , \nOut1_46[11] , \nOut1_46[10] , 
        \nOut1_46[9] , \nOut1_46[8] , \nOut1_46[7] , \nOut1_46[6] , 
        \nOut1_46[5] , \nOut1_46[4] , \nOut1_46[3] , \nOut1_46[2] , 
        \nOut1_46[1] , \nOut1_46[0] }), .SOUTH_EDGE({\nOut1_48[31] , 
        \nOut1_48[30] , \nOut1_48[29] , \nOut1_48[28] , \nOut1_48[27] , 
        \nOut1_48[26] , \nOut1_48[25] , \nOut1_48[24] , \nOut1_48[23] , 
        \nOut1_48[22] , \nOut1_48[21] , \nOut1_48[20] , \nOut1_48[19] , 
        \nOut1_48[18] , \nOut1_48[17] , \nOut1_48[16] , \nOut1_48[15] , 
        \nOut1_48[14] , \nOut1_48[13] , \nOut1_48[12] , \nOut1_48[11] , 
        \nOut1_48[10] , \nOut1_48[9] , \nOut1_48[8] , \nOut1_48[7] , 
        \nOut1_48[6] , \nOut1_48[5] , \nOut1_48[4] , \nOut1_48[3] , 
        \nOut1_48[2] , \nOut1_48[1] , \nOut1_48[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_47[0] ), .NW_EDGE(\nOut0_46[0] ), .SW_EDGE(
        \nOut0_48[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_39 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut40[31] , \nScanOut40[30] , \nScanOut40[29] , 
        \nScanOut40[28] , \nScanOut40[27] , \nScanOut40[26] , \nScanOut40[25] , 
        \nScanOut40[24] , \nScanOut40[23] , \nScanOut40[22] , \nScanOut40[21] , 
        \nScanOut40[20] , \nScanOut40[19] , \nScanOut40[18] , \nScanOut40[17] , 
        \nScanOut40[16] , \nScanOut40[15] , \nScanOut40[14] , \nScanOut40[13] , 
        \nScanOut40[12] , \nScanOut40[11] , \nScanOut40[10] , \nScanOut40[9] , 
        \nScanOut40[8] , \nScanOut40[7] , \nScanOut40[6] , \nScanOut40[5] , 
        \nScanOut40[4] , \nScanOut40[3] , \nScanOut40[2] , \nScanOut40[1] , 
        \nScanOut40[0] }), .ScanOut({\nScanOut39[31] , \nScanOut39[30] , 
        \nScanOut39[29] , \nScanOut39[28] , \nScanOut39[27] , \nScanOut39[26] , 
        \nScanOut39[25] , \nScanOut39[24] , \nScanOut39[23] , \nScanOut39[22] , 
        \nScanOut39[21] , \nScanOut39[20] , \nScanOut39[19] , \nScanOut39[18] , 
        \nScanOut39[17] , \nScanOut39[16] , \nScanOut39[15] , \nScanOut39[14] , 
        \nScanOut39[13] , \nScanOut39[12] , \nScanOut39[11] , \nScanOut39[10] , 
        \nScanOut39[9] , \nScanOut39[8] , \nScanOut39[7] , \nScanOut39[6] , 
        \nScanOut39[5] , \nScanOut39[4] , \nScanOut39[3] , \nScanOut39[2] , 
        \nScanOut39[1] , \nScanOut39[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_39[31] , 
        \nOut0_39[30] , \nOut0_39[29] , \nOut0_39[28] , \nOut0_39[27] , 
        \nOut0_39[26] , \nOut0_39[25] , \nOut0_39[24] , \nOut0_39[23] , 
        \nOut0_39[22] , \nOut0_39[21] , \nOut0_39[20] , \nOut0_39[19] , 
        \nOut0_39[18] , \nOut0_39[17] , \nOut0_39[16] , \nOut0_39[15] , 
        \nOut0_39[14] , \nOut0_39[13] , \nOut0_39[12] , \nOut0_39[11] , 
        \nOut0_39[10] , \nOut0_39[9] , \nOut0_39[8] , \nOut0_39[7] , 
        \nOut0_39[6] , \nOut0_39[5] , \nOut0_39[4] , \nOut0_39[3] , 
        \nOut0_39[2] , \nOut0_39[1] , \nOut0_39[0] }), .NORTH_EDGE({
        \nOut0_38[31] , \nOut0_38[30] , \nOut0_38[29] , \nOut0_38[28] , 
        \nOut0_38[27] , \nOut0_38[26] , \nOut0_38[25] , \nOut0_38[24] , 
        \nOut0_38[23] , \nOut0_38[22] , \nOut0_38[21] , \nOut0_38[20] , 
        \nOut0_38[19] , \nOut0_38[18] , \nOut0_38[17] , \nOut0_38[16] , 
        \nOut0_38[15] , \nOut0_38[14] , \nOut0_38[13] , \nOut0_38[12] , 
        \nOut0_38[11] , \nOut0_38[10] , \nOut0_38[9] , \nOut0_38[8] , 
        \nOut0_38[7] , \nOut0_38[6] , \nOut0_38[5] , \nOut0_38[4] , 
        \nOut0_38[3] , \nOut0_38[2] , \nOut0_38[1] , \nOut0_38[0] }), 
        .SOUTH_EDGE({\nOut0_40[31] , \nOut0_40[30] , \nOut0_40[29] , 
        \nOut0_40[28] , \nOut0_40[27] , \nOut0_40[26] , \nOut0_40[25] , 
        \nOut0_40[24] , \nOut0_40[23] , \nOut0_40[22] , \nOut0_40[21] , 
        \nOut0_40[20] , \nOut0_40[19] , \nOut0_40[18] , \nOut0_40[17] , 
        \nOut0_40[16] , \nOut0_40[15] , \nOut0_40[14] , \nOut0_40[13] , 
        \nOut0_40[12] , \nOut0_40[11] , \nOut0_40[10] , \nOut0_40[9] , 
        \nOut0_40[8] , \nOut0_40[7] , \nOut0_40[6] , \nOut0_40[5] , 
        \nOut0_40[4] , \nOut0_40[3] , \nOut0_40[2] , \nOut0_40[1] , 
        \nOut0_40[0] }), .EAST_EDGE(\nOut1_39[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_38[31] ), .SE_EDGE(
        \nOut1_40[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_95 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut96[31] , \nScanOut96[30] , \nScanOut96[29] , 
        \nScanOut96[28] , \nScanOut96[27] , \nScanOut96[26] , \nScanOut96[25] , 
        \nScanOut96[24] , \nScanOut96[23] , \nScanOut96[22] , \nScanOut96[21] , 
        \nScanOut96[20] , \nScanOut96[19] , \nScanOut96[18] , \nScanOut96[17] , 
        \nScanOut96[16] , \nScanOut96[15] , \nScanOut96[14] , \nScanOut96[13] , 
        \nScanOut96[12] , \nScanOut96[11] , \nScanOut96[10] , \nScanOut96[9] , 
        \nScanOut96[8] , \nScanOut96[7] , \nScanOut96[6] , \nScanOut96[5] , 
        \nScanOut96[4] , \nScanOut96[3] , \nScanOut96[2] , \nScanOut96[1] , 
        \nScanOut96[0] }), .ScanOut({\nScanOut95[31] , \nScanOut95[30] , 
        \nScanOut95[29] , \nScanOut95[28] , \nScanOut95[27] , \nScanOut95[26] , 
        \nScanOut95[25] , \nScanOut95[24] , \nScanOut95[23] , \nScanOut95[22] , 
        \nScanOut95[21] , \nScanOut95[20] , \nScanOut95[19] , \nScanOut95[18] , 
        \nScanOut95[17] , \nScanOut95[16] , \nScanOut95[15] , \nScanOut95[14] , 
        \nScanOut95[13] , \nScanOut95[12] , \nScanOut95[11] , \nScanOut95[10] , 
        \nScanOut95[9] , \nScanOut95[8] , \nScanOut95[7] , \nScanOut95[6] , 
        \nScanOut95[5] , \nScanOut95[4] , \nScanOut95[3] , \nScanOut95[2] , 
        \nScanOut95[1] , \nScanOut95[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_31[31] , 
        \nOut1_31[30] , \nOut1_31[29] , \nOut1_31[28] , \nOut1_31[27] , 
        \nOut1_31[26] , \nOut1_31[25] , \nOut1_31[24] , \nOut1_31[23] , 
        \nOut1_31[22] , \nOut1_31[21] , \nOut1_31[20] , \nOut1_31[19] , 
        \nOut1_31[18] , \nOut1_31[17] , \nOut1_31[16] , \nOut1_31[15] , 
        \nOut1_31[14] , \nOut1_31[13] , \nOut1_31[12] , \nOut1_31[11] , 
        \nOut1_31[10] , \nOut1_31[9] , \nOut1_31[8] , \nOut1_31[7] , 
        \nOut1_31[6] , \nOut1_31[5] , \nOut1_31[4] , \nOut1_31[3] , 
        \nOut1_31[2] , \nOut1_31[1] , \nOut1_31[0] }), .NORTH_EDGE({
        \nOut1_30[31] , \nOut1_30[30] , \nOut1_30[29] , \nOut1_30[28] , 
        \nOut1_30[27] , \nOut1_30[26] , \nOut1_30[25] , \nOut1_30[24] , 
        \nOut1_30[23] , \nOut1_30[22] , \nOut1_30[21] , \nOut1_30[20] , 
        \nOut1_30[19] , \nOut1_30[18] , \nOut1_30[17] , \nOut1_30[16] , 
        \nOut1_30[15] , \nOut1_30[14] , \nOut1_30[13] , \nOut1_30[12] , 
        \nOut1_30[11] , \nOut1_30[10] , \nOut1_30[9] , \nOut1_30[8] , 
        \nOut1_30[7] , \nOut1_30[6] , \nOut1_30[5] , \nOut1_30[4] , 
        \nOut1_30[3] , \nOut1_30[2] , \nOut1_30[1] , \nOut1_30[0] }), 
        .SOUTH_EDGE({\nOut1_32[31] , \nOut1_32[30] , \nOut1_32[29] , 
        \nOut1_32[28] , \nOut1_32[27] , \nOut1_32[26] , \nOut1_32[25] , 
        \nOut1_32[24] , \nOut1_32[23] , \nOut1_32[22] , \nOut1_32[21] , 
        \nOut1_32[20] , \nOut1_32[19] , \nOut1_32[18] , \nOut1_32[17] , 
        \nOut1_32[16] , \nOut1_32[15] , \nOut1_32[14] , \nOut1_32[13] , 
        \nOut1_32[12] , \nOut1_32[11] , \nOut1_32[10] , \nOut1_32[9] , 
        \nOut1_32[8] , \nOut1_32[7] , \nOut1_32[6] , \nOut1_32[5] , 
        \nOut1_32[4] , \nOut1_32[3] , \nOut1_32[2] , \nOut1_32[1] , 
        \nOut1_32[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_31[0] ), 
        .NW_EDGE(\nOut0_30[0] ), .SW_EDGE(\nOut0_32[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut2[31] , \nScanOut2[30] , \nScanOut2[29] , 
        \nScanOut2[28] , \nScanOut2[27] , \nScanOut2[26] , \nScanOut2[25] , 
        \nScanOut2[24] , \nScanOut2[23] , \nScanOut2[22] , \nScanOut2[21] , 
        \nScanOut2[20] , \nScanOut2[19] , \nScanOut2[18] , \nScanOut2[17] , 
        \nScanOut2[16] , \nScanOut2[15] , \nScanOut2[14] , \nScanOut2[13] , 
        \nScanOut2[12] , \nScanOut2[11] , \nScanOut2[10] , \nScanOut2[9] , 
        \nScanOut2[8] , \nScanOut2[7] , \nScanOut2[6] , \nScanOut2[5] , 
        \nScanOut2[4] , \nScanOut2[3] , \nScanOut2[2] , \nScanOut2[1] , 
        \nScanOut2[0] }), .ScanOut({\nScanOut1[31] , \nScanOut1[30] , 
        \nScanOut1[29] , \nScanOut1[28] , \nScanOut1[27] , \nScanOut1[26] , 
        \nScanOut1[25] , \nScanOut1[24] , \nScanOut1[23] , \nScanOut1[22] , 
        \nScanOut1[21] , \nScanOut1[20] , \nScanOut1[19] , \nScanOut1[18] , 
        \nScanOut1[17] , \nScanOut1[16] , \nScanOut1[15] , \nScanOut1[14] , 
        \nScanOut1[13] , \nScanOut1[12] , \nScanOut1[11] , \nScanOut1[10] , 
        \nScanOut1[9] , \nScanOut1[8] , \nScanOut1[7] , \nScanOut1[6] , 
        \nScanOut1[5] , \nScanOut1[4] , \nScanOut1[3] , \nScanOut1[2] , 
        \nScanOut1[1] , \nScanOut1[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_1[31] , 
        \nOut0_1[30] , \nOut0_1[29] , \nOut0_1[28] , \nOut0_1[27] , 
        \nOut0_1[26] , \nOut0_1[25] , \nOut0_1[24] , \nOut0_1[23] , 
        \nOut0_1[22] , \nOut0_1[21] , \nOut0_1[20] , \nOut0_1[19] , 
        \nOut0_1[18] , \nOut0_1[17] , \nOut0_1[16] , \nOut0_1[15] , 
        \nOut0_1[14] , \nOut0_1[13] , \nOut0_1[12] , \nOut0_1[11] , 
        \nOut0_1[10] , \nOut0_1[9] , \nOut0_1[8] , \nOut0_1[7] , \nOut0_1[6] , 
        \nOut0_1[5] , \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , 
        \nOut0_1[0] }), .NORTH_EDGE({\nOut0_0[31] , \nOut0_0[30] , 
        \nOut0_0[29] , \nOut0_0[28] , \nOut0_0[27] , \nOut0_0[26] , 
        \nOut0_0[25] , \nOut0_0[24] , \nOut0_0[23] , \nOut0_0[22] , 
        \nOut0_0[21] , \nOut0_0[20] , \nOut0_0[19] , \nOut0_0[18] , 
        \nOut0_0[17] , \nOut0_0[16] , \nOut0_0[15] , \nOut0_0[14] , 
        \nOut0_0[13] , \nOut0_0[12] , \nOut0_0[11] , \nOut0_0[10] , 
        \nOut0_0[9] , \nOut0_0[8] , \nOut0_0[7] , \nOut0_0[6] , \nOut0_0[5] , 
        \nOut0_0[4] , \nOut0_0[3] , \nOut0_0[2] , \nOut0_0[1] , \nOut0_0[0] }), 
        .SOUTH_EDGE({\nOut0_2[31] , \nOut0_2[30] , \nOut0_2[29] , 
        \nOut0_2[28] , \nOut0_2[27] , \nOut0_2[26] , \nOut0_2[25] , 
        \nOut0_2[24] , \nOut0_2[23] , \nOut0_2[22] , \nOut0_2[21] , 
        \nOut0_2[20] , \nOut0_2[19] , \nOut0_2[18] , \nOut0_2[17] , 
        \nOut0_2[16] , \nOut0_2[15] , \nOut0_2[14] , \nOut0_2[13] , 
        \nOut0_2[12] , \nOut0_2[11] , \nOut0_2[10] , \nOut0_2[9] , 
        \nOut0_2[8] , \nOut0_2[7] , \nOut0_2[6] , \nOut0_2[5] , \nOut0_2[4] , 
        \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , \nOut0_2[0] }), .EAST_EDGE(
        \nOut1_1[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_0[31] ), .SE_EDGE(\nOut1_2[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut7[31] , \nScanOut7[30] , \nScanOut7[29] , 
        \nScanOut7[28] , \nScanOut7[27] , \nScanOut7[26] , \nScanOut7[25] , 
        \nScanOut7[24] , \nScanOut7[23] , \nScanOut7[22] , \nScanOut7[21] , 
        \nScanOut7[20] , \nScanOut7[19] , \nScanOut7[18] , \nScanOut7[17] , 
        \nScanOut7[16] , \nScanOut7[15] , \nScanOut7[14] , \nScanOut7[13] , 
        \nScanOut7[12] , \nScanOut7[11] , \nScanOut7[10] , \nScanOut7[9] , 
        \nScanOut7[8] , \nScanOut7[7] , \nScanOut7[6] , \nScanOut7[5] , 
        \nScanOut7[4] , \nScanOut7[3] , \nScanOut7[2] , \nScanOut7[1] , 
        \nScanOut7[0] }), .ScanOut({\nScanOut6[31] , \nScanOut6[30] , 
        \nScanOut6[29] , \nScanOut6[28] , \nScanOut6[27] , \nScanOut6[26] , 
        \nScanOut6[25] , \nScanOut6[24] , \nScanOut6[23] , \nScanOut6[22] , 
        \nScanOut6[21] , \nScanOut6[20] , \nScanOut6[19] , \nScanOut6[18] , 
        \nScanOut6[17] , \nScanOut6[16] , \nScanOut6[15] , \nScanOut6[14] , 
        \nScanOut6[13] , \nScanOut6[12] , \nScanOut6[11] , \nScanOut6[10] , 
        \nScanOut6[9] , \nScanOut6[8] , \nScanOut6[7] , \nScanOut6[6] , 
        \nScanOut6[5] , \nScanOut6[4] , \nScanOut6[3] , \nScanOut6[2] , 
        \nScanOut6[1] , \nScanOut6[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_6[31] , 
        \nOut0_6[30] , \nOut0_6[29] , \nOut0_6[28] , \nOut0_6[27] , 
        \nOut0_6[26] , \nOut0_6[25] , \nOut0_6[24] , \nOut0_6[23] , 
        \nOut0_6[22] , \nOut0_6[21] , \nOut0_6[20] , \nOut0_6[19] , 
        \nOut0_6[18] , \nOut0_6[17] , \nOut0_6[16] , \nOut0_6[15] , 
        \nOut0_6[14] , \nOut0_6[13] , \nOut0_6[12] , \nOut0_6[11] , 
        \nOut0_6[10] , \nOut0_6[9] , \nOut0_6[8] , \nOut0_6[7] , \nOut0_6[6] , 
        \nOut0_6[5] , \nOut0_6[4] , \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , 
        \nOut0_6[0] }), .NORTH_EDGE({\nOut0_5[31] , \nOut0_5[30] , 
        \nOut0_5[29] , \nOut0_5[28] , \nOut0_5[27] , \nOut0_5[26] , 
        \nOut0_5[25] , \nOut0_5[24] , \nOut0_5[23] , \nOut0_5[22] , 
        \nOut0_5[21] , \nOut0_5[20] , \nOut0_5[19] , \nOut0_5[18] , 
        \nOut0_5[17] , \nOut0_5[16] , \nOut0_5[15] , \nOut0_5[14] , 
        \nOut0_5[13] , \nOut0_5[12] , \nOut0_5[11] , \nOut0_5[10] , 
        \nOut0_5[9] , \nOut0_5[8] , \nOut0_5[7] , \nOut0_5[6] , \nOut0_5[5] , 
        \nOut0_5[4] , \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , \nOut0_5[0] }), 
        .SOUTH_EDGE({\nOut0_7[31] , \nOut0_7[30] , \nOut0_7[29] , 
        \nOut0_7[28] , \nOut0_7[27] , \nOut0_7[26] , \nOut0_7[25] , 
        \nOut0_7[24] , \nOut0_7[23] , \nOut0_7[22] , \nOut0_7[21] , 
        \nOut0_7[20] , \nOut0_7[19] , \nOut0_7[18] , \nOut0_7[17] , 
        \nOut0_7[16] , \nOut0_7[15] , \nOut0_7[14] , \nOut0_7[13] , 
        \nOut0_7[12] , \nOut0_7[11] , \nOut0_7[10] , \nOut0_7[9] , 
        \nOut0_7[8] , \nOut0_7[7] , \nOut0_7[6] , \nOut0_7[5] , \nOut0_7[4] , 
        \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , \nOut0_7[0] }), .EAST_EDGE(
        \nOut1_6[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_5[31] ), .SE_EDGE(\nOut1_7[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut8[31] , \nScanOut8[30] , \nScanOut8[29] , 
        \nScanOut8[28] , \nScanOut8[27] , \nScanOut8[26] , \nScanOut8[25] , 
        \nScanOut8[24] , \nScanOut8[23] , \nScanOut8[22] , \nScanOut8[21] , 
        \nScanOut8[20] , \nScanOut8[19] , \nScanOut8[18] , \nScanOut8[17] , 
        \nScanOut8[16] , \nScanOut8[15] , \nScanOut8[14] , \nScanOut8[13] , 
        \nScanOut8[12] , \nScanOut8[11] , \nScanOut8[10] , \nScanOut8[9] , 
        \nScanOut8[8] , \nScanOut8[7] , \nScanOut8[6] , \nScanOut8[5] , 
        \nScanOut8[4] , \nScanOut8[3] , \nScanOut8[2] , \nScanOut8[1] , 
        \nScanOut8[0] }), .ScanOut({\nScanOut7[31] , \nScanOut7[30] , 
        \nScanOut7[29] , \nScanOut7[28] , \nScanOut7[27] , \nScanOut7[26] , 
        \nScanOut7[25] , \nScanOut7[24] , \nScanOut7[23] , \nScanOut7[22] , 
        \nScanOut7[21] , \nScanOut7[20] , \nScanOut7[19] , \nScanOut7[18] , 
        \nScanOut7[17] , \nScanOut7[16] , \nScanOut7[15] , \nScanOut7[14] , 
        \nScanOut7[13] , \nScanOut7[12] , \nScanOut7[11] , \nScanOut7[10] , 
        \nScanOut7[9] , \nScanOut7[8] , \nScanOut7[7] , \nScanOut7[6] , 
        \nScanOut7[5] , \nScanOut7[4] , \nScanOut7[3] , \nScanOut7[2] , 
        \nScanOut7[1] , \nScanOut7[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_7[31] , 
        \nOut0_7[30] , \nOut0_7[29] , \nOut0_7[28] , \nOut0_7[27] , 
        \nOut0_7[26] , \nOut0_7[25] , \nOut0_7[24] , \nOut0_7[23] , 
        \nOut0_7[22] , \nOut0_7[21] , \nOut0_7[20] , \nOut0_7[19] , 
        \nOut0_7[18] , \nOut0_7[17] , \nOut0_7[16] , \nOut0_7[15] , 
        \nOut0_7[14] , \nOut0_7[13] , \nOut0_7[12] , \nOut0_7[11] , 
        \nOut0_7[10] , \nOut0_7[9] , \nOut0_7[8] , \nOut0_7[7] , \nOut0_7[6] , 
        \nOut0_7[5] , \nOut0_7[4] , \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , 
        \nOut0_7[0] }), .NORTH_EDGE({\nOut0_6[31] , \nOut0_6[30] , 
        \nOut0_6[29] , \nOut0_6[28] , \nOut0_6[27] , \nOut0_6[26] , 
        \nOut0_6[25] , \nOut0_6[24] , \nOut0_6[23] , \nOut0_6[22] , 
        \nOut0_6[21] , \nOut0_6[20] , \nOut0_6[19] , \nOut0_6[18] , 
        \nOut0_6[17] , \nOut0_6[16] , \nOut0_6[15] , \nOut0_6[14] , 
        \nOut0_6[13] , \nOut0_6[12] , \nOut0_6[11] , \nOut0_6[10] , 
        \nOut0_6[9] , \nOut0_6[8] , \nOut0_6[7] , \nOut0_6[6] , \nOut0_6[5] , 
        \nOut0_6[4] , \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , \nOut0_6[0] }), 
        .SOUTH_EDGE({\nOut0_8[31] , \nOut0_8[30] , \nOut0_8[29] , 
        \nOut0_8[28] , \nOut0_8[27] , \nOut0_8[26] , \nOut0_8[25] , 
        \nOut0_8[24] , \nOut0_8[23] , \nOut0_8[22] , \nOut0_8[21] , 
        \nOut0_8[20] , \nOut0_8[19] , \nOut0_8[18] , \nOut0_8[17] , 
        \nOut0_8[16] , \nOut0_8[15] , \nOut0_8[14] , \nOut0_8[13] , 
        \nOut0_8[12] , \nOut0_8[11] , \nOut0_8[10] , \nOut0_8[9] , 
        \nOut0_8[8] , \nOut0_8[7] , \nOut0_8[6] , \nOut0_8[5] , \nOut0_8[4] , 
        \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , \nOut0_8[0] }), .EAST_EDGE(
        \nOut1_7[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_6[31] ), .SE_EDGE(\nOut1_8[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut10[31] , \nScanOut10[30] , \nScanOut10[29] , 
        \nScanOut10[28] , \nScanOut10[27] , \nScanOut10[26] , \nScanOut10[25] , 
        \nScanOut10[24] , \nScanOut10[23] , \nScanOut10[22] , \nScanOut10[21] , 
        \nScanOut10[20] , \nScanOut10[19] , \nScanOut10[18] , \nScanOut10[17] , 
        \nScanOut10[16] , \nScanOut10[15] , \nScanOut10[14] , \nScanOut10[13] , 
        \nScanOut10[12] , \nScanOut10[11] , \nScanOut10[10] , \nScanOut10[9] , 
        \nScanOut10[8] , \nScanOut10[7] , \nScanOut10[6] , \nScanOut10[5] , 
        \nScanOut10[4] , \nScanOut10[3] , \nScanOut10[2] , \nScanOut10[1] , 
        \nScanOut10[0] }), .ScanOut({\nScanOut9[31] , \nScanOut9[30] , 
        \nScanOut9[29] , \nScanOut9[28] , \nScanOut9[27] , \nScanOut9[26] , 
        \nScanOut9[25] , \nScanOut9[24] , \nScanOut9[23] , \nScanOut9[22] , 
        \nScanOut9[21] , \nScanOut9[20] , \nScanOut9[19] , \nScanOut9[18] , 
        \nScanOut9[17] , \nScanOut9[16] , \nScanOut9[15] , \nScanOut9[14] , 
        \nScanOut9[13] , \nScanOut9[12] , \nScanOut9[11] , \nScanOut9[10] , 
        \nScanOut9[9] , \nScanOut9[8] , \nScanOut9[7] , \nScanOut9[6] , 
        \nScanOut9[5] , \nScanOut9[4] , \nScanOut9[3] , \nScanOut9[2] , 
        \nScanOut9[1] , \nScanOut9[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_9[31] , 
        \nOut0_9[30] , \nOut0_9[29] , \nOut0_9[28] , \nOut0_9[27] , 
        \nOut0_9[26] , \nOut0_9[25] , \nOut0_9[24] , \nOut0_9[23] , 
        \nOut0_9[22] , \nOut0_9[21] , \nOut0_9[20] , \nOut0_9[19] , 
        \nOut0_9[18] , \nOut0_9[17] , \nOut0_9[16] , \nOut0_9[15] , 
        \nOut0_9[14] , \nOut0_9[13] , \nOut0_9[12] , \nOut0_9[11] , 
        \nOut0_9[10] , \nOut0_9[9] , \nOut0_9[8] , \nOut0_9[7] , \nOut0_9[6] , 
        \nOut0_9[5] , \nOut0_9[4] , \nOut0_9[3] , \nOut0_9[2] , \nOut0_9[1] , 
        \nOut0_9[0] }), .NORTH_EDGE({\nOut0_8[31] , \nOut0_8[30] , 
        \nOut0_8[29] , \nOut0_8[28] , \nOut0_8[27] , \nOut0_8[26] , 
        \nOut0_8[25] , \nOut0_8[24] , \nOut0_8[23] , \nOut0_8[22] , 
        \nOut0_8[21] , \nOut0_8[20] , \nOut0_8[19] , \nOut0_8[18] , 
        \nOut0_8[17] , \nOut0_8[16] , \nOut0_8[15] , \nOut0_8[14] , 
        \nOut0_8[13] , \nOut0_8[12] , \nOut0_8[11] , \nOut0_8[10] , 
        \nOut0_8[9] , \nOut0_8[8] , \nOut0_8[7] , \nOut0_8[6] , \nOut0_8[5] , 
        \nOut0_8[4] , \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , \nOut0_8[0] }), 
        .SOUTH_EDGE({\nOut0_10[31] , \nOut0_10[30] , \nOut0_10[29] , 
        \nOut0_10[28] , \nOut0_10[27] , \nOut0_10[26] , \nOut0_10[25] , 
        \nOut0_10[24] , \nOut0_10[23] , \nOut0_10[22] , \nOut0_10[21] , 
        \nOut0_10[20] , \nOut0_10[19] , \nOut0_10[18] , \nOut0_10[17] , 
        \nOut0_10[16] , \nOut0_10[15] , \nOut0_10[14] , \nOut0_10[13] , 
        \nOut0_10[12] , \nOut0_10[11] , \nOut0_10[10] , \nOut0_10[9] , 
        \nOut0_10[8] , \nOut0_10[7] , \nOut0_10[6] , \nOut0_10[5] , 
        \nOut0_10[4] , \nOut0_10[3] , \nOut0_10[2] , \nOut0_10[1] , 
        \nOut0_10[0] }), .EAST_EDGE(\nOut1_9[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_8[31] ), .SE_EDGE(
        \nOut1_10[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_17 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut18[31] , \nScanOut18[30] , \nScanOut18[29] , 
        \nScanOut18[28] , \nScanOut18[27] , \nScanOut18[26] , \nScanOut18[25] , 
        \nScanOut18[24] , \nScanOut18[23] , \nScanOut18[22] , \nScanOut18[21] , 
        \nScanOut18[20] , \nScanOut18[19] , \nScanOut18[18] , \nScanOut18[17] , 
        \nScanOut18[16] , \nScanOut18[15] , \nScanOut18[14] , \nScanOut18[13] , 
        \nScanOut18[12] , \nScanOut18[11] , \nScanOut18[10] , \nScanOut18[9] , 
        \nScanOut18[8] , \nScanOut18[7] , \nScanOut18[6] , \nScanOut18[5] , 
        \nScanOut18[4] , \nScanOut18[3] , \nScanOut18[2] , \nScanOut18[1] , 
        \nScanOut18[0] }), .ScanOut({\nScanOut17[31] , \nScanOut17[30] , 
        \nScanOut17[29] , \nScanOut17[28] , \nScanOut17[27] , \nScanOut17[26] , 
        \nScanOut17[25] , \nScanOut17[24] , \nScanOut17[23] , \nScanOut17[22] , 
        \nScanOut17[21] , \nScanOut17[20] , \nScanOut17[19] , \nScanOut17[18] , 
        \nScanOut17[17] , \nScanOut17[16] , \nScanOut17[15] , \nScanOut17[14] , 
        \nScanOut17[13] , \nScanOut17[12] , \nScanOut17[11] , \nScanOut17[10] , 
        \nScanOut17[9] , \nScanOut17[8] , \nScanOut17[7] , \nScanOut17[6] , 
        \nScanOut17[5] , \nScanOut17[4] , \nScanOut17[3] , \nScanOut17[2] , 
        \nScanOut17[1] , \nScanOut17[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_17[31] , 
        \nOut0_17[30] , \nOut0_17[29] , \nOut0_17[28] , \nOut0_17[27] , 
        \nOut0_17[26] , \nOut0_17[25] , \nOut0_17[24] , \nOut0_17[23] , 
        \nOut0_17[22] , \nOut0_17[21] , \nOut0_17[20] , \nOut0_17[19] , 
        \nOut0_17[18] , \nOut0_17[17] , \nOut0_17[16] , \nOut0_17[15] , 
        \nOut0_17[14] , \nOut0_17[13] , \nOut0_17[12] , \nOut0_17[11] , 
        \nOut0_17[10] , \nOut0_17[9] , \nOut0_17[8] , \nOut0_17[7] , 
        \nOut0_17[6] , \nOut0_17[5] , \nOut0_17[4] , \nOut0_17[3] , 
        \nOut0_17[2] , \nOut0_17[1] , \nOut0_17[0] }), .NORTH_EDGE({
        \nOut0_16[31] , \nOut0_16[30] , \nOut0_16[29] , \nOut0_16[28] , 
        \nOut0_16[27] , \nOut0_16[26] , \nOut0_16[25] , \nOut0_16[24] , 
        \nOut0_16[23] , \nOut0_16[22] , \nOut0_16[21] , \nOut0_16[20] , 
        \nOut0_16[19] , \nOut0_16[18] , \nOut0_16[17] , \nOut0_16[16] , 
        \nOut0_16[15] , \nOut0_16[14] , \nOut0_16[13] , \nOut0_16[12] , 
        \nOut0_16[11] , \nOut0_16[10] , \nOut0_16[9] , \nOut0_16[8] , 
        \nOut0_16[7] , \nOut0_16[6] , \nOut0_16[5] , \nOut0_16[4] , 
        \nOut0_16[3] , \nOut0_16[2] , \nOut0_16[1] , \nOut0_16[0] }), 
        .SOUTH_EDGE({\nOut0_18[31] , \nOut0_18[30] , \nOut0_18[29] , 
        \nOut0_18[28] , \nOut0_18[27] , \nOut0_18[26] , \nOut0_18[25] , 
        \nOut0_18[24] , \nOut0_18[23] , \nOut0_18[22] , \nOut0_18[21] , 
        \nOut0_18[20] , \nOut0_18[19] , \nOut0_18[18] , \nOut0_18[17] , 
        \nOut0_18[16] , \nOut0_18[15] , \nOut0_18[14] , \nOut0_18[13] , 
        \nOut0_18[12] , \nOut0_18[11] , \nOut0_18[10] , \nOut0_18[9] , 
        \nOut0_18[8] , \nOut0_18[7] , \nOut0_18[6] , \nOut0_18[5] , 
        \nOut0_18[4] , \nOut0_18[3] , \nOut0_18[2] , \nOut0_18[1] , 
        \nOut0_18[0] }), .EAST_EDGE(\nOut1_17[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_16[31] ), .SE_EDGE(
        \nOut1_18[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_22 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut23[31] , \nScanOut23[30] , \nScanOut23[29] , 
        \nScanOut23[28] , \nScanOut23[27] , \nScanOut23[26] , \nScanOut23[25] , 
        \nScanOut23[24] , \nScanOut23[23] , \nScanOut23[22] , \nScanOut23[21] , 
        \nScanOut23[20] , \nScanOut23[19] , \nScanOut23[18] , \nScanOut23[17] , 
        \nScanOut23[16] , \nScanOut23[15] , \nScanOut23[14] , \nScanOut23[13] , 
        \nScanOut23[12] , \nScanOut23[11] , \nScanOut23[10] , \nScanOut23[9] , 
        \nScanOut23[8] , \nScanOut23[7] , \nScanOut23[6] , \nScanOut23[5] , 
        \nScanOut23[4] , \nScanOut23[3] , \nScanOut23[2] , \nScanOut23[1] , 
        \nScanOut23[0] }), .ScanOut({\nScanOut22[31] , \nScanOut22[30] , 
        \nScanOut22[29] , \nScanOut22[28] , \nScanOut22[27] , \nScanOut22[26] , 
        \nScanOut22[25] , \nScanOut22[24] , \nScanOut22[23] , \nScanOut22[22] , 
        \nScanOut22[21] , \nScanOut22[20] , \nScanOut22[19] , \nScanOut22[18] , 
        \nScanOut22[17] , \nScanOut22[16] , \nScanOut22[15] , \nScanOut22[14] , 
        \nScanOut22[13] , \nScanOut22[12] , \nScanOut22[11] , \nScanOut22[10] , 
        \nScanOut22[9] , \nScanOut22[8] , \nScanOut22[7] , \nScanOut22[6] , 
        \nScanOut22[5] , \nScanOut22[4] , \nScanOut22[3] , \nScanOut22[2] , 
        \nScanOut22[1] , \nScanOut22[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_22[31] , 
        \nOut0_22[30] , \nOut0_22[29] , \nOut0_22[28] , \nOut0_22[27] , 
        \nOut0_22[26] , \nOut0_22[25] , \nOut0_22[24] , \nOut0_22[23] , 
        \nOut0_22[22] , \nOut0_22[21] , \nOut0_22[20] , \nOut0_22[19] , 
        \nOut0_22[18] , \nOut0_22[17] , \nOut0_22[16] , \nOut0_22[15] , 
        \nOut0_22[14] , \nOut0_22[13] , \nOut0_22[12] , \nOut0_22[11] , 
        \nOut0_22[10] , \nOut0_22[9] , \nOut0_22[8] , \nOut0_22[7] , 
        \nOut0_22[6] , \nOut0_22[5] , \nOut0_22[4] , \nOut0_22[3] , 
        \nOut0_22[2] , \nOut0_22[1] , \nOut0_22[0] }), .NORTH_EDGE({
        \nOut0_21[31] , \nOut0_21[30] , \nOut0_21[29] , \nOut0_21[28] , 
        \nOut0_21[27] , \nOut0_21[26] , \nOut0_21[25] , \nOut0_21[24] , 
        \nOut0_21[23] , \nOut0_21[22] , \nOut0_21[21] , \nOut0_21[20] , 
        \nOut0_21[19] , \nOut0_21[18] , \nOut0_21[17] , \nOut0_21[16] , 
        \nOut0_21[15] , \nOut0_21[14] , \nOut0_21[13] , \nOut0_21[12] , 
        \nOut0_21[11] , \nOut0_21[10] , \nOut0_21[9] , \nOut0_21[8] , 
        \nOut0_21[7] , \nOut0_21[6] , \nOut0_21[5] , \nOut0_21[4] , 
        \nOut0_21[3] , \nOut0_21[2] , \nOut0_21[1] , \nOut0_21[0] }), 
        .SOUTH_EDGE({\nOut0_23[31] , \nOut0_23[30] , \nOut0_23[29] , 
        \nOut0_23[28] , \nOut0_23[27] , \nOut0_23[26] , \nOut0_23[25] , 
        \nOut0_23[24] , \nOut0_23[23] , \nOut0_23[22] , \nOut0_23[21] , 
        \nOut0_23[20] , \nOut0_23[19] , \nOut0_23[18] , \nOut0_23[17] , 
        \nOut0_23[16] , \nOut0_23[15] , \nOut0_23[14] , \nOut0_23[13] , 
        \nOut0_23[12] , \nOut0_23[11] , \nOut0_23[10] , \nOut0_23[9] , 
        \nOut0_23[8] , \nOut0_23[7] , \nOut0_23[6] , \nOut0_23[5] , 
        \nOut0_23[4] , \nOut0_23[3] , \nOut0_23[2] , \nOut0_23[1] , 
        \nOut0_23[0] }), .EAST_EDGE(\nOut1_22[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_21[31] ), .SE_EDGE(
        \nOut1_23[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_57 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut58[31] , \nScanOut58[30] , \nScanOut58[29] , 
        \nScanOut58[28] , \nScanOut58[27] , \nScanOut58[26] , \nScanOut58[25] , 
        \nScanOut58[24] , \nScanOut58[23] , \nScanOut58[22] , \nScanOut58[21] , 
        \nScanOut58[20] , \nScanOut58[19] , \nScanOut58[18] , \nScanOut58[17] , 
        \nScanOut58[16] , \nScanOut58[15] , \nScanOut58[14] , \nScanOut58[13] , 
        \nScanOut58[12] , \nScanOut58[11] , \nScanOut58[10] , \nScanOut58[9] , 
        \nScanOut58[8] , \nScanOut58[7] , \nScanOut58[6] , \nScanOut58[5] , 
        \nScanOut58[4] , \nScanOut58[3] , \nScanOut58[2] , \nScanOut58[1] , 
        \nScanOut58[0] }), .ScanOut({\nScanOut57[31] , \nScanOut57[30] , 
        \nScanOut57[29] , \nScanOut57[28] , \nScanOut57[27] , \nScanOut57[26] , 
        \nScanOut57[25] , \nScanOut57[24] , \nScanOut57[23] , \nScanOut57[22] , 
        \nScanOut57[21] , \nScanOut57[20] , \nScanOut57[19] , \nScanOut57[18] , 
        \nScanOut57[17] , \nScanOut57[16] , \nScanOut57[15] , \nScanOut57[14] , 
        \nScanOut57[13] , \nScanOut57[12] , \nScanOut57[11] , \nScanOut57[10] , 
        \nScanOut57[9] , \nScanOut57[8] , \nScanOut57[7] , \nScanOut57[6] , 
        \nScanOut57[5] , \nScanOut57[4] , \nScanOut57[3] , \nScanOut57[2] , 
        \nScanOut57[1] , \nScanOut57[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_57[31] , 
        \nOut0_57[30] , \nOut0_57[29] , \nOut0_57[28] , \nOut0_57[27] , 
        \nOut0_57[26] , \nOut0_57[25] , \nOut0_57[24] , \nOut0_57[23] , 
        \nOut0_57[22] , \nOut0_57[21] , \nOut0_57[20] , \nOut0_57[19] , 
        \nOut0_57[18] , \nOut0_57[17] , \nOut0_57[16] , \nOut0_57[15] , 
        \nOut0_57[14] , \nOut0_57[13] , \nOut0_57[12] , \nOut0_57[11] , 
        \nOut0_57[10] , \nOut0_57[9] , \nOut0_57[8] , \nOut0_57[7] , 
        \nOut0_57[6] , \nOut0_57[5] , \nOut0_57[4] , \nOut0_57[3] , 
        \nOut0_57[2] , \nOut0_57[1] , \nOut0_57[0] }), .NORTH_EDGE({
        \nOut0_56[31] , \nOut0_56[30] , \nOut0_56[29] , \nOut0_56[28] , 
        \nOut0_56[27] , \nOut0_56[26] , \nOut0_56[25] , \nOut0_56[24] , 
        \nOut0_56[23] , \nOut0_56[22] , \nOut0_56[21] , \nOut0_56[20] , 
        \nOut0_56[19] , \nOut0_56[18] , \nOut0_56[17] , \nOut0_56[16] , 
        \nOut0_56[15] , \nOut0_56[14] , \nOut0_56[13] , \nOut0_56[12] , 
        \nOut0_56[11] , \nOut0_56[10] , \nOut0_56[9] , \nOut0_56[8] , 
        \nOut0_56[7] , \nOut0_56[6] , \nOut0_56[5] , \nOut0_56[4] , 
        \nOut0_56[3] , \nOut0_56[2] , \nOut0_56[1] , \nOut0_56[0] }), 
        .SOUTH_EDGE({\nOut0_58[31] , \nOut0_58[30] , \nOut0_58[29] , 
        \nOut0_58[28] , \nOut0_58[27] , \nOut0_58[26] , \nOut0_58[25] , 
        \nOut0_58[24] , \nOut0_58[23] , \nOut0_58[22] , \nOut0_58[21] , 
        \nOut0_58[20] , \nOut0_58[19] , \nOut0_58[18] , \nOut0_58[17] , 
        \nOut0_58[16] , \nOut0_58[15] , \nOut0_58[14] , \nOut0_58[13] , 
        \nOut0_58[12] , \nOut0_58[11] , \nOut0_58[10] , \nOut0_58[9] , 
        \nOut0_58[8] , \nOut0_58[7] , \nOut0_58[6] , \nOut0_58[5] , 
        \nOut0_58[4] , \nOut0_58[3] , \nOut0_58[2] , \nOut0_58[1] , 
        \nOut0_58[0] }), .EAST_EDGE(\nOut1_57[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_56[31] ), .SE_EDGE(
        \nOut1_58[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_70 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut71[31] , \nScanOut71[30] , \nScanOut71[29] , 
        \nScanOut71[28] , \nScanOut71[27] , \nScanOut71[26] , \nScanOut71[25] , 
        \nScanOut71[24] , \nScanOut71[23] , \nScanOut71[22] , \nScanOut71[21] , 
        \nScanOut71[20] , \nScanOut71[19] , \nScanOut71[18] , \nScanOut71[17] , 
        \nScanOut71[16] , \nScanOut71[15] , \nScanOut71[14] , \nScanOut71[13] , 
        \nScanOut71[12] , \nScanOut71[11] , \nScanOut71[10] , \nScanOut71[9] , 
        \nScanOut71[8] , \nScanOut71[7] , \nScanOut71[6] , \nScanOut71[5] , 
        \nScanOut71[4] , \nScanOut71[3] , \nScanOut71[2] , \nScanOut71[1] , 
        \nScanOut71[0] }), .ScanOut({\nScanOut70[31] , \nScanOut70[30] , 
        \nScanOut70[29] , \nScanOut70[28] , \nScanOut70[27] , \nScanOut70[26] , 
        \nScanOut70[25] , \nScanOut70[24] , \nScanOut70[23] , \nScanOut70[22] , 
        \nScanOut70[21] , \nScanOut70[20] , \nScanOut70[19] , \nScanOut70[18] , 
        \nScanOut70[17] , \nScanOut70[16] , \nScanOut70[15] , \nScanOut70[14] , 
        \nScanOut70[13] , \nScanOut70[12] , \nScanOut70[11] , \nScanOut70[10] , 
        \nScanOut70[9] , \nScanOut70[8] , \nScanOut70[7] , \nScanOut70[6] , 
        \nScanOut70[5] , \nScanOut70[4] , \nScanOut70[3] , \nScanOut70[2] , 
        \nScanOut70[1] , \nScanOut70[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_6[31] , 
        \nOut1_6[30] , \nOut1_6[29] , \nOut1_6[28] , \nOut1_6[27] , 
        \nOut1_6[26] , \nOut1_6[25] , \nOut1_6[24] , \nOut1_6[23] , 
        \nOut1_6[22] , \nOut1_6[21] , \nOut1_6[20] , \nOut1_6[19] , 
        \nOut1_6[18] , \nOut1_6[17] , \nOut1_6[16] , \nOut1_6[15] , 
        \nOut1_6[14] , \nOut1_6[13] , \nOut1_6[12] , \nOut1_6[11] , 
        \nOut1_6[10] , \nOut1_6[9] , \nOut1_6[8] , \nOut1_6[7] , \nOut1_6[6] , 
        \nOut1_6[5] , \nOut1_6[4] , \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , 
        \nOut1_6[0] }), .NORTH_EDGE({\nOut1_5[31] , \nOut1_5[30] , 
        \nOut1_5[29] , \nOut1_5[28] , \nOut1_5[27] , \nOut1_5[26] , 
        \nOut1_5[25] , \nOut1_5[24] , \nOut1_5[23] , \nOut1_5[22] , 
        \nOut1_5[21] , \nOut1_5[20] , \nOut1_5[19] , \nOut1_5[18] , 
        \nOut1_5[17] , \nOut1_5[16] , \nOut1_5[15] , \nOut1_5[14] , 
        \nOut1_5[13] , \nOut1_5[12] , \nOut1_5[11] , \nOut1_5[10] , 
        \nOut1_5[9] , \nOut1_5[8] , \nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , 
        \nOut1_5[4] , \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }), 
        .SOUTH_EDGE({\nOut1_7[31] , \nOut1_7[30] , \nOut1_7[29] , 
        \nOut1_7[28] , \nOut1_7[27] , \nOut1_7[26] , \nOut1_7[25] , 
        \nOut1_7[24] , \nOut1_7[23] , \nOut1_7[22] , \nOut1_7[21] , 
        \nOut1_7[20] , \nOut1_7[19] , \nOut1_7[18] , \nOut1_7[17] , 
        \nOut1_7[16] , \nOut1_7[15] , \nOut1_7[14] , \nOut1_7[13] , 
        \nOut1_7[12] , \nOut1_7[11] , \nOut1_7[10] , \nOut1_7[9] , 
        \nOut1_7[8] , \nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , \nOut1_7[4] , 
        \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_6[0] ), .NW_EDGE(\nOut0_5[0] ), .SW_EDGE(
        \nOut0_7[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_126 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut127[31] , \nScanOut127[30] , \nScanOut127[29] , 
        \nScanOut127[28] , \nScanOut127[27] , \nScanOut127[26] , 
        \nScanOut127[25] , \nScanOut127[24] , \nScanOut127[23] , 
        \nScanOut127[22] , \nScanOut127[21] , \nScanOut127[20] , 
        \nScanOut127[19] , \nScanOut127[18] , \nScanOut127[17] , 
        \nScanOut127[16] , \nScanOut127[15] , \nScanOut127[14] , 
        \nScanOut127[13] , \nScanOut127[12] , \nScanOut127[11] , 
        \nScanOut127[10] , \nScanOut127[9] , \nScanOut127[8] , 
        \nScanOut127[7] , \nScanOut127[6] , \nScanOut127[5] , \nScanOut127[4] , 
        \nScanOut127[3] , \nScanOut127[2] , \nScanOut127[1] , \nScanOut127[0] 
        }), .ScanOut({\nScanOut126[31] , \nScanOut126[30] , \nScanOut126[29] , 
        \nScanOut126[28] , \nScanOut126[27] , \nScanOut126[26] , 
        \nScanOut126[25] , \nScanOut126[24] , \nScanOut126[23] , 
        \nScanOut126[22] , \nScanOut126[21] , \nScanOut126[20] , 
        \nScanOut126[19] , \nScanOut126[18] , \nScanOut126[17] , 
        \nScanOut126[16] , \nScanOut126[15] , \nScanOut126[14] , 
        \nScanOut126[13] , \nScanOut126[12] , \nScanOut126[11] , 
        \nScanOut126[10] , \nScanOut126[9] , \nScanOut126[8] , 
        \nScanOut126[7] , \nScanOut126[6] , \nScanOut126[5] , \nScanOut126[4] , 
        \nScanOut126[3] , \nScanOut126[2] , \nScanOut126[1] , \nScanOut126[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_62[31] , \nOut1_62[30] , \nOut1_62[29] , 
        \nOut1_62[28] , \nOut1_62[27] , \nOut1_62[26] , \nOut1_62[25] , 
        \nOut1_62[24] , \nOut1_62[23] , \nOut1_62[22] , \nOut1_62[21] , 
        \nOut1_62[20] , \nOut1_62[19] , \nOut1_62[18] , \nOut1_62[17] , 
        \nOut1_62[16] , \nOut1_62[15] , \nOut1_62[14] , \nOut1_62[13] , 
        \nOut1_62[12] , \nOut1_62[11] , \nOut1_62[10] , \nOut1_62[9] , 
        \nOut1_62[8] , \nOut1_62[7] , \nOut1_62[6] , \nOut1_62[5] , 
        \nOut1_62[4] , \nOut1_62[3] , \nOut1_62[2] , \nOut1_62[1] , 
        \nOut1_62[0] }), .NORTH_EDGE({\nOut1_61[31] , \nOut1_61[30] , 
        \nOut1_61[29] , \nOut1_61[28] , \nOut1_61[27] , \nOut1_61[26] , 
        \nOut1_61[25] , \nOut1_61[24] , \nOut1_61[23] , \nOut1_61[22] , 
        \nOut1_61[21] , \nOut1_61[20] , \nOut1_61[19] , \nOut1_61[18] , 
        \nOut1_61[17] , \nOut1_61[16] , \nOut1_61[15] , \nOut1_61[14] , 
        \nOut1_61[13] , \nOut1_61[12] , \nOut1_61[11] , \nOut1_61[10] , 
        \nOut1_61[9] , \nOut1_61[8] , \nOut1_61[7] , \nOut1_61[6] , 
        \nOut1_61[5] , \nOut1_61[4] , \nOut1_61[3] , \nOut1_61[2] , 
        \nOut1_61[1] , \nOut1_61[0] }), .SOUTH_EDGE({\nOut1_63[31] , 
        \nOut1_63[30] , \nOut1_63[29] , \nOut1_63[28] , \nOut1_63[27] , 
        \nOut1_63[26] , \nOut1_63[25] , \nOut1_63[24] , \nOut1_63[23] , 
        \nOut1_63[22] , \nOut1_63[21] , \nOut1_63[20] , \nOut1_63[19] , 
        \nOut1_63[18] , \nOut1_63[17] , \nOut1_63[16] , \nOut1_63[15] , 
        \nOut1_63[14] , \nOut1_63[13] , \nOut1_63[12] , \nOut1_63[11] , 
        \nOut1_63[10] , \nOut1_63[9] , \nOut1_63[8] , \nOut1_63[7] , 
        \nOut1_63[6] , \nOut1_63[5] , \nOut1_63[4] , \nOut1_63[3] , 
        \nOut1_63[2] , \nOut1_63[1] , \nOut1_63[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_62[0] ), .NW_EDGE(\nOut0_61[0] ), .SW_EDGE(
        \nOut0_63[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_101 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut102[31] , \nScanOut102[30] , \nScanOut102[29] , 
        \nScanOut102[28] , \nScanOut102[27] , \nScanOut102[26] , 
        \nScanOut102[25] , \nScanOut102[24] , \nScanOut102[23] , 
        \nScanOut102[22] , \nScanOut102[21] , \nScanOut102[20] , 
        \nScanOut102[19] , \nScanOut102[18] , \nScanOut102[17] , 
        \nScanOut102[16] , \nScanOut102[15] , \nScanOut102[14] , 
        \nScanOut102[13] , \nScanOut102[12] , \nScanOut102[11] , 
        \nScanOut102[10] , \nScanOut102[9] , \nScanOut102[8] , 
        \nScanOut102[7] , \nScanOut102[6] , \nScanOut102[5] , \nScanOut102[4] , 
        \nScanOut102[3] , \nScanOut102[2] , \nScanOut102[1] , \nScanOut102[0] 
        }), .ScanOut({\nScanOut101[31] , \nScanOut101[30] , \nScanOut101[29] , 
        \nScanOut101[28] , \nScanOut101[27] , \nScanOut101[26] , 
        \nScanOut101[25] , \nScanOut101[24] , \nScanOut101[23] , 
        \nScanOut101[22] , \nScanOut101[21] , \nScanOut101[20] , 
        \nScanOut101[19] , \nScanOut101[18] , \nScanOut101[17] , 
        \nScanOut101[16] , \nScanOut101[15] , \nScanOut101[14] , 
        \nScanOut101[13] , \nScanOut101[12] , \nScanOut101[11] , 
        \nScanOut101[10] , \nScanOut101[9] , \nScanOut101[8] , 
        \nScanOut101[7] , \nScanOut101[6] , \nScanOut101[5] , \nScanOut101[4] , 
        \nScanOut101[3] , \nScanOut101[2] , \nScanOut101[1] , \nScanOut101[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_37[31] , \nOut1_37[30] , \nOut1_37[29] , 
        \nOut1_37[28] , \nOut1_37[27] , \nOut1_37[26] , \nOut1_37[25] , 
        \nOut1_37[24] , \nOut1_37[23] , \nOut1_37[22] , \nOut1_37[21] , 
        \nOut1_37[20] , \nOut1_37[19] , \nOut1_37[18] , \nOut1_37[17] , 
        \nOut1_37[16] , \nOut1_37[15] , \nOut1_37[14] , \nOut1_37[13] , 
        \nOut1_37[12] , \nOut1_37[11] , \nOut1_37[10] , \nOut1_37[9] , 
        \nOut1_37[8] , \nOut1_37[7] , \nOut1_37[6] , \nOut1_37[5] , 
        \nOut1_37[4] , \nOut1_37[3] , \nOut1_37[2] , \nOut1_37[1] , 
        \nOut1_37[0] }), .NORTH_EDGE({\nOut1_36[31] , \nOut1_36[30] , 
        \nOut1_36[29] , \nOut1_36[28] , \nOut1_36[27] , \nOut1_36[26] , 
        \nOut1_36[25] , \nOut1_36[24] , \nOut1_36[23] , \nOut1_36[22] , 
        \nOut1_36[21] , \nOut1_36[20] , \nOut1_36[19] , \nOut1_36[18] , 
        \nOut1_36[17] , \nOut1_36[16] , \nOut1_36[15] , \nOut1_36[14] , 
        \nOut1_36[13] , \nOut1_36[12] , \nOut1_36[11] , \nOut1_36[10] , 
        \nOut1_36[9] , \nOut1_36[8] , \nOut1_36[7] , \nOut1_36[6] , 
        \nOut1_36[5] , \nOut1_36[4] , \nOut1_36[3] , \nOut1_36[2] , 
        \nOut1_36[1] , \nOut1_36[0] }), .SOUTH_EDGE({\nOut1_38[31] , 
        \nOut1_38[30] , \nOut1_38[29] , \nOut1_38[28] , \nOut1_38[27] , 
        \nOut1_38[26] , \nOut1_38[25] , \nOut1_38[24] , \nOut1_38[23] , 
        \nOut1_38[22] , \nOut1_38[21] , \nOut1_38[20] , \nOut1_38[19] , 
        \nOut1_38[18] , \nOut1_38[17] , \nOut1_38[16] , \nOut1_38[15] , 
        \nOut1_38[14] , \nOut1_38[13] , \nOut1_38[12] , \nOut1_38[11] , 
        \nOut1_38[10] , \nOut1_38[9] , \nOut1_38[8] , \nOut1_38[7] , 
        \nOut1_38[6] , \nOut1_38[5] , \nOut1_38[4] , \nOut1_38[3] , 
        \nOut1_38[2] , \nOut1_38[1] , \nOut1_38[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_37[0] ), .NW_EDGE(\nOut0_36[0] ), .SW_EDGE(
        \nOut0_38[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_30 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut31[31] , \nScanOut31[30] , \nScanOut31[29] , 
        \nScanOut31[28] , \nScanOut31[27] , \nScanOut31[26] , \nScanOut31[25] , 
        \nScanOut31[24] , \nScanOut31[23] , \nScanOut31[22] , \nScanOut31[21] , 
        \nScanOut31[20] , \nScanOut31[19] , \nScanOut31[18] , \nScanOut31[17] , 
        \nScanOut31[16] , \nScanOut31[15] , \nScanOut31[14] , \nScanOut31[13] , 
        \nScanOut31[12] , \nScanOut31[11] , \nScanOut31[10] , \nScanOut31[9] , 
        \nScanOut31[8] , \nScanOut31[7] , \nScanOut31[6] , \nScanOut31[5] , 
        \nScanOut31[4] , \nScanOut31[3] , \nScanOut31[2] , \nScanOut31[1] , 
        \nScanOut31[0] }), .ScanOut({\nScanOut30[31] , \nScanOut30[30] , 
        \nScanOut30[29] , \nScanOut30[28] , \nScanOut30[27] , \nScanOut30[26] , 
        \nScanOut30[25] , \nScanOut30[24] , \nScanOut30[23] , \nScanOut30[22] , 
        \nScanOut30[21] , \nScanOut30[20] , \nScanOut30[19] , \nScanOut30[18] , 
        \nScanOut30[17] , \nScanOut30[16] , \nScanOut30[15] , \nScanOut30[14] , 
        \nScanOut30[13] , \nScanOut30[12] , \nScanOut30[11] , \nScanOut30[10] , 
        \nScanOut30[9] , \nScanOut30[8] , \nScanOut30[7] , \nScanOut30[6] , 
        \nScanOut30[5] , \nScanOut30[4] , \nScanOut30[3] , \nScanOut30[2] , 
        \nScanOut30[1] , \nScanOut30[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_30[31] , 
        \nOut0_30[30] , \nOut0_30[29] , \nOut0_30[28] , \nOut0_30[27] , 
        \nOut0_30[26] , \nOut0_30[25] , \nOut0_30[24] , \nOut0_30[23] , 
        \nOut0_30[22] , \nOut0_30[21] , \nOut0_30[20] , \nOut0_30[19] , 
        \nOut0_30[18] , \nOut0_30[17] , \nOut0_30[16] , \nOut0_30[15] , 
        \nOut0_30[14] , \nOut0_30[13] , \nOut0_30[12] , \nOut0_30[11] , 
        \nOut0_30[10] , \nOut0_30[9] , \nOut0_30[8] , \nOut0_30[7] , 
        \nOut0_30[6] , \nOut0_30[5] , \nOut0_30[4] , \nOut0_30[3] , 
        \nOut0_30[2] , \nOut0_30[1] , \nOut0_30[0] }), .NORTH_EDGE({
        \nOut0_29[31] , \nOut0_29[30] , \nOut0_29[29] , \nOut0_29[28] , 
        \nOut0_29[27] , \nOut0_29[26] , \nOut0_29[25] , \nOut0_29[24] , 
        \nOut0_29[23] , \nOut0_29[22] , \nOut0_29[21] , \nOut0_29[20] , 
        \nOut0_29[19] , \nOut0_29[18] , \nOut0_29[17] , \nOut0_29[16] , 
        \nOut0_29[15] , \nOut0_29[14] , \nOut0_29[13] , \nOut0_29[12] , 
        \nOut0_29[11] , \nOut0_29[10] , \nOut0_29[9] , \nOut0_29[8] , 
        \nOut0_29[7] , \nOut0_29[6] , \nOut0_29[5] , \nOut0_29[4] , 
        \nOut0_29[3] , \nOut0_29[2] , \nOut0_29[1] , \nOut0_29[0] }), 
        .SOUTH_EDGE({\nOut0_31[31] , \nOut0_31[30] , \nOut0_31[29] , 
        \nOut0_31[28] , \nOut0_31[27] , \nOut0_31[26] , \nOut0_31[25] , 
        \nOut0_31[24] , \nOut0_31[23] , \nOut0_31[22] , \nOut0_31[21] , 
        \nOut0_31[20] , \nOut0_31[19] , \nOut0_31[18] , \nOut0_31[17] , 
        \nOut0_31[16] , \nOut0_31[15] , \nOut0_31[14] , \nOut0_31[13] , 
        \nOut0_31[12] , \nOut0_31[11] , \nOut0_31[10] , \nOut0_31[9] , 
        \nOut0_31[8] , \nOut0_31[7] , \nOut0_31[6] , \nOut0_31[5] , 
        \nOut0_31[4] , \nOut0_31[3] , \nOut0_31[2] , \nOut0_31[1] , 
        \nOut0_31[0] }), .EAST_EDGE(\nOut1_30[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_29[31] ), .SE_EDGE(
        \nOut1_31[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut11[31] , \nScanOut11[30] , \nScanOut11[29] , 
        \nScanOut11[28] , \nScanOut11[27] , \nScanOut11[26] , \nScanOut11[25] , 
        \nScanOut11[24] , \nScanOut11[23] , \nScanOut11[22] , \nScanOut11[21] , 
        \nScanOut11[20] , \nScanOut11[19] , \nScanOut11[18] , \nScanOut11[17] , 
        \nScanOut11[16] , \nScanOut11[15] , \nScanOut11[14] , \nScanOut11[13] , 
        \nScanOut11[12] , \nScanOut11[11] , \nScanOut11[10] , \nScanOut11[9] , 
        \nScanOut11[8] , \nScanOut11[7] , \nScanOut11[6] , \nScanOut11[5] , 
        \nScanOut11[4] , \nScanOut11[3] , \nScanOut11[2] , \nScanOut11[1] , 
        \nScanOut11[0] }), .ScanOut({\nScanOut10[31] , \nScanOut10[30] , 
        \nScanOut10[29] , \nScanOut10[28] , \nScanOut10[27] , \nScanOut10[26] , 
        \nScanOut10[25] , \nScanOut10[24] , \nScanOut10[23] , \nScanOut10[22] , 
        \nScanOut10[21] , \nScanOut10[20] , \nScanOut10[19] , \nScanOut10[18] , 
        \nScanOut10[17] , \nScanOut10[16] , \nScanOut10[15] , \nScanOut10[14] , 
        \nScanOut10[13] , \nScanOut10[12] , \nScanOut10[11] , \nScanOut10[10] , 
        \nScanOut10[9] , \nScanOut10[8] , \nScanOut10[7] , \nScanOut10[6] , 
        \nScanOut10[5] , \nScanOut10[4] , \nScanOut10[3] , \nScanOut10[2] , 
        \nScanOut10[1] , \nScanOut10[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_10[31] , 
        \nOut0_10[30] , \nOut0_10[29] , \nOut0_10[28] , \nOut0_10[27] , 
        \nOut0_10[26] , \nOut0_10[25] , \nOut0_10[24] , \nOut0_10[23] , 
        \nOut0_10[22] , \nOut0_10[21] , \nOut0_10[20] , \nOut0_10[19] , 
        \nOut0_10[18] , \nOut0_10[17] , \nOut0_10[16] , \nOut0_10[15] , 
        \nOut0_10[14] , \nOut0_10[13] , \nOut0_10[12] , \nOut0_10[11] , 
        \nOut0_10[10] , \nOut0_10[9] , \nOut0_10[8] , \nOut0_10[7] , 
        \nOut0_10[6] , \nOut0_10[5] , \nOut0_10[4] , \nOut0_10[3] , 
        \nOut0_10[2] , \nOut0_10[1] , \nOut0_10[0] }), .NORTH_EDGE({
        \nOut0_9[31] , \nOut0_9[30] , \nOut0_9[29] , \nOut0_9[28] , 
        \nOut0_9[27] , \nOut0_9[26] , \nOut0_9[25] , \nOut0_9[24] , 
        \nOut0_9[23] , \nOut0_9[22] , \nOut0_9[21] , \nOut0_9[20] , 
        \nOut0_9[19] , \nOut0_9[18] , \nOut0_9[17] , \nOut0_9[16] , 
        \nOut0_9[15] , \nOut0_9[14] , \nOut0_9[13] , \nOut0_9[12] , 
        \nOut0_9[11] , \nOut0_9[10] , \nOut0_9[9] , \nOut0_9[8] , \nOut0_9[7] , 
        \nOut0_9[6] , \nOut0_9[5] , \nOut0_9[4] , \nOut0_9[3] , \nOut0_9[2] , 
        \nOut0_9[1] , \nOut0_9[0] }), .SOUTH_EDGE({\nOut0_11[31] , 
        \nOut0_11[30] , \nOut0_11[29] , \nOut0_11[28] , \nOut0_11[27] , 
        \nOut0_11[26] , \nOut0_11[25] , \nOut0_11[24] , \nOut0_11[23] , 
        \nOut0_11[22] , \nOut0_11[21] , \nOut0_11[20] , \nOut0_11[19] , 
        \nOut0_11[18] , \nOut0_11[17] , \nOut0_11[16] , \nOut0_11[15] , 
        \nOut0_11[14] , \nOut0_11[13] , \nOut0_11[12] , \nOut0_11[11] , 
        \nOut0_11[10] , \nOut0_11[9] , \nOut0_11[8] , \nOut0_11[7] , 
        \nOut0_11[6] , \nOut0_11[5] , \nOut0_11[4] , \nOut0_11[3] , 
        \nOut0_11[2] , \nOut0_11[1] , \nOut0_11[0] }), .EAST_EDGE(
        \nOut1_10[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_9[31] ), .SE_EDGE(\nOut1_11[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_37 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut38[31] , \nScanOut38[30] , \nScanOut38[29] , 
        \nScanOut38[28] , \nScanOut38[27] , \nScanOut38[26] , \nScanOut38[25] , 
        \nScanOut38[24] , \nScanOut38[23] , \nScanOut38[22] , \nScanOut38[21] , 
        \nScanOut38[20] , \nScanOut38[19] , \nScanOut38[18] , \nScanOut38[17] , 
        \nScanOut38[16] , \nScanOut38[15] , \nScanOut38[14] , \nScanOut38[13] , 
        \nScanOut38[12] , \nScanOut38[11] , \nScanOut38[10] , \nScanOut38[9] , 
        \nScanOut38[8] , \nScanOut38[7] , \nScanOut38[6] , \nScanOut38[5] , 
        \nScanOut38[4] , \nScanOut38[3] , \nScanOut38[2] , \nScanOut38[1] , 
        \nScanOut38[0] }), .ScanOut({\nScanOut37[31] , \nScanOut37[30] , 
        \nScanOut37[29] , \nScanOut37[28] , \nScanOut37[27] , \nScanOut37[26] , 
        \nScanOut37[25] , \nScanOut37[24] , \nScanOut37[23] , \nScanOut37[22] , 
        \nScanOut37[21] , \nScanOut37[20] , \nScanOut37[19] , \nScanOut37[18] , 
        \nScanOut37[17] , \nScanOut37[16] , \nScanOut37[15] , \nScanOut37[14] , 
        \nScanOut37[13] , \nScanOut37[12] , \nScanOut37[11] , \nScanOut37[10] , 
        \nScanOut37[9] , \nScanOut37[8] , \nScanOut37[7] , \nScanOut37[6] , 
        \nScanOut37[5] , \nScanOut37[4] , \nScanOut37[3] , \nScanOut37[2] , 
        \nScanOut37[1] , \nScanOut37[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_37[31] , 
        \nOut0_37[30] , \nOut0_37[29] , \nOut0_37[28] , \nOut0_37[27] , 
        \nOut0_37[26] , \nOut0_37[25] , \nOut0_37[24] , \nOut0_37[23] , 
        \nOut0_37[22] , \nOut0_37[21] , \nOut0_37[20] , \nOut0_37[19] , 
        \nOut0_37[18] , \nOut0_37[17] , \nOut0_37[16] , \nOut0_37[15] , 
        \nOut0_37[14] , \nOut0_37[13] , \nOut0_37[12] , \nOut0_37[11] , 
        \nOut0_37[10] , \nOut0_37[9] , \nOut0_37[8] , \nOut0_37[7] , 
        \nOut0_37[6] , \nOut0_37[5] , \nOut0_37[4] , \nOut0_37[3] , 
        \nOut0_37[2] , \nOut0_37[1] , \nOut0_37[0] }), .NORTH_EDGE({
        \nOut0_36[31] , \nOut0_36[30] , \nOut0_36[29] , \nOut0_36[28] , 
        \nOut0_36[27] , \nOut0_36[26] , \nOut0_36[25] , \nOut0_36[24] , 
        \nOut0_36[23] , \nOut0_36[22] , \nOut0_36[21] , \nOut0_36[20] , 
        \nOut0_36[19] , \nOut0_36[18] , \nOut0_36[17] , \nOut0_36[16] , 
        \nOut0_36[15] , \nOut0_36[14] , \nOut0_36[13] , \nOut0_36[12] , 
        \nOut0_36[11] , \nOut0_36[10] , \nOut0_36[9] , \nOut0_36[8] , 
        \nOut0_36[7] , \nOut0_36[6] , \nOut0_36[5] , \nOut0_36[4] , 
        \nOut0_36[3] , \nOut0_36[2] , \nOut0_36[1] , \nOut0_36[0] }), 
        .SOUTH_EDGE({\nOut0_38[31] , \nOut0_38[30] , \nOut0_38[29] , 
        \nOut0_38[28] , \nOut0_38[27] , \nOut0_38[26] , \nOut0_38[25] , 
        \nOut0_38[24] , \nOut0_38[23] , \nOut0_38[22] , \nOut0_38[21] , 
        \nOut0_38[20] , \nOut0_38[19] , \nOut0_38[18] , \nOut0_38[17] , 
        \nOut0_38[16] , \nOut0_38[15] , \nOut0_38[14] , \nOut0_38[13] , 
        \nOut0_38[12] , \nOut0_38[11] , \nOut0_38[10] , \nOut0_38[9] , 
        \nOut0_38[8] , \nOut0_38[7] , \nOut0_38[6] , \nOut0_38[5] , 
        \nOut0_38[4] , \nOut0_38[3] , \nOut0_38[2] , \nOut0_38[1] , 
        \nOut0_38[0] }), .EAST_EDGE(\nOut1_37[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_36[31] ), .SE_EDGE(
        \nOut1_38[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_42 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut43[31] , \nScanOut43[30] , \nScanOut43[29] , 
        \nScanOut43[28] , \nScanOut43[27] , \nScanOut43[26] , \nScanOut43[25] , 
        \nScanOut43[24] , \nScanOut43[23] , \nScanOut43[22] , \nScanOut43[21] , 
        \nScanOut43[20] , \nScanOut43[19] , \nScanOut43[18] , \nScanOut43[17] , 
        \nScanOut43[16] , \nScanOut43[15] , \nScanOut43[14] , \nScanOut43[13] , 
        \nScanOut43[12] , \nScanOut43[11] , \nScanOut43[10] , \nScanOut43[9] , 
        \nScanOut43[8] , \nScanOut43[7] , \nScanOut43[6] , \nScanOut43[5] , 
        \nScanOut43[4] , \nScanOut43[3] , \nScanOut43[2] , \nScanOut43[1] , 
        \nScanOut43[0] }), .ScanOut({\nScanOut42[31] , \nScanOut42[30] , 
        \nScanOut42[29] , \nScanOut42[28] , \nScanOut42[27] , \nScanOut42[26] , 
        \nScanOut42[25] , \nScanOut42[24] , \nScanOut42[23] , \nScanOut42[22] , 
        \nScanOut42[21] , \nScanOut42[20] , \nScanOut42[19] , \nScanOut42[18] , 
        \nScanOut42[17] , \nScanOut42[16] , \nScanOut42[15] , \nScanOut42[14] , 
        \nScanOut42[13] , \nScanOut42[12] , \nScanOut42[11] , \nScanOut42[10] , 
        \nScanOut42[9] , \nScanOut42[8] , \nScanOut42[7] , \nScanOut42[6] , 
        \nScanOut42[5] , \nScanOut42[4] , \nScanOut42[3] , \nScanOut42[2] , 
        \nScanOut42[1] , \nScanOut42[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_42[31] , 
        \nOut0_42[30] , \nOut0_42[29] , \nOut0_42[28] , \nOut0_42[27] , 
        \nOut0_42[26] , \nOut0_42[25] , \nOut0_42[24] , \nOut0_42[23] , 
        \nOut0_42[22] , \nOut0_42[21] , \nOut0_42[20] , \nOut0_42[19] , 
        \nOut0_42[18] , \nOut0_42[17] , \nOut0_42[16] , \nOut0_42[15] , 
        \nOut0_42[14] , \nOut0_42[13] , \nOut0_42[12] , \nOut0_42[11] , 
        \nOut0_42[10] , \nOut0_42[9] , \nOut0_42[8] , \nOut0_42[7] , 
        \nOut0_42[6] , \nOut0_42[5] , \nOut0_42[4] , \nOut0_42[3] , 
        \nOut0_42[2] , \nOut0_42[1] , \nOut0_42[0] }), .NORTH_EDGE({
        \nOut0_41[31] , \nOut0_41[30] , \nOut0_41[29] , \nOut0_41[28] , 
        \nOut0_41[27] , \nOut0_41[26] , \nOut0_41[25] , \nOut0_41[24] , 
        \nOut0_41[23] , \nOut0_41[22] , \nOut0_41[21] , \nOut0_41[20] , 
        \nOut0_41[19] , \nOut0_41[18] , \nOut0_41[17] , \nOut0_41[16] , 
        \nOut0_41[15] , \nOut0_41[14] , \nOut0_41[13] , \nOut0_41[12] , 
        \nOut0_41[11] , \nOut0_41[10] , \nOut0_41[9] , \nOut0_41[8] , 
        \nOut0_41[7] , \nOut0_41[6] , \nOut0_41[5] , \nOut0_41[4] , 
        \nOut0_41[3] , \nOut0_41[2] , \nOut0_41[1] , \nOut0_41[0] }), 
        .SOUTH_EDGE({\nOut0_43[31] , \nOut0_43[30] , \nOut0_43[29] , 
        \nOut0_43[28] , \nOut0_43[27] , \nOut0_43[26] , \nOut0_43[25] , 
        \nOut0_43[24] , \nOut0_43[23] , \nOut0_43[22] , \nOut0_43[21] , 
        \nOut0_43[20] , \nOut0_43[19] , \nOut0_43[18] , \nOut0_43[17] , 
        \nOut0_43[16] , \nOut0_43[15] , \nOut0_43[14] , \nOut0_43[13] , 
        \nOut0_43[12] , \nOut0_43[11] , \nOut0_43[10] , \nOut0_43[9] , 
        \nOut0_43[8] , \nOut0_43[7] , \nOut0_43[6] , \nOut0_43[5] , 
        \nOut0_43[4] , \nOut0_43[3] , \nOut0_43[2] , \nOut0_43[1] , 
        \nOut0_43[0] }), .EAST_EDGE(\nOut1_42[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_41[31] ), .SE_EDGE(
        \nOut1_43[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_45 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut46[31] , \nScanOut46[30] , \nScanOut46[29] , 
        \nScanOut46[28] , \nScanOut46[27] , \nScanOut46[26] , \nScanOut46[25] , 
        \nScanOut46[24] , \nScanOut46[23] , \nScanOut46[22] , \nScanOut46[21] , 
        \nScanOut46[20] , \nScanOut46[19] , \nScanOut46[18] , \nScanOut46[17] , 
        \nScanOut46[16] , \nScanOut46[15] , \nScanOut46[14] , \nScanOut46[13] , 
        \nScanOut46[12] , \nScanOut46[11] , \nScanOut46[10] , \nScanOut46[9] , 
        \nScanOut46[8] , \nScanOut46[7] , \nScanOut46[6] , \nScanOut46[5] , 
        \nScanOut46[4] , \nScanOut46[3] , \nScanOut46[2] , \nScanOut46[1] , 
        \nScanOut46[0] }), .ScanOut({\nScanOut45[31] , \nScanOut45[30] , 
        \nScanOut45[29] , \nScanOut45[28] , \nScanOut45[27] , \nScanOut45[26] , 
        \nScanOut45[25] , \nScanOut45[24] , \nScanOut45[23] , \nScanOut45[22] , 
        \nScanOut45[21] , \nScanOut45[20] , \nScanOut45[19] , \nScanOut45[18] , 
        \nScanOut45[17] , \nScanOut45[16] , \nScanOut45[15] , \nScanOut45[14] , 
        \nScanOut45[13] , \nScanOut45[12] , \nScanOut45[11] , \nScanOut45[10] , 
        \nScanOut45[9] , \nScanOut45[8] , \nScanOut45[7] , \nScanOut45[6] , 
        \nScanOut45[5] , \nScanOut45[4] , \nScanOut45[3] , \nScanOut45[2] , 
        \nScanOut45[1] , \nScanOut45[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_45[31] , 
        \nOut0_45[30] , \nOut0_45[29] , \nOut0_45[28] , \nOut0_45[27] , 
        \nOut0_45[26] , \nOut0_45[25] , \nOut0_45[24] , \nOut0_45[23] , 
        \nOut0_45[22] , \nOut0_45[21] , \nOut0_45[20] , \nOut0_45[19] , 
        \nOut0_45[18] , \nOut0_45[17] , \nOut0_45[16] , \nOut0_45[15] , 
        \nOut0_45[14] , \nOut0_45[13] , \nOut0_45[12] , \nOut0_45[11] , 
        \nOut0_45[10] , \nOut0_45[9] , \nOut0_45[8] , \nOut0_45[7] , 
        \nOut0_45[6] , \nOut0_45[5] , \nOut0_45[4] , \nOut0_45[3] , 
        \nOut0_45[2] , \nOut0_45[1] , \nOut0_45[0] }), .NORTH_EDGE({
        \nOut0_44[31] , \nOut0_44[30] , \nOut0_44[29] , \nOut0_44[28] , 
        \nOut0_44[27] , \nOut0_44[26] , \nOut0_44[25] , \nOut0_44[24] , 
        \nOut0_44[23] , \nOut0_44[22] , \nOut0_44[21] , \nOut0_44[20] , 
        \nOut0_44[19] , \nOut0_44[18] , \nOut0_44[17] , \nOut0_44[16] , 
        \nOut0_44[15] , \nOut0_44[14] , \nOut0_44[13] , \nOut0_44[12] , 
        \nOut0_44[11] , \nOut0_44[10] , \nOut0_44[9] , \nOut0_44[8] , 
        \nOut0_44[7] , \nOut0_44[6] , \nOut0_44[5] , \nOut0_44[4] , 
        \nOut0_44[3] , \nOut0_44[2] , \nOut0_44[1] , \nOut0_44[0] }), 
        .SOUTH_EDGE({\nOut0_46[31] , \nOut0_46[30] , \nOut0_46[29] , 
        \nOut0_46[28] , \nOut0_46[27] , \nOut0_46[26] , \nOut0_46[25] , 
        \nOut0_46[24] , \nOut0_46[23] , \nOut0_46[22] , \nOut0_46[21] , 
        \nOut0_46[20] , \nOut0_46[19] , \nOut0_46[18] , \nOut0_46[17] , 
        \nOut0_46[16] , \nOut0_46[15] , \nOut0_46[14] , \nOut0_46[13] , 
        \nOut0_46[12] , \nOut0_46[11] , \nOut0_46[10] , \nOut0_46[9] , 
        \nOut0_46[8] , \nOut0_46[7] , \nOut0_46[6] , \nOut0_46[5] , 
        \nOut0_46[4] , \nOut0_46[3] , \nOut0_46[2] , \nOut0_46[1] , 
        \nOut0_46[0] }), .EAST_EDGE(\nOut1_45[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_44[31] ), .SE_EDGE(
        \nOut1_46[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_62 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut63[31] , \nScanOut63[30] , \nScanOut63[29] , 
        \nScanOut63[28] , \nScanOut63[27] , \nScanOut63[26] , \nScanOut63[25] , 
        \nScanOut63[24] , \nScanOut63[23] , \nScanOut63[22] , \nScanOut63[21] , 
        \nScanOut63[20] , \nScanOut63[19] , \nScanOut63[18] , \nScanOut63[17] , 
        \nScanOut63[16] , \nScanOut63[15] , \nScanOut63[14] , \nScanOut63[13] , 
        \nScanOut63[12] , \nScanOut63[11] , \nScanOut63[10] , \nScanOut63[9] , 
        \nScanOut63[8] , \nScanOut63[7] , \nScanOut63[6] , \nScanOut63[5] , 
        \nScanOut63[4] , \nScanOut63[3] , \nScanOut63[2] , \nScanOut63[1] , 
        \nScanOut63[0] }), .ScanOut({\nScanOut62[31] , \nScanOut62[30] , 
        \nScanOut62[29] , \nScanOut62[28] , \nScanOut62[27] , \nScanOut62[26] , 
        \nScanOut62[25] , \nScanOut62[24] , \nScanOut62[23] , \nScanOut62[22] , 
        \nScanOut62[21] , \nScanOut62[20] , \nScanOut62[19] , \nScanOut62[18] , 
        \nScanOut62[17] , \nScanOut62[16] , \nScanOut62[15] , \nScanOut62[14] , 
        \nScanOut62[13] , \nScanOut62[12] , \nScanOut62[11] , \nScanOut62[10] , 
        \nScanOut62[9] , \nScanOut62[8] , \nScanOut62[7] , \nScanOut62[6] , 
        \nScanOut62[5] , \nScanOut62[4] , \nScanOut62[3] , \nScanOut62[2] , 
        \nScanOut62[1] , \nScanOut62[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_62[31] , 
        \nOut0_62[30] , \nOut0_62[29] , \nOut0_62[28] , \nOut0_62[27] , 
        \nOut0_62[26] , \nOut0_62[25] , \nOut0_62[24] , \nOut0_62[23] , 
        \nOut0_62[22] , \nOut0_62[21] , \nOut0_62[20] , \nOut0_62[19] , 
        \nOut0_62[18] , \nOut0_62[17] , \nOut0_62[16] , \nOut0_62[15] , 
        \nOut0_62[14] , \nOut0_62[13] , \nOut0_62[12] , \nOut0_62[11] , 
        \nOut0_62[10] , \nOut0_62[9] , \nOut0_62[8] , \nOut0_62[7] , 
        \nOut0_62[6] , \nOut0_62[5] , \nOut0_62[4] , \nOut0_62[3] , 
        \nOut0_62[2] , \nOut0_62[1] , \nOut0_62[0] }), .NORTH_EDGE({
        \nOut0_61[31] , \nOut0_61[30] , \nOut0_61[29] , \nOut0_61[28] , 
        \nOut0_61[27] , \nOut0_61[26] , \nOut0_61[25] , \nOut0_61[24] , 
        \nOut0_61[23] , \nOut0_61[22] , \nOut0_61[21] , \nOut0_61[20] , 
        \nOut0_61[19] , \nOut0_61[18] , \nOut0_61[17] , \nOut0_61[16] , 
        \nOut0_61[15] , \nOut0_61[14] , \nOut0_61[13] , \nOut0_61[12] , 
        \nOut0_61[11] , \nOut0_61[10] , \nOut0_61[9] , \nOut0_61[8] , 
        \nOut0_61[7] , \nOut0_61[6] , \nOut0_61[5] , \nOut0_61[4] , 
        \nOut0_61[3] , \nOut0_61[2] , \nOut0_61[1] , \nOut0_61[0] }), 
        .SOUTH_EDGE({\nOut0_63[31] , \nOut0_63[30] , \nOut0_63[29] , 
        \nOut0_63[28] , \nOut0_63[27] , \nOut0_63[26] , \nOut0_63[25] , 
        \nOut0_63[24] , \nOut0_63[23] , \nOut0_63[22] , \nOut0_63[21] , 
        \nOut0_63[20] , \nOut0_63[19] , \nOut0_63[18] , \nOut0_63[17] , 
        \nOut0_63[16] , \nOut0_63[15] , \nOut0_63[14] , \nOut0_63[13] , 
        \nOut0_63[12] , \nOut0_63[11] , \nOut0_63[10] , \nOut0_63[9] , 
        \nOut0_63[8] , \nOut0_63[7] , \nOut0_63[6] , \nOut0_63[5] , 
        \nOut0_63[4] , \nOut0_63[3] , \nOut0_63[2] , \nOut0_63[1] , 
        \nOut0_63[0] }), .EAST_EDGE(\nOut1_62[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_61[31] ), .SE_EDGE(
        \nOut1_63[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_79 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut80[31] , \nScanOut80[30] , \nScanOut80[29] , 
        \nScanOut80[28] , \nScanOut80[27] , \nScanOut80[26] , \nScanOut80[25] , 
        \nScanOut80[24] , \nScanOut80[23] , \nScanOut80[22] , \nScanOut80[21] , 
        \nScanOut80[20] , \nScanOut80[19] , \nScanOut80[18] , \nScanOut80[17] , 
        \nScanOut80[16] , \nScanOut80[15] , \nScanOut80[14] , \nScanOut80[13] , 
        \nScanOut80[12] , \nScanOut80[11] , \nScanOut80[10] , \nScanOut80[9] , 
        \nScanOut80[8] , \nScanOut80[7] , \nScanOut80[6] , \nScanOut80[5] , 
        \nScanOut80[4] , \nScanOut80[3] , \nScanOut80[2] , \nScanOut80[1] , 
        \nScanOut80[0] }), .ScanOut({\nScanOut79[31] , \nScanOut79[30] , 
        \nScanOut79[29] , \nScanOut79[28] , \nScanOut79[27] , \nScanOut79[26] , 
        \nScanOut79[25] , \nScanOut79[24] , \nScanOut79[23] , \nScanOut79[22] , 
        \nScanOut79[21] , \nScanOut79[20] , \nScanOut79[19] , \nScanOut79[18] , 
        \nScanOut79[17] , \nScanOut79[16] , \nScanOut79[15] , \nScanOut79[14] , 
        \nScanOut79[13] , \nScanOut79[12] , \nScanOut79[11] , \nScanOut79[10] , 
        \nScanOut79[9] , \nScanOut79[8] , \nScanOut79[7] , \nScanOut79[6] , 
        \nScanOut79[5] , \nScanOut79[4] , \nScanOut79[3] , \nScanOut79[2] , 
        \nScanOut79[1] , \nScanOut79[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_15[31] , 
        \nOut1_15[30] , \nOut1_15[29] , \nOut1_15[28] , \nOut1_15[27] , 
        \nOut1_15[26] , \nOut1_15[25] , \nOut1_15[24] , \nOut1_15[23] , 
        \nOut1_15[22] , \nOut1_15[21] , \nOut1_15[20] , \nOut1_15[19] , 
        \nOut1_15[18] , \nOut1_15[17] , \nOut1_15[16] , \nOut1_15[15] , 
        \nOut1_15[14] , \nOut1_15[13] , \nOut1_15[12] , \nOut1_15[11] , 
        \nOut1_15[10] , \nOut1_15[9] , \nOut1_15[8] , \nOut1_15[7] , 
        \nOut1_15[6] , \nOut1_15[5] , \nOut1_15[4] , \nOut1_15[3] , 
        \nOut1_15[2] , \nOut1_15[1] , \nOut1_15[0] }), .NORTH_EDGE({
        \nOut1_14[31] , \nOut1_14[30] , \nOut1_14[29] , \nOut1_14[28] , 
        \nOut1_14[27] , \nOut1_14[26] , \nOut1_14[25] , \nOut1_14[24] , 
        \nOut1_14[23] , \nOut1_14[22] , \nOut1_14[21] , \nOut1_14[20] , 
        \nOut1_14[19] , \nOut1_14[18] , \nOut1_14[17] , \nOut1_14[16] , 
        \nOut1_14[15] , \nOut1_14[14] , \nOut1_14[13] , \nOut1_14[12] , 
        \nOut1_14[11] , \nOut1_14[10] , \nOut1_14[9] , \nOut1_14[8] , 
        \nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), 
        .SOUTH_EDGE({\nOut1_16[31] , \nOut1_16[30] , \nOut1_16[29] , 
        \nOut1_16[28] , \nOut1_16[27] , \nOut1_16[26] , \nOut1_16[25] , 
        \nOut1_16[24] , \nOut1_16[23] , \nOut1_16[22] , \nOut1_16[21] , 
        \nOut1_16[20] , \nOut1_16[19] , \nOut1_16[18] , \nOut1_16[17] , 
        \nOut1_16[16] , \nOut1_16[15] , \nOut1_16[14] , \nOut1_16[13] , 
        \nOut1_16[12] , \nOut1_16[11] , \nOut1_16[10] , \nOut1_16[9] , 
        \nOut1_16[8] , \nOut1_16[7] , \nOut1_16[6] , \nOut1_16[5] , 
        \nOut1_16[4] , \nOut1_16[3] , \nOut1_16[2] , \nOut1_16[1] , 
        \nOut1_16[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_15[0] ), 
        .NW_EDGE(\nOut0_14[0] ), .SW_EDGE(\nOut0_16[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_108 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut109[31] , \nScanOut109[30] , \nScanOut109[29] , 
        \nScanOut109[28] , \nScanOut109[27] , \nScanOut109[26] , 
        \nScanOut109[25] , \nScanOut109[24] , \nScanOut109[23] , 
        \nScanOut109[22] , \nScanOut109[21] , \nScanOut109[20] , 
        \nScanOut109[19] , \nScanOut109[18] , \nScanOut109[17] , 
        \nScanOut109[16] , \nScanOut109[15] , \nScanOut109[14] , 
        \nScanOut109[13] , \nScanOut109[12] , \nScanOut109[11] , 
        \nScanOut109[10] , \nScanOut109[9] , \nScanOut109[8] , 
        \nScanOut109[7] , \nScanOut109[6] , \nScanOut109[5] , \nScanOut109[4] , 
        \nScanOut109[3] , \nScanOut109[2] , \nScanOut109[1] , \nScanOut109[0] 
        }), .ScanOut({\nScanOut108[31] , \nScanOut108[30] , \nScanOut108[29] , 
        \nScanOut108[28] , \nScanOut108[27] , \nScanOut108[26] , 
        \nScanOut108[25] , \nScanOut108[24] , \nScanOut108[23] , 
        \nScanOut108[22] , \nScanOut108[21] , \nScanOut108[20] , 
        \nScanOut108[19] , \nScanOut108[18] , \nScanOut108[17] , 
        \nScanOut108[16] , \nScanOut108[15] , \nScanOut108[14] , 
        \nScanOut108[13] , \nScanOut108[12] , \nScanOut108[11] , 
        \nScanOut108[10] , \nScanOut108[9] , \nScanOut108[8] , 
        \nScanOut108[7] , \nScanOut108[6] , \nScanOut108[5] , \nScanOut108[4] , 
        \nScanOut108[3] , \nScanOut108[2] , \nScanOut108[1] , \nScanOut108[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_44[31] , \nOut1_44[30] , \nOut1_44[29] , 
        \nOut1_44[28] , \nOut1_44[27] , \nOut1_44[26] , \nOut1_44[25] , 
        \nOut1_44[24] , \nOut1_44[23] , \nOut1_44[22] , \nOut1_44[21] , 
        \nOut1_44[20] , \nOut1_44[19] , \nOut1_44[18] , \nOut1_44[17] , 
        \nOut1_44[16] , \nOut1_44[15] , \nOut1_44[14] , \nOut1_44[13] , 
        \nOut1_44[12] , \nOut1_44[11] , \nOut1_44[10] , \nOut1_44[9] , 
        \nOut1_44[8] , \nOut1_44[7] , \nOut1_44[6] , \nOut1_44[5] , 
        \nOut1_44[4] , \nOut1_44[3] , \nOut1_44[2] , \nOut1_44[1] , 
        \nOut1_44[0] }), .NORTH_EDGE({\nOut1_43[31] , \nOut1_43[30] , 
        \nOut1_43[29] , \nOut1_43[28] , \nOut1_43[27] , \nOut1_43[26] , 
        \nOut1_43[25] , \nOut1_43[24] , \nOut1_43[23] , \nOut1_43[22] , 
        \nOut1_43[21] , \nOut1_43[20] , \nOut1_43[19] , \nOut1_43[18] , 
        \nOut1_43[17] , \nOut1_43[16] , \nOut1_43[15] , \nOut1_43[14] , 
        \nOut1_43[13] , \nOut1_43[12] , \nOut1_43[11] , \nOut1_43[10] , 
        \nOut1_43[9] , \nOut1_43[8] , \nOut1_43[7] , \nOut1_43[6] , 
        \nOut1_43[5] , \nOut1_43[4] , \nOut1_43[3] , \nOut1_43[2] , 
        \nOut1_43[1] , \nOut1_43[0] }), .SOUTH_EDGE({\nOut1_45[31] , 
        \nOut1_45[30] , \nOut1_45[29] , \nOut1_45[28] , \nOut1_45[27] , 
        \nOut1_45[26] , \nOut1_45[25] , \nOut1_45[24] , \nOut1_45[23] , 
        \nOut1_45[22] , \nOut1_45[21] , \nOut1_45[20] , \nOut1_45[19] , 
        \nOut1_45[18] , \nOut1_45[17] , \nOut1_45[16] , \nOut1_45[15] , 
        \nOut1_45[14] , \nOut1_45[13] , \nOut1_45[12] , \nOut1_45[11] , 
        \nOut1_45[10] , \nOut1_45[9] , \nOut1_45[8] , \nOut1_45[7] , 
        \nOut1_45[6] , \nOut1_45[5] , \nOut1_45[4] , \nOut1_45[3] , 
        \nOut1_45[2] , \nOut1_45[1] , \nOut1_45[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_44[0] ), .NW_EDGE(\nOut0_43[0] ), .SW_EDGE(
        \nOut0_45[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_80 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut81[31] , \nScanOut81[30] , \nScanOut81[29] , 
        \nScanOut81[28] , \nScanOut81[27] , \nScanOut81[26] , \nScanOut81[25] , 
        \nScanOut81[24] , \nScanOut81[23] , \nScanOut81[22] , \nScanOut81[21] , 
        \nScanOut81[20] , \nScanOut81[19] , \nScanOut81[18] , \nScanOut81[17] , 
        \nScanOut81[16] , \nScanOut81[15] , \nScanOut81[14] , \nScanOut81[13] , 
        \nScanOut81[12] , \nScanOut81[11] , \nScanOut81[10] , \nScanOut81[9] , 
        \nScanOut81[8] , \nScanOut81[7] , \nScanOut81[6] , \nScanOut81[5] , 
        \nScanOut81[4] , \nScanOut81[3] , \nScanOut81[2] , \nScanOut81[1] , 
        \nScanOut81[0] }), .ScanOut({\nScanOut80[31] , \nScanOut80[30] , 
        \nScanOut80[29] , \nScanOut80[28] , \nScanOut80[27] , \nScanOut80[26] , 
        \nScanOut80[25] , \nScanOut80[24] , \nScanOut80[23] , \nScanOut80[22] , 
        \nScanOut80[21] , \nScanOut80[20] , \nScanOut80[19] , \nScanOut80[18] , 
        \nScanOut80[17] , \nScanOut80[16] , \nScanOut80[15] , \nScanOut80[14] , 
        \nScanOut80[13] , \nScanOut80[12] , \nScanOut80[11] , \nScanOut80[10] , 
        \nScanOut80[9] , \nScanOut80[8] , \nScanOut80[7] , \nScanOut80[6] , 
        \nScanOut80[5] , \nScanOut80[4] , \nScanOut80[3] , \nScanOut80[2] , 
        \nScanOut80[1] , \nScanOut80[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_16[31] , 
        \nOut1_16[30] , \nOut1_16[29] , \nOut1_16[28] , \nOut1_16[27] , 
        \nOut1_16[26] , \nOut1_16[25] , \nOut1_16[24] , \nOut1_16[23] , 
        \nOut1_16[22] , \nOut1_16[21] , \nOut1_16[20] , \nOut1_16[19] , 
        \nOut1_16[18] , \nOut1_16[17] , \nOut1_16[16] , \nOut1_16[15] , 
        \nOut1_16[14] , \nOut1_16[13] , \nOut1_16[12] , \nOut1_16[11] , 
        \nOut1_16[10] , \nOut1_16[9] , \nOut1_16[8] , \nOut1_16[7] , 
        \nOut1_16[6] , \nOut1_16[5] , \nOut1_16[4] , \nOut1_16[3] , 
        \nOut1_16[2] , \nOut1_16[1] , \nOut1_16[0] }), .NORTH_EDGE({
        \nOut1_15[31] , \nOut1_15[30] , \nOut1_15[29] , \nOut1_15[28] , 
        \nOut1_15[27] , \nOut1_15[26] , \nOut1_15[25] , \nOut1_15[24] , 
        \nOut1_15[23] , \nOut1_15[22] , \nOut1_15[21] , \nOut1_15[20] , 
        \nOut1_15[19] , \nOut1_15[18] , \nOut1_15[17] , \nOut1_15[16] , 
        \nOut1_15[15] , \nOut1_15[14] , \nOut1_15[13] , \nOut1_15[12] , 
        \nOut1_15[11] , \nOut1_15[10] , \nOut1_15[9] , \nOut1_15[8] , 
        \nOut1_15[7] , \nOut1_15[6] , \nOut1_15[5] , \nOut1_15[4] , 
        \nOut1_15[3] , \nOut1_15[2] , \nOut1_15[1] , \nOut1_15[0] }), 
        .SOUTH_EDGE({\nOut1_17[31] , \nOut1_17[30] , \nOut1_17[29] , 
        \nOut1_17[28] , \nOut1_17[27] , \nOut1_17[26] , \nOut1_17[25] , 
        \nOut1_17[24] , \nOut1_17[23] , \nOut1_17[22] , \nOut1_17[21] , 
        \nOut1_17[20] , \nOut1_17[19] , \nOut1_17[18] , \nOut1_17[17] , 
        \nOut1_17[16] , \nOut1_17[15] , \nOut1_17[14] , \nOut1_17[13] , 
        \nOut1_17[12] , \nOut1_17[11] , \nOut1_17[10] , \nOut1_17[9] , 
        \nOut1_17[8] , \nOut1_17[7] , \nOut1_17[6] , \nOut1_17[5] , 
        \nOut1_17[4] , \nOut1_17[3] , \nOut1_17[2] , \nOut1_17[1] , 
        \nOut1_17[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_16[0] ), 
        .NW_EDGE(\nOut0_15[0] ), .SW_EDGE(\nOut0_17[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_87 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut88[31] , \nScanOut88[30] , \nScanOut88[29] , 
        \nScanOut88[28] , \nScanOut88[27] , \nScanOut88[26] , \nScanOut88[25] , 
        \nScanOut88[24] , \nScanOut88[23] , \nScanOut88[22] , \nScanOut88[21] , 
        \nScanOut88[20] , \nScanOut88[19] , \nScanOut88[18] , \nScanOut88[17] , 
        \nScanOut88[16] , \nScanOut88[15] , \nScanOut88[14] , \nScanOut88[13] , 
        \nScanOut88[12] , \nScanOut88[11] , \nScanOut88[10] , \nScanOut88[9] , 
        \nScanOut88[8] , \nScanOut88[7] , \nScanOut88[6] , \nScanOut88[5] , 
        \nScanOut88[4] , \nScanOut88[3] , \nScanOut88[2] , \nScanOut88[1] , 
        \nScanOut88[0] }), .ScanOut({\nScanOut87[31] , \nScanOut87[30] , 
        \nScanOut87[29] , \nScanOut87[28] , \nScanOut87[27] , \nScanOut87[26] , 
        \nScanOut87[25] , \nScanOut87[24] , \nScanOut87[23] , \nScanOut87[22] , 
        \nScanOut87[21] , \nScanOut87[20] , \nScanOut87[19] , \nScanOut87[18] , 
        \nScanOut87[17] , \nScanOut87[16] , \nScanOut87[15] , \nScanOut87[14] , 
        \nScanOut87[13] , \nScanOut87[12] , \nScanOut87[11] , \nScanOut87[10] , 
        \nScanOut87[9] , \nScanOut87[8] , \nScanOut87[7] , \nScanOut87[6] , 
        \nScanOut87[5] , \nScanOut87[4] , \nScanOut87[3] , \nScanOut87[2] , 
        \nScanOut87[1] , \nScanOut87[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_23[31] , 
        \nOut1_23[30] , \nOut1_23[29] , \nOut1_23[28] , \nOut1_23[27] , 
        \nOut1_23[26] , \nOut1_23[25] , \nOut1_23[24] , \nOut1_23[23] , 
        \nOut1_23[22] , \nOut1_23[21] , \nOut1_23[20] , \nOut1_23[19] , 
        \nOut1_23[18] , \nOut1_23[17] , \nOut1_23[16] , \nOut1_23[15] , 
        \nOut1_23[14] , \nOut1_23[13] , \nOut1_23[12] , \nOut1_23[11] , 
        \nOut1_23[10] , \nOut1_23[9] , \nOut1_23[8] , \nOut1_23[7] , 
        \nOut1_23[6] , \nOut1_23[5] , \nOut1_23[4] , \nOut1_23[3] , 
        \nOut1_23[2] , \nOut1_23[1] , \nOut1_23[0] }), .NORTH_EDGE({
        \nOut1_22[31] , \nOut1_22[30] , \nOut1_22[29] , \nOut1_22[28] , 
        \nOut1_22[27] , \nOut1_22[26] , \nOut1_22[25] , \nOut1_22[24] , 
        \nOut1_22[23] , \nOut1_22[22] , \nOut1_22[21] , \nOut1_22[20] , 
        \nOut1_22[19] , \nOut1_22[18] , \nOut1_22[17] , \nOut1_22[16] , 
        \nOut1_22[15] , \nOut1_22[14] , \nOut1_22[13] , \nOut1_22[12] , 
        \nOut1_22[11] , \nOut1_22[10] , \nOut1_22[9] , \nOut1_22[8] , 
        \nOut1_22[7] , \nOut1_22[6] , \nOut1_22[5] , \nOut1_22[4] , 
        \nOut1_22[3] , \nOut1_22[2] , \nOut1_22[1] , \nOut1_22[0] }), 
        .SOUTH_EDGE({\nOut1_24[31] , \nOut1_24[30] , \nOut1_24[29] , 
        \nOut1_24[28] , \nOut1_24[27] , \nOut1_24[26] , \nOut1_24[25] , 
        \nOut1_24[24] , \nOut1_24[23] , \nOut1_24[22] , \nOut1_24[21] , 
        \nOut1_24[20] , \nOut1_24[19] , \nOut1_24[18] , \nOut1_24[17] , 
        \nOut1_24[16] , \nOut1_24[15] , \nOut1_24[14] , \nOut1_24[13] , 
        \nOut1_24[12] , \nOut1_24[11] , \nOut1_24[10] , \nOut1_24[9] , 
        \nOut1_24[8] , \nOut1_24[7] , \nOut1_24[6] , \nOut1_24[5] , 
        \nOut1_24[4] , \nOut1_24[3] , \nOut1_24[2] , \nOut1_24[1] , 
        \nOut1_24[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_23[0] ), 
        .NW_EDGE(\nOut0_22[0] ), .SW_EDGE(\nOut0_24[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_113 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut114[31] , \nScanOut114[30] , \nScanOut114[29] , 
        \nScanOut114[28] , \nScanOut114[27] , \nScanOut114[26] , 
        \nScanOut114[25] , \nScanOut114[24] , \nScanOut114[23] , 
        \nScanOut114[22] , \nScanOut114[21] , \nScanOut114[20] , 
        \nScanOut114[19] , \nScanOut114[18] , \nScanOut114[17] , 
        \nScanOut114[16] , \nScanOut114[15] , \nScanOut114[14] , 
        \nScanOut114[13] , \nScanOut114[12] , \nScanOut114[11] , 
        \nScanOut114[10] , \nScanOut114[9] , \nScanOut114[8] , 
        \nScanOut114[7] , \nScanOut114[6] , \nScanOut114[5] , \nScanOut114[4] , 
        \nScanOut114[3] , \nScanOut114[2] , \nScanOut114[1] , \nScanOut114[0] 
        }), .ScanOut({\nScanOut113[31] , \nScanOut113[30] , \nScanOut113[29] , 
        \nScanOut113[28] , \nScanOut113[27] , \nScanOut113[26] , 
        \nScanOut113[25] , \nScanOut113[24] , \nScanOut113[23] , 
        \nScanOut113[22] , \nScanOut113[21] , \nScanOut113[20] , 
        \nScanOut113[19] , \nScanOut113[18] , \nScanOut113[17] , 
        \nScanOut113[16] , \nScanOut113[15] , \nScanOut113[14] , 
        \nScanOut113[13] , \nScanOut113[12] , \nScanOut113[11] , 
        \nScanOut113[10] , \nScanOut113[9] , \nScanOut113[8] , 
        \nScanOut113[7] , \nScanOut113[6] , \nScanOut113[5] , \nScanOut113[4] , 
        \nScanOut113[3] , \nScanOut113[2] , \nScanOut113[1] , \nScanOut113[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_49[31] , \nOut1_49[30] , \nOut1_49[29] , 
        \nOut1_49[28] , \nOut1_49[27] , \nOut1_49[26] , \nOut1_49[25] , 
        \nOut1_49[24] , \nOut1_49[23] , \nOut1_49[22] , \nOut1_49[21] , 
        \nOut1_49[20] , \nOut1_49[19] , \nOut1_49[18] , \nOut1_49[17] , 
        \nOut1_49[16] , \nOut1_49[15] , \nOut1_49[14] , \nOut1_49[13] , 
        \nOut1_49[12] , \nOut1_49[11] , \nOut1_49[10] , \nOut1_49[9] , 
        \nOut1_49[8] , \nOut1_49[7] , \nOut1_49[6] , \nOut1_49[5] , 
        \nOut1_49[4] , \nOut1_49[3] , \nOut1_49[2] , \nOut1_49[1] , 
        \nOut1_49[0] }), .NORTH_EDGE({\nOut1_48[31] , \nOut1_48[30] , 
        \nOut1_48[29] , \nOut1_48[28] , \nOut1_48[27] , \nOut1_48[26] , 
        \nOut1_48[25] , \nOut1_48[24] , \nOut1_48[23] , \nOut1_48[22] , 
        \nOut1_48[21] , \nOut1_48[20] , \nOut1_48[19] , \nOut1_48[18] , 
        \nOut1_48[17] , \nOut1_48[16] , \nOut1_48[15] , \nOut1_48[14] , 
        \nOut1_48[13] , \nOut1_48[12] , \nOut1_48[11] , \nOut1_48[10] , 
        \nOut1_48[9] , \nOut1_48[8] , \nOut1_48[7] , \nOut1_48[6] , 
        \nOut1_48[5] , \nOut1_48[4] , \nOut1_48[3] , \nOut1_48[2] , 
        \nOut1_48[1] , \nOut1_48[0] }), .SOUTH_EDGE({\nOut1_50[31] , 
        \nOut1_50[30] , \nOut1_50[29] , \nOut1_50[28] , \nOut1_50[27] , 
        \nOut1_50[26] , \nOut1_50[25] , \nOut1_50[24] , \nOut1_50[23] , 
        \nOut1_50[22] , \nOut1_50[21] , \nOut1_50[20] , \nOut1_50[19] , 
        \nOut1_50[18] , \nOut1_50[17] , \nOut1_50[16] , \nOut1_50[15] , 
        \nOut1_50[14] , \nOut1_50[13] , \nOut1_50[12] , \nOut1_50[11] , 
        \nOut1_50[10] , \nOut1_50[9] , \nOut1_50[8] , \nOut1_50[7] , 
        \nOut1_50[6] , \nOut1_50[5] , \nOut1_50[4] , \nOut1_50[3] , 
        \nOut1_50[2] , \nOut1_50[1] , \nOut1_50[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_49[0] ), .NW_EDGE(\nOut0_48[0] ), .SW_EDGE(
        \nOut0_50[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_114 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut115[31] , \nScanOut115[30] , \nScanOut115[29] , 
        \nScanOut115[28] , \nScanOut115[27] , \nScanOut115[26] , 
        \nScanOut115[25] , \nScanOut115[24] , \nScanOut115[23] , 
        \nScanOut115[22] , \nScanOut115[21] , \nScanOut115[20] , 
        \nScanOut115[19] , \nScanOut115[18] , \nScanOut115[17] , 
        \nScanOut115[16] , \nScanOut115[15] , \nScanOut115[14] , 
        \nScanOut115[13] , \nScanOut115[12] , \nScanOut115[11] , 
        \nScanOut115[10] , \nScanOut115[9] , \nScanOut115[8] , 
        \nScanOut115[7] , \nScanOut115[6] , \nScanOut115[5] , \nScanOut115[4] , 
        \nScanOut115[3] , \nScanOut115[2] , \nScanOut115[1] , \nScanOut115[0] 
        }), .ScanOut({\nScanOut114[31] , \nScanOut114[30] , \nScanOut114[29] , 
        \nScanOut114[28] , \nScanOut114[27] , \nScanOut114[26] , 
        \nScanOut114[25] , \nScanOut114[24] , \nScanOut114[23] , 
        \nScanOut114[22] , \nScanOut114[21] , \nScanOut114[20] , 
        \nScanOut114[19] , \nScanOut114[18] , \nScanOut114[17] , 
        \nScanOut114[16] , \nScanOut114[15] , \nScanOut114[14] , 
        \nScanOut114[13] , \nScanOut114[12] , \nScanOut114[11] , 
        \nScanOut114[10] , \nScanOut114[9] , \nScanOut114[8] , 
        \nScanOut114[7] , \nScanOut114[6] , \nScanOut114[5] , \nScanOut114[4] , 
        \nScanOut114[3] , \nScanOut114[2] , \nScanOut114[1] , \nScanOut114[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_50[31] , \nOut1_50[30] , \nOut1_50[29] , 
        \nOut1_50[28] , \nOut1_50[27] , \nOut1_50[26] , \nOut1_50[25] , 
        \nOut1_50[24] , \nOut1_50[23] , \nOut1_50[22] , \nOut1_50[21] , 
        \nOut1_50[20] , \nOut1_50[19] , \nOut1_50[18] , \nOut1_50[17] , 
        \nOut1_50[16] , \nOut1_50[15] , \nOut1_50[14] , \nOut1_50[13] , 
        \nOut1_50[12] , \nOut1_50[11] , \nOut1_50[10] , \nOut1_50[9] , 
        \nOut1_50[8] , \nOut1_50[7] , \nOut1_50[6] , \nOut1_50[5] , 
        \nOut1_50[4] , \nOut1_50[3] , \nOut1_50[2] , \nOut1_50[1] , 
        \nOut1_50[0] }), .NORTH_EDGE({\nOut1_49[31] , \nOut1_49[30] , 
        \nOut1_49[29] , \nOut1_49[28] , \nOut1_49[27] , \nOut1_49[26] , 
        \nOut1_49[25] , \nOut1_49[24] , \nOut1_49[23] , \nOut1_49[22] , 
        \nOut1_49[21] , \nOut1_49[20] , \nOut1_49[19] , \nOut1_49[18] , 
        \nOut1_49[17] , \nOut1_49[16] , \nOut1_49[15] , \nOut1_49[14] , 
        \nOut1_49[13] , \nOut1_49[12] , \nOut1_49[11] , \nOut1_49[10] , 
        \nOut1_49[9] , \nOut1_49[8] , \nOut1_49[7] , \nOut1_49[6] , 
        \nOut1_49[5] , \nOut1_49[4] , \nOut1_49[3] , \nOut1_49[2] , 
        \nOut1_49[1] , \nOut1_49[0] }), .SOUTH_EDGE({\nOut1_51[31] , 
        \nOut1_51[30] , \nOut1_51[29] , \nOut1_51[28] , \nOut1_51[27] , 
        \nOut1_51[26] , \nOut1_51[25] , \nOut1_51[24] , \nOut1_51[23] , 
        \nOut1_51[22] , \nOut1_51[21] , \nOut1_51[20] , \nOut1_51[19] , 
        \nOut1_51[18] , \nOut1_51[17] , \nOut1_51[16] , \nOut1_51[15] , 
        \nOut1_51[14] , \nOut1_51[13] , \nOut1_51[12] , \nOut1_51[11] , 
        \nOut1_51[10] , \nOut1_51[9] , \nOut1_51[8] , \nOut1_51[7] , 
        \nOut1_51[6] , \nOut1_51[5] , \nOut1_51[4] , \nOut1_51[3] , 
        \nOut1_51[2] , \nOut1_51[1] , \nOut1_51[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_50[0] ), .NW_EDGE(\nOut0_49[0] ), .SW_EDGE(
        \nOut0_51[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_59 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut60[31] , \nScanOut60[30] , \nScanOut60[29] , 
        \nScanOut60[28] , \nScanOut60[27] , \nScanOut60[26] , \nScanOut60[25] , 
        \nScanOut60[24] , \nScanOut60[23] , \nScanOut60[22] , \nScanOut60[21] , 
        \nScanOut60[20] , \nScanOut60[19] , \nScanOut60[18] , \nScanOut60[17] , 
        \nScanOut60[16] , \nScanOut60[15] , \nScanOut60[14] , \nScanOut60[13] , 
        \nScanOut60[12] , \nScanOut60[11] , \nScanOut60[10] , \nScanOut60[9] , 
        \nScanOut60[8] , \nScanOut60[7] , \nScanOut60[6] , \nScanOut60[5] , 
        \nScanOut60[4] , \nScanOut60[3] , \nScanOut60[2] , \nScanOut60[1] , 
        \nScanOut60[0] }), .ScanOut({\nScanOut59[31] , \nScanOut59[30] , 
        \nScanOut59[29] , \nScanOut59[28] , \nScanOut59[27] , \nScanOut59[26] , 
        \nScanOut59[25] , \nScanOut59[24] , \nScanOut59[23] , \nScanOut59[22] , 
        \nScanOut59[21] , \nScanOut59[20] , \nScanOut59[19] , \nScanOut59[18] , 
        \nScanOut59[17] , \nScanOut59[16] , \nScanOut59[15] , \nScanOut59[14] , 
        \nScanOut59[13] , \nScanOut59[12] , \nScanOut59[11] , \nScanOut59[10] , 
        \nScanOut59[9] , \nScanOut59[8] , \nScanOut59[7] , \nScanOut59[6] , 
        \nScanOut59[5] , \nScanOut59[4] , \nScanOut59[3] , \nScanOut59[2] , 
        \nScanOut59[1] , \nScanOut59[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_59[31] , 
        \nOut0_59[30] , \nOut0_59[29] , \nOut0_59[28] , \nOut0_59[27] , 
        \nOut0_59[26] , \nOut0_59[25] , \nOut0_59[24] , \nOut0_59[23] , 
        \nOut0_59[22] , \nOut0_59[21] , \nOut0_59[20] , \nOut0_59[19] , 
        \nOut0_59[18] , \nOut0_59[17] , \nOut0_59[16] , \nOut0_59[15] , 
        \nOut0_59[14] , \nOut0_59[13] , \nOut0_59[12] , \nOut0_59[11] , 
        \nOut0_59[10] , \nOut0_59[9] , \nOut0_59[8] , \nOut0_59[7] , 
        \nOut0_59[6] , \nOut0_59[5] , \nOut0_59[4] , \nOut0_59[3] , 
        \nOut0_59[2] , \nOut0_59[1] , \nOut0_59[0] }), .NORTH_EDGE({
        \nOut0_58[31] , \nOut0_58[30] , \nOut0_58[29] , \nOut0_58[28] , 
        \nOut0_58[27] , \nOut0_58[26] , \nOut0_58[25] , \nOut0_58[24] , 
        \nOut0_58[23] , \nOut0_58[22] , \nOut0_58[21] , \nOut0_58[20] , 
        \nOut0_58[19] , \nOut0_58[18] , \nOut0_58[17] , \nOut0_58[16] , 
        \nOut0_58[15] , \nOut0_58[14] , \nOut0_58[13] , \nOut0_58[12] , 
        \nOut0_58[11] , \nOut0_58[10] , \nOut0_58[9] , \nOut0_58[8] , 
        \nOut0_58[7] , \nOut0_58[6] , \nOut0_58[5] , \nOut0_58[4] , 
        \nOut0_58[3] , \nOut0_58[2] , \nOut0_58[1] , \nOut0_58[0] }), 
        .SOUTH_EDGE({\nOut0_60[31] , \nOut0_60[30] , \nOut0_60[29] , 
        \nOut0_60[28] , \nOut0_60[27] , \nOut0_60[26] , \nOut0_60[25] , 
        \nOut0_60[24] , \nOut0_60[23] , \nOut0_60[22] , \nOut0_60[21] , 
        \nOut0_60[20] , \nOut0_60[19] , \nOut0_60[18] , \nOut0_60[17] , 
        \nOut0_60[16] , \nOut0_60[15] , \nOut0_60[14] , \nOut0_60[13] , 
        \nOut0_60[12] , \nOut0_60[11] , \nOut0_60[10] , \nOut0_60[9] , 
        \nOut0_60[8] , \nOut0_60[7] , \nOut0_60[6] , \nOut0_60[5] , 
        \nOut0_60[4] , \nOut0_60[3] , \nOut0_60[2] , \nOut0_60[1] , 
        \nOut0_60[0] }), .EAST_EDGE(\nOut1_59[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_58[31] ), .SE_EDGE(
        \nOut1_60[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_65 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut66[31] , \nScanOut66[30] , \nScanOut66[29] , 
        \nScanOut66[28] , \nScanOut66[27] , \nScanOut66[26] , \nScanOut66[25] , 
        \nScanOut66[24] , \nScanOut66[23] , \nScanOut66[22] , \nScanOut66[21] , 
        \nScanOut66[20] , \nScanOut66[19] , \nScanOut66[18] , \nScanOut66[17] , 
        \nScanOut66[16] , \nScanOut66[15] , \nScanOut66[14] , \nScanOut66[13] , 
        \nScanOut66[12] , \nScanOut66[11] , \nScanOut66[10] , \nScanOut66[9] , 
        \nScanOut66[8] , \nScanOut66[7] , \nScanOut66[6] , \nScanOut66[5] , 
        \nScanOut66[4] , \nScanOut66[3] , \nScanOut66[2] , \nScanOut66[1] , 
        \nScanOut66[0] }), .ScanOut({\nScanOut65[31] , \nScanOut65[30] , 
        \nScanOut65[29] , \nScanOut65[28] , \nScanOut65[27] , \nScanOut65[26] , 
        \nScanOut65[25] , \nScanOut65[24] , \nScanOut65[23] , \nScanOut65[22] , 
        \nScanOut65[21] , \nScanOut65[20] , \nScanOut65[19] , \nScanOut65[18] , 
        \nScanOut65[17] , \nScanOut65[16] , \nScanOut65[15] , \nScanOut65[14] , 
        \nScanOut65[13] , \nScanOut65[12] , \nScanOut65[11] , \nScanOut65[10] , 
        \nScanOut65[9] , \nScanOut65[8] , \nScanOut65[7] , \nScanOut65[6] , 
        \nScanOut65[5] , \nScanOut65[4] , \nScanOut65[3] , \nScanOut65[2] , 
        \nScanOut65[1] , \nScanOut65[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_1[31] , 
        \nOut1_1[30] , \nOut1_1[29] , \nOut1_1[28] , \nOut1_1[27] , 
        \nOut1_1[26] , \nOut1_1[25] , \nOut1_1[24] , \nOut1_1[23] , 
        \nOut1_1[22] , \nOut1_1[21] , \nOut1_1[20] , \nOut1_1[19] , 
        \nOut1_1[18] , \nOut1_1[17] , \nOut1_1[16] , \nOut1_1[15] , 
        \nOut1_1[14] , \nOut1_1[13] , \nOut1_1[12] , \nOut1_1[11] , 
        \nOut1_1[10] , \nOut1_1[9] , \nOut1_1[8] , \nOut1_1[7] , \nOut1_1[6] , 
        \nOut1_1[5] , \nOut1_1[4] , \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , 
        \nOut1_1[0] }), .NORTH_EDGE({\nOut1_0[31] , \nOut1_0[30] , 
        \nOut1_0[29] , \nOut1_0[28] , \nOut1_0[27] , \nOut1_0[26] , 
        \nOut1_0[25] , \nOut1_0[24] , \nOut1_0[23] , \nOut1_0[22] , 
        \nOut1_0[21] , \nOut1_0[20] , \nOut1_0[19] , \nOut1_0[18] , 
        \nOut1_0[17] , \nOut1_0[16] , \nOut1_0[15] , \nOut1_0[14] , 
        \nOut1_0[13] , \nOut1_0[12] , \nOut1_0[11] , \nOut1_0[10] , 
        \nOut1_0[9] , \nOut1_0[8] , \nOut1_0[7] , \nOut1_0[6] , \nOut1_0[5] , 
        \nOut1_0[4] , \nOut1_0[3] , \nOut1_0[2] , \nOut1_0[1] , \nOut1_0[0] }), 
        .SOUTH_EDGE({\nOut1_2[31] , \nOut1_2[30] , \nOut1_2[29] , 
        \nOut1_2[28] , \nOut1_2[27] , \nOut1_2[26] , \nOut1_2[25] , 
        \nOut1_2[24] , \nOut1_2[23] , \nOut1_2[22] , \nOut1_2[21] , 
        \nOut1_2[20] , \nOut1_2[19] , \nOut1_2[18] , \nOut1_2[17] , 
        \nOut1_2[16] , \nOut1_2[15] , \nOut1_2[14] , \nOut1_2[13] , 
        \nOut1_2[12] , \nOut1_2[11] , \nOut1_2[10] , \nOut1_2[9] , 
        \nOut1_2[8] , \nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , 
        \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_1[0] ), .NW_EDGE(\nOut0_0[0] ), .SW_EDGE(
        \nOut0_2[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_25 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut26[31] , \nScanOut26[30] , \nScanOut26[29] , 
        \nScanOut26[28] , \nScanOut26[27] , \nScanOut26[26] , \nScanOut26[25] , 
        \nScanOut26[24] , \nScanOut26[23] , \nScanOut26[22] , \nScanOut26[21] , 
        \nScanOut26[20] , \nScanOut26[19] , \nScanOut26[18] , \nScanOut26[17] , 
        \nScanOut26[16] , \nScanOut26[15] , \nScanOut26[14] , \nScanOut26[13] , 
        \nScanOut26[12] , \nScanOut26[11] , \nScanOut26[10] , \nScanOut26[9] , 
        \nScanOut26[8] , \nScanOut26[7] , \nScanOut26[6] , \nScanOut26[5] , 
        \nScanOut26[4] , \nScanOut26[3] , \nScanOut26[2] , \nScanOut26[1] , 
        \nScanOut26[0] }), .ScanOut({\nScanOut25[31] , \nScanOut25[30] , 
        \nScanOut25[29] , \nScanOut25[28] , \nScanOut25[27] , \nScanOut25[26] , 
        \nScanOut25[25] , \nScanOut25[24] , \nScanOut25[23] , \nScanOut25[22] , 
        \nScanOut25[21] , \nScanOut25[20] , \nScanOut25[19] , \nScanOut25[18] , 
        \nScanOut25[17] , \nScanOut25[16] , \nScanOut25[15] , \nScanOut25[14] , 
        \nScanOut25[13] , \nScanOut25[12] , \nScanOut25[11] , \nScanOut25[10] , 
        \nScanOut25[9] , \nScanOut25[8] , \nScanOut25[7] , \nScanOut25[6] , 
        \nScanOut25[5] , \nScanOut25[4] , \nScanOut25[3] , \nScanOut25[2] , 
        \nScanOut25[1] , \nScanOut25[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_25[31] , 
        \nOut0_25[30] , \nOut0_25[29] , \nOut0_25[28] , \nOut0_25[27] , 
        \nOut0_25[26] , \nOut0_25[25] , \nOut0_25[24] , \nOut0_25[23] , 
        \nOut0_25[22] , \nOut0_25[21] , \nOut0_25[20] , \nOut0_25[19] , 
        \nOut0_25[18] , \nOut0_25[17] , \nOut0_25[16] , \nOut0_25[15] , 
        \nOut0_25[14] , \nOut0_25[13] , \nOut0_25[12] , \nOut0_25[11] , 
        \nOut0_25[10] , \nOut0_25[9] , \nOut0_25[8] , \nOut0_25[7] , 
        \nOut0_25[6] , \nOut0_25[5] , \nOut0_25[4] , \nOut0_25[3] , 
        \nOut0_25[2] , \nOut0_25[1] , \nOut0_25[0] }), .NORTH_EDGE({
        \nOut0_24[31] , \nOut0_24[30] , \nOut0_24[29] , \nOut0_24[28] , 
        \nOut0_24[27] , \nOut0_24[26] , \nOut0_24[25] , \nOut0_24[24] , 
        \nOut0_24[23] , \nOut0_24[22] , \nOut0_24[21] , \nOut0_24[20] , 
        \nOut0_24[19] , \nOut0_24[18] , \nOut0_24[17] , \nOut0_24[16] , 
        \nOut0_24[15] , \nOut0_24[14] , \nOut0_24[13] , \nOut0_24[12] , 
        \nOut0_24[11] , \nOut0_24[10] , \nOut0_24[9] , \nOut0_24[8] , 
        \nOut0_24[7] , \nOut0_24[6] , \nOut0_24[5] , \nOut0_24[4] , 
        \nOut0_24[3] , \nOut0_24[2] , \nOut0_24[1] , \nOut0_24[0] }), 
        .SOUTH_EDGE({\nOut0_26[31] , \nOut0_26[30] , \nOut0_26[29] , 
        \nOut0_26[28] , \nOut0_26[27] , \nOut0_26[26] , \nOut0_26[25] , 
        \nOut0_26[24] , \nOut0_26[23] , \nOut0_26[22] , \nOut0_26[21] , 
        \nOut0_26[20] , \nOut0_26[19] , \nOut0_26[18] , \nOut0_26[17] , 
        \nOut0_26[16] , \nOut0_26[15] , \nOut0_26[14] , \nOut0_26[13] , 
        \nOut0_26[12] , \nOut0_26[11] , \nOut0_26[10] , \nOut0_26[9] , 
        \nOut0_26[8] , \nOut0_26[7] , \nOut0_26[6] , \nOut0_26[5] , 
        \nOut0_26[4] , \nOut0_26[3] , \nOut0_26[2] , \nOut0_26[1] , 
        \nOut0_26[0] }), .EAST_EDGE(\nOut1_25[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_24[31] ), .SE_EDGE(
        \nOut1_26[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_89 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut90[31] , \nScanOut90[30] , \nScanOut90[29] , 
        \nScanOut90[28] , \nScanOut90[27] , \nScanOut90[26] , \nScanOut90[25] , 
        \nScanOut90[24] , \nScanOut90[23] , \nScanOut90[22] , \nScanOut90[21] , 
        \nScanOut90[20] , \nScanOut90[19] , \nScanOut90[18] , \nScanOut90[17] , 
        \nScanOut90[16] , \nScanOut90[15] , \nScanOut90[14] , \nScanOut90[13] , 
        \nScanOut90[12] , \nScanOut90[11] , \nScanOut90[10] , \nScanOut90[9] , 
        \nScanOut90[8] , \nScanOut90[7] , \nScanOut90[6] , \nScanOut90[5] , 
        \nScanOut90[4] , \nScanOut90[3] , \nScanOut90[2] , \nScanOut90[1] , 
        \nScanOut90[0] }), .ScanOut({\nScanOut89[31] , \nScanOut89[30] , 
        \nScanOut89[29] , \nScanOut89[28] , \nScanOut89[27] , \nScanOut89[26] , 
        \nScanOut89[25] , \nScanOut89[24] , \nScanOut89[23] , \nScanOut89[22] , 
        \nScanOut89[21] , \nScanOut89[20] , \nScanOut89[19] , \nScanOut89[18] , 
        \nScanOut89[17] , \nScanOut89[16] , \nScanOut89[15] , \nScanOut89[14] , 
        \nScanOut89[13] , \nScanOut89[12] , \nScanOut89[11] , \nScanOut89[10] , 
        \nScanOut89[9] , \nScanOut89[8] , \nScanOut89[7] , \nScanOut89[6] , 
        \nScanOut89[5] , \nScanOut89[4] , \nScanOut89[3] , \nScanOut89[2] , 
        \nScanOut89[1] , \nScanOut89[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_25[31] , 
        \nOut1_25[30] , \nOut1_25[29] , \nOut1_25[28] , \nOut1_25[27] , 
        \nOut1_25[26] , \nOut1_25[25] , \nOut1_25[24] , \nOut1_25[23] , 
        \nOut1_25[22] , \nOut1_25[21] , \nOut1_25[20] , \nOut1_25[19] , 
        \nOut1_25[18] , \nOut1_25[17] , \nOut1_25[16] , \nOut1_25[15] , 
        \nOut1_25[14] , \nOut1_25[13] , \nOut1_25[12] , \nOut1_25[11] , 
        \nOut1_25[10] , \nOut1_25[9] , \nOut1_25[8] , \nOut1_25[7] , 
        \nOut1_25[6] , \nOut1_25[5] , \nOut1_25[4] , \nOut1_25[3] , 
        \nOut1_25[2] , \nOut1_25[1] , \nOut1_25[0] }), .NORTH_EDGE({
        \nOut1_24[31] , \nOut1_24[30] , \nOut1_24[29] , \nOut1_24[28] , 
        \nOut1_24[27] , \nOut1_24[26] , \nOut1_24[25] , \nOut1_24[24] , 
        \nOut1_24[23] , \nOut1_24[22] , \nOut1_24[21] , \nOut1_24[20] , 
        \nOut1_24[19] , \nOut1_24[18] , \nOut1_24[17] , \nOut1_24[16] , 
        \nOut1_24[15] , \nOut1_24[14] , \nOut1_24[13] , \nOut1_24[12] , 
        \nOut1_24[11] , \nOut1_24[10] , \nOut1_24[9] , \nOut1_24[8] , 
        \nOut1_24[7] , \nOut1_24[6] , \nOut1_24[5] , \nOut1_24[4] , 
        \nOut1_24[3] , \nOut1_24[2] , \nOut1_24[1] , \nOut1_24[0] }), 
        .SOUTH_EDGE({\nOut1_26[31] , \nOut1_26[30] , \nOut1_26[29] , 
        \nOut1_26[28] , \nOut1_26[27] , \nOut1_26[26] , \nOut1_26[25] , 
        \nOut1_26[24] , \nOut1_26[23] , \nOut1_26[22] , \nOut1_26[21] , 
        \nOut1_26[20] , \nOut1_26[19] , \nOut1_26[18] , \nOut1_26[17] , 
        \nOut1_26[16] , \nOut1_26[15] , \nOut1_26[14] , \nOut1_26[13] , 
        \nOut1_26[12] , \nOut1_26[11] , \nOut1_26[10] , \nOut1_26[9] , 
        \nOut1_26[8] , \nOut1_26[7] , \nOut1_26[6] , \nOut1_26[5] , 
        \nOut1_26[4] , \nOut1_26[3] , \nOut1_26[2] , \nOut1_26[1] , 
        \nOut1_26[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_25[0] ), 
        .NW_EDGE(\nOut0_24[0] ), .SW_EDGE(\nOut0_26[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut12[31] , \nScanOut12[30] , \nScanOut12[29] , 
        \nScanOut12[28] , \nScanOut12[27] , \nScanOut12[26] , \nScanOut12[25] , 
        \nScanOut12[24] , \nScanOut12[23] , \nScanOut12[22] , \nScanOut12[21] , 
        \nScanOut12[20] , \nScanOut12[19] , \nScanOut12[18] , \nScanOut12[17] , 
        \nScanOut12[16] , \nScanOut12[15] , \nScanOut12[14] , \nScanOut12[13] , 
        \nScanOut12[12] , \nScanOut12[11] , \nScanOut12[10] , \nScanOut12[9] , 
        \nScanOut12[8] , \nScanOut12[7] , \nScanOut12[6] , \nScanOut12[5] , 
        \nScanOut12[4] , \nScanOut12[3] , \nScanOut12[2] , \nScanOut12[1] , 
        \nScanOut12[0] }), .ScanOut({\nScanOut11[31] , \nScanOut11[30] , 
        \nScanOut11[29] , \nScanOut11[28] , \nScanOut11[27] , \nScanOut11[26] , 
        \nScanOut11[25] , \nScanOut11[24] , \nScanOut11[23] , \nScanOut11[22] , 
        \nScanOut11[21] , \nScanOut11[20] , \nScanOut11[19] , \nScanOut11[18] , 
        \nScanOut11[17] , \nScanOut11[16] , \nScanOut11[15] , \nScanOut11[14] , 
        \nScanOut11[13] , \nScanOut11[12] , \nScanOut11[11] , \nScanOut11[10] , 
        \nScanOut11[9] , \nScanOut11[8] , \nScanOut11[7] , \nScanOut11[6] , 
        \nScanOut11[5] , \nScanOut11[4] , \nScanOut11[3] , \nScanOut11[2] , 
        \nScanOut11[1] , \nScanOut11[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_11[31] , 
        \nOut0_11[30] , \nOut0_11[29] , \nOut0_11[28] , \nOut0_11[27] , 
        \nOut0_11[26] , \nOut0_11[25] , \nOut0_11[24] , \nOut0_11[23] , 
        \nOut0_11[22] , \nOut0_11[21] , \nOut0_11[20] , \nOut0_11[19] , 
        \nOut0_11[18] , \nOut0_11[17] , \nOut0_11[16] , \nOut0_11[15] , 
        \nOut0_11[14] , \nOut0_11[13] , \nOut0_11[12] , \nOut0_11[11] , 
        \nOut0_11[10] , \nOut0_11[9] , \nOut0_11[8] , \nOut0_11[7] , 
        \nOut0_11[6] , \nOut0_11[5] , \nOut0_11[4] , \nOut0_11[3] , 
        \nOut0_11[2] , \nOut0_11[1] , \nOut0_11[0] }), .NORTH_EDGE({
        \nOut0_10[31] , \nOut0_10[30] , \nOut0_10[29] , \nOut0_10[28] , 
        \nOut0_10[27] , \nOut0_10[26] , \nOut0_10[25] , \nOut0_10[24] , 
        \nOut0_10[23] , \nOut0_10[22] , \nOut0_10[21] , \nOut0_10[20] , 
        \nOut0_10[19] , \nOut0_10[18] , \nOut0_10[17] , \nOut0_10[16] , 
        \nOut0_10[15] , \nOut0_10[14] , \nOut0_10[13] , \nOut0_10[12] , 
        \nOut0_10[11] , \nOut0_10[10] , \nOut0_10[9] , \nOut0_10[8] , 
        \nOut0_10[7] , \nOut0_10[6] , \nOut0_10[5] , \nOut0_10[4] , 
        \nOut0_10[3] , \nOut0_10[2] , \nOut0_10[1] , \nOut0_10[0] }), 
        .SOUTH_EDGE({\nOut0_12[31] , \nOut0_12[30] , \nOut0_12[29] , 
        \nOut0_12[28] , \nOut0_12[27] , \nOut0_12[26] , \nOut0_12[25] , 
        \nOut0_12[24] , \nOut0_12[23] , \nOut0_12[22] , \nOut0_12[21] , 
        \nOut0_12[20] , \nOut0_12[19] , \nOut0_12[18] , \nOut0_12[17] , 
        \nOut0_12[16] , \nOut0_12[15] , \nOut0_12[14] , \nOut0_12[13] , 
        \nOut0_12[12] , \nOut0_12[11] , \nOut0_12[10] , \nOut0_12[9] , 
        \nOut0_12[8] , \nOut0_12[7] , \nOut0_12[6] , \nOut0_12[5] , 
        \nOut0_12[4] , \nOut0_12[3] , \nOut0_12[2] , \nOut0_12[1] , 
        \nOut0_12[0] }), .EAST_EDGE(\nOut1_11[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_10[31] ), .SE_EDGE(
        \nOut1_12[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_19 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut20[31] , \nScanOut20[30] , \nScanOut20[29] , 
        \nScanOut20[28] , \nScanOut20[27] , \nScanOut20[26] , \nScanOut20[25] , 
        \nScanOut20[24] , \nScanOut20[23] , \nScanOut20[22] , \nScanOut20[21] , 
        \nScanOut20[20] , \nScanOut20[19] , \nScanOut20[18] , \nScanOut20[17] , 
        \nScanOut20[16] , \nScanOut20[15] , \nScanOut20[14] , \nScanOut20[13] , 
        \nScanOut20[12] , \nScanOut20[11] , \nScanOut20[10] , \nScanOut20[9] , 
        \nScanOut20[8] , \nScanOut20[7] , \nScanOut20[6] , \nScanOut20[5] , 
        \nScanOut20[4] , \nScanOut20[3] , \nScanOut20[2] , \nScanOut20[1] , 
        \nScanOut20[0] }), .ScanOut({\nScanOut19[31] , \nScanOut19[30] , 
        \nScanOut19[29] , \nScanOut19[28] , \nScanOut19[27] , \nScanOut19[26] , 
        \nScanOut19[25] , \nScanOut19[24] , \nScanOut19[23] , \nScanOut19[22] , 
        \nScanOut19[21] , \nScanOut19[20] , \nScanOut19[19] , \nScanOut19[18] , 
        \nScanOut19[17] , \nScanOut19[16] , \nScanOut19[15] , \nScanOut19[14] , 
        \nScanOut19[13] , \nScanOut19[12] , \nScanOut19[11] , \nScanOut19[10] , 
        \nScanOut19[9] , \nScanOut19[8] , \nScanOut19[7] , \nScanOut19[6] , 
        \nScanOut19[5] , \nScanOut19[4] , \nScanOut19[3] , \nScanOut19[2] , 
        \nScanOut19[1] , \nScanOut19[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_19[31] , 
        \nOut0_19[30] , \nOut0_19[29] , \nOut0_19[28] , \nOut0_19[27] , 
        \nOut0_19[26] , \nOut0_19[25] , \nOut0_19[24] , \nOut0_19[23] , 
        \nOut0_19[22] , \nOut0_19[21] , \nOut0_19[20] , \nOut0_19[19] , 
        \nOut0_19[18] , \nOut0_19[17] , \nOut0_19[16] , \nOut0_19[15] , 
        \nOut0_19[14] , \nOut0_19[13] , \nOut0_19[12] , \nOut0_19[11] , 
        \nOut0_19[10] , \nOut0_19[9] , \nOut0_19[8] , \nOut0_19[7] , 
        \nOut0_19[6] , \nOut0_19[5] , \nOut0_19[4] , \nOut0_19[3] , 
        \nOut0_19[2] , \nOut0_19[1] , \nOut0_19[0] }), .NORTH_EDGE({
        \nOut0_18[31] , \nOut0_18[30] , \nOut0_18[29] , \nOut0_18[28] , 
        \nOut0_18[27] , \nOut0_18[26] , \nOut0_18[25] , \nOut0_18[24] , 
        \nOut0_18[23] , \nOut0_18[22] , \nOut0_18[21] , \nOut0_18[20] , 
        \nOut0_18[19] , \nOut0_18[18] , \nOut0_18[17] , \nOut0_18[16] , 
        \nOut0_18[15] , \nOut0_18[14] , \nOut0_18[13] , \nOut0_18[12] , 
        \nOut0_18[11] , \nOut0_18[10] , \nOut0_18[9] , \nOut0_18[8] , 
        \nOut0_18[7] , \nOut0_18[6] , \nOut0_18[5] , \nOut0_18[4] , 
        \nOut0_18[3] , \nOut0_18[2] , \nOut0_18[1] , \nOut0_18[0] }), 
        .SOUTH_EDGE({\nOut0_20[31] , \nOut0_20[30] , \nOut0_20[29] , 
        \nOut0_20[28] , \nOut0_20[27] , \nOut0_20[26] , \nOut0_20[25] , 
        \nOut0_20[24] , \nOut0_20[23] , \nOut0_20[22] , \nOut0_20[21] , 
        \nOut0_20[20] , \nOut0_20[19] , \nOut0_20[18] , \nOut0_20[17] , 
        \nOut0_20[16] , \nOut0_20[15] , \nOut0_20[14] , \nOut0_20[13] , 
        \nOut0_20[12] , \nOut0_20[11] , \nOut0_20[10] , \nOut0_20[9] , 
        \nOut0_20[8] , \nOut0_20[7] , \nOut0_20[6] , \nOut0_20[5] , 
        \nOut0_20[4] , \nOut0_20[3] , \nOut0_20[2] , \nOut0_20[1] , 
        \nOut0_20[0] }), .EAST_EDGE(\nOut1_19[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_18[31] ), .SE_EDGE(
        \nOut1_20[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_50 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut51[31] , \nScanOut51[30] , \nScanOut51[29] , 
        \nScanOut51[28] , \nScanOut51[27] , \nScanOut51[26] , \nScanOut51[25] , 
        \nScanOut51[24] , \nScanOut51[23] , \nScanOut51[22] , \nScanOut51[21] , 
        \nScanOut51[20] , \nScanOut51[19] , \nScanOut51[18] , \nScanOut51[17] , 
        \nScanOut51[16] , \nScanOut51[15] , \nScanOut51[14] , \nScanOut51[13] , 
        \nScanOut51[12] , \nScanOut51[11] , \nScanOut51[10] , \nScanOut51[9] , 
        \nScanOut51[8] , \nScanOut51[7] , \nScanOut51[6] , \nScanOut51[5] , 
        \nScanOut51[4] , \nScanOut51[3] , \nScanOut51[2] , \nScanOut51[1] , 
        \nScanOut51[0] }), .ScanOut({\nScanOut50[31] , \nScanOut50[30] , 
        \nScanOut50[29] , \nScanOut50[28] , \nScanOut50[27] , \nScanOut50[26] , 
        \nScanOut50[25] , \nScanOut50[24] , \nScanOut50[23] , \nScanOut50[22] , 
        \nScanOut50[21] , \nScanOut50[20] , \nScanOut50[19] , \nScanOut50[18] , 
        \nScanOut50[17] , \nScanOut50[16] , \nScanOut50[15] , \nScanOut50[14] , 
        \nScanOut50[13] , \nScanOut50[12] , \nScanOut50[11] , \nScanOut50[10] , 
        \nScanOut50[9] , \nScanOut50[8] , \nScanOut50[7] , \nScanOut50[6] , 
        \nScanOut50[5] , \nScanOut50[4] , \nScanOut50[3] , \nScanOut50[2] , 
        \nScanOut50[1] , \nScanOut50[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_50[31] , 
        \nOut0_50[30] , \nOut0_50[29] , \nOut0_50[28] , \nOut0_50[27] , 
        \nOut0_50[26] , \nOut0_50[25] , \nOut0_50[24] , \nOut0_50[23] , 
        \nOut0_50[22] , \nOut0_50[21] , \nOut0_50[20] , \nOut0_50[19] , 
        \nOut0_50[18] , \nOut0_50[17] , \nOut0_50[16] , \nOut0_50[15] , 
        \nOut0_50[14] , \nOut0_50[13] , \nOut0_50[12] , \nOut0_50[11] , 
        \nOut0_50[10] , \nOut0_50[9] , \nOut0_50[8] , \nOut0_50[7] , 
        \nOut0_50[6] , \nOut0_50[5] , \nOut0_50[4] , \nOut0_50[3] , 
        \nOut0_50[2] , \nOut0_50[1] , \nOut0_50[0] }), .NORTH_EDGE({
        \nOut0_49[31] , \nOut0_49[30] , \nOut0_49[29] , \nOut0_49[28] , 
        \nOut0_49[27] , \nOut0_49[26] , \nOut0_49[25] , \nOut0_49[24] , 
        \nOut0_49[23] , \nOut0_49[22] , \nOut0_49[21] , \nOut0_49[20] , 
        \nOut0_49[19] , \nOut0_49[18] , \nOut0_49[17] , \nOut0_49[16] , 
        \nOut0_49[15] , \nOut0_49[14] , \nOut0_49[13] , \nOut0_49[12] , 
        \nOut0_49[11] , \nOut0_49[10] , \nOut0_49[9] , \nOut0_49[8] , 
        \nOut0_49[7] , \nOut0_49[6] , \nOut0_49[5] , \nOut0_49[4] , 
        \nOut0_49[3] , \nOut0_49[2] , \nOut0_49[1] , \nOut0_49[0] }), 
        .SOUTH_EDGE({\nOut0_51[31] , \nOut0_51[30] , \nOut0_51[29] , 
        \nOut0_51[28] , \nOut0_51[27] , \nOut0_51[26] , \nOut0_51[25] , 
        \nOut0_51[24] , \nOut0_51[23] , \nOut0_51[22] , \nOut0_51[21] , 
        \nOut0_51[20] , \nOut0_51[19] , \nOut0_51[18] , \nOut0_51[17] , 
        \nOut0_51[16] , \nOut0_51[15] , \nOut0_51[14] , \nOut0_51[13] , 
        \nOut0_51[12] , \nOut0_51[11] , \nOut0_51[10] , \nOut0_51[9] , 
        \nOut0_51[8] , \nOut0_51[7] , \nOut0_51[6] , \nOut0_51[5] , 
        \nOut0_51[4] , \nOut0_51[3] , \nOut0_51[2] , \nOut0_51[1] , 
        \nOut0_51[0] }), .EAST_EDGE(\nOut1_50[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_49[31] ), .SE_EDGE(
        \nOut1_51[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_106 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut107[31] , \nScanOut107[30] , \nScanOut107[29] , 
        \nScanOut107[28] , \nScanOut107[27] , \nScanOut107[26] , 
        \nScanOut107[25] , \nScanOut107[24] , \nScanOut107[23] , 
        \nScanOut107[22] , \nScanOut107[21] , \nScanOut107[20] , 
        \nScanOut107[19] , \nScanOut107[18] , \nScanOut107[17] , 
        \nScanOut107[16] , \nScanOut107[15] , \nScanOut107[14] , 
        \nScanOut107[13] , \nScanOut107[12] , \nScanOut107[11] , 
        \nScanOut107[10] , \nScanOut107[9] , \nScanOut107[8] , 
        \nScanOut107[7] , \nScanOut107[6] , \nScanOut107[5] , \nScanOut107[4] , 
        \nScanOut107[3] , \nScanOut107[2] , \nScanOut107[1] , \nScanOut107[0] 
        }), .ScanOut({\nScanOut106[31] , \nScanOut106[30] , \nScanOut106[29] , 
        \nScanOut106[28] , \nScanOut106[27] , \nScanOut106[26] , 
        \nScanOut106[25] , \nScanOut106[24] , \nScanOut106[23] , 
        \nScanOut106[22] , \nScanOut106[21] , \nScanOut106[20] , 
        \nScanOut106[19] , \nScanOut106[18] , \nScanOut106[17] , 
        \nScanOut106[16] , \nScanOut106[15] , \nScanOut106[14] , 
        \nScanOut106[13] , \nScanOut106[12] , \nScanOut106[11] , 
        \nScanOut106[10] , \nScanOut106[9] , \nScanOut106[8] , 
        \nScanOut106[7] , \nScanOut106[6] , \nScanOut106[5] , \nScanOut106[4] , 
        \nScanOut106[3] , \nScanOut106[2] , \nScanOut106[1] , \nScanOut106[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_42[31] , \nOut1_42[30] , \nOut1_42[29] , 
        \nOut1_42[28] , \nOut1_42[27] , \nOut1_42[26] , \nOut1_42[25] , 
        \nOut1_42[24] , \nOut1_42[23] , \nOut1_42[22] , \nOut1_42[21] , 
        \nOut1_42[20] , \nOut1_42[19] , \nOut1_42[18] , \nOut1_42[17] , 
        \nOut1_42[16] , \nOut1_42[15] , \nOut1_42[14] , \nOut1_42[13] , 
        \nOut1_42[12] , \nOut1_42[11] , \nOut1_42[10] , \nOut1_42[9] , 
        \nOut1_42[8] , \nOut1_42[7] , \nOut1_42[6] , \nOut1_42[5] , 
        \nOut1_42[4] , \nOut1_42[3] , \nOut1_42[2] , \nOut1_42[1] , 
        \nOut1_42[0] }), .NORTH_EDGE({\nOut1_41[31] , \nOut1_41[30] , 
        \nOut1_41[29] , \nOut1_41[28] , \nOut1_41[27] , \nOut1_41[26] , 
        \nOut1_41[25] , \nOut1_41[24] , \nOut1_41[23] , \nOut1_41[22] , 
        \nOut1_41[21] , \nOut1_41[20] , \nOut1_41[19] , \nOut1_41[18] , 
        \nOut1_41[17] , \nOut1_41[16] , \nOut1_41[15] , \nOut1_41[14] , 
        \nOut1_41[13] , \nOut1_41[12] , \nOut1_41[11] , \nOut1_41[10] , 
        \nOut1_41[9] , \nOut1_41[8] , \nOut1_41[7] , \nOut1_41[6] , 
        \nOut1_41[5] , \nOut1_41[4] , \nOut1_41[3] , \nOut1_41[2] , 
        \nOut1_41[1] , \nOut1_41[0] }), .SOUTH_EDGE({\nOut1_43[31] , 
        \nOut1_43[30] , \nOut1_43[29] , \nOut1_43[28] , \nOut1_43[27] , 
        \nOut1_43[26] , \nOut1_43[25] , \nOut1_43[24] , \nOut1_43[23] , 
        \nOut1_43[22] , \nOut1_43[21] , \nOut1_43[20] , \nOut1_43[19] , 
        \nOut1_43[18] , \nOut1_43[17] , \nOut1_43[16] , \nOut1_43[15] , 
        \nOut1_43[14] , \nOut1_43[13] , \nOut1_43[12] , \nOut1_43[11] , 
        \nOut1_43[10] , \nOut1_43[9] , \nOut1_43[8] , \nOut1_43[7] , 
        \nOut1_43[6] , \nOut1_43[5] , \nOut1_43[4] , \nOut1_43[3] , 
        \nOut1_43[2] , \nOut1_43[1] , \nOut1_43[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_42[0] ), .NW_EDGE(\nOut0_41[0] ), .SW_EDGE(
        \nOut0_43[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_77 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut78[31] , \nScanOut78[30] , \nScanOut78[29] , 
        \nScanOut78[28] , \nScanOut78[27] , \nScanOut78[26] , \nScanOut78[25] , 
        \nScanOut78[24] , \nScanOut78[23] , \nScanOut78[22] , \nScanOut78[21] , 
        \nScanOut78[20] , \nScanOut78[19] , \nScanOut78[18] , \nScanOut78[17] , 
        \nScanOut78[16] , \nScanOut78[15] , \nScanOut78[14] , \nScanOut78[13] , 
        \nScanOut78[12] , \nScanOut78[11] , \nScanOut78[10] , \nScanOut78[9] , 
        \nScanOut78[8] , \nScanOut78[7] , \nScanOut78[6] , \nScanOut78[5] , 
        \nScanOut78[4] , \nScanOut78[3] , \nScanOut78[2] , \nScanOut78[1] , 
        \nScanOut78[0] }), .ScanOut({\nScanOut77[31] , \nScanOut77[30] , 
        \nScanOut77[29] , \nScanOut77[28] , \nScanOut77[27] , \nScanOut77[26] , 
        \nScanOut77[25] , \nScanOut77[24] , \nScanOut77[23] , \nScanOut77[22] , 
        \nScanOut77[21] , \nScanOut77[20] , \nScanOut77[19] , \nScanOut77[18] , 
        \nScanOut77[17] , \nScanOut77[16] , \nScanOut77[15] , \nScanOut77[14] , 
        \nScanOut77[13] , \nScanOut77[12] , \nScanOut77[11] , \nScanOut77[10] , 
        \nScanOut77[9] , \nScanOut77[8] , \nScanOut77[7] , \nScanOut77[6] , 
        \nScanOut77[5] , \nScanOut77[4] , \nScanOut77[3] , \nScanOut77[2] , 
        \nScanOut77[1] , \nScanOut77[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_13[31] , 
        \nOut1_13[30] , \nOut1_13[29] , \nOut1_13[28] , \nOut1_13[27] , 
        \nOut1_13[26] , \nOut1_13[25] , \nOut1_13[24] , \nOut1_13[23] , 
        \nOut1_13[22] , \nOut1_13[21] , \nOut1_13[20] , \nOut1_13[19] , 
        \nOut1_13[18] , \nOut1_13[17] , \nOut1_13[16] , \nOut1_13[15] , 
        \nOut1_13[14] , \nOut1_13[13] , \nOut1_13[12] , \nOut1_13[11] , 
        \nOut1_13[10] , \nOut1_13[9] , \nOut1_13[8] , \nOut1_13[7] , 
        \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , \nOut1_13[3] , 
        \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), .NORTH_EDGE({
        \nOut1_12[31] , \nOut1_12[30] , \nOut1_12[29] , \nOut1_12[28] , 
        \nOut1_12[27] , \nOut1_12[26] , \nOut1_12[25] , \nOut1_12[24] , 
        \nOut1_12[23] , \nOut1_12[22] , \nOut1_12[21] , \nOut1_12[20] , 
        \nOut1_12[19] , \nOut1_12[18] , \nOut1_12[17] , \nOut1_12[16] , 
        \nOut1_12[15] , \nOut1_12[14] , \nOut1_12[13] , \nOut1_12[12] , 
        \nOut1_12[11] , \nOut1_12[10] , \nOut1_12[9] , \nOut1_12[8] , 
        \nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), 
        .SOUTH_EDGE({\nOut1_14[31] , \nOut1_14[30] , \nOut1_14[29] , 
        \nOut1_14[28] , \nOut1_14[27] , \nOut1_14[26] , \nOut1_14[25] , 
        \nOut1_14[24] , \nOut1_14[23] , \nOut1_14[22] , \nOut1_14[21] , 
        \nOut1_14[20] , \nOut1_14[19] , \nOut1_14[18] , \nOut1_14[17] , 
        \nOut1_14[16] , \nOut1_14[15] , \nOut1_14[14] , \nOut1_14[13] , 
        \nOut1_14[12] , \nOut1_14[11] , \nOut1_14[10] , \nOut1_14[9] , 
        \nOut1_14[8] , \nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , 
        \nOut1_14[4] , \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , 
        \nOut1_14[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_13[0] ), 
        .NW_EDGE(\nOut0_12[0] ), .SW_EDGE(\nOut0_14[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_121 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut122[31] , \nScanOut122[30] , \nScanOut122[29] , 
        \nScanOut122[28] , \nScanOut122[27] , \nScanOut122[26] , 
        \nScanOut122[25] , \nScanOut122[24] , \nScanOut122[23] , 
        \nScanOut122[22] , \nScanOut122[21] , \nScanOut122[20] , 
        \nScanOut122[19] , \nScanOut122[18] , \nScanOut122[17] , 
        \nScanOut122[16] , \nScanOut122[15] , \nScanOut122[14] , 
        \nScanOut122[13] , \nScanOut122[12] , \nScanOut122[11] , 
        \nScanOut122[10] , \nScanOut122[9] , \nScanOut122[8] , 
        \nScanOut122[7] , \nScanOut122[6] , \nScanOut122[5] , \nScanOut122[4] , 
        \nScanOut122[3] , \nScanOut122[2] , \nScanOut122[1] , \nScanOut122[0] 
        }), .ScanOut({\nScanOut121[31] , \nScanOut121[30] , \nScanOut121[29] , 
        \nScanOut121[28] , \nScanOut121[27] , \nScanOut121[26] , 
        \nScanOut121[25] , \nScanOut121[24] , \nScanOut121[23] , 
        \nScanOut121[22] , \nScanOut121[21] , \nScanOut121[20] , 
        \nScanOut121[19] , \nScanOut121[18] , \nScanOut121[17] , 
        \nScanOut121[16] , \nScanOut121[15] , \nScanOut121[14] , 
        \nScanOut121[13] , \nScanOut121[12] , \nScanOut121[11] , 
        \nScanOut121[10] , \nScanOut121[9] , \nScanOut121[8] , 
        \nScanOut121[7] , \nScanOut121[6] , \nScanOut121[5] , \nScanOut121[4] , 
        \nScanOut121[3] , \nScanOut121[2] , \nScanOut121[1] , \nScanOut121[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_57[31] , \nOut1_57[30] , \nOut1_57[29] , 
        \nOut1_57[28] , \nOut1_57[27] , \nOut1_57[26] , \nOut1_57[25] , 
        \nOut1_57[24] , \nOut1_57[23] , \nOut1_57[22] , \nOut1_57[21] , 
        \nOut1_57[20] , \nOut1_57[19] , \nOut1_57[18] , \nOut1_57[17] , 
        \nOut1_57[16] , \nOut1_57[15] , \nOut1_57[14] , \nOut1_57[13] , 
        \nOut1_57[12] , \nOut1_57[11] , \nOut1_57[10] , \nOut1_57[9] , 
        \nOut1_57[8] , \nOut1_57[7] , \nOut1_57[6] , \nOut1_57[5] , 
        \nOut1_57[4] , \nOut1_57[3] , \nOut1_57[2] , \nOut1_57[1] , 
        \nOut1_57[0] }), .NORTH_EDGE({\nOut1_56[31] , \nOut1_56[30] , 
        \nOut1_56[29] , \nOut1_56[28] , \nOut1_56[27] , \nOut1_56[26] , 
        \nOut1_56[25] , \nOut1_56[24] , \nOut1_56[23] , \nOut1_56[22] , 
        \nOut1_56[21] , \nOut1_56[20] , \nOut1_56[19] , \nOut1_56[18] , 
        \nOut1_56[17] , \nOut1_56[16] , \nOut1_56[15] , \nOut1_56[14] , 
        \nOut1_56[13] , \nOut1_56[12] , \nOut1_56[11] , \nOut1_56[10] , 
        \nOut1_56[9] , \nOut1_56[8] , \nOut1_56[7] , \nOut1_56[6] , 
        \nOut1_56[5] , \nOut1_56[4] , \nOut1_56[3] , \nOut1_56[2] , 
        \nOut1_56[1] , \nOut1_56[0] }), .SOUTH_EDGE({\nOut1_58[31] , 
        \nOut1_58[30] , \nOut1_58[29] , \nOut1_58[28] , \nOut1_58[27] , 
        \nOut1_58[26] , \nOut1_58[25] , \nOut1_58[24] , \nOut1_58[23] , 
        \nOut1_58[22] , \nOut1_58[21] , \nOut1_58[20] , \nOut1_58[19] , 
        \nOut1_58[18] , \nOut1_58[17] , \nOut1_58[16] , \nOut1_58[15] , 
        \nOut1_58[14] , \nOut1_58[13] , \nOut1_58[12] , \nOut1_58[11] , 
        \nOut1_58[10] , \nOut1_58[9] , \nOut1_58[8] , \nOut1_58[7] , 
        \nOut1_58[6] , \nOut1_58[5] , \nOut1_58[4] , \nOut1_58[3] , 
        \nOut1_58[2] , \nOut1_58[1] , \nOut1_58[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_57[0] ), .NW_EDGE(\nOut0_56[0] ), .SW_EDGE(
        \nOut0_58[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_36 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut37[31] , \nScanOut37[30] , \nScanOut37[29] , 
        \nScanOut37[28] , \nScanOut37[27] , \nScanOut37[26] , \nScanOut37[25] , 
        \nScanOut37[24] , \nScanOut37[23] , \nScanOut37[22] , \nScanOut37[21] , 
        \nScanOut37[20] , \nScanOut37[19] , \nScanOut37[18] , \nScanOut37[17] , 
        \nScanOut37[16] , \nScanOut37[15] , \nScanOut37[14] , \nScanOut37[13] , 
        \nScanOut37[12] , \nScanOut37[11] , \nScanOut37[10] , \nScanOut37[9] , 
        \nScanOut37[8] , \nScanOut37[7] , \nScanOut37[6] , \nScanOut37[5] , 
        \nScanOut37[4] , \nScanOut37[3] , \nScanOut37[2] , \nScanOut37[1] , 
        \nScanOut37[0] }), .ScanOut({\nScanOut36[31] , \nScanOut36[30] , 
        \nScanOut36[29] , \nScanOut36[28] , \nScanOut36[27] , \nScanOut36[26] , 
        \nScanOut36[25] , \nScanOut36[24] , \nScanOut36[23] , \nScanOut36[22] , 
        \nScanOut36[21] , \nScanOut36[20] , \nScanOut36[19] , \nScanOut36[18] , 
        \nScanOut36[17] , \nScanOut36[16] , \nScanOut36[15] , \nScanOut36[14] , 
        \nScanOut36[13] , \nScanOut36[12] , \nScanOut36[11] , \nScanOut36[10] , 
        \nScanOut36[9] , \nScanOut36[8] , \nScanOut36[7] , \nScanOut36[6] , 
        \nScanOut36[5] , \nScanOut36[4] , \nScanOut36[3] , \nScanOut36[2] , 
        \nScanOut36[1] , \nScanOut36[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_36[31] , 
        \nOut0_36[30] , \nOut0_36[29] , \nOut0_36[28] , \nOut0_36[27] , 
        \nOut0_36[26] , \nOut0_36[25] , \nOut0_36[24] , \nOut0_36[23] , 
        \nOut0_36[22] , \nOut0_36[21] , \nOut0_36[20] , \nOut0_36[19] , 
        \nOut0_36[18] , \nOut0_36[17] , \nOut0_36[16] , \nOut0_36[15] , 
        \nOut0_36[14] , \nOut0_36[13] , \nOut0_36[12] , \nOut0_36[11] , 
        \nOut0_36[10] , \nOut0_36[9] , \nOut0_36[8] , \nOut0_36[7] , 
        \nOut0_36[6] , \nOut0_36[5] , \nOut0_36[4] , \nOut0_36[3] , 
        \nOut0_36[2] , \nOut0_36[1] , \nOut0_36[0] }), .NORTH_EDGE({
        \nOut0_35[31] , \nOut0_35[30] , \nOut0_35[29] , \nOut0_35[28] , 
        \nOut0_35[27] , \nOut0_35[26] , \nOut0_35[25] , \nOut0_35[24] , 
        \nOut0_35[23] , \nOut0_35[22] , \nOut0_35[21] , \nOut0_35[20] , 
        \nOut0_35[19] , \nOut0_35[18] , \nOut0_35[17] , \nOut0_35[16] , 
        \nOut0_35[15] , \nOut0_35[14] , \nOut0_35[13] , \nOut0_35[12] , 
        \nOut0_35[11] , \nOut0_35[10] , \nOut0_35[9] , \nOut0_35[8] , 
        \nOut0_35[7] , \nOut0_35[6] , \nOut0_35[5] , \nOut0_35[4] , 
        \nOut0_35[3] , \nOut0_35[2] , \nOut0_35[1] , \nOut0_35[0] }), 
        .SOUTH_EDGE({\nOut0_37[31] , \nOut0_37[30] , \nOut0_37[29] , 
        \nOut0_37[28] , \nOut0_37[27] , \nOut0_37[26] , \nOut0_37[25] , 
        \nOut0_37[24] , \nOut0_37[23] , \nOut0_37[22] , \nOut0_37[21] , 
        \nOut0_37[20] , \nOut0_37[19] , \nOut0_37[18] , \nOut0_37[17] , 
        \nOut0_37[16] , \nOut0_37[15] , \nOut0_37[14] , \nOut0_37[13] , 
        \nOut0_37[12] , \nOut0_37[11] , \nOut0_37[10] , \nOut0_37[9] , 
        \nOut0_37[8] , \nOut0_37[7] , \nOut0_37[6] , \nOut0_37[5] , 
        \nOut0_37[4] , \nOut0_37[3] , \nOut0_37[2] , \nOut0_37[1] , 
        \nOut0_37[0] }), .EAST_EDGE(\nOut1_36[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_35[31] ), .SE_EDGE(
        \nOut1_37[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_92 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut93[31] , \nScanOut93[30] , \nScanOut93[29] , 
        \nScanOut93[28] , \nScanOut93[27] , \nScanOut93[26] , \nScanOut93[25] , 
        \nScanOut93[24] , \nScanOut93[23] , \nScanOut93[22] , \nScanOut93[21] , 
        \nScanOut93[20] , \nScanOut93[19] , \nScanOut93[18] , \nScanOut93[17] , 
        \nScanOut93[16] , \nScanOut93[15] , \nScanOut93[14] , \nScanOut93[13] , 
        \nScanOut93[12] , \nScanOut93[11] , \nScanOut93[10] , \nScanOut93[9] , 
        \nScanOut93[8] , \nScanOut93[7] , \nScanOut93[6] , \nScanOut93[5] , 
        \nScanOut93[4] , \nScanOut93[3] , \nScanOut93[2] , \nScanOut93[1] , 
        \nScanOut93[0] }), .ScanOut({\nScanOut92[31] , \nScanOut92[30] , 
        \nScanOut92[29] , \nScanOut92[28] , \nScanOut92[27] , \nScanOut92[26] , 
        \nScanOut92[25] , \nScanOut92[24] , \nScanOut92[23] , \nScanOut92[22] , 
        \nScanOut92[21] , \nScanOut92[20] , \nScanOut92[19] , \nScanOut92[18] , 
        \nScanOut92[17] , \nScanOut92[16] , \nScanOut92[15] , \nScanOut92[14] , 
        \nScanOut92[13] , \nScanOut92[12] , \nScanOut92[11] , \nScanOut92[10] , 
        \nScanOut92[9] , \nScanOut92[8] , \nScanOut92[7] , \nScanOut92[6] , 
        \nScanOut92[5] , \nScanOut92[4] , \nScanOut92[3] , \nScanOut92[2] , 
        \nScanOut92[1] , \nScanOut92[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_28[31] , 
        \nOut1_28[30] , \nOut1_28[29] , \nOut1_28[28] , \nOut1_28[27] , 
        \nOut1_28[26] , \nOut1_28[25] , \nOut1_28[24] , \nOut1_28[23] , 
        \nOut1_28[22] , \nOut1_28[21] , \nOut1_28[20] , \nOut1_28[19] , 
        \nOut1_28[18] , \nOut1_28[17] , \nOut1_28[16] , \nOut1_28[15] , 
        \nOut1_28[14] , \nOut1_28[13] , \nOut1_28[12] , \nOut1_28[11] , 
        \nOut1_28[10] , \nOut1_28[9] , \nOut1_28[8] , \nOut1_28[7] , 
        \nOut1_28[6] , \nOut1_28[5] , \nOut1_28[4] , \nOut1_28[3] , 
        \nOut1_28[2] , \nOut1_28[1] , \nOut1_28[0] }), .NORTH_EDGE({
        \nOut1_27[31] , \nOut1_27[30] , \nOut1_27[29] , \nOut1_27[28] , 
        \nOut1_27[27] , \nOut1_27[26] , \nOut1_27[25] , \nOut1_27[24] , 
        \nOut1_27[23] , \nOut1_27[22] , \nOut1_27[21] , \nOut1_27[20] , 
        \nOut1_27[19] , \nOut1_27[18] , \nOut1_27[17] , \nOut1_27[16] , 
        \nOut1_27[15] , \nOut1_27[14] , \nOut1_27[13] , \nOut1_27[12] , 
        \nOut1_27[11] , \nOut1_27[10] , \nOut1_27[9] , \nOut1_27[8] , 
        \nOut1_27[7] , \nOut1_27[6] , \nOut1_27[5] , \nOut1_27[4] , 
        \nOut1_27[3] , \nOut1_27[2] , \nOut1_27[1] , \nOut1_27[0] }), 
        .SOUTH_EDGE({\nOut1_29[31] , \nOut1_29[30] , \nOut1_29[29] , 
        \nOut1_29[28] , \nOut1_29[27] , \nOut1_29[26] , \nOut1_29[25] , 
        \nOut1_29[24] , \nOut1_29[23] , \nOut1_29[22] , \nOut1_29[21] , 
        \nOut1_29[20] , \nOut1_29[19] , \nOut1_29[18] , \nOut1_29[17] , 
        \nOut1_29[16] , \nOut1_29[15] , \nOut1_29[14] , \nOut1_29[13] , 
        \nOut1_29[12] , \nOut1_29[11] , \nOut1_29[10] , \nOut1_29[9] , 
        \nOut1_29[8] , \nOut1_29[7] , \nOut1_29[6] , \nOut1_29[5] , 
        \nOut1_29[4] , \nOut1_29[3] , \nOut1_29[2] , \nOut1_29[1] , 
        \nOut1_29[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_28[0] ), 
        .NW_EDGE(\nOut0_27[0] ), .SW_EDGE(\nOut0_29[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_18 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut19[31] , \nScanOut19[30] , \nScanOut19[29] , 
        \nScanOut19[28] , \nScanOut19[27] , \nScanOut19[26] , \nScanOut19[25] , 
        \nScanOut19[24] , \nScanOut19[23] , \nScanOut19[22] , \nScanOut19[21] , 
        \nScanOut19[20] , \nScanOut19[19] , \nScanOut19[18] , \nScanOut19[17] , 
        \nScanOut19[16] , \nScanOut19[15] , \nScanOut19[14] , \nScanOut19[13] , 
        \nScanOut19[12] , \nScanOut19[11] , \nScanOut19[10] , \nScanOut19[9] , 
        \nScanOut19[8] , \nScanOut19[7] , \nScanOut19[6] , \nScanOut19[5] , 
        \nScanOut19[4] , \nScanOut19[3] , \nScanOut19[2] , \nScanOut19[1] , 
        \nScanOut19[0] }), .ScanOut({\nScanOut18[31] , \nScanOut18[30] , 
        \nScanOut18[29] , \nScanOut18[28] , \nScanOut18[27] , \nScanOut18[26] , 
        \nScanOut18[25] , \nScanOut18[24] , \nScanOut18[23] , \nScanOut18[22] , 
        \nScanOut18[21] , \nScanOut18[20] , \nScanOut18[19] , \nScanOut18[18] , 
        \nScanOut18[17] , \nScanOut18[16] , \nScanOut18[15] , \nScanOut18[14] , 
        \nScanOut18[13] , \nScanOut18[12] , \nScanOut18[11] , \nScanOut18[10] , 
        \nScanOut18[9] , \nScanOut18[8] , \nScanOut18[7] , \nScanOut18[6] , 
        \nScanOut18[5] , \nScanOut18[4] , \nScanOut18[3] , \nScanOut18[2] , 
        \nScanOut18[1] , \nScanOut18[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_18[31] , 
        \nOut0_18[30] , \nOut0_18[29] , \nOut0_18[28] , \nOut0_18[27] , 
        \nOut0_18[26] , \nOut0_18[25] , \nOut0_18[24] , \nOut0_18[23] , 
        \nOut0_18[22] , \nOut0_18[21] , \nOut0_18[20] , \nOut0_18[19] , 
        \nOut0_18[18] , \nOut0_18[17] , \nOut0_18[16] , \nOut0_18[15] , 
        \nOut0_18[14] , \nOut0_18[13] , \nOut0_18[12] , \nOut0_18[11] , 
        \nOut0_18[10] , \nOut0_18[9] , \nOut0_18[8] , \nOut0_18[7] , 
        \nOut0_18[6] , \nOut0_18[5] , \nOut0_18[4] , \nOut0_18[3] , 
        \nOut0_18[2] , \nOut0_18[1] , \nOut0_18[0] }), .NORTH_EDGE({
        \nOut0_17[31] , \nOut0_17[30] , \nOut0_17[29] , \nOut0_17[28] , 
        \nOut0_17[27] , \nOut0_17[26] , \nOut0_17[25] , \nOut0_17[24] , 
        \nOut0_17[23] , \nOut0_17[22] , \nOut0_17[21] , \nOut0_17[20] , 
        \nOut0_17[19] , \nOut0_17[18] , \nOut0_17[17] , \nOut0_17[16] , 
        \nOut0_17[15] , \nOut0_17[14] , \nOut0_17[13] , \nOut0_17[12] , 
        \nOut0_17[11] , \nOut0_17[10] , \nOut0_17[9] , \nOut0_17[8] , 
        \nOut0_17[7] , \nOut0_17[6] , \nOut0_17[5] , \nOut0_17[4] , 
        \nOut0_17[3] , \nOut0_17[2] , \nOut0_17[1] , \nOut0_17[0] }), 
        .SOUTH_EDGE({\nOut0_19[31] , \nOut0_19[30] , \nOut0_19[29] , 
        \nOut0_19[28] , \nOut0_19[27] , \nOut0_19[26] , \nOut0_19[25] , 
        \nOut0_19[24] , \nOut0_19[23] , \nOut0_19[22] , \nOut0_19[21] , 
        \nOut0_19[20] , \nOut0_19[19] , \nOut0_19[18] , \nOut0_19[17] , 
        \nOut0_19[16] , \nOut0_19[15] , \nOut0_19[14] , \nOut0_19[13] , 
        \nOut0_19[12] , \nOut0_19[11] , \nOut0_19[10] , \nOut0_19[9] , 
        \nOut0_19[8] , \nOut0_19[7] , \nOut0_19[6] , \nOut0_19[5] , 
        \nOut0_19[4] , \nOut0_19[3] , \nOut0_19[2] , \nOut0_19[1] , 
        \nOut0_19[0] }), .EAST_EDGE(\nOut1_18[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_17[31] ), .SE_EDGE(
        \nOut1_19[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_43 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut44[31] , \nScanOut44[30] , \nScanOut44[29] , 
        \nScanOut44[28] , \nScanOut44[27] , \nScanOut44[26] , \nScanOut44[25] , 
        \nScanOut44[24] , \nScanOut44[23] , \nScanOut44[22] , \nScanOut44[21] , 
        \nScanOut44[20] , \nScanOut44[19] , \nScanOut44[18] , \nScanOut44[17] , 
        \nScanOut44[16] , \nScanOut44[15] , \nScanOut44[14] , \nScanOut44[13] , 
        \nScanOut44[12] , \nScanOut44[11] , \nScanOut44[10] , \nScanOut44[9] , 
        \nScanOut44[8] , \nScanOut44[7] , \nScanOut44[6] , \nScanOut44[5] , 
        \nScanOut44[4] , \nScanOut44[3] , \nScanOut44[2] , \nScanOut44[1] , 
        \nScanOut44[0] }), .ScanOut({\nScanOut43[31] , \nScanOut43[30] , 
        \nScanOut43[29] , \nScanOut43[28] , \nScanOut43[27] , \nScanOut43[26] , 
        \nScanOut43[25] , \nScanOut43[24] , \nScanOut43[23] , \nScanOut43[22] , 
        \nScanOut43[21] , \nScanOut43[20] , \nScanOut43[19] , \nScanOut43[18] , 
        \nScanOut43[17] , \nScanOut43[16] , \nScanOut43[15] , \nScanOut43[14] , 
        \nScanOut43[13] , \nScanOut43[12] , \nScanOut43[11] , \nScanOut43[10] , 
        \nScanOut43[9] , \nScanOut43[8] , \nScanOut43[7] , \nScanOut43[6] , 
        \nScanOut43[5] , \nScanOut43[4] , \nScanOut43[3] , \nScanOut43[2] , 
        \nScanOut43[1] , \nScanOut43[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_43[31] , 
        \nOut0_43[30] , \nOut0_43[29] , \nOut0_43[28] , \nOut0_43[27] , 
        \nOut0_43[26] , \nOut0_43[25] , \nOut0_43[24] , \nOut0_43[23] , 
        \nOut0_43[22] , \nOut0_43[21] , \nOut0_43[20] , \nOut0_43[19] , 
        \nOut0_43[18] , \nOut0_43[17] , \nOut0_43[16] , \nOut0_43[15] , 
        \nOut0_43[14] , \nOut0_43[13] , \nOut0_43[12] , \nOut0_43[11] , 
        \nOut0_43[10] , \nOut0_43[9] , \nOut0_43[8] , \nOut0_43[7] , 
        \nOut0_43[6] , \nOut0_43[5] , \nOut0_43[4] , \nOut0_43[3] , 
        \nOut0_43[2] , \nOut0_43[1] , \nOut0_43[0] }), .NORTH_EDGE({
        \nOut0_42[31] , \nOut0_42[30] , \nOut0_42[29] , \nOut0_42[28] , 
        \nOut0_42[27] , \nOut0_42[26] , \nOut0_42[25] , \nOut0_42[24] , 
        \nOut0_42[23] , \nOut0_42[22] , \nOut0_42[21] , \nOut0_42[20] , 
        \nOut0_42[19] , \nOut0_42[18] , \nOut0_42[17] , \nOut0_42[16] , 
        \nOut0_42[15] , \nOut0_42[14] , \nOut0_42[13] , \nOut0_42[12] , 
        \nOut0_42[11] , \nOut0_42[10] , \nOut0_42[9] , \nOut0_42[8] , 
        \nOut0_42[7] , \nOut0_42[6] , \nOut0_42[5] , \nOut0_42[4] , 
        \nOut0_42[3] , \nOut0_42[2] , \nOut0_42[1] , \nOut0_42[0] }), 
        .SOUTH_EDGE({\nOut0_44[31] , \nOut0_44[30] , \nOut0_44[29] , 
        \nOut0_44[28] , \nOut0_44[27] , \nOut0_44[26] , \nOut0_44[25] , 
        \nOut0_44[24] , \nOut0_44[23] , \nOut0_44[22] , \nOut0_44[21] , 
        \nOut0_44[20] , \nOut0_44[19] , \nOut0_44[18] , \nOut0_44[17] , 
        \nOut0_44[16] , \nOut0_44[15] , \nOut0_44[14] , \nOut0_44[13] , 
        \nOut0_44[12] , \nOut0_44[11] , \nOut0_44[10] , \nOut0_44[9] , 
        \nOut0_44[8] , \nOut0_44[7] , \nOut0_44[6] , \nOut0_44[5] , 
        \nOut0_44[4] , \nOut0_44[3] , \nOut0_44[2] , \nOut0_44[1] , 
        \nOut0_44[0] }), .EAST_EDGE(\nOut1_43[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_42[31] ), .SE_EDGE(
        \nOut1_44[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_58 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut59[31] , \nScanOut59[30] , \nScanOut59[29] , 
        \nScanOut59[28] , \nScanOut59[27] , \nScanOut59[26] , \nScanOut59[25] , 
        \nScanOut59[24] , \nScanOut59[23] , \nScanOut59[22] , \nScanOut59[21] , 
        \nScanOut59[20] , \nScanOut59[19] , \nScanOut59[18] , \nScanOut59[17] , 
        \nScanOut59[16] , \nScanOut59[15] , \nScanOut59[14] , \nScanOut59[13] , 
        \nScanOut59[12] , \nScanOut59[11] , \nScanOut59[10] , \nScanOut59[9] , 
        \nScanOut59[8] , \nScanOut59[7] , \nScanOut59[6] , \nScanOut59[5] , 
        \nScanOut59[4] , \nScanOut59[3] , \nScanOut59[2] , \nScanOut59[1] , 
        \nScanOut59[0] }), .ScanOut({\nScanOut58[31] , \nScanOut58[30] , 
        \nScanOut58[29] , \nScanOut58[28] , \nScanOut58[27] , \nScanOut58[26] , 
        \nScanOut58[25] , \nScanOut58[24] , \nScanOut58[23] , \nScanOut58[22] , 
        \nScanOut58[21] , \nScanOut58[20] , \nScanOut58[19] , \nScanOut58[18] , 
        \nScanOut58[17] , \nScanOut58[16] , \nScanOut58[15] , \nScanOut58[14] , 
        \nScanOut58[13] , \nScanOut58[12] , \nScanOut58[11] , \nScanOut58[10] , 
        \nScanOut58[9] , \nScanOut58[8] , \nScanOut58[7] , \nScanOut58[6] , 
        \nScanOut58[5] , \nScanOut58[4] , \nScanOut58[3] , \nScanOut58[2] , 
        \nScanOut58[1] , \nScanOut58[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_58[31] , 
        \nOut0_58[30] , \nOut0_58[29] , \nOut0_58[28] , \nOut0_58[27] , 
        \nOut0_58[26] , \nOut0_58[25] , \nOut0_58[24] , \nOut0_58[23] , 
        \nOut0_58[22] , \nOut0_58[21] , \nOut0_58[20] , \nOut0_58[19] , 
        \nOut0_58[18] , \nOut0_58[17] , \nOut0_58[16] , \nOut0_58[15] , 
        \nOut0_58[14] , \nOut0_58[13] , \nOut0_58[12] , \nOut0_58[11] , 
        \nOut0_58[10] , \nOut0_58[9] , \nOut0_58[8] , \nOut0_58[7] , 
        \nOut0_58[6] , \nOut0_58[5] , \nOut0_58[4] , \nOut0_58[3] , 
        \nOut0_58[2] , \nOut0_58[1] , \nOut0_58[0] }), .NORTH_EDGE({
        \nOut0_57[31] , \nOut0_57[30] , \nOut0_57[29] , \nOut0_57[28] , 
        \nOut0_57[27] , \nOut0_57[26] , \nOut0_57[25] , \nOut0_57[24] , 
        \nOut0_57[23] , \nOut0_57[22] , \nOut0_57[21] , \nOut0_57[20] , 
        \nOut0_57[19] , \nOut0_57[18] , \nOut0_57[17] , \nOut0_57[16] , 
        \nOut0_57[15] , \nOut0_57[14] , \nOut0_57[13] , \nOut0_57[12] , 
        \nOut0_57[11] , \nOut0_57[10] , \nOut0_57[9] , \nOut0_57[8] , 
        \nOut0_57[7] , \nOut0_57[6] , \nOut0_57[5] , \nOut0_57[4] , 
        \nOut0_57[3] , \nOut0_57[2] , \nOut0_57[1] , \nOut0_57[0] }), 
        .SOUTH_EDGE({\nOut0_59[31] , \nOut0_59[30] , \nOut0_59[29] , 
        \nOut0_59[28] , \nOut0_59[27] , \nOut0_59[26] , \nOut0_59[25] , 
        \nOut0_59[24] , \nOut0_59[23] , \nOut0_59[22] , \nOut0_59[21] , 
        \nOut0_59[20] , \nOut0_59[19] , \nOut0_59[18] , \nOut0_59[17] , 
        \nOut0_59[16] , \nOut0_59[15] , \nOut0_59[14] , \nOut0_59[13] , 
        \nOut0_59[12] , \nOut0_59[11] , \nOut0_59[10] , \nOut0_59[9] , 
        \nOut0_59[8] , \nOut0_59[7] , \nOut0_59[6] , \nOut0_59[5] , 
        \nOut0_59[4] , \nOut0_59[3] , \nOut0_59[2] , \nOut0_59[1] , 
        \nOut0_59[0] }), .EAST_EDGE(\nOut1_58[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_57[31] ), .SE_EDGE(
        \nOut1_59[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_115 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut116[31] , \nScanOut116[30] , \nScanOut116[29] , 
        \nScanOut116[28] , \nScanOut116[27] , \nScanOut116[26] , 
        \nScanOut116[25] , \nScanOut116[24] , \nScanOut116[23] , 
        \nScanOut116[22] , \nScanOut116[21] , \nScanOut116[20] , 
        \nScanOut116[19] , \nScanOut116[18] , \nScanOut116[17] , 
        \nScanOut116[16] , \nScanOut116[15] , \nScanOut116[14] , 
        \nScanOut116[13] , \nScanOut116[12] , \nScanOut116[11] , 
        \nScanOut116[10] , \nScanOut116[9] , \nScanOut116[8] , 
        \nScanOut116[7] , \nScanOut116[6] , \nScanOut116[5] , \nScanOut116[4] , 
        \nScanOut116[3] , \nScanOut116[2] , \nScanOut116[1] , \nScanOut116[0] 
        }), .ScanOut({\nScanOut115[31] , \nScanOut115[30] , \nScanOut115[29] , 
        \nScanOut115[28] , \nScanOut115[27] , \nScanOut115[26] , 
        \nScanOut115[25] , \nScanOut115[24] , \nScanOut115[23] , 
        \nScanOut115[22] , \nScanOut115[21] , \nScanOut115[20] , 
        \nScanOut115[19] , \nScanOut115[18] , \nScanOut115[17] , 
        \nScanOut115[16] , \nScanOut115[15] , \nScanOut115[14] , 
        \nScanOut115[13] , \nScanOut115[12] , \nScanOut115[11] , 
        \nScanOut115[10] , \nScanOut115[9] , \nScanOut115[8] , 
        \nScanOut115[7] , \nScanOut115[6] , \nScanOut115[5] , \nScanOut115[4] , 
        \nScanOut115[3] , \nScanOut115[2] , \nScanOut115[1] , \nScanOut115[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_51[31] , \nOut1_51[30] , \nOut1_51[29] , 
        \nOut1_51[28] , \nOut1_51[27] , \nOut1_51[26] , \nOut1_51[25] , 
        \nOut1_51[24] , \nOut1_51[23] , \nOut1_51[22] , \nOut1_51[21] , 
        \nOut1_51[20] , \nOut1_51[19] , \nOut1_51[18] , \nOut1_51[17] , 
        \nOut1_51[16] , \nOut1_51[15] , \nOut1_51[14] , \nOut1_51[13] , 
        \nOut1_51[12] , \nOut1_51[11] , \nOut1_51[10] , \nOut1_51[9] , 
        \nOut1_51[8] , \nOut1_51[7] , \nOut1_51[6] , \nOut1_51[5] , 
        \nOut1_51[4] , \nOut1_51[3] , \nOut1_51[2] , \nOut1_51[1] , 
        \nOut1_51[0] }), .NORTH_EDGE({\nOut1_50[31] , \nOut1_50[30] , 
        \nOut1_50[29] , \nOut1_50[28] , \nOut1_50[27] , \nOut1_50[26] , 
        \nOut1_50[25] , \nOut1_50[24] , \nOut1_50[23] , \nOut1_50[22] , 
        \nOut1_50[21] , \nOut1_50[20] , \nOut1_50[19] , \nOut1_50[18] , 
        \nOut1_50[17] , \nOut1_50[16] , \nOut1_50[15] , \nOut1_50[14] , 
        \nOut1_50[13] , \nOut1_50[12] , \nOut1_50[11] , \nOut1_50[10] , 
        \nOut1_50[9] , \nOut1_50[8] , \nOut1_50[7] , \nOut1_50[6] , 
        \nOut1_50[5] , \nOut1_50[4] , \nOut1_50[3] , \nOut1_50[2] , 
        \nOut1_50[1] , \nOut1_50[0] }), .SOUTH_EDGE({\nOut1_52[31] , 
        \nOut1_52[30] , \nOut1_52[29] , \nOut1_52[28] , \nOut1_52[27] , 
        \nOut1_52[26] , \nOut1_52[25] , \nOut1_52[24] , \nOut1_52[23] , 
        \nOut1_52[22] , \nOut1_52[21] , \nOut1_52[20] , \nOut1_52[19] , 
        \nOut1_52[18] , \nOut1_52[17] , \nOut1_52[16] , \nOut1_52[15] , 
        \nOut1_52[14] , \nOut1_52[13] , \nOut1_52[12] , \nOut1_52[11] , 
        \nOut1_52[10] , \nOut1_52[9] , \nOut1_52[8] , \nOut1_52[7] , 
        \nOut1_52[6] , \nOut1_52[5] , \nOut1_52[4] , \nOut1_52[3] , 
        \nOut1_52[2] , \nOut1_52[1] , \nOut1_52[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_51[0] ), .NW_EDGE(\nOut0_50[0] ), .SW_EDGE(
        \nOut0_52[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_64 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut65[31] , \nScanOut65[30] , \nScanOut65[29] , 
        \nScanOut65[28] , \nScanOut65[27] , \nScanOut65[26] , \nScanOut65[25] , 
        \nScanOut65[24] , \nScanOut65[23] , \nScanOut65[22] , \nScanOut65[21] , 
        \nScanOut65[20] , \nScanOut65[19] , \nScanOut65[18] , \nScanOut65[17] , 
        \nScanOut65[16] , \nScanOut65[15] , \nScanOut65[14] , \nScanOut65[13] , 
        \nScanOut65[12] , \nScanOut65[11] , \nScanOut65[10] , \nScanOut65[9] , 
        \nScanOut65[8] , \nScanOut65[7] , \nScanOut65[6] , \nScanOut65[5] , 
        \nScanOut65[4] , \nScanOut65[3] , \nScanOut65[2] , \nScanOut65[1] , 
        \nScanOut65[0] }), .ScanOut({\nScanOut64[31] , \nScanOut64[30] , 
        \nScanOut64[29] , \nScanOut64[28] , \nScanOut64[27] , \nScanOut64[26] , 
        \nScanOut64[25] , \nScanOut64[24] , \nScanOut64[23] , \nScanOut64[22] , 
        \nScanOut64[21] , \nScanOut64[20] , \nScanOut64[19] , \nScanOut64[18] , 
        \nScanOut64[17] , \nScanOut64[16] , \nScanOut64[15] , \nScanOut64[14] , 
        \nScanOut64[13] , \nScanOut64[12] , \nScanOut64[11] , \nScanOut64[10] , 
        \nScanOut64[9] , \nScanOut64[8] , \nScanOut64[7] , \nScanOut64[6] , 
        \nScanOut64[5] , \nScanOut64[4] , \nScanOut64[3] , \nScanOut64[2] , 
        \nScanOut64[1] , \nScanOut64[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_0[31] , 
        \nOut1_0[30] , \nOut1_0[29] , \nOut1_0[28] , \nOut1_0[27] , 
        \nOut1_0[26] , \nOut1_0[25] , \nOut1_0[24] , \nOut1_0[23] , 
        \nOut1_0[22] , \nOut1_0[21] , \nOut1_0[20] , \nOut1_0[19] , 
        \nOut1_0[18] , \nOut1_0[17] , \nOut1_0[16] , \nOut1_0[15] , 
        \nOut1_0[14] , \nOut1_0[13] , \nOut1_0[12] , \nOut1_0[11] , 
        \nOut1_0[10] , \nOut1_0[9] , \nOut1_0[8] , \nOut1_0[7] , \nOut1_0[6] , 
        \nOut1_0[5] , \nOut1_0[4] , \nOut1_0[3] , \nOut1_0[2] , \nOut1_0[1] , 
        \nOut1_0[0] }), .NORTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .SOUTH_EDGE({\nOut1_1[31] , \nOut1_1[30] , \nOut1_1[29] , 
        \nOut1_1[28] , \nOut1_1[27] , \nOut1_1[26] , \nOut1_1[25] , 
        \nOut1_1[24] , \nOut1_1[23] , \nOut1_1[22] , \nOut1_1[21] , 
        \nOut1_1[20] , \nOut1_1[19] , \nOut1_1[18] , \nOut1_1[17] , 
        \nOut1_1[16] , \nOut1_1[15] , \nOut1_1[14] , \nOut1_1[13] , 
        \nOut1_1[12] , \nOut1_1[11] , \nOut1_1[10] , \nOut1_1[9] , 
        \nOut1_1[8] , \nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , \nOut1_1[4] , 
        \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_0[0] ), .NW_EDGE(1'b0), .SW_EDGE(\nOut0_1[0] 
        ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_81 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut82[31] , \nScanOut82[30] , \nScanOut82[29] , 
        \nScanOut82[28] , \nScanOut82[27] , \nScanOut82[26] , \nScanOut82[25] , 
        \nScanOut82[24] , \nScanOut82[23] , \nScanOut82[22] , \nScanOut82[21] , 
        \nScanOut82[20] , \nScanOut82[19] , \nScanOut82[18] , \nScanOut82[17] , 
        \nScanOut82[16] , \nScanOut82[15] , \nScanOut82[14] , \nScanOut82[13] , 
        \nScanOut82[12] , \nScanOut82[11] , \nScanOut82[10] , \nScanOut82[9] , 
        \nScanOut82[8] , \nScanOut82[7] , \nScanOut82[6] , \nScanOut82[5] , 
        \nScanOut82[4] , \nScanOut82[3] , \nScanOut82[2] , \nScanOut82[1] , 
        \nScanOut82[0] }), .ScanOut({\nScanOut81[31] , \nScanOut81[30] , 
        \nScanOut81[29] , \nScanOut81[28] , \nScanOut81[27] , \nScanOut81[26] , 
        \nScanOut81[25] , \nScanOut81[24] , \nScanOut81[23] , \nScanOut81[22] , 
        \nScanOut81[21] , \nScanOut81[20] , \nScanOut81[19] , \nScanOut81[18] , 
        \nScanOut81[17] , \nScanOut81[16] , \nScanOut81[15] , \nScanOut81[14] , 
        \nScanOut81[13] , \nScanOut81[12] , \nScanOut81[11] , \nScanOut81[10] , 
        \nScanOut81[9] , \nScanOut81[8] , \nScanOut81[7] , \nScanOut81[6] , 
        \nScanOut81[5] , \nScanOut81[4] , \nScanOut81[3] , \nScanOut81[2] , 
        \nScanOut81[1] , \nScanOut81[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_17[31] , 
        \nOut1_17[30] , \nOut1_17[29] , \nOut1_17[28] , \nOut1_17[27] , 
        \nOut1_17[26] , \nOut1_17[25] , \nOut1_17[24] , \nOut1_17[23] , 
        \nOut1_17[22] , \nOut1_17[21] , \nOut1_17[20] , \nOut1_17[19] , 
        \nOut1_17[18] , \nOut1_17[17] , \nOut1_17[16] , \nOut1_17[15] , 
        \nOut1_17[14] , \nOut1_17[13] , \nOut1_17[12] , \nOut1_17[11] , 
        \nOut1_17[10] , \nOut1_17[9] , \nOut1_17[8] , \nOut1_17[7] , 
        \nOut1_17[6] , \nOut1_17[5] , \nOut1_17[4] , \nOut1_17[3] , 
        \nOut1_17[2] , \nOut1_17[1] , \nOut1_17[0] }), .NORTH_EDGE({
        \nOut1_16[31] , \nOut1_16[30] , \nOut1_16[29] , \nOut1_16[28] , 
        \nOut1_16[27] , \nOut1_16[26] , \nOut1_16[25] , \nOut1_16[24] , 
        \nOut1_16[23] , \nOut1_16[22] , \nOut1_16[21] , \nOut1_16[20] , 
        \nOut1_16[19] , \nOut1_16[18] , \nOut1_16[17] , \nOut1_16[16] , 
        \nOut1_16[15] , \nOut1_16[14] , \nOut1_16[13] , \nOut1_16[12] , 
        \nOut1_16[11] , \nOut1_16[10] , \nOut1_16[9] , \nOut1_16[8] , 
        \nOut1_16[7] , \nOut1_16[6] , \nOut1_16[5] , \nOut1_16[4] , 
        \nOut1_16[3] , \nOut1_16[2] , \nOut1_16[1] , \nOut1_16[0] }), 
        .SOUTH_EDGE({\nOut1_18[31] , \nOut1_18[30] , \nOut1_18[29] , 
        \nOut1_18[28] , \nOut1_18[27] , \nOut1_18[26] , \nOut1_18[25] , 
        \nOut1_18[24] , \nOut1_18[23] , \nOut1_18[22] , \nOut1_18[21] , 
        \nOut1_18[20] , \nOut1_18[19] , \nOut1_18[18] , \nOut1_18[17] , 
        \nOut1_18[16] , \nOut1_18[15] , \nOut1_18[14] , \nOut1_18[13] , 
        \nOut1_18[12] , \nOut1_18[11] , \nOut1_18[10] , \nOut1_18[9] , 
        \nOut1_18[8] , \nOut1_18[7] , \nOut1_18[6] , \nOut1_18[5] , 
        \nOut1_18[4] , \nOut1_18[3] , \nOut1_18[2] , \nOut1_18[1] , 
        \nOut1_18[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_17[0] ), 
        .NW_EDGE(\nOut0_16[0] ), .SW_EDGE(\nOut0_18[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_93 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut94[31] , \nScanOut94[30] , \nScanOut94[29] , 
        \nScanOut94[28] , \nScanOut94[27] , \nScanOut94[26] , \nScanOut94[25] , 
        \nScanOut94[24] , \nScanOut94[23] , \nScanOut94[22] , \nScanOut94[21] , 
        \nScanOut94[20] , \nScanOut94[19] , \nScanOut94[18] , \nScanOut94[17] , 
        \nScanOut94[16] , \nScanOut94[15] , \nScanOut94[14] , \nScanOut94[13] , 
        \nScanOut94[12] , \nScanOut94[11] , \nScanOut94[10] , \nScanOut94[9] , 
        \nScanOut94[8] , \nScanOut94[7] , \nScanOut94[6] , \nScanOut94[5] , 
        \nScanOut94[4] , \nScanOut94[3] , \nScanOut94[2] , \nScanOut94[1] , 
        \nScanOut94[0] }), .ScanOut({\nScanOut93[31] , \nScanOut93[30] , 
        \nScanOut93[29] , \nScanOut93[28] , \nScanOut93[27] , \nScanOut93[26] , 
        \nScanOut93[25] , \nScanOut93[24] , \nScanOut93[23] , \nScanOut93[22] , 
        \nScanOut93[21] , \nScanOut93[20] , \nScanOut93[19] , \nScanOut93[18] , 
        \nScanOut93[17] , \nScanOut93[16] , \nScanOut93[15] , \nScanOut93[14] , 
        \nScanOut93[13] , \nScanOut93[12] , \nScanOut93[11] , \nScanOut93[10] , 
        \nScanOut93[9] , \nScanOut93[8] , \nScanOut93[7] , \nScanOut93[6] , 
        \nScanOut93[5] , \nScanOut93[4] , \nScanOut93[3] , \nScanOut93[2] , 
        \nScanOut93[1] , \nScanOut93[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_29[31] , 
        \nOut1_29[30] , \nOut1_29[29] , \nOut1_29[28] , \nOut1_29[27] , 
        \nOut1_29[26] , \nOut1_29[25] , \nOut1_29[24] , \nOut1_29[23] , 
        \nOut1_29[22] , \nOut1_29[21] , \nOut1_29[20] , \nOut1_29[19] , 
        \nOut1_29[18] , \nOut1_29[17] , \nOut1_29[16] , \nOut1_29[15] , 
        \nOut1_29[14] , \nOut1_29[13] , \nOut1_29[12] , \nOut1_29[11] , 
        \nOut1_29[10] , \nOut1_29[9] , \nOut1_29[8] , \nOut1_29[7] , 
        \nOut1_29[6] , \nOut1_29[5] , \nOut1_29[4] , \nOut1_29[3] , 
        \nOut1_29[2] , \nOut1_29[1] , \nOut1_29[0] }), .NORTH_EDGE({
        \nOut1_28[31] , \nOut1_28[30] , \nOut1_28[29] , \nOut1_28[28] , 
        \nOut1_28[27] , \nOut1_28[26] , \nOut1_28[25] , \nOut1_28[24] , 
        \nOut1_28[23] , \nOut1_28[22] , \nOut1_28[21] , \nOut1_28[20] , 
        \nOut1_28[19] , \nOut1_28[18] , \nOut1_28[17] , \nOut1_28[16] , 
        \nOut1_28[15] , \nOut1_28[14] , \nOut1_28[13] , \nOut1_28[12] , 
        \nOut1_28[11] , \nOut1_28[10] , \nOut1_28[9] , \nOut1_28[8] , 
        \nOut1_28[7] , \nOut1_28[6] , \nOut1_28[5] , \nOut1_28[4] , 
        \nOut1_28[3] , \nOut1_28[2] , \nOut1_28[1] , \nOut1_28[0] }), 
        .SOUTH_EDGE({\nOut1_30[31] , \nOut1_30[30] , \nOut1_30[29] , 
        \nOut1_30[28] , \nOut1_30[27] , \nOut1_30[26] , \nOut1_30[25] , 
        \nOut1_30[24] , \nOut1_30[23] , \nOut1_30[22] , \nOut1_30[21] , 
        \nOut1_30[20] , \nOut1_30[19] , \nOut1_30[18] , \nOut1_30[17] , 
        \nOut1_30[16] , \nOut1_30[15] , \nOut1_30[14] , \nOut1_30[13] , 
        \nOut1_30[12] , \nOut1_30[11] , \nOut1_30[10] , \nOut1_30[9] , 
        \nOut1_30[8] , \nOut1_30[7] , \nOut1_30[6] , \nOut1_30[5] , 
        \nOut1_30[4] , \nOut1_30[3] , \nOut1_30[2] , \nOut1_30[1] , 
        \nOut1_30[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_29[0] ), 
        .NW_EDGE(\nOut0_28[0] ), .SW_EDGE(\nOut0_30[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_23 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut24[31] , \nScanOut24[30] , \nScanOut24[29] , 
        \nScanOut24[28] , \nScanOut24[27] , \nScanOut24[26] , \nScanOut24[25] , 
        \nScanOut24[24] , \nScanOut24[23] , \nScanOut24[22] , \nScanOut24[21] , 
        \nScanOut24[20] , \nScanOut24[19] , \nScanOut24[18] , \nScanOut24[17] , 
        \nScanOut24[16] , \nScanOut24[15] , \nScanOut24[14] , \nScanOut24[13] , 
        \nScanOut24[12] , \nScanOut24[11] , \nScanOut24[10] , \nScanOut24[9] , 
        \nScanOut24[8] , \nScanOut24[7] , \nScanOut24[6] , \nScanOut24[5] , 
        \nScanOut24[4] , \nScanOut24[3] , \nScanOut24[2] , \nScanOut24[1] , 
        \nScanOut24[0] }), .ScanOut({\nScanOut23[31] , \nScanOut23[30] , 
        \nScanOut23[29] , \nScanOut23[28] , \nScanOut23[27] , \nScanOut23[26] , 
        \nScanOut23[25] , \nScanOut23[24] , \nScanOut23[23] , \nScanOut23[22] , 
        \nScanOut23[21] , \nScanOut23[20] , \nScanOut23[19] , \nScanOut23[18] , 
        \nScanOut23[17] , \nScanOut23[16] , \nScanOut23[15] , \nScanOut23[14] , 
        \nScanOut23[13] , \nScanOut23[12] , \nScanOut23[11] , \nScanOut23[10] , 
        \nScanOut23[9] , \nScanOut23[8] , \nScanOut23[7] , \nScanOut23[6] , 
        \nScanOut23[5] , \nScanOut23[4] , \nScanOut23[3] , \nScanOut23[2] , 
        \nScanOut23[1] , \nScanOut23[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_23[31] , 
        \nOut0_23[30] , \nOut0_23[29] , \nOut0_23[28] , \nOut0_23[27] , 
        \nOut0_23[26] , \nOut0_23[25] , \nOut0_23[24] , \nOut0_23[23] , 
        \nOut0_23[22] , \nOut0_23[21] , \nOut0_23[20] , \nOut0_23[19] , 
        \nOut0_23[18] , \nOut0_23[17] , \nOut0_23[16] , \nOut0_23[15] , 
        \nOut0_23[14] , \nOut0_23[13] , \nOut0_23[12] , \nOut0_23[11] , 
        \nOut0_23[10] , \nOut0_23[9] , \nOut0_23[8] , \nOut0_23[7] , 
        \nOut0_23[6] , \nOut0_23[5] , \nOut0_23[4] , \nOut0_23[3] , 
        \nOut0_23[2] , \nOut0_23[1] , \nOut0_23[0] }), .NORTH_EDGE({
        \nOut0_22[31] , \nOut0_22[30] , \nOut0_22[29] , \nOut0_22[28] , 
        \nOut0_22[27] , \nOut0_22[26] , \nOut0_22[25] , \nOut0_22[24] , 
        \nOut0_22[23] , \nOut0_22[22] , \nOut0_22[21] , \nOut0_22[20] , 
        \nOut0_22[19] , \nOut0_22[18] , \nOut0_22[17] , \nOut0_22[16] , 
        \nOut0_22[15] , \nOut0_22[14] , \nOut0_22[13] , \nOut0_22[12] , 
        \nOut0_22[11] , \nOut0_22[10] , \nOut0_22[9] , \nOut0_22[8] , 
        \nOut0_22[7] , \nOut0_22[6] , \nOut0_22[5] , \nOut0_22[4] , 
        \nOut0_22[3] , \nOut0_22[2] , \nOut0_22[1] , \nOut0_22[0] }), 
        .SOUTH_EDGE({\nOut0_24[31] , \nOut0_24[30] , \nOut0_24[29] , 
        \nOut0_24[28] , \nOut0_24[27] , \nOut0_24[26] , \nOut0_24[25] , 
        \nOut0_24[24] , \nOut0_24[23] , \nOut0_24[22] , \nOut0_24[21] , 
        \nOut0_24[20] , \nOut0_24[19] , \nOut0_24[18] , \nOut0_24[17] , 
        \nOut0_24[16] , \nOut0_24[15] , \nOut0_24[14] , \nOut0_24[13] , 
        \nOut0_24[12] , \nOut0_24[11] , \nOut0_24[10] , \nOut0_24[9] , 
        \nOut0_24[8] , \nOut0_24[7] , \nOut0_24[6] , \nOut0_24[5] , 
        \nOut0_24[4] , \nOut0_24[3] , \nOut0_24[2] , \nOut0_24[1] , 
        \nOut0_24[0] }), .EAST_EDGE(\nOut1_23[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_22[31] ), .SE_EDGE(
        \nOut1_24[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_24 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut25[31] , \nScanOut25[30] , \nScanOut25[29] , 
        \nScanOut25[28] , \nScanOut25[27] , \nScanOut25[26] , \nScanOut25[25] , 
        \nScanOut25[24] , \nScanOut25[23] , \nScanOut25[22] , \nScanOut25[21] , 
        \nScanOut25[20] , \nScanOut25[19] , \nScanOut25[18] , \nScanOut25[17] , 
        \nScanOut25[16] , \nScanOut25[15] , \nScanOut25[14] , \nScanOut25[13] , 
        \nScanOut25[12] , \nScanOut25[11] , \nScanOut25[10] , \nScanOut25[9] , 
        \nScanOut25[8] , \nScanOut25[7] , \nScanOut25[6] , \nScanOut25[5] , 
        \nScanOut25[4] , \nScanOut25[3] , \nScanOut25[2] , \nScanOut25[1] , 
        \nScanOut25[0] }), .ScanOut({\nScanOut24[31] , \nScanOut24[30] , 
        \nScanOut24[29] , \nScanOut24[28] , \nScanOut24[27] , \nScanOut24[26] , 
        \nScanOut24[25] , \nScanOut24[24] , \nScanOut24[23] , \nScanOut24[22] , 
        \nScanOut24[21] , \nScanOut24[20] , \nScanOut24[19] , \nScanOut24[18] , 
        \nScanOut24[17] , \nScanOut24[16] , \nScanOut24[15] , \nScanOut24[14] , 
        \nScanOut24[13] , \nScanOut24[12] , \nScanOut24[11] , \nScanOut24[10] , 
        \nScanOut24[9] , \nScanOut24[8] , \nScanOut24[7] , \nScanOut24[6] , 
        \nScanOut24[5] , \nScanOut24[4] , \nScanOut24[3] , \nScanOut24[2] , 
        \nScanOut24[1] , \nScanOut24[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_24[31] , 
        \nOut0_24[30] , \nOut0_24[29] , \nOut0_24[28] , \nOut0_24[27] , 
        \nOut0_24[26] , \nOut0_24[25] , \nOut0_24[24] , \nOut0_24[23] , 
        \nOut0_24[22] , \nOut0_24[21] , \nOut0_24[20] , \nOut0_24[19] , 
        \nOut0_24[18] , \nOut0_24[17] , \nOut0_24[16] , \nOut0_24[15] , 
        \nOut0_24[14] , \nOut0_24[13] , \nOut0_24[12] , \nOut0_24[11] , 
        \nOut0_24[10] , \nOut0_24[9] , \nOut0_24[8] , \nOut0_24[7] , 
        \nOut0_24[6] , \nOut0_24[5] , \nOut0_24[4] , \nOut0_24[3] , 
        \nOut0_24[2] , \nOut0_24[1] , \nOut0_24[0] }), .NORTH_EDGE({
        \nOut0_23[31] , \nOut0_23[30] , \nOut0_23[29] , \nOut0_23[28] , 
        \nOut0_23[27] , \nOut0_23[26] , \nOut0_23[25] , \nOut0_23[24] , 
        \nOut0_23[23] , \nOut0_23[22] , \nOut0_23[21] , \nOut0_23[20] , 
        \nOut0_23[19] , \nOut0_23[18] , \nOut0_23[17] , \nOut0_23[16] , 
        \nOut0_23[15] , \nOut0_23[14] , \nOut0_23[13] , \nOut0_23[12] , 
        \nOut0_23[11] , \nOut0_23[10] , \nOut0_23[9] , \nOut0_23[8] , 
        \nOut0_23[7] , \nOut0_23[6] , \nOut0_23[5] , \nOut0_23[4] , 
        \nOut0_23[3] , \nOut0_23[2] , \nOut0_23[1] , \nOut0_23[0] }), 
        .SOUTH_EDGE({\nOut0_25[31] , \nOut0_25[30] , \nOut0_25[29] , 
        \nOut0_25[28] , \nOut0_25[27] , \nOut0_25[26] , \nOut0_25[25] , 
        \nOut0_25[24] , \nOut0_25[23] , \nOut0_25[22] , \nOut0_25[21] , 
        \nOut0_25[20] , \nOut0_25[19] , \nOut0_25[18] , \nOut0_25[17] , 
        \nOut0_25[16] , \nOut0_25[15] , \nOut0_25[14] , \nOut0_25[13] , 
        \nOut0_25[12] , \nOut0_25[11] , \nOut0_25[10] , \nOut0_25[9] , 
        \nOut0_25[8] , \nOut0_25[7] , \nOut0_25[6] , \nOut0_25[5] , 
        \nOut0_25[4] , \nOut0_25[3] , \nOut0_25[2] , \nOut0_25[1] , 
        \nOut0_25[0] }), .EAST_EDGE(\nOut1_24[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_23[31] ), .SE_EDGE(
        \nOut1_25[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_51 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut52[31] , \nScanOut52[30] , \nScanOut52[29] , 
        \nScanOut52[28] , \nScanOut52[27] , \nScanOut52[26] , \nScanOut52[25] , 
        \nScanOut52[24] , \nScanOut52[23] , \nScanOut52[22] , \nScanOut52[21] , 
        \nScanOut52[20] , \nScanOut52[19] , \nScanOut52[18] , \nScanOut52[17] , 
        \nScanOut52[16] , \nScanOut52[15] , \nScanOut52[14] , \nScanOut52[13] , 
        \nScanOut52[12] , \nScanOut52[11] , \nScanOut52[10] , \nScanOut52[9] , 
        \nScanOut52[8] , \nScanOut52[7] , \nScanOut52[6] , \nScanOut52[5] , 
        \nScanOut52[4] , \nScanOut52[3] , \nScanOut52[2] , \nScanOut52[1] , 
        \nScanOut52[0] }), .ScanOut({\nScanOut51[31] , \nScanOut51[30] , 
        \nScanOut51[29] , \nScanOut51[28] , \nScanOut51[27] , \nScanOut51[26] , 
        \nScanOut51[25] , \nScanOut51[24] , \nScanOut51[23] , \nScanOut51[22] , 
        \nScanOut51[21] , \nScanOut51[20] , \nScanOut51[19] , \nScanOut51[18] , 
        \nScanOut51[17] , \nScanOut51[16] , \nScanOut51[15] , \nScanOut51[14] , 
        \nScanOut51[13] , \nScanOut51[12] , \nScanOut51[11] , \nScanOut51[10] , 
        \nScanOut51[9] , \nScanOut51[8] , \nScanOut51[7] , \nScanOut51[6] , 
        \nScanOut51[5] , \nScanOut51[4] , \nScanOut51[3] , \nScanOut51[2] , 
        \nScanOut51[1] , \nScanOut51[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_51[31] , 
        \nOut0_51[30] , \nOut0_51[29] , \nOut0_51[28] , \nOut0_51[27] , 
        \nOut0_51[26] , \nOut0_51[25] , \nOut0_51[24] , \nOut0_51[23] , 
        \nOut0_51[22] , \nOut0_51[21] , \nOut0_51[20] , \nOut0_51[19] , 
        \nOut0_51[18] , \nOut0_51[17] , \nOut0_51[16] , \nOut0_51[15] , 
        \nOut0_51[14] , \nOut0_51[13] , \nOut0_51[12] , \nOut0_51[11] , 
        \nOut0_51[10] , \nOut0_51[9] , \nOut0_51[8] , \nOut0_51[7] , 
        \nOut0_51[6] , \nOut0_51[5] , \nOut0_51[4] , \nOut0_51[3] , 
        \nOut0_51[2] , \nOut0_51[1] , \nOut0_51[0] }), .NORTH_EDGE({
        \nOut0_50[31] , \nOut0_50[30] , \nOut0_50[29] , \nOut0_50[28] , 
        \nOut0_50[27] , \nOut0_50[26] , \nOut0_50[25] , \nOut0_50[24] , 
        \nOut0_50[23] , \nOut0_50[22] , \nOut0_50[21] , \nOut0_50[20] , 
        \nOut0_50[19] , \nOut0_50[18] , \nOut0_50[17] , \nOut0_50[16] , 
        \nOut0_50[15] , \nOut0_50[14] , \nOut0_50[13] , \nOut0_50[12] , 
        \nOut0_50[11] , \nOut0_50[10] , \nOut0_50[9] , \nOut0_50[8] , 
        \nOut0_50[7] , \nOut0_50[6] , \nOut0_50[5] , \nOut0_50[4] , 
        \nOut0_50[3] , \nOut0_50[2] , \nOut0_50[1] , \nOut0_50[0] }), 
        .SOUTH_EDGE({\nOut0_52[31] , \nOut0_52[30] , \nOut0_52[29] , 
        \nOut0_52[28] , \nOut0_52[27] , \nOut0_52[26] , \nOut0_52[25] , 
        \nOut0_52[24] , \nOut0_52[23] , \nOut0_52[22] , \nOut0_52[21] , 
        \nOut0_52[20] , \nOut0_52[19] , \nOut0_52[18] , \nOut0_52[17] , 
        \nOut0_52[16] , \nOut0_52[15] , \nOut0_52[14] , \nOut0_52[13] , 
        \nOut0_52[12] , \nOut0_52[11] , \nOut0_52[10] , \nOut0_52[9] , 
        \nOut0_52[8] , \nOut0_52[7] , \nOut0_52[6] , \nOut0_52[5] , 
        \nOut0_52[4] , \nOut0_52[3] , \nOut0_52[2] , \nOut0_52[1] , 
        \nOut0_52[0] }), .EAST_EDGE(\nOut1_51[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_50[31] ), .SE_EDGE(
        \nOut1_52[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_107 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut108[31] , \nScanOut108[30] , \nScanOut108[29] , 
        \nScanOut108[28] , \nScanOut108[27] , \nScanOut108[26] , 
        \nScanOut108[25] , \nScanOut108[24] , \nScanOut108[23] , 
        \nScanOut108[22] , \nScanOut108[21] , \nScanOut108[20] , 
        \nScanOut108[19] , \nScanOut108[18] , \nScanOut108[17] , 
        \nScanOut108[16] , \nScanOut108[15] , \nScanOut108[14] , 
        \nScanOut108[13] , \nScanOut108[12] , \nScanOut108[11] , 
        \nScanOut108[10] , \nScanOut108[9] , \nScanOut108[8] , 
        \nScanOut108[7] , \nScanOut108[6] , \nScanOut108[5] , \nScanOut108[4] , 
        \nScanOut108[3] , \nScanOut108[2] , \nScanOut108[1] , \nScanOut108[0] 
        }), .ScanOut({\nScanOut107[31] , \nScanOut107[30] , \nScanOut107[29] , 
        \nScanOut107[28] , \nScanOut107[27] , \nScanOut107[26] , 
        \nScanOut107[25] , \nScanOut107[24] , \nScanOut107[23] , 
        \nScanOut107[22] , \nScanOut107[21] , \nScanOut107[20] , 
        \nScanOut107[19] , \nScanOut107[18] , \nScanOut107[17] , 
        \nScanOut107[16] , \nScanOut107[15] , \nScanOut107[14] , 
        \nScanOut107[13] , \nScanOut107[12] , \nScanOut107[11] , 
        \nScanOut107[10] , \nScanOut107[9] , \nScanOut107[8] , 
        \nScanOut107[7] , \nScanOut107[6] , \nScanOut107[5] , \nScanOut107[4] , 
        \nScanOut107[3] , \nScanOut107[2] , \nScanOut107[1] , \nScanOut107[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_43[31] , \nOut1_43[30] , \nOut1_43[29] , 
        \nOut1_43[28] , \nOut1_43[27] , \nOut1_43[26] , \nOut1_43[25] , 
        \nOut1_43[24] , \nOut1_43[23] , \nOut1_43[22] , \nOut1_43[21] , 
        \nOut1_43[20] , \nOut1_43[19] , \nOut1_43[18] , \nOut1_43[17] , 
        \nOut1_43[16] , \nOut1_43[15] , \nOut1_43[14] , \nOut1_43[13] , 
        \nOut1_43[12] , \nOut1_43[11] , \nOut1_43[10] , \nOut1_43[9] , 
        \nOut1_43[8] , \nOut1_43[7] , \nOut1_43[6] , \nOut1_43[5] , 
        \nOut1_43[4] , \nOut1_43[3] , \nOut1_43[2] , \nOut1_43[1] , 
        \nOut1_43[0] }), .NORTH_EDGE({\nOut1_42[31] , \nOut1_42[30] , 
        \nOut1_42[29] , \nOut1_42[28] , \nOut1_42[27] , \nOut1_42[26] , 
        \nOut1_42[25] , \nOut1_42[24] , \nOut1_42[23] , \nOut1_42[22] , 
        \nOut1_42[21] , \nOut1_42[20] , \nOut1_42[19] , \nOut1_42[18] , 
        \nOut1_42[17] , \nOut1_42[16] , \nOut1_42[15] , \nOut1_42[14] , 
        \nOut1_42[13] , \nOut1_42[12] , \nOut1_42[11] , \nOut1_42[10] , 
        \nOut1_42[9] , \nOut1_42[8] , \nOut1_42[7] , \nOut1_42[6] , 
        \nOut1_42[5] , \nOut1_42[4] , \nOut1_42[3] , \nOut1_42[2] , 
        \nOut1_42[1] , \nOut1_42[0] }), .SOUTH_EDGE({\nOut1_44[31] , 
        \nOut1_44[30] , \nOut1_44[29] , \nOut1_44[28] , \nOut1_44[27] , 
        \nOut1_44[26] , \nOut1_44[25] , \nOut1_44[24] , \nOut1_44[23] , 
        \nOut1_44[22] , \nOut1_44[21] , \nOut1_44[20] , \nOut1_44[19] , 
        \nOut1_44[18] , \nOut1_44[17] , \nOut1_44[16] , \nOut1_44[15] , 
        \nOut1_44[14] , \nOut1_44[13] , \nOut1_44[12] , \nOut1_44[11] , 
        \nOut1_44[10] , \nOut1_44[9] , \nOut1_44[8] , \nOut1_44[7] , 
        \nOut1_44[6] , \nOut1_44[5] , \nOut1_44[4] , \nOut1_44[3] , 
        \nOut1_44[2] , \nOut1_44[1] , \nOut1_44[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_43[0] ), .NW_EDGE(\nOut0_42[0] ), .SW_EDGE(
        \nOut0_44[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_76 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut77[31] , \nScanOut77[30] , \nScanOut77[29] , 
        \nScanOut77[28] , \nScanOut77[27] , \nScanOut77[26] , \nScanOut77[25] , 
        \nScanOut77[24] , \nScanOut77[23] , \nScanOut77[22] , \nScanOut77[21] , 
        \nScanOut77[20] , \nScanOut77[19] , \nScanOut77[18] , \nScanOut77[17] , 
        \nScanOut77[16] , \nScanOut77[15] , \nScanOut77[14] , \nScanOut77[13] , 
        \nScanOut77[12] , \nScanOut77[11] , \nScanOut77[10] , \nScanOut77[9] , 
        \nScanOut77[8] , \nScanOut77[7] , \nScanOut77[6] , \nScanOut77[5] , 
        \nScanOut77[4] , \nScanOut77[3] , \nScanOut77[2] , \nScanOut77[1] , 
        \nScanOut77[0] }), .ScanOut({\nScanOut76[31] , \nScanOut76[30] , 
        \nScanOut76[29] , \nScanOut76[28] , \nScanOut76[27] , \nScanOut76[26] , 
        \nScanOut76[25] , \nScanOut76[24] , \nScanOut76[23] , \nScanOut76[22] , 
        \nScanOut76[21] , \nScanOut76[20] , \nScanOut76[19] , \nScanOut76[18] , 
        \nScanOut76[17] , \nScanOut76[16] , \nScanOut76[15] , \nScanOut76[14] , 
        \nScanOut76[13] , \nScanOut76[12] , \nScanOut76[11] , \nScanOut76[10] , 
        \nScanOut76[9] , \nScanOut76[8] , \nScanOut76[7] , \nScanOut76[6] , 
        \nScanOut76[5] , \nScanOut76[4] , \nScanOut76[3] , \nScanOut76[2] , 
        \nScanOut76[1] , \nScanOut76[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_12[31] , 
        \nOut1_12[30] , \nOut1_12[29] , \nOut1_12[28] , \nOut1_12[27] , 
        \nOut1_12[26] , \nOut1_12[25] , \nOut1_12[24] , \nOut1_12[23] , 
        \nOut1_12[22] , \nOut1_12[21] , \nOut1_12[20] , \nOut1_12[19] , 
        \nOut1_12[18] , \nOut1_12[17] , \nOut1_12[16] , \nOut1_12[15] , 
        \nOut1_12[14] , \nOut1_12[13] , \nOut1_12[12] , \nOut1_12[11] , 
        \nOut1_12[10] , \nOut1_12[9] , \nOut1_12[8] , \nOut1_12[7] , 
        \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , \nOut1_12[3] , 
        \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), .NORTH_EDGE({
        \nOut1_11[31] , \nOut1_11[30] , \nOut1_11[29] , \nOut1_11[28] , 
        \nOut1_11[27] , \nOut1_11[26] , \nOut1_11[25] , \nOut1_11[24] , 
        \nOut1_11[23] , \nOut1_11[22] , \nOut1_11[21] , \nOut1_11[20] , 
        \nOut1_11[19] , \nOut1_11[18] , \nOut1_11[17] , \nOut1_11[16] , 
        \nOut1_11[15] , \nOut1_11[14] , \nOut1_11[13] , \nOut1_11[12] , 
        \nOut1_11[11] , \nOut1_11[10] , \nOut1_11[9] , \nOut1_11[8] , 
        \nOut1_11[7] , \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , 
        \nOut1_11[3] , \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), 
        .SOUTH_EDGE({\nOut1_13[31] , \nOut1_13[30] , \nOut1_13[29] , 
        \nOut1_13[28] , \nOut1_13[27] , \nOut1_13[26] , \nOut1_13[25] , 
        \nOut1_13[24] , \nOut1_13[23] , \nOut1_13[22] , \nOut1_13[21] , 
        \nOut1_13[20] , \nOut1_13[19] , \nOut1_13[18] , \nOut1_13[17] , 
        \nOut1_13[16] , \nOut1_13[15] , \nOut1_13[14] , \nOut1_13[13] , 
        \nOut1_13[12] , \nOut1_13[11] , \nOut1_13[10] , \nOut1_13[9] , 
        \nOut1_13[8] , \nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , 
        \nOut1_13[4] , \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , 
        \nOut1_13[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_12[0] ), 
        .NW_EDGE(\nOut0_11[0] ), .SW_EDGE(\nOut0_13[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_88 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut89[31] , \nScanOut89[30] , \nScanOut89[29] , 
        \nScanOut89[28] , \nScanOut89[27] , \nScanOut89[26] , \nScanOut89[25] , 
        \nScanOut89[24] , \nScanOut89[23] , \nScanOut89[22] , \nScanOut89[21] , 
        \nScanOut89[20] , \nScanOut89[19] , \nScanOut89[18] , \nScanOut89[17] , 
        \nScanOut89[16] , \nScanOut89[15] , \nScanOut89[14] , \nScanOut89[13] , 
        \nScanOut89[12] , \nScanOut89[11] , \nScanOut89[10] , \nScanOut89[9] , 
        \nScanOut89[8] , \nScanOut89[7] , \nScanOut89[6] , \nScanOut89[5] , 
        \nScanOut89[4] , \nScanOut89[3] , \nScanOut89[2] , \nScanOut89[1] , 
        \nScanOut89[0] }), .ScanOut({\nScanOut88[31] , \nScanOut88[30] , 
        \nScanOut88[29] , \nScanOut88[28] , \nScanOut88[27] , \nScanOut88[26] , 
        \nScanOut88[25] , \nScanOut88[24] , \nScanOut88[23] , \nScanOut88[22] , 
        \nScanOut88[21] , \nScanOut88[20] , \nScanOut88[19] , \nScanOut88[18] , 
        \nScanOut88[17] , \nScanOut88[16] , \nScanOut88[15] , \nScanOut88[14] , 
        \nScanOut88[13] , \nScanOut88[12] , \nScanOut88[11] , \nScanOut88[10] , 
        \nScanOut88[9] , \nScanOut88[8] , \nScanOut88[7] , \nScanOut88[6] , 
        \nScanOut88[5] , \nScanOut88[4] , \nScanOut88[3] , \nScanOut88[2] , 
        \nScanOut88[1] , \nScanOut88[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_24[31] , 
        \nOut1_24[30] , \nOut1_24[29] , \nOut1_24[28] , \nOut1_24[27] , 
        \nOut1_24[26] , \nOut1_24[25] , \nOut1_24[24] , \nOut1_24[23] , 
        \nOut1_24[22] , \nOut1_24[21] , \nOut1_24[20] , \nOut1_24[19] , 
        \nOut1_24[18] , \nOut1_24[17] , \nOut1_24[16] , \nOut1_24[15] , 
        \nOut1_24[14] , \nOut1_24[13] , \nOut1_24[12] , \nOut1_24[11] , 
        \nOut1_24[10] , \nOut1_24[9] , \nOut1_24[8] , \nOut1_24[7] , 
        \nOut1_24[6] , \nOut1_24[5] , \nOut1_24[4] , \nOut1_24[3] , 
        \nOut1_24[2] , \nOut1_24[1] , \nOut1_24[0] }), .NORTH_EDGE({
        \nOut1_23[31] , \nOut1_23[30] , \nOut1_23[29] , \nOut1_23[28] , 
        \nOut1_23[27] , \nOut1_23[26] , \nOut1_23[25] , \nOut1_23[24] , 
        \nOut1_23[23] , \nOut1_23[22] , \nOut1_23[21] , \nOut1_23[20] , 
        \nOut1_23[19] , \nOut1_23[18] , \nOut1_23[17] , \nOut1_23[16] , 
        \nOut1_23[15] , \nOut1_23[14] , \nOut1_23[13] , \nOut1_23[12] , 
        \nOut1_23[11] , \nOut1_23[10] , \nOut1_23[9] , \nOut1_23[8] , 
        \nOut1_23[7] , \nOut1_23[6] , \nOut1_23[5] , \nOut1_23[4] , 
        \nOut1_23[3] , \nOut1_23[2] , \nOut1_23[1] , \nOut1_23[0] }), 
        .SOUTH_EDGE({\nOut1_25[31] , \nOut1_25[30] , \nOut1_25[29] , 
        \nOut1_25[28] , \nOut1_25[27] , \nOut1_25[26] , \nOut1_25[25] , 
        \nOut1_25[24] , \nOut1_25[23] , \nOut1_25[22] , \nOut1_25[21] , 
        \nOut1_25[20] , \nOut1_25[19] , \nOut1_25[18] , \nOut1_25[17] , 
        \nOut1_25[16] , \nOut1_25[15] , \nOut1_25[14] , \nOut1_25[13] , 
        \nOut1_25[12] , \nOut1_25[11] , \nOut1_25[10] , \nOut1_25[9] , 
        \nOut1_25[8] , \nOut1_25[7] , \nOut1_25[6] , \nOut1_25[5] , 
        \nOut1_25[4] , \nOut1_25[3] , \nOut1_25[2] , \nOut1_25[1] , 
        \nOut1_25[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_24[0] ), 
        .NW_EDGE(\nOut0_23[0] ), .SW_EDGE(\nOut0_25[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_120 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut121[31] , \nScanOut121[30] , \nScanOut121[29] , 
        \nScanOut121[28] , \nScanOut121[27] , \nScanOut121[26] , 
        \nScanOut121[25] , \nScanOut121[24] , \nScanOut121[23] , 
        \nScanOut121[22] , \nScanOut121[21] , \nScanOut121[20] , 
        \nScanOut121[19] , \nScanOut121[18] , \nScanOut121[17] , 
        \nScanOut121[16] , \nScanOut121[15] , \nScanOut121[14] , 
        \nScanOut121[13] , \nScanOut121[12] , \nScanOut121[11] , 
        \nScanOut121[10] , \nScanOut121[9] , \nScanOut121[8] , 
        \nScanOut121[7] , \nScanOut121[6] , \nScanOut121[5] , \nScanOut121[4] , 
        \nScanOut121[3] , \nScanOut121[2] , \nScanOut121[1] , \nScanOut121[0] 
        }), .ScanOut({\nScanOut120[31] , \nScanOut120[30] , \nScanOut120[29] , 
        \nScanOut120[28] , \nScanOut120[27] , \nScanOut120[26] , 
        \nScanOut120[25] , \nScanOut120[24] , \nScanOut120[23] , 
        \nScanOut120[22] , \nScanOut120[21] , \nScanOut120[20] , 
        \nScanOut120[19] , \nScanOut120[18] , \nScanOut120[17] , 
        \nScanOut120[16] , \nScanOut120[15] , \nScanOut120[14] , 
        \nScanOut120[13] , \nScanOut120[12] , \nScanOut120[11] , 
        \nScanOut120[10] , \nScanOut120[9] , \nScanOut120[8] , 
        \nScanOut120[7] , \nScanOut120[6] , \nScanOut120[5] , \nScanOut120[4] , 
        \nScanOut120[3] , \nScanOut120[2] , \nScanOut120[1] , \nScanOut120[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_56[31] , \nOut1_56[30] , \nOut1_56[29] , 
        \nOut1_56[28] , \nOut1_56[27] , \nOut1_56[26] , \nOut1_56[25] , 
        \nOut1_56[24] , \nOut1_56[23] , \nOut1_56[22] , \nOut1_56[21] , 
        \nOut1_56[20] , \nOut1_56[19] , \nOut1_56[18] , \nOut1_56[17] , 
        \nOut1_56[16] , \nOut1_56[15] , \nOut1_56[14] , \nOut1_56[13] , 
        \nOut1_56[12] , \nOut1_56[11] , \nOut1_56[10] , \nOut1_56[9] , 
        \nOut1_56[8] , \nOut1_56[7] , \nOut1_56[6] , \nOut1_56[5] , 
        \nOut1_56[4] , \nOut1_56[3] , \nOut1_56[2] , \nOut1_56[1] , 
        \nOut1_56[0] }), .NORTH_EDGE({\nOut1_55[31] , \nOut1_55[30] , 
        \nOut1_55[29] , \nOut1_55[28] , \nOut1_55[27] , \nOut1_55[26] , 
        \nOut1_55[25] , \nOut1_55[24] , \nOut1_55[23] , \nOut1_55[22] , 
        \nOut1_55[21] , \nOut1_55[20] , \nOut1_55[19] , \nOut1_55[18] , 
        \nOut1_55[17] , \nOut1_55[16] , \nOut1_55[15] , \nOut1_55[14] , 
        \nOut1_55[13] , \nOut1_55[12] , \nOut1_55[11] , \nOut1_55[10] , 
        \nOut1_55[9] , \nOut1_55[8] , \nOut1_55[7] , \nOut1_55[6] , 
        \nOut1_55[5] , \nOut1_55[4] , \nOut1_55[3] , \nOut1_55[2] , 
        \nOut1_55[1] , \nOut1_55[0] }), .SOUTH_EDGE({\nOut1_57[31] , 
        \nOut1_57[30] , \nOut1_57[29] , \nOut1_57[28] , \nOut1_57[27] , 
        \nOut1_57[26] , \nOut1_57[25] , \nOut1_57[24] , \nOut1_57[23] , 
        \nOut1_57[22] , \nOut1_57[21] , \nOut1_57[20] , \nOut1_57[19] , 
        \nOut1_57[18] , \nOut1_57[17] , \nOut1_57[16] , \nOut1_57[15] , 
        \nOut1_57[14] , \nOut1_57[13] , \nOut1_57[12] , \nOut1_57[11] , 
        \nOut1_57[10] , \nOut1_57[9] , \nOut1_57[8] , \nOut1_57[7] , 
        \nOut1_57[6] , \nOut1_57[5] , \nOut1_57[4] , \nOut1_57[3] , 
        \nOut1_57[2] , \nOut1_57[1] , \nOut1_57[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_56[0] ), .NW_EDGE(\nOut0_55[0] ), .SW_EDGE(
        \nOut0_57[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut9[31] , \nScanOut9[30] , \nScanOut9[29] , 
        \nScanOut9[28] , \nScanOut9[27] , \nScanOut9[26] , \nScanOut9[25] , 
        \nScanOut9[24] , \nScanOut9[23] , \nScanOut9[22] , \nScanOut9[21] , 
        \nScanOut9[20] , \nScanOut9[19] , \nScanOut9[18] , \nScanOut9[17] , 
        \nScanOut9[16] , \nScanOut9[15] , \nScanOut9[14] , \nScanOut9[13] , 
        \nScanOut9[12] , \nScanOut9[11] , \nScanOut9[10] , \nScanOut9[9] , 
        \nScanOut9[8] , \nScanOut9[7] , \nScanOut9[6] , \nScanOut9[5] , 
        \nScanOut9[4] , \nScanOut9[3] , \nScanOut9[2] , \nScanOut9[1] , 
        \nScanOut9[0] }), .ScanOut({\nScanOut8[31] , \nScanOut8[30] , 
        \nScanOut8[29] , \nScanOut8[28] , \nScanOut8[27] , \nScanOut8[26] , 
        \nScanOut8[25] , \nScanOut8[24] , \nScanOut8[23] , \nScanOut8[22] , 
        \nScanOut8[21] , \nScanOut8[20] , \nScanOut8[19] , \nScanOut8[18] , 
        \nScanOut8[17] , \nScanOut8[16] , \nScanOut8[15] , \nScanOut8[14] , 
        \nScanOut8[13] , \nScanOut8[12] , \nScanOut8[11] , \nScanOut8[10] , 
        \nScanOut8[9] , \nScanOut8[8] , \nScanOut8[7] , \nScanOut8[6] , 
        \nScanOut8[5] , \nScanOut8[4] , \nScanOut8[3] , \nScanOut8[2] , 
        \nScanOut8[1] , \nScanOut8[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_8[31] , 
        \nOut0_8[30] , \nOut0_8[29] , \nOut0_8[28] , \nOut0_8[27] , 
        \nOut0_8[26] , \nOut0_8[25] , \nOut0_8[24] , \nOut0_8[23] , 
        \nOut0_8[22] , \nOut0_8[21] , \nOut0_8[20] , \nOut0_8[19] , 
        \nOut0_8[18] , \nOut0_8[17] , \nOut0_8[16] , \nOut0_8[15] , 
        \nOut0_8[14] , \nOut0_8[13] , \nOut0_8[12] , \nOut0_8[11] , 
        \nOut0_8[10] , \nOut0_8[9] , \nOut0_8[8] , \nOut0_8[7] , \nOut0_8[6] , 
        \nOut0_8[5] , \nOut0_8[4] , \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , 
        \nOut0_8[0] }), .NORTH_EDGE({\nOut0_7[31] , \nOut0_7[30] , 
        \nOut0_7[29] , \nOut0_7[28] , \nOut0_7[27] , \nOut0_7[26] , 
        \nOut0_7[25] , \nOut0_7[24] , \nOut0_7[23] , \nOut0_7[22] , 
        \nOut0_7[21] , \nOut0_7[20] , \nOut0_7[19] , \nOut0_7[18] , 
        \nOut0_7[17] , \nOut0_7[16] , \nOut0_7[15] , \nOut0_7[14] , 
        \nOut0_7[13] , \nOut0_7[12] , \nOut0_7[11] , \nOut0_7[10] , 
        \nOut0_7[9] , \nOut0_7[8] , \nOut0_7[7] , \nOut0_7[6] , \nOut0_7[5] , 
        \nOut0_7[4] , \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , \nOut0_7[0] }), 
        .SOUTH_EDGE({\nOut0_9[31] , \nOut0_9[30] , \nOut0_9[29] , 
        \nOut0_9[28] , \nOut0_9[27] , \nOut0_9[26] , \nOut0_9[25] , 
        \nOut0_9[24] , \nOut0_9[23] , \nOut0_9[22] , \nOut0_9[21] , 
        \nOut0_9[20] , \nOut0_9[19] , \nOut0_9[18] , \nOut0_9[17] , 
        \nOut0_9[16] , \nOut0_9[15] , \nOut0_9[14] , \nOut0_9[13] , 
        \nOut0_9[12] , \nOut0_9[11] , \nOut0_9[10] , \nOut0_9[9] , 
        \nOut0_9[8] , \nOut0_9[7] , \nOut0_9[6] , \nOut0_9[5] , \nOut0_9[4] , 
        \nOut0_9[3] , \nOut0_9[2] , \nOut0_9[1] , \nOut0_9[0] }), .EAST_EDGE(
        \nOut1_8[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_7[31] ), .SE_EDGE(\nOut1_9[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_38 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut39[31] , \nScanOut39[30] , \nScanOut39[29] , 
        \nScanOut39[28] , \nScanOut39[27] , \nScanOut39[26] , \nScanOut39[25] , 
        \nScanOut39[24] , \nScanOut39[23] , \nScanOut39[22] , \nScanOut39[21] , 
        \nScanOut39[20] , \nScanOut39[19] , \nScanOut39[18] , \nScanOut39[17] , 
        \nScanOut39[16] , \nScanOut39[15] , \nScanOut39[14] , \nScanOut39[13] , 
        \nScanOut39[12] , \nScanOut39[11] , \nScanOut39[10] , \nScanOut39[9] , 
        \nScanOut39[8] , \nScanOut39[7] , \nScanOut39[6] , \nScanOut39[5] , 
        \nScanOut39[4] , \nScanOut39[3] , \nScanOut39[2] , \nScanOut39[1] , 
        \nScanOut39[0] }), .ScanOut({\nScanOut38[31] , \nScanOut38[30] , 
        \nScanOut38[29] , \nScanOut38[28] , \nScanOut38[27] , \nScanOut38[26] , 
        \nScanOut38[25] , \nScanOut38[24] , \nScanOut38[23] , \nScanOut38[22] , 
        \nScanOut38[21] , \nScanOut38[20] , \nScanOut38[19] , \nScanOut38[18] , 
        \nScanOut38[17] , \nScanOut38[16] , \nScanOut38[15] , \nScanOut38[14] , 
        \nScanOut38[13] , \nScanOut38[12] , \nScanOut38[11] , \nScanOut38[10] , 
        \nScanOut38[9] , \nScanOut38[8] , \nScanOut38[7] , \nScanOut38[6] , 
        \nScanOut38[5] , \nScanOut38[4] , \nScanOut38[3] , \nScanOut38[2] , 
        \nScanOut38[1] , \nScanOut38[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_38[31] , 
        \nOut0_38[30] , \nOut0_38[29] , \nOut0_38[28] , \nOut0_38[27] , 
        \nOut0_38[26] , \nOut0_38[25] , \nOut0_38[24] , \nOut0_38[23] , 
        \nOut0_38[22] , \nOut0_38[21] , \nOut0_38[20] , \nOut0_38[19] , 
        \nOut0_38[18] , \nOut0_38[17] , \nOut0_38[16] , \nOut0_38[15] , 
        \nOut0_38[14] , \nOut0_38[13] , \nOut0_38[12] , \nOut0_38[11] , 
        \nOut0_38[10] , \nOut0_38[9] , \nOut0_38[8] , \nOut0_38[7] , 
        \nOut0_38[6] , \nOut0_38[5] , \nOut0_38[4] , \nOut0_38[3] , 
        \nOut0_38[2] , \nOut0_38[1] , \nOut0_38[0] }), .NORTH_EDGE({
        \nOut0_37[31] , \nOut0_37[30] , \nOut0_37[29] , \nOut0_37[28] , 
        \nOut0_37[27] , \nOut0_37[26] , \nOut0_37[25] , \nOut0_37[24] , 
        \nOut0_37[23] , \nOut0_37[22] , \nOut0_37[21] , \nOut0_37[20] , 
        \nOut0_37[19] , \nOut0_37[18] , \nOut0_37[17] , \nOut0_37[16] , 
        \nOut0_37[15] , \nOut0_37[14] , \nOut0_37[13] , \nOut0_37[12] , 
        \nOut0_37[11] , \nOut0_37[10] , \nOut0_37[9] , \nOut0_37[8] , 
        \nOut0_37[7] , \nOut0_37[6] , \nOut0_37[5] , \nOut0_37[4] , 
        \nOut0_37[3] , \nOut0_37[2] , \nOut0_37[1] , \nOut0_37[0] }), 
        .SOUTH_EDGE({\nOut0_39[31] , \nOut0_39[30] , \nOut0_39[29] , 
        \nOut0_39[28] , \nOut0_39[27] , \nOut0_39[26] , \nOut0_39[25] , 
        \nOut0_39[24] , \nOut0_39[23] , \nOut0_39[22] , \nOut0_39[21] , 
        \nOut0_39[20] , \nOut0_39[19] , \nOut0_39[18] , \nOut0_39[17] , 
        \nOut0_39[16] , \nOut0_39[15] , \nOut0_39[14] , \nOut0_39[13] , 
        \nOut0_39[12] , \nOut0_39[11] , \nOut0_39[10] , \nOut0_39[9] , 
        \nOut0_39[8] , \nOut0_39[7] , \nOut0_39[6] , \nOut0_39[5] , 
        \nOut0_39[4] , \nOut0_39[3] , \nOut0_39[2] , \nOut0_39[1] , 
        \nOut0_39[0] }), .EAST_EDGE(\nOut1_38[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_37[31] ), .SE_EDGE(
        \nOut1_39[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_56 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut57[31] , \nScanOut57[30] , \nScanOut57[29] , 
        \nScanOut57[28] , \nScanOut57[27] , \nScanOut57[26] , \nScanOut57[25] , 
        \nScanOut57[24] , \nScanOut57[23] , \nScanOut57[22] , \nScanOut57[21] , 
        \nScanOut57[20] , \nScanOut57[19] , \nScanOut57[18] , \nScanOut57[17] , 
        \nScanOut57[16] , \nScanOut57[15] , \nScanOut57[14] , \nScanOut57[13] , 
        \nScanOut57[12] , \nScanOut57[11] , \nScanOut57[10] , \nScanOut57[9] , 
        \nScanOut57[8] , \nScanOut57[7] , \nScanOut57[6] , \nScanOut57[5] , 
        \nScanOut57[4] , \nScanOut57[3] , \nScanOut57[2] , \nScanOut57[1] , 
        \nScanOut57[0] }), .ScanOut({\nScanOut56[31] , \nScanOut56[30] , 
        \nScanOut56[29] , \nScanOut56[28] , \nScanOut56[27] , \nScanOut56[26] , 
        \nScanOut56[25] , \nScanOut56[24] , \nScanOut56[23] , \nScanOut56[22] , 
        \nScanOut56[21] , \nScanOut56[20] , \nScanOut56[19] , \nScanOut56[18] , 
        \nScanOut56[17] , \nScanOut56[16] , \nScanOut56[15] , \nScanOut56[14] , 
        \nScanOut56[13] , \nScanOut56[12] , \nScanOut56[11] , \nScanOut56[10] , 
        \nScanOut56[9] , \nScanOut56[8] , \nScanOut56[7] , \nScanOut56[6] , 
        \nScanOut56[5] , \nScanOut56[4] , \nScanOut56[3] , \nScanOut56[2] , 
        \nScanOut56[1] , \nScanOut56[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_56[31] , 
        \nOut0_56[30] , \nOut0_56[29] , \nOut0_56[28] , \nOut0_56[27] , 
        \nOut0_56[26] , \nOut0_56[25] , \nOut0_56[24] , \nOut0_56[23] , 
        \nOut0_56[22] , \nOut0_56[21] , \nOut0_56[20] , \nOut0_56[19] , 
        \nOut0_56[18] , \nOut0_56[17] , \nOut0_56[16] , \nOut0_56[15] , 
        \nOut0_56[14] , \nOut0_56[13] , \nOut0_56[12] , \nOut0_56[11] , 
        \nOut0_56[10] , \nOut0_56[9] , \nOut0_56[8] , \nOut0_56[7] , 
        \nOut0_56[6] , \nOut0_56[5] , \nOut0_56[4] , \nOut0_56[3] , 
        \nOut0_56[2] , \nOut0_56[1] , \nOut0_56[0] }), .NORTH_EDGE({
        \nOut0_55[31] , \nOut0_55[30] , \nOut0_55[29] , \nOut0_55[28] , 
        \nOut0_55[27] , \nOut0_55[26] , \nOut0_55[25] , \nOut0_55[24] , 
        \nOut0_55[23] , \nOut0_55[22] , \nOut0_55[21] , \nOut0_55[20] , 
        \nOut0_55[19] , \nOut0_55[18] , \nOut0_55[17] , \nOut0_55[16] , 
        \nOut0_55[15] , \nOut0_55[14] , \nOut0_55[13] , \nOut0_55[12] , 
        \nOut0_55[11] , \nOut0_55[10] , \nOut0_55[9] , \nOut0_55[8] , 
        \nOut0_55[7] , \nOut0_55[6] , \nOut0_55[5] , \nOut0_55[4] , 
        \nOut0_55[3] , \nOut0_55[2] , \nOut0_55[1] , \nOut0_55[0] }), 
        .SOUTH_EDGE({\nOut0_57[31] , \nOut0_57[30] , \nOut0_57[29] , 
        \nOut0_57[28] , \nOut0_57[27] , \nOut0_57[26] , \nOut0_57[25] , 
        \nOut0_57[24] , \nOut0_57[23] , \nOut0_57[22] , \nOut0_57[21] , 
        \nOut0_57[20] , \nOut0_57[19] , \nOut0_57[18] , \nOut0_57[17] , 
        \nOut0_57[16] , \nOut0_57[15] , \nOut0_57[14] , \nOut0_57[13] , 
        \nOut0_57[12] , \nOut0_57[11] , \nOut0_57[10] , \nOut0_57[9] , 
        \nOut0_57[8] , \nOut0_57[7] , \nOut0_57[6] , \nOut0_57[5] , 
        \nOut0_57[4] , \nOut0_57[3] , \nOut0_57[2] , \nOut0_57[1] , 
        \nOut0_57[0] }), .EAST_EDGE(\nOut1_56[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_55[31] ), .SE_EDGE(
        \nOut1_57[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_71 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut72[31] , \nScanOut72[30] , \nScanOut72[29] , 
        \nScanOut72[28] , \nScanOut72[27] , \nScanOut72[26] , \nScanOut72[25] , 
        \nScanOut72[24] , \nScanOut72[23] , \nScanOut72[22] , \nScanOut72[21] , 
        \nScanOut72[20] , \nScanOut72[19] , \nScanOut72[18] , \nScanOut72[17] , 
        \nScanOut72[16] , \nScanOut72[15] , \nScanOut72[14] , \nScanOut72[13] , 
        \nScanOut72[12] , \nScanOut72[11] , \nScanOut72[10] , \nScanOut72[9] , 
        \nScanOut72[8] , \nScanOut72[7] , \nScanOut72[6] , \nScanOut72[5] , 
        \nScanOut72[4] , \nScanOut72[3] , \nScanOut72[2] , \nScanOut72[1] , 
        \nScanOut72[0] }), .ScanOut({\nScanOut71[31] , \nScanOut71[30] , 
        \nScanOut71[29] , \nScanOut71[28] , \nScanOut71[27] , \nScanOut71[26] , 
        \nScanOut71[25] , \nScanOut71[24] , \nScanOut71[23] , \nScanOut71[22] , 
        \nScanOut71[21] , \nScanOut71[20] , \nScanOut71[19] , \nScanOut71[18] , 
        \nScanOut71[17] , \nScanOut71[16] , \nScanOut71[15] , \nScanOut71[14] , 
        \nScanOut71[13] , \nScanOut71[12] , \nScanOut71[11] , \nScanOut71[10] , 
        \nScanOut71[9] , \nScanOut71[8] , \nScanOut71[7] , \nScanOut71[6] , 
        \nScanOut71[5] , \nScanOut71[4] , \nScanOut71[3] , \nScanOut71[2] , 
        \nScanOut71[1] , \nScanOut71[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_7[31] , 
        \nOut1_7[30] , \nOut1_7[29] , \nOut1_7[28] , \nOut1_7[27] , 
        \nOut1_7[26] , \nOut1_7[25] , \nOut1_7[24] , \nOut1_7[23] , 
        \nOut1_7[22] , \nOut1_7[21] , \nOut1_7[20] , \nOut1_7[19] , 
        \nOut1_7[18] , \nOut1_7[17] , \nOut1_7[16] , \nOut1_7[15] , 
        \nOut1_7[14] , \nOut1_7[13] , \nOut1_7[12] , \nOut1_7[11] , 
        \nOut1_7[10] , \nOut1_7[9] , \nOut1_7[8] , \nOut1_7[7] , \nOut1_7[6] , 
        \nOut1_7[5] , \nOut1_7[4] , \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , 
        \nOut1_7[0] }), .NORTH_EDGE({\nOut1_6[31] , \nOut1_6[30] , 
        \nOut1_6[29] , \nOut1_6[28] , \nOut1_6[27] , \nOut1_6[26] , 
        \nOut1_6[25] , \nOut1_6[24] , \nOut1_6[23] , \nOut1_6[22] , 
        \nOut1_6[21] , \nOut1_6[20] , \nOut1_6[19] , \nOut1_6[18] , 
        \nOut1_6[17] , \nOut1_6[16] , \nOut1_6[15] , \nOut1_6[14] , 
        \nOut1_6[13] , \nOut1_6[12] , \nOut1_6[11] , \nOut1_6[10] , 
        \nOut1_6[9] , \nOut1_6[8] , \nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , 
        \nOut1_6[4] , \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }), 
        .SOUTH_EDGE({\nOut1_8[31] , \nOut1_8[30] , \nOut1_8[29] , 
        \nOut1_8[28] , \nOut1_8[27] , \nOut1_8[26] , \nOut1_8[25] , 
        \nOut1_8[24] , \nOut1_8[23] , \nOut1_8[22] , \nOut1_8[21] , 
        \nOut1_8[20] , \nOut1_8[19] , \nOut1_8[18] , \nOut1_8[17] , 
        \nOut1_8[16] , \nOut1_8[15] , \nOut1_8[14] , \nOut1_8[13] , 
        \nOut1_8[12] , \nOut1_8[11] , \nOut1_8[10] , \nOut1_8[9] , 
        \nOut1_8[8] , \nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , \nOut1_8[4] , 
        \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut0_7[0] ), .NW_EDGE(\nOut0_6[0] ), .SW_EDGE(
        \nOut0_8[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_127 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut128[31] , \nScanOut128[30] , \nScanOut128[29] , 
        \nScanOut128[28] , \nScanOut128[27] , \nScanOut128[26] , 
        \nScanOut128[25] , \nScanOut128[24] , \nScanOut128[23] , 
        \nScanOut128[22] , \nScanOut128[21] , \nScanOut128[20] , 
        \nScanOut128[19] , \nScanOut128[18] , \nScanOut128[17] , 
        \nScanOut128[16] , \nScanOut128[15] , \nScanOut128[14] , 
        \nScanOut128[13] , \nScanOut128[12] , \nScanOut128[11] , 
        \nScanOut128[10] , \nScanOut128[9] , \nScanOut128[8] , 
        \nScanOut128[7] , \nScanOut128[6] , \nScanOut128[5] , \nScanOut128[4] , 
        \nScanOut128[3] , \nScanOut128[2] , \nScanOut128[1] , \nScanOut128[0] 
        }), .ScanOut({\nScanOut127[31] , \nScanOut127[30] , \nScanOut127[29] , 
        \nScanOut127[28] , \nScanOut127[27] , \nScanOut127[26] , 
        \nScanOut127[25] , \nScanOut127[24] , \nScanOut127[23] , 
        \nScanOut127[22] , \nScanOut127[21] , \nScanOut127[20] , 
        \nScanOut127[19] , \nScanOut127[18] , \nScanOut127[17] , 
        \nScanOut127[16] , \nScanOut127[15] , \nScanOut127[14] , 
        \nScanOut127[13] , \nScanOut127[12] , \nScanOut127[11] , 
        \nScanOut127[10] , \nScanOut127[9] , \nScanOut127[8] , 
        \nScanOut127[7] , \nScanOut127[6] , \nScanOut127[5] , \nScanOut127[4] , 
        \nScanOut127[3] , \nScanOut127[2] , \nScanOut127[1] , \nScanOut127[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_63[31] , \nOut1_63[30] , \nOut1_63[29] , 
        \nOut1_63[28] , \nOut1_63[27] , \nOut1_63[26] , \nOut1_63[25] , 
        \nOut1_63[24] , \nOut1_63[23] , \nOut1_63[22] , \nOut1_63[21] , 
        \nOut1_63[20] , \nOut1_63[19] , \nOut1_63[18] , \nOut1_63[17] , 
        \nOut1_63[16] , \nOut1_63[15] , \nOut1_63[14] , \nOut1_63[13] , 
        \nOut1_63[12] , \nOut1_63[11] , \nOut1_63[10] , \nOut1_63[9] , 
        \nOut1_63[8] , \nOut1_63[7] , \nOut1_63[6] , \nOut1_63[5] , 
        \nOut1_63[4] , \nOut1_63[3] , \nOut1_63[2] , \nOut1_63[1] , 
        \nOut1_63[0] }), .NORTH_EDGE({\nOut1_62[31] , \nOut1_62[30] , 
        \nOut1_62[29] , \nOut1_62[28] , \nOut1_62[27] , \nOut1_62[26] , 
        \nOut1_62[25] , \nOut1_62[24] , \nOut1_62[23] , \nOut1_62[22] , 
        \nOut1_62[21] , \nOut1_62[20] , \nOut1_62[19] , \nOut1_62[18] , 
        \nOut1_62[17] , \nOut1_62[16] , \nOut1_62[15] , \nOut1_62[14] , 
        \nOut1_62[13] , \nOut1_62[12] , \nOut1_62[11] , \nOut1_62[10] , 
        \nOut1_62[9] , \nOut1_62[8] , \nOut1_62[7] , \nOut1_62[6] , 
        \nOut1_62[5] , \nOut1_62[4] , \nOut1_62[3] , \nOut1_62[2] , 
        \nOut1_62[1] , \nOut1_62[0] }), .SOUTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_63[0] ), 
        .NW_EDGE(\nOut0_62[0] ), .SW_EDGE(1'b0), .NE_EDGE(1'b0), .SE_EDGE(1'b0
        ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_100 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut101[31] , \nScanOut101[30] , \nScanOut101[29] , 
        \nScanOut101[28] , \nScanOut101[27] , \nScanOut101[26] , 
        \nScanOut101[25] , \nScanOut101[24] , \nScanOut101[23] , 
        \nScanOut101[22] , \nScanOut101[21] , \nScanOut101[20] , 
        \nScanOut101[19] , \nScanOut101[18] , \nScanOut101[17] , 
        \nScanOut101[16] , \nScanOut101[15] , \nScanOut101[14] , 
        \nScanOut101[13] , \nScanOut101[12] , \nScanOut101[11] , 
        \nScanOut101[10] , \nScanOut101[9] , \nScanOut101[8] , 
        \nScanOut101[7] , \nScanOut101[6] , \nScanOut101[5] , \nScanOut101[4] , 
        \nScanOut101[3] , \nScanOut101[2] , \nScanOut101[1] , \nScanOut101[0] 
        }), .ScanOut({\nScanOut100[31] , \nScanOut100[30] , \nScanOut100[29] , 
        \nScanOut100[28] , \nScanOut100[27] , \nScanOut100[26] , 
        \nScanOut100[25] , \nScanOut100[24] , \nScanOut100[23] , 
        \nScanOut100[22] , \nScanOut100[21] , \nScanOut100[20] , 
        \nScanOut100[19] , \nScanOut100[18] , \nScanOut100[17] , 
        \nScanOut100[16] , \nScanOut100[15] , \nScanOut100[14] , 
        \nScanOut100[13] , \nScanOut100[12] , \nScanOut100[11] , 
        \nScanOut100[10] , \nScanOut100[9] , \nScanOut100[8] , 
        \nScanOut100[7] , \nScanOut100[6] , \nScanOut100[5] , \nScanOut100[4] , 
        \nScanOut100[3] , \nScanOut100[2] , \nScanOut100[1] , \nScanOut100[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_36[31] , \nOut1_36[30] , \nOut1_36[29] , 
        \nOut1_36[28] , \nOut1_36[27] , \nOut1_36[26] , \nOut1_36[25] , 
        \nOut1_36[24] , \nOut1_36[23] , \nOut1_36[22] , \nOut1_36[21] , 
        \nOut1_36[20] , \nOut1_36[19] , \nOut1_36[18] , \nOut1_36[17] , 
        \nOut1_36[16] , \nOut1_36[15] , \nOut1_36[14] , \nOut1_36[13] , 
        \nOut1_36[12] , \nOut1_36[11] , \nOut1_36[10] , \nOut1_36[9] , 
        \nOut1_36[8] , \nOut1_36[7] , \nOut1_36[6] , \nOut1_36[5] , 
        \nOut1_36[4] , \nOut1_36[3] , \nOut1_36[2] , \nOut1_36[1] , 
        \nOut1_36[0] }), .NORTH_EDGE({\nOut1_35[31] , \nOut1_35[30] , 
        \nOut1_35[29] , \nOut1_35[28] , \nOut1_35[27] , \nOut1_35[26] , 
        \nOut1_35[25] , \nOut1_35[24] , \nOut1_35[23] , \nOut1_35[22] , 
        \nOut1_35[21] , \nOut1_35[20] , \nOut1_35[19] , \nOut1_35[18] , 
        \nOut1_35[17] , \nOut1_35[16] , \nOut1_35[15] , \nOut1_35[14] , 
        \nOut1_35[13] , \nOut1_35[12] , \nOut1_35[11] , \nOut1_35[10] , 
        \nOut1_35[9] , \nOut1_35[8] , \nOut1_35[7] , \nOut1_35[6] , 
        \nOut1_35[5] , \nOut1_35[4] , \nOut1_35[3] , \nOut1_35[2] , 
        \nOut1_35[1] , \nOut1_35[0] }), .SOUTH_EDGE({\nOut1_37[31] , 
        \nOut1_37[30] , \nOut1_37[29] , \nOut1_37[28] , \nOut1_37[27] , 
        \nOut1_37[26] , \nOut1_37[25] , \nOut1_37[24] , \nOut1_37[23] , 
        \nOut1_37[22] , \nOut1_37[21] , \nOut1_37[20] , \nOut1_37[19] , 
        \nOut1_37[18] , \nOut1_37[17] , \nOut1_37[16] , \nOut1_37[15] , 
        \nOut1_37[14] , \nOut1_37[13] , \nOut1_37[12] , \nOut1_37[11] , 
        \nOut1_37[10] , \nOut1_37[9] , \nOut1_37[8] , \nOut1_37[7] , 
        \nOut1_37[6] , \nOut1_37[5] , \nOut1_37[4] , \nOut1_37[3] , 
        \nOut1_37[2] , \nOut1_37[1] , \nOut1_37[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_36[0] ), .NW_EDGE(\nOut0_35[0] ), .SW_EDGE(
        \nOut0_37[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_44 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut45[31] , \nScanOut45[30] , \nScanOut45[29] , 
        \nScanOut45[28] , \nScanOut45[27] , \nScanOut45[26] , \nScanOut45[25] , 
        \nScanOut45[24] , \nScanOut45[23] , \nScanOut45[22] , \nScanOut45[21] , 
        \nScanOut45[20] , \nScanOut45[19] , \nScanOut45[18] , \nScanOut45[17] , 
        \nScanOut45[16] , \nScanOut45[15] , \nScanOut45[14] , \nScanOut45[13] , 
        \nScanOut45[12] , \nScanOut45[11] , \nScanOut45[10] , \nScanOut45[9] , 
        \nScanOut45[8] , \nScanOut45[7] , \nScanOut45[6] , \nScanOut45[5] , 
        \nScanOut45[4] , \nScanOut45[3] , \nScanOut45[2] , \nScanOut45[1] , 
        \nScanOut45[0] }), .ScanOut({\nScanOut44[31] , \nScanOut44[30] , 
        \nScanOut44[29] , \nScanOut44[28] , \nScanOut44[27] , \nScanOut44[26] , 
        \nScanOut44[25] , \nScanOut44[24] , \nScanOut44[23] , \nScanOut44[22] , 
        \nScanOut44[21] , \nScanOut44[20] , \nScanOut44[19] , \nScanOut44[18] , 
        \nScanOut44[17] , \nScanOut44[16] , \nScanOut44[15] , \nScanOut44[14] , 
        \nScanOut44[13] , \nScanOut44[12] , \nScanOut44[11] , \nScanOut44[10] , 
        \nScanOut44[9] , \nScanOut44[8] , \nScanOut44[7] , \nScanOut44[6] , 
        \nScanOut44[5] , \nScanOut44[4] , \nScanOut44[3] , \nScanOut44[2] , 
        \nScanOut44[1] , \nScanOut44[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_44[31] , 
        \nOut0_44[30] , \nOut0_44[29] , \nOut0_44[28] , \nOut0_44[27] , 
        \nOut0_44[26] , \nOut0_44[25] , \nOut0_44[24] , \nOut0_44[23] , 
        \nOut0_44[22] , \nOut0_44[21] , \nOut0_44[20] , \nOut0_44[19] , 
        \nOut0_44[18] , \nOut0_44[17] , \nOut0_44[16] , \nOut0_44[15] , 
        \nOut0_44[14] , \nOut0_44[13] , \nOut0_44[12] , \nOut0_44[11] , 
        \nOut0_44[10] , \nOut0_44[9] , \nOut0_44[8] , \nOut0_44[7] , 
        \nOut0_44[6] , \nOut0_44[5] , \nOut0_44[4] , \nOut0_44[3] , 
        \nOut0_44[2] , \nOut0_44[1] , \nOut0_44[0] }), .NORTH_EDGE({
        \nOut0_43[31] , \nOut0_43[30] , \nOut0_43[29] , \nOut0_43[28] , 
        \nOut0_43[27] , \nOut0_43[26] , \nOut0_43[25] , \nOut0_43[24] , 
        \nOut0_43[23] , \nOut0_43[22] , \nOut0_43[21] , \nOut0_43[20] , 
        \nOut0_43[19] , \nOut0_43[18] , \nOut0_43[17] , \nOut0_43[16] , 
        \nOut0_43[15] , \nOut0_43[14] , \nOut0_43[13] , \nOut0_43[12] , 
        \nOut0_43[11] , \nOut0_43[10] , \nOut0_43[9] , \nOut0_43[8] , 
        \nOut0_43[7] , \nOut0_43[6] , \nOut0_43[5] , \nOut0_43[4] , 
        \nOut0_43[3] , \nOut0_43[2] , \nOut0_43[1] , \nOut0_43[0] }), 
        .SOUTH_EDGE({\nOut0_45[31] , \nOut0_45[30] , \nOut0_45[29] , 
        \nOut0_45[28] , \nOut0_45[27] , \nOut0_45[26] , \nOut0_45[25] , 
        \nOut0_45[24] , \nOut0_45[23] , \nOut0_45[22] , \nOut0_45[21] , 
        \nOut0_45[20] , \nOut0_45[19] , \nOut0_45[18] , \nOut0_45[17] , 
        \nOut0_45[16] , \nOut0_45[15] , \nOut0_45[14] , \nOut0_45[13] , 
        \nOut0_45[12] , \nOut0_45[11] , \nOut0_45[10] , \nOut0_45[9] , 
        \nOut0_45[8] , \nOut0_45[7] , \nOut0_45[6] , \nOut0_45[5] , 
        \nOut0_45[4] , \nOut0_45[3] , \nOut0_45[2] , \nOut0_45[1] , 
        \nOut0_45[0] }), .EAST_EDGE(\nOut1_44[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_43[31] ), .SE_EDGE(
        \nOut1_45[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_63 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut64[31] , \nScanOut64[30] , \nScanOut64[29] , 
        \nScanOut64[28] , \nScanOut64[27] , \nScanOut64[26] , \nScanOut64[25] , 
        \nScanOut64[24] , \nScanOut64[23] , \nScanOut64[22] , \nScanOut64[21] , 
        \nScanOut64[20] , \nScanOut64[19] , \nScanOut64[18] , \nScanOut64[17] , 
        \nScanOut64[16] , \nScanOut64[15] , \nScanOut64[14] , \nScanOut64[13] , 
        \nScanOut64[12] , \nScanOut64[11] , \nScanOut64[10] , \nScanOut64[9] , 
        \nScanOut64[8] , \nScanOut64[7] , \nScanOut64[6] , \nScanOut64[5] , 
        \nScanOut64[4] , \nScanOut64[3] , \nScanOut64[2] , \nScanOut64[1] , 
        \nScanOut64[0] }), .ScanOut({\nScanOut63[31] , \nScanOut63[30] , 
        \nScanOut63[29] , \nScanOut63[28] , \nScanOut63[27] , \nScanOut63[26] , 
        \nScanOut63[25] , \nScanOut63[24] , \nScanOut63[23] , \nScanOut63[22] , 
        \nScanOut63[21] , \nScanOut63[20] , \nScanOut63[19] , \nScanOut63[18] , 
        \nScanOut63[17] , \nScanOut63[16] , \nScanOut63[15] , \nScanOut63[14] , 
        \nScanOut63[13] , \nScanOut63[12] , \nScanOut63[11] , \nScanOut63[10] , 
        \nScanOut63[9] , \nScanOut63[8] , \nScanOut63[7] , \nScanOut63[6] , 
        \nScanOut63[5] , \nScanOut63[4] , \nScanOut63[3] , \nScanOut63[2] , 
        \nScanOut63[1] , \nScanOut63[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_63[31] , 
        \nOut0_63[30] , \nOut0_63[29] , \nOut0_63[28] , \nOut0_63[27] , 
        \nOut0_63[26] , \nOut0_63[25] , \nOut0_63[24] , \nOut0_63[23] , 
        \nOut0_63[22] , \nOut0_63[21] , \nOut0_63[20] , \nOut0_63[19] , 
        \nOut0_63[18] , \nOut0_63[17] , \nOut0_63[16] , \nOut0_63[15] , 
        \nOut0_63[14] , \nOut0_63[13] , \nOut0_63[12] , \nOut0_63[11] , 
        \nOut0_63[10] , \nOut0_63[9] , \nOut0_63[8] , \nOut0_63[7] , 
        \nOut0_63[6] , \nOut0_63[5] , \nOut0_63[4] , \nOut0_63[3] , 
        \nOut0_63[2] , \nOut0_63[1] , \nOut0_63[0] }), .NORTH_EDGE({
        \nOut0_62[31] , \nOut0_62[30] , \nOut0_62[29] , \nOut0_62[28] , 
        \nOut0_62[27] , \nOut0_62[26] , \nOut0_62[25] , \nOut0_62[24] , 
        \nOut0_62[23] , \nOut0_62[22] , \nOut0_62[21] , \nOut0_62[20] , 
        \nOut0_62[19] , \nOut0_62[18] , \nOut0_62[17] , \nOut0_62[16] , 
        \nOut0_62[15] , \nOut0_62[14] , \nOut0_62[13] , \nOut0_62[12] , 
        \nOut0_62[11] , \nOut0_62[10] , \nOut0_62[9] , \nOut0_62[8] , 
        \nOut0_62[7] , \nOut0_62[6] , \nOut0_62[5] , \nOut0_62[4] , 
        \nOut0_62[3] , \nOut0_62[2] , \nOut0_62[1] , \nOut0_62[0] }), 
        .SOUTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .EAST_EDGE(\nOut1_63[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), 
        .SW_EDGE(1'b0), .NE_EDGE(\nOut1_62[31] ), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_86 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut87[31] , \nScanOut87[30] , \nScanOut87[29] , 
        \nScanOut87[28] , \nScanOut87[27] , \nScanOut87[26] , \nScanOut87[25] , 
        \nScanOut87[24] , \nScanOut87[23] , \nScanOut87[22] , \nScanOut87[21] , 
        \nScanOut87[20] , \nScanOut87[19] , \nScanOut87[18] , \nScanOut87[17] , 
        \nScanOut87[16] , \nScanOut87[15] , \nScanOut87[14] , \nScanOut87[13] , 
        \nScanOut87[12] , \nScanOut87[11] , \nScanOut87[10] , \nScanOut87[9] , 
        \nScanOut87[8] , \nScanOut87[7] , \nScanOut87[6] , \nScanOut87[5] , 
        \nScanOut87[4] , \nScanOut87[3] , \nScanOut87[2] , \nScanOut87[1] , 
        \nScanOut87[0] }), .ScanOut({\nScanOut86[31] , \nScanOut86[30] , 
        \nScanOut86[29] , \nScanOut86[28] , \nScanOut86[27] , \nScanOut86[26] , 
        \nScanOut86[25] , \nScanOut86[24] , \nScanOut86[23] , \nScanOut86[22] , 
        \nScanOut86[21] , \nScanOut86[20] , \nScanOut86[19] , \nScanOut86[18] , 
        \nScanOut86[17] , \nScanOut86[16] , \nScanOut86[15] , \nScanOut86[14] , 
        \nScanOut86[13] , \nScanOut86[12] , \nScanOut86[11] , \nScanOut86[10] , 
        \nScanOut86[9] , \nScanOut86[8] , \nScanOut86[7] , \nScanOut86[6] , 
        \nScanOut86[5] , \nScanOut86[4] , \nScanOut86[3] , \nScanOut86[2] , 
        \nScanOut86[1] , \nScanOut86[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_22[31] , 
        \nOut1_22[30] , \nOut1_22[29] , \nOut1_22[28] , \nOut1_22[27] , 
        \nOut1_22[26] , \nOut1_22[25] , \nOut1_22[24] , \nOut1_22[23] , 
        \nOut1_22[22] , \nOut1_22[21] , \nOut1_22[20] , \nOut1_22[19] , 
        \nOut1_22[18] , \nOut1_22[17] , \nOut1_22[16] , \nOut1_22[15] , 
        \nOut1_22[14] , \nOut1_22[13] , \nOut1_22[12] , \nOut1_22[11] , 
        \nOut1_22[10] , \nOut1_22[9] , \nOut1_22[8] , \nOut1_22[7] , 
        \nOut1_22[6] , \nOut1_22[5] , \nOut1_22[4] , \nOut1_22[3] , 
        \nOut1_22[2] , \nOut1_22[1] , \nOut1_22[0] }), .NORTH_EDGE({
        \nOut1_21[31] , \nOut1_21[30] , \nOut1_21[29] , \nOut1_21[28] , 
        \nOut1_21[27] , \nOut1_21[26] , \nOut1_21[25] , \nOut1_21[24] , 
        \nOut1_21[23] , \nOut1_21[22] , \nOut1_21[21] , \nOut1_21[20] , 
        \nOut1_21[19] , \nOut1_21[18] , \nOut1_21[17] , \nOut1_21[16] , 
        \nOut1_21[15] , \nOut1_21[14] , \nOut1_21[13] , \nOut1_21[12] , 
        \nOut1_21[11] , \nOut1_21[10] , \nOut1_21[9] , \nOut1_21[8] , 
        \nOut1_21[7] , \nOut1_21[6] , \nOut1_21[5] , \nOut1_21[4] , 
        \nOut1_21[3] , \nOut1_21[2] , \nOut1_21[1] , \nOut1_21[0] }), 
        .SOUTH_EDGE({\nOut1_23[31] , \nOut1_23[30] , \nOut1_23[29] , 
        \nOut1_23[28] , \nOut1_23[27] , \nOut1_23[26] , \nOut1_23[25] , 
        \nOut1_23[24] , \nOut1_23[23] , \nOut1_23[22] , \nOut1_23[21] , 
        \nOut1_23[20] , \nOut1_23[19] , \nOut1_23[18] , \nOut1_23[17] , 
        \nOut1_23[16] , \nOut1_23[15] , \nOut1_23[14] , \nOut1_23[13] , 
        \nOut1_23[12] , \nOut1_23[11] , \nOut1_23[10] , \nOut1_23[9] , 
        \nOut1_23[8] , \nOut1_23[7] , \nOut1_23[6] , \nOut1_23[5] , 
        \nOut1_23[4] , \nOut1_23[3] , \nOut1_23[2] , \nOut1_23[1] , 
        \nOut1_23[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_22[0] ), 
        .NW_EDGE(\nOut0_21[0] ), .SW_EDGE(\nOut0_23[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_94 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut95[31] , \nScanOut95[30] , \nScanOut95[29] , 
        \nScanOut95[28] , \nScanOut95[27] , \nScanOut95[26] , \nScanOut95[25] , 
        \nScanOut95[24] , \nScanOut95[23] , \nScanOut95[22] , \nScanOut95[21] , 
        \nScanOut95[20] , \nScanOut95[19] , \nScanOut95[18] , \nScanOut95[17] , 
        \nScanOut95[16] , \nScanOut95[15] , \nScanOut95[14] , \nScanOut95[13] , 
        \nScanOut95[12] , \nScanOut95[11] , \nScanOut95[10] , \nScanOut95[9] , 
        \nScanOut95[8] , \nScanOut95[7] , \nScanOut95[6] , \nScanOut95[5] , 
        \nScanOut95[4] , \nScanOut95[3] , \nScanOut95[2] , \nScanOut95[1] , 
        \nScanOut95[0] }), .ScanOut({\nScanOut94[31] , \nScanOut94[30] , 
        \nScanOut94[29] , \nScanOut94[28] , \nScanOut94[27] , \nScanOut94[26] , 
        \nScanOut94[25] , \nScanOut94[24] , \nScanOut94[23] , \nScanOut94[22] , 
        \nScanOut94[21] , \nScanOut94[20] , \nScanOut94[19] , \nScanOut94[18] , 
        \nScanOut94[17] , \nScanOut94[16] , \nScanOut94[15] , \nScanOut94[14] , 
        \nScanOut94[13] , \nScanOut94[12] , \nScanOut94[11] , \nScanOut94[10] , 
        \nScanOut94[9] , \nScanOut94[8] , \nScanOut94[7] , \nScanOut94[6] , 
        \nScanOut94[5] , \nScanOut94[4] , \nScanOut94[3] , \nScanOut94[2] , 
        \nScanOut94[1] , \nScanOut94[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_30[31] , 
        \nOut1_30[30] , \nOut1_30[29] , \nOut1_30[28] , \nOut1_30[27] , 
        \nOut1_30[26] , \nOut1_30[25] , \nOut1_30[24] , \nOut1_30[23] , 
        \nOut1_30[22] , \nOut1_30[21] , \nOut1_30[20] , \nOut1_30[19] , 
        \nOut1_30[18] , \nOut1_30[17] , \nOut1_30[16] , \nOut1_30[15] , 
        \nOut1_30[14] , \nOut1_30[13] , \nOut1_30[12] , \nOut1_30[11] , 
        \nOut1_30[10] , \nOut1_30[9] , \nOut1_30[8] , \nOut1_30[7] , 
        \nOut1_30[6] , \nOut1_30[5] , \nOut1_30[4] , \nOut1_30[3] , 
        \nOut1_30[2] , \nOut1_30[1] , \nOut1_30[0] }), .NORTH_EDGE({
        \nOut1_29[31] , \nOut1_29[30] , \nOut1_29[29] , \nOut1_29[28] , 
        \nOut1_29[27] , \nOut1_29[26] , \nOut1_29[25] , \nOut1_29[24] , 
        \nOut1_29[23] , \nOut1_29[22] , \nOut1_29[21] , \nOut1_29[20] , 
        \nOut1_29[19] , \nOut1_29[18] , \nOut1_29[17] , \nOut1_29[16] , 
        \nOut1_29[15] , \nOut1_29[14] , \nOut1_29[13] , \nOut1_29[12] , 
        \nOut1_29[11] , \nOut1_29[10] , \nOut1_29[9] , \nOut1_29[8] , 
        \nOut1_29[7] , \nOut1_29[6] , \nOut1_29[5] , \nOut1_29[4] , 
        \nOut1_29[3] , \nOut1_29[2] , \nOut1_29[1] , \nOut1_29[0] }), 
        .SOUTH_EDGE({\nOut1_31[31] , \nOut1_31[30] , \nOut1_31[29] , 
        \nOut1_31[28] , \nOut1_31[27] , \nOut1_31[26] , \nOut1_31[25] , 
        \nOut1_31[24] , \nOut1_31[23] , \nOut1_31[22] , \nOut1_31[21] , 
        \nOut1_31[20] , \nOut1_31[19] , \nOut1_31[18] , \nOut1_31[17] , 
        \nOut1_31[16] , \nOut1_31[15] , \nOut1_31[14] , \nOut1_31[13] , 
        \nOut1_31[12] , \nOut1_31[11] , \nOut1_31[10] , \nOut1_31[9] , 
        \nOut1_31[8] , \nOut1_31[7] , \nOut1_31[6] , \nOut1_31[5] , 
        \nOut1_31[4] , \nOut1_31[3] , \nOut1_31[2] , \nOut1_31[1] , 
        \nOut1_31[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_30[0] ), 
        .NW_EDGE(\nOut0_29[0] ), .SW_EDGE(\nOut0_31[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_112 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut113[31] , \nScanOut113[30] , \nScanOut113[29] , 
        \nScanOut113[28] , \nScanOut113[27] , \nScanOut113[26] , 
        \nScanOut113[25] , \nScanOut113[24] , \nScanOut113[23] , 
        \nScanOut113[22] , \nScanOut113[21] , \nScanOut113[20] , 
        \nScanOut113[19] , \nScanOut113[18] , \nScanOut113[17] , 
        \nScanOut113[16] , \nScanOut113[15] , \nScanOut113[14] , 
        \nScanOut113[13] , \nScanOut113[12] , \nScanOut113[11] , 
        \nScanOut113[10] , \nScanOut113[9] , \nScanOut113[8] , 
        \nScanOut113[7] , \nScanOut113[6] , \nScanOut113[5] , \nScanOut113[4] , 
        \nScanOut113[3] , \nScanOut113[2] , \nScanOut113[1] , \nScanOut113[0] 
        }), .ScanOut({\nScanOut112[31] , \nScanOut112[30] , \nScanOut112[29] , 
        \nScanOut112[28] , \nScanOut112[27] , \nScanOut112[26] , 
        \nScanOut112[25] , \nScanOut112[24] , \nScanOut112[23] , 
        \nScanOut112[22] , \nScanOut112[21] , \nScanOut112[20] , 
        \nScanOut112[19] , \nScanOut112[18] , \nScanOut112[17] , 
        \nScanOut112[16] , \nScanOut112[15] , \nScanOut112[14] , 
        \nScanOut112[13] , \nScanOut112[12] , \nScanOut112[11] , 
        \nScanOut112[10] , \nScanOut112[9] , \nScanOut112[8] , 
        \nScanOut112[7] , \nScanOut112[6] , \nScanOut112[5] , \nScanOut112[4] , 
        \nScanOut112[3] , \nScanOut112[2] , \nScanOut112[1] , \nScanOut112[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_48[31] , \nOut1_48[30] , \nOut1_48[29] , 
        \nOut1_48[28] , \nOut1_48[27] , \nOut1_48[26] , \nOut1_48[25] , 
        \nOut1_48[24] , \nOut1_48[23] , \nOut1_48[22] , \nOut1_48[21] , 
        \nOut1_48[20] , \nOut1_48[19] , \nOut1_48[18] , \nOut1_48[17] , 
        \nOut1_48[16] , \nOut1_48[15] , \nOut1_48[14] , \nOut1_48[13] , 
        \nOut1_48[12] , \nOut1_48[11] , \nOut1_48[10] , \nOut1_48[9] , 
        \nOut1_48[8] , \nOut1_48[7] , \nOut1_48[6] , \nOut1_48[5] , 
        \nOut1_48[4] , \nOut1_48[3] , \nOut1_48[2] , \nOut1_48[1] , 
        \nOut1_48[0] }), .NORTH_EDGE({\nOut1_47[31] , \nOut1_47[30] , 
        \nOut1_47[29] , \nOut1_47[28] , \nOut1_47[27] , \nOut1_47[26] , 
        \nOut1_47[25] , \nOut1_47[24] , \nOut1_47[23] , \nOut1_47[22] , 
        \nOut1_47[21] , \nOut1_47[20] , \nOut1_47[19] , \nOut1_47[18] , 
        \nOut1_47[17] , \nOut1_47[16] , \nOut1_47[15] , \nOut1_47[14] , 
        \nOut1_47[13] , \nOut1_47[12] , \nOut1_47[11] , \nOut1_47[10] , 
        \nOut1_47[9] , \nOut1_47[8] , \nOut1_47[7] , \nOut1_47[6] , 
        \nOut1_47[5] , \nOut1_47[4] , \nOut1_47[3] , \nOut1_47[2] , 
        \nOut1_47[1] , \nOut1_47[0] }), .SOUTH_EDGE({\nOut1_49[31] , 
        \nOut1_49[30] , \nOut1_49[29] , \nOut1_49[28] , \nOut1_49[27] , 
        \nOut1_49[26] , \nOut1_49[25] , \nOut1_49[24] , \nOut1_49[23] , 
        \nOut1_49[22] , \nOut1_49[21] , \nOut1_49[20] , \nOut1_49[19] , 
        \nOut1_49[18] , \nOut1_49[17] , \nOut1_49[16] , \nOut1_49[15] , 
        \nOut1_49[14] , \nOut1_49[13] , \nOut1_49[12] , \nOut1_49[11] , 
        \nOut1_49[10] , \nOut1_49[9] , \nOut1_49[8] , \nOut1_49[7] , 
        \nOut1_49[6] , \nOut1_49[5] , \nOut1_49[4] , \nOut1_49[3] , 
        \nOut1_49[2] , \nOut1_49[1] , \nOut1_49[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_48[0] ), .NW_EDGE(\nOut0_47[0] ), .SW_EDGE(
        \nOut0_49[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Control_WIDTH32_CWIDTH7_IDWIDTH1_SCAN1 U_Life_Control ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut0[31] , \nScanOut0[30] , 
        \nScanOut0[29] , \nScanOut0[28] , \nScanOut0[27] , \nScanOut0[26] , 
        \nScanOut0[25] , \nScanOut0[24] , \nScanOut0[23] , \nScanOut0[22] , 
        \nScanOut0[21] , \nScanOut0[20] , \nScanOut0[19] , \nScanOut0[18] , 
        \nScanOut0[17] , \nScanOut0[16] , \nScanOut0[15] , \nScanOut0[14] , 
        \nScanOut0[13] , \nScanOut0[12] , \nScanOut0[11] , \nScanOut0[10] , 
        \nScanOut0[9] , \nScanOut0[8] , \nScanOut0[7] , \nScanOut0[6] , 
        \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , \nScanOut0[2] , 
        \nScanOut0[1] , \nScanOut0[0] }), .ScanOut({\nScanOut128[31] , 
        \nScanOut128[30] , \nScanOut128[29] , \nScanOut128[28] , 
        \nScanOut128[27] , \nScanOut128[26] , \nScanOut128[25] , 
        \nScanOut128[24] , \nScanOut128[23] , \nScanOut128[22] , 
        \nScanOut128[21] , \nScanOut128[20] , \nScanOut128[19] , 
        \nScanOut128[18] , \nScanOut128[17] , \nScanOut128[16] , 
        \nScanOut128[15] , \nScanOut128[14] , \nScanOut128[13] , 
        \nScanOut128[12] , \nScanOut128[11] , \nScanOut128[10] , 
        \nScanOut128[9] , \nScanOut128[8] , \nScanOut128[7] , \nScanOut128[6] , 
        \nScanOut128[5] , \nScanOut128[4] , \nScanOut128[3] , \nScanOut128[2] , 
        \nScanOut128[1] , \nScanOut128[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b1), .ScanId(1'b0), .Enable(\nEnable[0] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_16 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut17[31] , \nScanOut17[30] , \nScanOut17[29] , 
        \nScanOut17[28] , \nScanOut17[27] , \nScanOut17[26] , \nScanOut17[25] , 
        \nScanOut17[24] , \nScanOut17[23] , \nScanOut17[22] , \nScanOut17[21] , 
        \nScanOut17[20] , \nScanOut17[19] , \nScanOut17[18] , \nScanOut17[17] , 
        \nScanOut17[16] , \nScanOut17[15] , \nScanOut17[14] , \nScanOut17[13] , 
        \nScanOut17[12] , \nScanOut17[11] , \nScanOut17[10] , \nScanOut17[9] , 
        \nScanOut17[8] , \nScanOut17[7] , \nScanOut17[6] , \nScanOut17[5] , 
        \nScanOut17[4] , \nScanOut17[3] , \nScanOut17[2] , \nScanOut17[1] , 
        \nScanOut17[0] }), .ScanOut({\nScanOut16[31] , \nScanOut16[30] , 
        \nScanOut16[29] , \nScanOut16[28] , \nScanOut16[27] , \nScanOut16[26] , 
        \nScanOut16[25] , \nScanOut16[24] , \nScanOut16[23] , \nScanOut16[22] , 
        \nScanOut16[21] , \nScanOut16[20] , \nScanOut16[19] , \nScanOut16[18] , 
        \nScanOut16[17] , \nScanOut16[16] , \nScanOut16[15] , \nScanOut16[14] , 
        \nScanOut16[13] , \nScanOut16[12] , \nScanOut16[11] , \nScanOut16[10] , 
        \nScanOut16[9] , \nScanOut16[8] , \nScanOut16[7] , \nScanOut16[6] , 
        \nScanOut16[5] , \nScanOut16[4] , \nScanOut16[3] , \nScanOut16[2] , 
        \nScanOut16[1] , \nScanOut16[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_16[31] , 
        \nOut0_16[30] , \nOut0_16[29] , \nOut0_16[28] , \nOut0_16[27] , 
        \nOut0_16[26] , \nOut0_16[25] , \nOut0_16[24] , \nOut0_16[23] , 
        \nOut0_16[22] , \nOut0_16[21] , \nOut0_16[20] , \nOut0_16[19] , 
        \nOut0_16[18] , \nOut0_16[17] , \nOut0_16[16] , \nOut0_16[15] , 
        \nOut0_16[14] , \nOut0_16[13] , \nOut0_16[12] , \nOut0_16[11] , 
        \nOut0_16[10] , \nOut0_16[9] , \nOut0_16[8] , \nOut0_16[7] , 
        \nOut0_16[6] , \nOut0_16[5] , \nOut0_16[4] , \nOut0_16[3] , 
        \nOut0_16[2] , \nOut0_16[1] , \nOut0_16[0] }), .NORTH_EDGE({
        \nOut0_15[31] , \nOut0_15[30] , \nOut0_15[29] , \nOut0_15[28] , 
        \nOut0_15[27] , \nOut0_15[26] , \nOut0_15[25] , \nOut0_15[24] , 
        \nOut0_15[23] , \nOut0_15[22] , \nOut0_15[21] , \nOut0_15[20] , 
        \nOut0_15[19] , \nOut0_15[18] , \nOut0_15[17] , \nOut0_15[16] , 
        \nOut0_15[15] , \nOut0_15[14] , \nOut0_15[13] , \nOut0_15[12] , 
        \nOut0_15[11] , \nOut0_15[10] , \nOut0_15[9] , \nOut0_15[8] , 
        \nOut0_15[7] , \nOut0_15[6] , \nOut0_15[5] , \nOut0_15[4] , 
        \nOut0_15[3] , \nOut0_15[2] , \nOut0_15[1] , \nOut0_15[0] }), 
        .SOUTH_EDGE({\nOut0_17[31] , \nOut0_17[30] , \nOut0_17[29] , 
        \nOut0_17[28] , \nOut0_17[27] , \nOut0_17[26] , \nOut0_17[25] , 
        \nOut0_17[24] , \nOut0_17[23] , \nOut0_17[22] , \nOut0_17[21] , 
        \nOut0_17[20] , \nOut0_17[19] , \nOut0_17[18] , \nOut0_17[17] , 
        \nOut0_17[16] , \nOut0_17[15] , \nOut0_17[14] , \nOut0_17[13] , 
        \nOut0_17[12] , \nOut0_17[11] , \nOut0_17[10] , \nOut0_17[9] , 
        \nOut0_17[8] , \nOut0_17[7] , \nOut0_17[6] , \nOut0_17[5] , 
        \nOut0_17[4] , \nOut0_17[3] , \nOut0_17[2] , \nOut0_17[1] , 
        \nOut0_17[0] }), .EAST_EDGE(\nOut1_16[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_15[31] ), .SE_EDGE(
        \nOut1_17[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_78 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut79[31] , \nScanOut79[30] , \nScanOut79[29] , 
        \nScanOut79[28] , \nScanOut79[27] , \nScanOut79[26] , \nScanOut79[25] , 
        \nScanOut79[24] , \nScanOut79[23] , \nScanOut79[22] , \nScanOut79[21] , 
        \nScanOut79[20] , \nScanOut79[19] , \nScanOut79[18] , \nScanOut79[17] , 
        \nScanOut79[16] , \nScanOut79[15] , \nScanOut79[14] , \nScanOut79[13] , 
        \nScanOut79[12] , \nScanOut79[11] , \nScanOut79[10] , \nScanOut79[9] , 
        \nScanOut79[8] , \nScanOut79[7] , \nScanOut79[6] , \nScanOut79[5] , 
        \nScanOut79[4] , \nScanOut79[3] , \nScanOut79[2] , \nScanOut79[1] , 
        \nScanOut79[0] }), .ScanOut({\nScanOut78[31] , \nScanOut78[30] , 
        \nScanOut78[29] , \nScanOut78[28] , \nScanOut78[27] , \nScanOut78[26] , 
        \nScanOut78[25] , \nScanOut78[24] , \nScanOut78[23] , \nScanOut78[22] , 
        \nScanOut78[21] , \nScanOut78[20] , \nScanOut78[19] , \nScanOut78[18] , 
        \nScanOut78[17] , \nScanOut78[16] , \nScanOut78[15] , \nScanOut78[14] , 
        \nScanOut78[13] , \nScanOut78[12] , \nScanOut78[11] , \nScanOut78[10] , 
        \nScanOut78[9] , \nScanOut78[8] , \nScanOut78[7] , \nScanOut78[6] , 
        \nScanOut78[5] , \nScanOut78[4] , \nScanOut78[3] , \nScanOut78[2] , 
        \nScanOut78[1] , \nScanOut78[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_14[31] , 
        \nOut1_14[30] , \nOut1_14[29] , \nOut1_14[28] , \nOut1_14[27] , 
        \nOut1_14[26] , \nOut1_14[25] , \nOut1_14[24] , \nOut1_14[23] , 
        \nOut1_14[22] , \nOut1_14[21] , \nOut1_14[20] , \nOut1_14[19] , 
        \nOut1_14[18] , \nOut1_14[17] , \nOut1_14[16] , \nOut1_14[15] , 
        \nOut1_14[14] , \nOut1_14[13] , \nOut1_14[12] , \nOut1_14[11] , 
        \nOut1_14[10] , \nOut1_14[9] , \nOut1_14[8] , \nOut1_14[7] , 
        \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , \nOut1_14[3] , 
        \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), .NORTH_EDGE({
        \nOut1_13[31] , \nOut1_13[30] , \nOut1_13[29] , \nOut1_13[28] , 
        \nOut1_13[27] , \nOut1_13[26] , \nOut1_13[25] , \nOut1_13[24] , 
        \nOut1_13[23] , \nOut1_13[22] , \nOut1_13[21] , \nOut1_13[20] , 
        \nOut1_13[19] , \nOut1_13[18] , \nOut1_13[17] , \nOut1_13[16] , 
        \nOut1_13[15] , \nOut1_13[14] , \nOut1_13[13] , \nOut1_13[12] , 
        \nOut1_13[11] , \nOut1_13[10] , \nOut1_13[9] , \nOut1_13[8] , 
        \nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), 
        .SOUTH_EDGE({\nOut1_15[31] , \nOut1_15[30] , \nOut1_15[29] , 
        \nOut1_15[28] , \nOut1_15[27] , \nOut1_15[26] , \nOut1_15[25] , 
        \nOut1_15[24] , \nOut1_15[23] , \nOut1_15[22] , \nOut1_15[21] , 
        \nOut1_15[20] , \nOut1_15[19] , \nOut1_15[18] , \nOut1_15[17] , 
        \nOut1_15[16] , \nOut1_15[15] , \nOut1_15[14] , \nOut1_15[13] , 
        \nOut1_15[12] , \nOut1_15[11] , \nOut1_15[10] , \nOut1_15[9] , 
        \nOut1_15[8] , \nOut1_15[7] , \nOut1_15[6] , \nOut1_15[5] , 
        \nOut1_15[4] , \nOut1_15[3] , \nOut1_15[2] , \nOut1_15[1] , 
        \nOut1_15[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut0_14[0] ), 
        .NW_EDGE(\nOut0_13[0] ), .SW_EDGE(\nOut0_15[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_109 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut110[31] , \nScanOut110[30] , \nScanOut110[29] , 
        \nScanOut110[28] , \nScanOut110[27] , \nScanOut110[26] , 
        \nScanOut110[25] , \nScanOut110[24] , \nScanOut110[23] , 
        \nScanOut110[22] , \nScanOut110[21] , \nScanOut110[20] , 
        \nScanOut110[19] , \nScanOut110[18] , \nScanOut110[17] , 
        \nScanOut110[16] , \nScanOut110[15] , \nScanOut110[14] , 
        \nScanOut110[13] , \nScanOut110[12] , \nScanOut110[11] , 
        \nScanOut110[10] , \nScanOut110[9] , \nScanOut110[8] , 
        \nScanOut110[7] , \nScanOut110[6] , \nScanOut110[5] , \nScanOut110[4] , 
        \nScanOut110[3] , \nScanOut110[2] , \nScanOut110[1] , \nScanOut110[0] 
        }), .ScanOut({\nScanOut109[31] , \nScanOut109[30] , \nScanOut109[29] , 
        \nScanOut109[28] , \nScanOut109[27] , \nScanOut109[26] , 
        \nScanOut109[25] , \nScanOut109[24] , \nScanOut109[23] , 
        \nScanOut109[22] , \nScanOut109[21] , \nScanOut109[20] , 
        \nScanOut109[19] , \nScanOut109[18] , \nScanOut109[17] , 
        \nScanOut109[16] , \nScanOut109[15] , \nScanOut109[14] , 
        \nScanOut109[13] , \nScanOut109[12] , \nScanOut109[11] , 
        \nScanOut109[10] , \nScanOut109[9] , \nScanOut109[8] , 
        \nScanOut109[7] , \nScanOut109[6] , \nScanOut109[5] , \nScanOut109[4] , 
        \nScanOut109[3] , \nScanOut109[2] , \nScanOut109[1] , \nScanOut109[0] 
        }), .ScanEnable(\nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), 
        .BLOCK_VALUE({\nOut1_45[31] , \nOut1_45[30] , \nOut1_45[29] , 
        \nOut1_45[28] , \nOut1_45[27] , \nOut1_45[26] , \nOut1_45[25] , 
        \nOut1_45[24] , \nOut1_45[23] , \nOut1_45[22] , \nOut1_45[21] , 
        \nOut1_45[20] , \nOut1_45[19] , \nOut1_45[18] , \nOut1_45[17] , 
        \nOut1_45[16] , \nOut1_45[15] , \nOut1_45[14] , \nOut1_45[13] , 
        \nOut1_45[12] , \nOut1_45[11] , \nOut1_45[10] , \nOut1_45[9] , 
        \nOut1_45[8] , \nOut1_45[7] , \nOut1_45[6] , \nOut1_45[5] , 
        \nOut1_45[4] , \nOut1_45[3] , \nOut1_45[2] , \nOut1_45[1] , 
        \nOut1_45[0] }), .NORTH_EDGE({\nOut1_44[31] , \nOut1_44[30] , 
        \nOut1_44[29] , \nOut1_44[28] , \nOut1_44[27] , \nOut1_44[26] , 
        \nOut1_44[25] , \nOut1_44[24] , \nOut1_44[23] , \nOut1_44[22] , 
        \nOut1_44[21] , \nOut1_44[20] , \nOut1_44[19] , \nOut1_44[18] , 
        \nOut1_44[17] , \nOut1_44[16] , \nOut1_44[15] , \nOut1_44[14] , 
        \nOut1_44[13] , \nOut1_44[12] , \nOut1_44[11] , \nOut1_44[10] , 
        \nOut1_44[9] , \nOut1_44[8] , \nOut1_44[7] , \nOut1_44[6] , 
        \nOut1_44[5] , \nOut1_44[4] , \nOut1_44[3] , \nOut1_44[2] , 
        \nOut1_44[1] , \nOut1_44[0] }), .SOUTH_EDGE({\nOut1_46[31] , 
        \nOut1_46[30] , \nOut1_46[29] , \nOut1_46[28] , \nOut1_46[27] , 
        \nOut1_46[26] , \nOut1_46[25] , \nOut1_46[24] , \nOut1_46[23] , 
        \nOut1_46[22] , \nOut1_46[21] , \nOut1_46[20] , \nOut1_46[19] , 
        \nOut1_46[18] , \nOut1_46[17] , \nOut1_46[16] , \nOut1_46[15] , 
        \nOut1_46[14] , \nOut1_46[13] , \nOut1_46[12] , \nOut1_46[11] , 
        \nOut1_46[10] , \nOut1_46[9] , \nOut1_46[8] , \nOut1_46[7] , 
        \nOut1_46[6] , \nOut1_46[5] , \nOut1_46[4] , \nOut1_46[3] , 
        \nOut1_46[2] , \nOut1_46[1] , \nOut1_46[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut0_45[0] ), .NW_EDGE(\nOut0_44[0] ), .SW_EDGE(
        \nOut0_46[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_31 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut32[31] , \nScanOut32[30] , \nScanOut32[29] , 
        \nScanOut32[28] , \nScanOut32[27] , \nScanOut32[26] , \nScanOut32[25] , 
        \nScanOut32[24] , \nScanOut32[23] , \nScanOut32[22] , \nScanOut32[21] , 
        \nScanOut32[20] , \nScanOut32[19] , \nScanOut32[18] , \nScanOut32[17] , 
        \nScanOut32[16] , \nScanOut32[15] , \nScanOut32[14] , \nScanOut32[13] , 
        \nScanOut32[12] , \nScanOut32[11] , \nScanOut32[10] , \nScanOut32[9] , 
        \nScanOut32[8] , \nScanOut32[7] , \nScanOut32[6] , \nScanOut32[5] , 
        \nScanOut32[4] , \nScanOut32[3] , \nScanOut32[2] , \nScanOut32[1] , 
        \nScanOut32[0] }), .ScanOut({\nScanOut31[31] , \nScanOut31[30] , 
        \nScanOut31[29] , \nScanOut31[28] , \nScanOut31[27] , \nScanOut31[26] , 
        \nScanOut31[25] , \nScanOut31[24] , \nScanOut31[23] , \nScanOut31[22] , 
        \nScanOut31[21] , \nScanOut31[20] , \nScanOut31[19] , \nScanOut31[18] , 
        \nScanOut31[17] , \nScanOut31[16] , \nScanOut31[15] , \nScanOut31[14] , 
        \nScanOut31[13] , \nScanOut31[12] , \nScanOut31[11] , \nScanOut31[10] , 
        \nScanOut31[9] , \nScanOut31[8] , \nScanOut31[7] , \nScanOut31[6] , 
        \nScanOut31[5] , \nScanOut31[4] , \nScanOut31[3] , \nScanOut31[2] , 
        \nScanOut31[1] , \nScanOut31[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_31[31] , 
        \nOut0_31[30] , \nOut0_31[29] , \nOut0_31[28] , \nOut0_31[27] , 
        \nOut0_31[26] , \nOut0_31[25] , \nOut0_31[24] , \nOut0_31[23] , 
        \nOut0_31[22] , \nOut0_31[21] , \nOut0_31[20] , \nOut0_31[19] , 
        \nOut0_31[18] , \nOut0_31[17] , \nOut0_31[16] , \nOut0_31[15] , 
        \nOut0_31[14] , \nOut0_31[13] , \nOut0_31[12] , \nOut0_31[11] , 
        \nOut0_31[10] , \nOut0_31[9] , \nOut0_31[8] , \nOut0_31[7] , 
        \nOut0_31[6] , \nOut0_31[5] , \nOut0_31[4] , \nOut0_31[3] , 
        \nOut0_31[2] , \nOut0_31[1] , \nOut0_31[0] }), .NORTH_EDGE({
        \nOut0_30[31] , \nOut0_30[30] , \nOut0_30[29] , \nOut0_30[28] , 
        \nOut0_30[27] , \nOut0_30[26] , \nOut0_30[25] , \nOut0_30[24] , 
        \nOut0_30[23] , \nOut0_30[22] , \nOut0_30[21] , \nOut0_30[20] , 
        \nOut0_30[19] , \nOut0_30[18] , \nOut0_30[17] , \nOut0_30[16] , 
        \nOut0_30[15] , \nOut0_30[14] , \nOut0_30[13] , \nOut0_30[12] , 
        \nOut0_30[11] , \nOut0_30[10] , \nOut0_30[9] , \nOut0_30[8] , 
        \nOut0_30[7] , \nOut0_30[6] , \nOut0_30[5] , \nOut0_30[4] , 
        \nOut0_30[3] , \nOut0_30[2] , \nOut0_30[1] , \nOut0_30[0] }), 
        .SOUTH_EDGE({\nOut0_32[31] , \nOut0_32[30] , \nOut0_32[29] , 
        \nOut0_32[28] , \nOut0_32[27] , \nOut0_32[26] , \nOut0_32[25] , 
        \nOut0_32[24] , \nOut0_32[23] , \nOut0_32[22] , \nOut0_32[21] , 
        \nOut0_32[20] , \nOut0_32[19] , \nOut0_32[18] , \nOut0_32[17] , 
        \nOut0_32[16] , \nOut0_32[15] , \nOut0_32[14] , \nOut0_32[13] , 
        \nOut0_32[12] , \nOut0_32[11] , \nOut0_32[10] , \nOut0_32[9] , 
        \nOut0_32[8] , \nOut0_32[7] , \nOut0_32[6] , \nOut0_32[5] , 
        \nOut0_32[4] , \nOut0_32[3] , \nOut0_32[2] , \nOut0_32[1] , 
        \nOut0_32[0] }), .EAST_EDGE(\nOut1_31[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_30[31] ), .SE_EDGE(
        \nOut1_32[31] ) );
endmodule

