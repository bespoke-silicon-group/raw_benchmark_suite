
module BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, Out, Enable1, Enable2, In1, In2
     );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] In1;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In2;
input  Clk, Reset, RD, WR, ScanEnable, Enable1, Enable2;
    wire \ScanOut[31] , n288, \ScanOut[5]1 , \ScanOut[4]1 , n245, n287, n262, 
        n279, n217, n230, \ScanOut[10]1 , n302, n222, n305, n257, n270, n295, 
        n239, n292, \ScanOut[23]1 , \ScanOut[8]1 , n219, n225, n250, n277, 
        n289, n237, n259, \ScanOut[22]1 , \ScanOut[11]1 , n265, n242, 
        \ScanOut[9]1 , n310, n280, n224, n276, n303, n251, n293, 
        \ScanOut[19]1 , n218, n311, n281, \ScanOut[26]1 , \ScanOut[18]1 , 
        \ScanOut[1]1 , n264, \ScanOut[0]1 , n243, n258, \ScanOut[15]1 , n236, 
        n216, n231, n278, \ScanOut[27]1 , n244, \ScanOut[14]1 , n263, n316, 
        n286, n304, n294, n271, n238, n256, n223, n233, n228, n314, n284, n214, 
        n246, n261, \ScanOut[28]1 , n221, \ScanOut[3]1 , n268, \ScanOut[30]1 , 
        \ScanOut[29]1 , \ScanOut[2]1 , n254, n273, n306, n296, n301, n291, 
        \ScanOut[25]1 , \ScanOut[24]1 , \ScanOut[17]1 , n253, n248, n274, 
        \ScanOut[16]1 , n226, n234, n308, n298, n241, n313, n266, n283, 
        \ScanOut[6]1 , n227, n249, \ScanOut[7]1 , n312, n300, n252, n290, n275, 
        n282, n215, n309, n235, n240, n267, n299, \ScanOut[13]1 , n232, n247, 
        n260, \ScanOut[21]1 , n315, n285, n229, n307, n297, \ScanOut[12]1 , 
        n272, n255, n269, \ScanOut[20]1 , n220;
    assign ScanOut[31] = \ScanOut[31] ;
    assign ScanOut[30] = \ScanOut[30]1 ;
    assign ScanOut[29] = \ScanOut[29]1 ;
    assign ScanOut[28] = \ScanOut[28]1 ;
    assign ScanOut[27] = \ScanOut[27]1 ;
    assign ScanOut[26] = \ScanOut[26]1 ;
    assign ScanOut[25] = \ScanOut[25]1 ;
    assign ScanOut[24] = \ScanOut[24]1 ;
    assign ScanOut[23] = \ScanOut[23]1 ;
    assign ScanOut[22] = \ScanOut[22]1 ;
    assign ScanOut[21] = \ScanOut[21]1 ;
    assign ScanOut[20] = \ScanOut[20]1 ;
    assign ScanOut[19] = \ScanOut[19]1 ;
    assign ScanOut[18] = \ScanOut[18]1 ;
    assign ScanOut[17] = \ScanOut[17]1 ;
    assign ScanOut[16] = \ScanOut[16]1 ;
    assign ScanOut[15] = \ScanOut[15]1 ;
    assign ScanOut[14] = \ScanOut[14]1 ;
    assign ScanOut[13] = \ScanOut[13]1 ;
    assign ScanOut[12] = \ScanOut[12]1 ;
    assign ScanOut[11] = \ScanOut[11]1 ;
    assign ScanOut[10] = \ScanOut[10]1 ;
    assign ScanOut[9] = \ScanOut[9]1 ;
    assign ScanOut[8] = \ScanOut[8]1 ;
    assign ScanOut[7] = \ScanOut[7]1 ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[31] = \ScanOut[31] ;
    assign Out[30] = \ScanOut[30]1 ;
    assign Out[29] = \ScanOut[29]1 ;
    assign Out[28] = \ScanOut[28]1 ;
    assign Out[27] = \ScanOut[27]1 ;
    assign Out[26] = \ScanOut[26]1 ;
    assign Out[25] = \ScanOut[25]1 ;
    assign Out[24] = \ScanOut[24]1 ;
    assign Out[23] = \ScanOut[23]1 ;
    assign Out[22] = \ScanOut[22]1 ;
    assign Out[21] = \ScanOut[21]1 ;
    assign Out[20] = \ScanOut[20]1 ;
    assign Out[19] = \ScanOut[19]1 ;
    assign Out[18] = \ScanOut[18]1 ;
    assign Out[17] = \ScanOut[17]1 ;
    assign Out[16] = \ScanOut[16]1 ;
    assign Out[15] = \ScanOut[15]1 ;
    assign Out[14] = \ScanOut[14]1 ;
    assign Out[13] = \ScanOut[13]1 ;
    assign Out[12] = \ScanOut[12]1 ;
    assign Out[11] = \ScanOut[11]1 ;
    assign Out[10] = \ScanOut[10]1 ;
    assign Out[9] = \ScanOut[9]1 ;
    assign Out[8] = \ScanOut[8]1 ;
    assign Out[7] = \ScanOut[7]1 ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_OR2 U54 ( .A(n258), .B(n259), .Z(n294) );
    VMW_AO22 U73 ( .A(In1[7]), .B(n281), .C(In2[7]), .D(n280), .Z(n228) );
    VMW_AO22 U113 ( .A(In1[18]), .B(n281), .C(In2[18]), .D(n280), .Z(n250) );
    VMW_INV U134 ( .A(Enable1), .Z(n282) );
    VMW_NOR4 U68 ( .A(Enable1), .B(Enable2), .C(ScanEnable), .D(Reset), .Z(
        n279) );
    VMW_AO22 U96 ( .A(\ScanOut[26]1 ), .B(n279), .C(ScanIn[26]), .D(n283), .Z(
        n267) );
    VMW_AO22 U108 ( .A(\ScanOut[20]1 ), .B(n279), .C(ScanIn[20]), .D(n283), 
        .Z(n255) );
    VMW_OR2 U33 ( .A(n216), .B(n217), .Z(n315) );
    VMW_OR2 U34 ( .A(n218), .B(n219), .Z(n314) );
    VMW_OR2 U41 ( .A(n232), .B(n233), .Z(n307) );
    VMW_OR2 U46 ( .A(n242), .B(n243), .Z(n302) );
    VMW_OR2 U61 ( .A(n272), .B(n273), .Z(n287) );
    VMW_AO22 U84 ( .A(\ScanOut[31] ), .B(n279), .C(ScanIn[31]), .D(n283), .Z(
        n277) );
    VMW_AO22 U101 ( .A(In1[23]), .B(n281), .C(In2[23]), .D(n280), .Z(n260) );
    VMW_AO22 U126 ( .A(\ScanOut[12]1 ), .B(n279), .C(ScanIn[12]), .D(n283), 
        .Z(n239) );
    VMW_NOR2 U66 ( .A(n278), .B(n282), .Z(n281) );
    VMW_AO22 U106 ( .A(\ScanOut[21]1 ), .B(n279), .C(ScanIn[21]), .D(n283), 
        .Z(n257) );
    VMW_AO22 U121 ( .A(In1[14]), .B(n281), .C(In2[14]), .D(n280), .Z(n242) );
    VMW_AO22 U83 ( .A(In1[31]), .B(n281), .C(In2[31]), .D(n280), .Z(n276) );
    VMW_AO22 U98 ( .A(\ScanOut[25]1 ), .B(n279), .C(ScanIn[25]), .D(n283), .Z(
        n265) );
    VMW_OR2 U35 ( .A(n220), .B(n221), .Z(n313) );
    VMW_OR2 U48 ( .A(n246), .B(n247), .Z(n300) );
    VMW_AO22 U128 ( .A(\ScanOut[11]1 ), .B(n279), .C(ScanIn[11]), .D(n283), 
        .Z(n237) );
    VMW_OR2 U53 ( .A(n256), .B(n257), .Z(n295) );
    VMW_AO22 U91 ( .A(In1[28]), .B(n281), .C(In2[28]), .D(n280), .Z(n270) );
    VMW_AO22 U74 ( .A(\ScanOut[7]1 ), .B(n279), .C(ScanIn[7]), .D(n283), .Z(
        n229) );
    VMW_AO22 U114 ( .A(\ScanOut[18]1 ), .B(n279), .C(ScanIn[18]), .D(n283), 
        .Z(n251) );
    VMW_INV U133 ( .A(ScanEnable), .Z(n284) );
    VMW_AO22 U99 ( .A(In1[24]), .B(n281), .C(In2[24]), .D(n280), .Z(n262) );
    VMW_FD \Out_reg[25]  ( .D(n291), .CP(Clk), .Q(\ScanOut[25]1 ) );
    VMW_FD \Out_reg[16]  ( .D(n300), .CP(Clk), .Q(\ScanOut[16]1 ) );
    VMW_OR2 U32 ( .A(n214), .B(n215), .Z(n316) );
    VMW_OR2 U40 ( .A(n230), .B(n231), .Z(n308) );
    VMW_AO22 U82 ( .A(\ScanOut[3]1 ), .B(n279), .C(ScanIn[3]), .D(n283), .Z(
        n221) );
    VMW_FD \Out_reg[5]  ( .D(n311), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_OR2 U47 ( .A(n244), .B(n245), .Z(n301) );
    VMW_OR2 U49 ( .A(n248), .B(n249), .Z(n299) );
    VMW_OR2 U52 ( .A(n254), .B(n255), .Z(n296) );
    VMW_NOR2 U67 ( .A(n284), .B(Reset), .Z(n283) );
    VMW_AO22 U107 ( .A(In1[20]), .B(n281), .C(In2[20]), .D(n280), .Z(n254) );
    VMW_AO22 U120 ( .A(\ScanOut[15]1 ), .B(n279), .C(ScanIn[15]), .D(n283), 
        .Z(n245) );
    VMW_AO22 U75 ( .A(In1[6]), .B(n281), .C(In2[6]), .D(n280), .Z(n226) );
    VMW_AO22 U115 ( .A(In1[17]), .B(n281), .C(In2[17]), .D(n280), .Z(n248) );
    VMW_AO22 U132 ( .A(\ScanOut[0]1 ), .B(n279), .C(ScanIn[0]), .D(n283), .Z(
        n215) );
    VMW_FD \Out_reg[12]  ( .D(n304), .CP(Clk), .Q(\ScanOut[12]1 ) );
    VMW_AO22 U90 ( .A(\ScanOut[29]1 ), .B(n279), .C(ScanIn[29]), .D(n283), .Z(
        n273) );
    VMW_FD \Out_reg[21]  ( .D(n295), .CP(Clk), .Q(\ScanOut[21]1 ) );
    VMW_AO22 U129 ( .A(In1[10]), .B(n281), .C(In2[10]), .D(n280), .Z(n234) );
    VMW_FD \Out_reg[31]  ( .D(n285), .CP(Clk), .Q(\ScanOut[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n288), .CP(Clk), .Q(\ScanOut[28]1 ) );
    VMW_FD \Out_reg[8]  ( .D(n308), .CP(Clk), .Q(\ScanOut[8]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n315), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_OR2 U55 ( .A(n260), .B(n261), .Z(n293) );
    VMW_AO22 U69 ( .A(In1[9]), .B(n281), .C(In2[9]), .D(n280), .Z(n232) );
    VMW_AO22 U109 ( .A(In1[1]), .B(n281), .C(In2[1]), .D(n280), .Z(n216) );
    VMW_FD \Out_reg[19]  ( .D(n297), .CP(Clk), .Q(\ScanOut[19]1 ) );
    VMW_AO22 U72 ( .A(\ScanOut[8]1 ), .B(n279), .C(ScanIn[8]), .D(n283), .Z(
        n231) );
    VMW_AO22 U97 ( .A(In1[25]), .B(n281), .C(In2[25]), .D(n280), .Z(n264) );
    VMW_FD \Out_reg[3]  ( .D(n313), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_AO22 U112 ( .A(\ScanOut[19]1 ), .B(n279), .C(ScanIn[19]), .D(n283), 
        .Z(n253) );
    VMW_FD \Out_reg[23]  ( .D(n293), .CP(Clk), .Q(\ScanOut[23]1 ) );
    VMW_FD \Out_reg[10]  ( .D(n306), .CP(Clk), .Q(\ScanOut[10]1 ) );
    VMW_OR2 U60 ( .A(n270), .B(n271), .Z(n288) );
    VMW_FD \Out_reg[7]  ( .D(n309), .CP(Clk), .Q(\ScanOut[7]1 ) );
    VMW_AO22 U100 ( .A(\ScanOut[24]1 ), .B(n279), .C(ScanIn[24]), .D(n283), 
        .Z(n263) );
    VMW_AO22 U127 ( .A(In1[11]), .B(n281), .C(In2[11]), .D(n280), .Z(n236) );
    VMW_AO22 U85 ( .A(In1[30]), .B(n281), .C(In2[30]), .D(n280), .Z(n274) );
    VMW_FD \Out_reg[27]  ( .D(n289), .CP(Clk), .Q(\ScanOut[27]1 ) );
    VMW_FD \Out_reg[14]  ( .D(n302), .CP(Clk), .Q(\ScanOut[14]1 ) );
    VMW_OR2 U36 ( .A(n222), .B(n223), .Z(n312) );
    VMW_OR2 U37 ( .A(n224), .B(n225), .Z(n311) );
    VMW_OR2 U39 ( .A(n228), .B(n229), .Z(n309) );
    VMW_OR2 U57 ( .A(n264), .B(n265), .Z(n291) );
    VMW_FD \Out_reg[6]  ( .D(n310), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U70 ( .A(\ScanOut[9]1 ), .B(n279), .C(ScanIn[9]), .D(n283), .Z(
        n233) );
    VMW_AO22 U110 ( .A(\ScanOut[1]1 ), .B(n279), .C(ScanIn[1]), .D(n283), .Z(
        n217) );
    VMW_OR2 U42 ( .A(n234), .B(n235), .Z(n306) );
    VMW_OR2 U45 ( .A(n240), .B(n241), .Z(n303) );
    VMW_AO22 U79 ( .A(In1[4]), .B(n281), .C(In2[4]), .D(n280), .Z(n222) );
    VMW_AO22 U95 ( .A(In1[26]), .B(n281), .C(In2[26]), .D(n280), .Z(n266) );
    VMW_AO22 U119 ( .A(In1[15]), .B(n281), .C(In2[15]), .D(n280), .Z(n244) );
    VMW_FD \Out_reg[26]  ( .D(n290), .CP(Clk), .Q(\ScanOut[26]1 ) );
    VMW_FD \Out_reg[15]  ( .D(n301), .CP(Clk), .Q(\ScanOut[15]1 ) );
    VMW_FD \Out_reg[18]  ( .D(n298), .CP(Clk), .Q(\ScanOut[18]1 ) );
    VMW_AO22 U87 ( .A(In1[2]), .B(n281), .C(In2[2]), .D(n280), .Z(n218) );
    VMW_FD \Out_reg[2]  ( .D(n314), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_AO22 U125 ( .A(In1[12]), .B(n281), .C(In2[12]), .D(n280), .Z(n238) );
    VMW_FD \Out_reg[11]  ( .D(n305), .CP(Clk), .Q(\ScanOut[11]1 ) );
    VMW_OR2 U62 ( .A(n274), .B(n275), .Z(n286) );
    VMW_FD \Out_reg[22]  ( .D(n294), .CP(Clk), .Q(\ScanOut[22]1 ) );
    VMW_NOR2 U65 ( .A(Enable1), .B(n278), .Z(n280) );
    VMW_AO22 U102 ( .A(\ScanOut[23]1 ), .B(n279), .C(ScanIn[23]), .D(n283), 
        .Z(n261) );
    VMW_AO22 U105 ( .A(In1[21]), .B(n281), .C(In2[21]), .D(n280), .Z(n256) );
    VMW_FD \Out_reg[20]  ( .D(n296), .CP(Clk), .Q(\ScanOut[20]1 ) );
    VMW_FD \Out_reg[13]  ( .D(n303), .CP(Clk), .Q(\ScanOut[13]1 ) );
    VMW_AO22 U80 ( .A(\ScanOut[4]1 ), .B(n279), .C(ScanIn[4]), .D(n283), .Z(
        n223) );
    VMW_AO22 U122 ( .A(\ScanOut[14]1 ), .B(n279), .C(ScanIn[14]), .D(n283), 
        .Z(n243) );
    VMW_FD \Out_reg[9]  ( .D(n307), .CP(Clk), .Q(\ScanOut[9]1 ) );
    VMW_OR2 U50 ( .A(n250), .B(n251), .Z(n298) );
    VMW_OR2 U59 ( .A(n268), .B(n269), .Z(n289) );
    VMW_FD \Out_reg[30]  ( .D(n286), .CP(Clk), .Q(\ScanOut[30]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n316), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_FD \Out_reg[29]  ( .D(n287), .CP(Clk), .Q(\ScanOut[29]1 ) );
    VMW_AO22 U77 ( .A(In1[5]), .B(n281), .C(In2[5]), .D(n280), .Z(n224) );
    VMW_AO22 U89 ( .A(In1[29]), .B(n281), .C(In2[29]), .D(n280), .Z(n272) );
    VMW_AO22 U92 ( .A(\ScanOut[28]1 ), .B(n279), .C(ScanIn[28]), .D(n283), .Z(
        n271) );
    VMW_FD \Out_reg[24]  ( .D(n292), .CP(Clk), .Q(\ScanOut[24]1 ) );
    VMW_FD \Out_reg[17]  ( .D(n299), .CP(Clk), .Q(\ScanOut[17]1 ) );
    VMW_AO22 U117 ( .A(In1[16]), .B(n281), .C(In2[16]), .D(n280), .Z(n246) );
    VMW_FD \Out_reg[4]  ( .D(n312), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_OR2 U58 ( .A(n266), .B(n267), .Z(n290) );
    VMW_AO22 U130 ( .A(\ScanOut[10]1 ), .B(n279), .C(ScanIn[10]), .D(n283), 
        .Z(n235) );
    VMW_OR2 U38 ( .A(n226), .B(n227), .Z(n310) );
    VMW_OR2 U43 ( .A(n236), .B(n237), .Z(n305) );
    VMW_OR3 U64 ( .A(Reset), .B(ScanEnable), .C(n279), .Z(n278) );
    VMW_AO22 U81 ( .A(In1[3]), .B(n281), .C(In2[3]), .D(n280), .Z(n220) );
    VMW_AO22 U104 ( .A(\ScanOut[22]1 ), .B(n279), .C(ScanIn[22]), .D(n283), 
        .Z(n259) );
    VMW_OR2 U51 ( .A(n252), .B(n253), .Z(n297) );
    VMW_AO22 U76 ( .A(\ScanOut[6]1 ), .B(n279), .C(ScanIn[6]), .D(n283), .Z(
        n227) );
    VMW_AO22 U116 ( .A(\ScanOut[17]1 ), .B(n279), .C(ScanIn[17]), .D(n283), 
        .Z(n249) );
    VMW_AO22 U123 ( .A(In1[13]), .B(n281), .C(In2[13]), .D(n280), .Z(n240) );
    VMW_AO22 U88 ( .A(\ScanOut[2]1 ), .B(n279), .C(ScanIn[2]), .D(n283), .Z(
        n219) );
    VMW_AO22 U93 ( .A(In1[27]), .B(n281), .C(In2[27]), .D(n280), .Z(n268) );
    VMW_AO22 U131 ( .A(In1[0]), .B(n281), .C(In2[0]), .D(n280), .Z(n214) );
    VMW_OR2 U44 ( .A(n238), .B(n239), .Z(n304) );
    VMW_OR2 U56 ( .A(n262), .B(n263), .Z(n292) );
    VMW_AO22 U94 ( .A(\ScanOut[27]1 ), .B(n279), .C(ScanIn[27]), .D(n283), .Z(
        n269) );
    VMW_AO22 U71 ( .A(In1[8]), .B(n281), .C(In2[8]), .D(n280), .Z(n230) );
    VMW_AO22 U111 ( .A(In1[19]), .B(n281), .C(In2[19]), .D(n280), .Z(n252) );
    VMW_AO22 U124 ( .A(\ScanOut[13]1 ), .B(n279), .C(ScanIn[13]), .D(n283), 
        .Z(n241) );
    VMW_OR2 U63 ( .A(n276), .B(n277), .Z(n285) );
    VMW_AO22 U78 ( .A(\ScanOut[5]1 ), .B(n279), .C(ScanIn[5]), .D(n283), .Z(
        n225) );
    VMW_AO22 U86 ( .A(\ScanOut[30]1 ), .B(n279), .C(ScanIn[30]), .D(n283), .Z(
        n275) );
    VMW_AO22 U103 ( .A(In1[22]), .B(n281), .C(In2[22]), .D(n280), .Z(n258) );
    VMW_AO22 U118 ( .A(\ScanOut[16]1 ), .B(n279), .C(ScanIn[16]), .D(n283), 
        .Z(n247) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_3 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n112, n32, n29, n85, n47, n60, n109, 
        n40, n67, n82, n99, n27, n35, n49, n115, n107, n52, n75, n114, n34, 
        n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, n21, n46, n54, 
        n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, n113, n118, n94, 
        n23, n103, n16, n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, n58, 
        n116, n104, n18, n24, n88, n37, n51, n93, n59, n76, n117, n80, n42, 
        n65, n19, n50, n77, n89, n25, n102, n105, n22, n39, n95, n45, n57, n70, 
        n62, n87, n17, n30, n79, n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_OR2 U54 ( .A(B[26]), .B(n99), .Z(n103) );
    VMW_INV U73 ( .A(B[27]), .Z(n109) );
    VMW_INV U96 ( .A(B[31]), .Z(n15) );
    VMW_INV U68 ( .A(A[30]), .Z(n117) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n66), .C(n62), .D(n57), .Z(n65) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U34 ( .A(B[16]), .B(n64), .Z(n67) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n75), .D(n70), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_NAND2 U61 ( .A(n114), .B(A[29]), .Z(n115) );
    VMW_INV U84 ( .A(B[15]), .Z(n66) );
    VMW_INV U101 ( .A(A[6]), .Z(n32) );
    VMW_INV U66 ( .A(B[7]), .Z(n41) );
    VMW_INV U83 ( .A(A[15]), .Z(n69) );
    VMW_INV U98 ( .A(B[13]), .Z(n60) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_NAND2 U48 ( .A(n91), .B(B[24]), .Z(n89) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n69), .C(n67), .D(n65), .Z(n68) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n102), .C(n96), .D(n89), .Z(n101) );
    VMW_INV U91 ( .A(B[11]), .Z(n54) );
    VMW_INV U74 ( .A(A[3]), .Z(n30) );
    VMW_INV U99 ( .A(A[26]), .Z(n99) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U40 ( .A(n78), .B(B[20]), .Z(n77) );
    VMW_INV U82 ( .A(B[29]), .Z(n114) );
    VMW_NAND2 U52 ( .A(n99), .B(B[26]), .Z(n97) );
    VMW_INV U67 ( .A(A[7]), .Z(n44) );
    VMW_INV U75 ( .A(B[3]), .Z(n27) );
    VMW_INV U90 ( .A(A[14]), .Z(n58) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n94), .C(n88), .D(n83), .Z(n93) );
    VMW_INV U69 ( .A(B[17]), .Z(n73) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n105), .C(n103), .D(n101), .Z(n104) );
    VMW_INV U72 ( .A(A[27]), .Z(n112) );
    VMW_INV U97 ( .A(A[16]), .Z(n64) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n114), .C(n111), .D(n106), .Z(n113) );
    VMW_INV U100 ( .A(B[23]), .Z(n94) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_INV U85 ( .A(A[4]), .Z(n25) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_NAND2 U32 ( .A(n64), .B(B[16]), .Z(n63) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n76), .C(n74), .D(n72), .Z(n75) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n109), .C(n104), .D(n97), .Z(n108) );
    VMW_INV U70 ( .A(A[17]), .Z(n76) );
    VMW_INV U95 ( .A(A[1]), .Z(n21) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_INV U79 ( .A(B[19]), .Z(n80) );
    VMW_INV U87 ( .A(A[8]), .Z(n39) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n77), .Z(n85) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n117), .C(n115), .D(n113), .Z(n116) );
    VMW_INV U65 ( .A(A[12]), .Z(n52) );
    VMW_INV U102 ( .A(A[2]), .Z(n18) );
    VMW_INV U80 ( .A(A[10]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n73), .C(n68), .D(n63), .Z(n72) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n112), .C(n110), .D(n108), .Z(n111) );
    VMW_INV U89 ( .A(A[18]), .Z(n71) );
    VMW_NAND2 U50 ( .A(n94), .B(A[23]), .Z(n95) );
    VMW_INV U77 ( .A(A[25]), .Z(n105) );
    VMW_INV U92 ( .A(A[28]), .Z(n107) );
    VMW_OR2 U58 ( .A(B[28]), .B(n107), .Z(n110) );
    VMW_NAND2 U36 ( .A(n71), .B(B[18]), .Z(n70) );
    VMW_INV U81 ( .A(B[9]), .Z(n48) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n78), .C(n81), .D(n79), .Z(n82) );
    VMW_AO22 U64 ( .A(n116), .B(n118), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n91), .C(n95), .D(n93), .Z(n96) );
    VMW_INV U76 ( .A(B[25]), .Z(n102) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_INV U88 ( .A(B[21]), .Z(n86) );
    VMW_INV U93 ( .A(A[5]), .Z(n37) );
    VMW_OR2 U38 ( .A(B[18]), .B(n71), .Z(n74) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n107), .B(B[28]), .Z(n106) );
    VMW_INV U94 ( .A(B[5]), .Z(n34) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_NAND2 U63 ( .A(n117), .B(B[30]), .Z(n118) );
    VMW_INV U86 ( .A(A[24]), .Z(n91) );
    VMW_INV U103 ( .A(A[0]), .Z(n20) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_INV U78 ( .A(A[20]), .Z(n78) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_2 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n190, n149, n152, n175, n127, n217, n135, n205, n199, n140, n167, 
        n182, n120, n129, n185, n147, n160, n132, n202, n169, n210, n155, n172, 
        n197, n133, n203, n146, n161, n121, n128, n184, n218, n154, n196, n168, 
        n173, n211, n216, n126, n148, n153, n174, n183, n191, n166, n141, n134, 
        n204, n151, n193, n198, n176, n124, n214, n188, n206, n136, n143, n158, 
        n144, n164, n163, n181, n186, n178, n123, n131, n201, n213, n171, n156, 
        n130, n138, n194, n208, n179, n200, n145, n162, n187, n195, n122, n139, 
        n209, n170, n157, n125, n212, n215, n189, n150, n177, n192, n119, n142, 
        n180, n165, n159, n137, n207;
    VMW_OAI21 U3 ( .A(A[31]), .B(n119), .C(n120), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n124), .B(B[0]), .C(n125), .D(B[1]), .Z(n123) );
    VMW_OR2 U6 ( .A(B[2]), .B(n122), .Z(n126) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n152), .C(n147), .D(n142), .Z(n151) );
    VMW_OR2 U54 ( .A(B[26]), .B(n200), .Z(n203) );
    VMW_INV U73 ( .A(B[27]), .Z(n209) );
    VMW_INV U96 ( .A(B[31]), .Z(n119) );
    VMW_INV U68 ( .A(A[30]), .Z(n217) );
    VMW_NAND2 U28 ( .A(n162), .B(B[14]), .Z(n161) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n170), .C(n166), .D(n161), .Z(n169) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n125), .C(n126), .D(n123), .Z(n127) );
    VMW_NAND2 U8 ( .A(n129), .B(B[4]), .Z(n128) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n133), .D(n128), .Z(n137) );
    VMW_OR2 U34 ( .A(B[16]), .B(n168), .Z(n171) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n184), .C(n179), .D(n174), .Z(n183) );
    VMW_NAND2 U46 ( .A(n190), .B(A[21]), .Z(n191) );
    VMW_NAND2 U61 ( .A(n214), .B(A[29]), .Z(n215) );
    VMW_INV U84 ( .A(B[15]), .Z(n170) );
    VMW_INV U101 ( .A(A[6]), .Z(n136) );
    VMW_INV U66 ( .A(B[7]), .Z(n145) );
    VMW_INV U83 ( .A(A[15]), .Z(n173) );
    VMW_INV U98 ( .A(B[13]), .Z(n164) );
    VMW_NAND2 U26 ( .A(n158), .B(A[11]), .Z(n159) );
    VMW_NAND2 U48 ( .A(n194), .B(B[24]), .Z(n193) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n131), .C(n127), .D(n121), .Z(n130) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n173), .C(n171), .D(n169), .Z(n172) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n202), .C(n198), .D(n193), .Z(n201) );
    VMW_INV U91 ( .A(B[11]), .Z(n158) );
    VMW_INV U74 ( .A(A[3]), .Z(n134) );
    VMW_INV U99 ( .A(A[26]), .Z(n200) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_NAND2 U40 ( .A(n182), .B(B[20]), .Z(n181) );
    VMW_INV U82 ( .A(B[29]), .Z(n214) );
    VMW_NAND2 U52 ( .A(n200), .B(B[26]), .Z(n199) );
    VMW_INV U67 ( .A(A[7]), .Z(n148) );
    VMW_INV U75 ( .A(B[3]), .Z(n131) );
    VMW_INV U90 ( .A(A[14]), .Z(n162) );
    VMW_NAND2 U20 ( .A(n150), .B(B[10]), .Z(n149) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n196), .C(n192), .D(n187), .Z(n195) );
    VMW_INV U69 ( .A(B[17]), .Z(n177) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n188), .C(n191), .D(n189), .Z(n192) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n205), .C(n203), .D(n201), .Z(n204) );
    VMW_INV U72 ( .A(A[27]), .Z(n212) );
    VMW_INV U97 ( .A(A[16]), .Z(n168) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n214), .C(n211), .D(n206), .Z(n213) );
    VMW_INV U100 ( .A(B[23]), .Z(n196) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_INV U85 ( .A(A[4]), .Z(n129) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n145), .C(n140), .D(n135), .Z(n144) );
    VMW_NAND2 U22 ( .A(n152), .B(A[9]), .Z(n153) );
    VMW_NAND2 U32 ( .A(n168), .B(B[16]), .Z(n167) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n180), .C(n178), .D(n176), .Z(n179) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n209), .C(n204), .D(n199), .Z(n208) );
    VMW_INV U70 ( .A(A[17]), .Z(n180) );
    VMW_INV U95 ( .A(A[1]), .Z(n125) );
    VMW_NAND2 U30 ( .A(n164), .B(A[13]), .Z(n165) );
    VMW_INV U79 ( .A(B[19]), .Z(n184) );
    VMW_INV U87 ( .A(A[8]), .Z(n143) );
    VMW_OR2 U10 ( .A(B[4]), .B(n129), .Z(n132) );
    VMW_NAND2 U42 ( .A(n184), .B(A[19]), .Z(n185) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n190), .C(n186), .D(n181), .Z(n189) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n217), .C(n215), .D(n213), .Z(n216) );
    VMW_INV U65 ( .A(A[12]), .Z(n156) );
    VMW_INV U102 ( .A(A[2]), .Z(n122) );
    VMW_INV U80 ( .A(A[10]), .Z(n150) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n134), .C(n132), .D(n130), .Z(n133) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n148), .C(n146), .D(n144), .Z(n147) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n177), .C(n172), .D(n167), .Z(n176) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n212), .C(n210), .D(n208), .Z(n211) );
    VMW_INV U89 ( .A(A[18]), .Z(n175) );
    VMW_NAND2 U50 ( .A(n196), .B(A[23]), .Z(n197) );
    VMW_INV U77 ( .A(A[25]), .Z(n205) );
    VMW_INV U92 ( .A(A[28]), .Z(n207) );
    VMW_OR2 U58 ( .A(B[28]), .B(n207), .Z(n210) );
    VMW_NAND2 U36 ( .A(n175), .B(B[18]), .Z(n174) );
    VMW_INV U81 ( .A(B[9]), .Z(n152) );
    VMW_NAND2 U4 ( .A(n122), .B(B[2]), .Z(n121) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n146) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n182), .C(n185), .D(n183), .Z(n186) );
    VMW_AO22 U64 ( .A(n216), .B(n218), .C(A[31]), .D(n119), .Z(n120) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n194), .C(n197), .D(n195), .Z(n198) );
    VMW_INV U76 ( .A(B[25]), .Z(n202) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U24 ( .A(n156), .B(B[12]), .Z(n155) );
    VMW_INV U88 ( .A(B[21]), .Z(n190) );
    VMW_INV U93 ( .A(A[5]), .Z(n141) );
    VMW_OR2 U38 ( .A(B[18]), .B(n175), .Z(n178) );
    VMW_NAND2 U44 ( .A(n188), .B(B[22]), .Z(n187) );
    VMW_NAND2 U56 ( .A(n207), .B(B[28]), .Z(n206) );
    VMW_INV U94 ( .A(B[5]), .Z(n138) );
    VMW_INV U71 ( .A(A[22]), .Z(n188) );
    VMW_NAND2 U63 ( .A(n217), .B(B[30]), .Z(n218) );
    VMW_INV U86 ( .A(A[24]), .Z(n194) );
    VMW_INV U103 ( .A(A[0]), .Z(n124) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n162), .C(n165), .D(n163), .Z(n166) );
    VMW_INV U78 ( .A(A[20]), .Z(n182) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n287, n317, n245, n262, n279, n222, n230, n257, n270, n239, n295, 
        n305, n219, n292, n302, n250, n277, n225, n237, n289, n259, n265, n242, 
        n280, n310, n224, n288, n318, n276, n236, n243, n251, n264, n281, n293, 
        n303, n311, n258, n231, n238, n244, n278, n263, n286, n316, n294, n304, 
        n256, n271, n223, n228, n284, n314, n261, n246, n233, n221, n248, n253, 
        n254, n268, n273, n291, n296, n301, n306, n274, n226, n234, n298, n308, 
        n241, n266, n227, n283, n313, n249, n252, n275, n290, n300, n282, n312, 
        n240, n267, n232, n235, n299, n309, n247, n260, n229, n285, n315, n255, 
        n272, n297, n307, n269, n220;
    VMW_OAI21 U3 ( .A(A[31]), .B(n219), .C(n220), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n224), .B(B[0]), .C(n225), .D(B[1]), .Z(n223) );
    VMW_OR2 U6 ( .A(B[2]), .B(n222), .Z(n226) );
    VMW_OR2 U14 ( .A(B[6]), .B(n236), .Z(n239) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n252), .C(n247), .D(n242), .Z(n251) );
    VMW_OR2 U54 ( .A(B[26]), .B(n300), .Z(n303) );
    VMW_INV U73 ( .A(B[27]), .Z(n309) );
    VMW_INV U96 ( .A(B[31]), .Z(n219) );
    VMW_INV U68 ( .A(A[30]), .Z(n317) );
    VMW_NAND2 U28 ( .A(n262), .B(B[14]), .Z(n261) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n270), .C(n266), .D(n261), .Z(n269) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n225), .C(n226), .D(n223), .Z(n227) );
    VMW_NAND2 U8 ( .A(n229), .B(B[4]), .Z(n228) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n238), .C(n233), .D(n228), .Z(n237) );
    VMW_OR2 U34 ( .A(B[16]), .B(n268), .Z(n271) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n284), .C(n279), .D(n274), .Z(n283) );
    VMW_NAND2 U46 ( .A(n290), .B(A[21]), .Z(n291) );
    VMW_NAND2 U61 ( .A(n314), .B(A[29]), .Z(n315) );
    VMW_INV U84 ( .A(B[15]), .Z(n270) );
    VMW_INV U101 ( .A(A[6]), .Z(n236) );
    VMW_INV U66 ( .A(B[7]), .Z(n245) );
    VMW_INV U83 ( .A(A[15]), .Z(n273) );
    VMW_INV U98 ( .A(B[13]), .Z(n264) );
    VMW_NAND2 U26 ( .A(n258), .B(A[11]), .Z(n259) );
    VMW_NAND2 U48 ( .A(n294), .B(B[24]), .Z(n293) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n231), .C(n227), .D(n221), .Z(n230) );
    VMW_NAND2 U12 ( .A(n236), .B(B[6]), .Z(n235) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n273), .C(n271), .D(n269), .Z(n272) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n302), .C(n298), .D(n293), .Z(n301) );
    VMW_INV U91 ( .A(B[11]), .Z(n258) );
    VMW_INV U74 ( .A(A[3]), .Z(n234) );
    VMW_INV U99 ( .A(A[26]), .Z(n300) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n256), .C(n259), .D(n257), .Z(n260) );
    VMW_NAND2 U40 ( .A(n282), .B(B[20]), .Z(n281) );
    VMW_INV U82 ( .A(B[29]), .Z(n314) );
    VMW_NAND2 U52 ( .A(n300), .B(B[26]), .Z(n299) );
    VMW_INV U67 ( .A(A[7]), .Z(n248) );
    VMW_INV U75 ( .A(B[3]), .Z(n231) );
    VMW_INV U90 ( .A(A[14]), .Z(n262) );
    VMW_NAND2 U20 ( .A(n250), .B(B[10]), .Z(n249) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n296), .C(n292), .D(n287), .Z(n295) );
    VMW_INV U69 ( .A(B[17]), .Z(n277) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n264), .C(n260), .D(n255), .Z(n263) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n288), .C(n291), .D(n289), .Z(n292) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n305), .C(n303), .D(n301), .Z(n304) );
    VMW_INV U72 ( .A(A[27]), .Z(n312) );
    VMW_INV U97 ( .A(A[16]), .Z(n268) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n314), .C(n311), .D(n306), .Z(n313) );
    VMW_INV U100 ( .A(B[23]), .Z(n296) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n241), .C(n239), .D(n237), .Z(n240) );
    VMW_INV U85 ( .A(A[4]), .Z(n229) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n245), .C(n240), .D(n235), .Z(n244) );
    VMW_NAND2 U22 ( .A(n252), .B(A[9]), .Z(n253) );
    VMW_NAND2 U32 ( .A(n268), .B(B[16]), .Z(n267) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n280), .C(n278), .D(n276), .Z(n279) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n309), .C(n304), .D(n299), .Z(n308) );
    VMW_INV U70 ( .A(A[17]), .Z(n280) );
    VMW_INV U95 ( .A(A[1]), .Z(n225) );
    VMW_NAND2 U30 ( .A(n264), .B(A[13]), .Z(n265) );
    VMW_INV U79 ( .A(B[19]), .Z(n284) );
    VMW_INV U87 ( .A(A[8]), .Z(n243) );
    VMW_OR2 U10 ( .A(B[4]), .B(n229), .Z(n232) );
    VMW_NAND2 U42 ( .A(n284), .B(A[19]), .Z(n285) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n290), .C(n286), .D(n281), .Z(n289) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n317), .C(n315), .D(n313), .Z(n316) );
    VMW_INV U65 ( .A(A[12]), .Z(n256) );
    VMW_INV U102 ( .A(A[2]), .Z(n222) );
    VMW_INV U80 ( .A(A[10]), .Z(n250) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n234), .C(n232), .D(n230), .Z(n233) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n248), .C(n246), .D(n244), .Z(n247) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n258), .C(n254), .D(n249), .Z(n257) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n277), .C(n272), .D(n267), .Z(n276) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n312), .C(n310), .D(n308), .Z(n311) );
    VMW_INV U89 ( .A(A[18]), .Z(n275) );
    VMW_NAND2 U50 ( .A(n296), .B(A[23]), .Z(n297) );
    VMW_INV U77 ( .A(A[25]), .Z(n305) );
    VMW_INV U92 ( .A(A[28]), .Z(n307) );
    VMW_OR2 U58 ( .A(B[28]), .B(n307), .Z(n310) );
    VMW_NAND2 U36 ( .A(n275), .B(B[18]), .Z(n274) );
    VMW_INV U81 ( .A(B[9]), .Z(n252) );
    VMW_NAND2 U4 ( .A(n222), .B(B[2]), .Z(n221) );
    VMW_OR2 U18 ( .A(B[8]), .B(n243), .Z(n246) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n282), .C(n285), .D(n283), .Z(n286) );
    VMW_AO22 U64 ( .A(n316), .B(n318), .C(A[31]), .D(n219), .Z(n220) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n294), .C(n297), .D(n295), .Z(n298) );
    VMW_INV U76 ( .A(B[25]), .Z(n302) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n250), .C(n253), .D(n251), .Z(n254) );
    VMW_NAND2 U24 ( .A(n256), .B(B[12]), .Z(n255) );
    VMW_INV U88 ( .A(B[21]), .Z(n290) );
    VMW_INV U93 ( .A(A[5]), .Z(n241) );
    VMW_OR2 U38 ( .A(B[18]), .B(n275), .Z(n278) );
    VMW_NAND2 U44 ( .A(n288), .B(B[22]), .Z(n287) );
    VMW_NAND2 U56 ( .A(n307), .B(B[28]), .Z(n306) );
    VMW_INV U94 ( .A(B[5]), .Z(n238) );
    VMW_INV U71 ( .A(A[22]), .Z(n288) );
    VMW_NAND2 U63 ( .A(n317), .B(B[30]), .Z(n318) );
    VMW_INV U86 ( .A(A[24]), .Z(n294) );
    VMW_INV U103 ( .A(A[0]), .Z(n224) );
    VMW_NAND2 U16 ( .A(n243), .B(B[8]), .Z(n242) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n262), .C(n265), .D(n263), .Z(n266) );
    VMW_INV U78 ( .A(A[20]), .Z(n282) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n330, n379, n362, n339, n345, n387, n395, n406, n414, n370, n357, 
        n322, n319, n325, n389, n408, n350, n377, n392, n413, n342, n380, n401, 
        n359, n365, n337, n351, n393, n412, n376, n324, n336, n388, n409, n343, 
        n358, n364, n381, n400, n386, n407, n323, n331, n344, n363, n378, n356, 
        n371, n333, n338, n394, n415, n328, n346, n361, n384, n405, n396, n321, 
        n354, n368, n373, n326, n348, n353, n374, n383, n391, n410, n402, n341, 
        n366, n334, n390, n398, n411, n349, n352, n375, n327, n335, n399, n340, 
        n367, n329, n382, n403, n385, n404, n347, n360, n332, n320, n369, n355, 
        n372, n397, n416;
    VMW_OAI21 U3 ( .A(A[31]), .B(n319), .C(n320), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n322), .C(B[0]), .Z(n323) );
    VMW_AO22 U6 ( .A(A[2]), .B(n325), .C(n323), .D(A[0]), .Z(n324) );
    VMW_OR2 U14 ( .A(B[6]), .B(n334), .Z(n337) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n350), .C(n345), .D(n340), .Z(n349) );
    VMW_OR2 U54 ( .A(B[26]), .B(n398), .Z(n401) );
    VMW_INV U73 ( .A(B[27]), .Z(n407) );
    VMW_INV U96 ( .A(A[16]), .Z(n366) );
    VMW_INV U68 ( .A(A[30]), .Z(n415) );
    VMW_NAND2 U28 ( .A(n360), .B(B[14]), .Z(n359) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n368), .C(n364), .D(n359), .Z(n367) );
    VMW_OAI22 U7 ( .A(n321), .B(n324), .C(A[2]), .D(n325), .Z(n326) );
    VMW_NAND2 U8 ( .A(n328), .B(B[4]), .Z(n327) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n336), .C(n332), .D(n327), .Z(n335) );
    VMW_OR2 U34 ( .A(B[16]), .B(n366), .Z(n369) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n382), .C(n377), .D(n372), .Z(n381) );
    VMW_NAND2 U46 ( .A(n388), .B(A[21]), .Z(n389) );
    VMW_NAND2 U61 ( .A(n412), .B(A[29]), .Z(n413) );
    VMW_INV U84 ( .A(A[4]), .Z(n328) );
    VMW_INV U101 ( .A(B[2]), .Z(n325) );
    VMW_INV U66 ( .A(B[7]), .Z(n343) );
    VMW_INV U83 ( .A(B[15]), .Z(n368) );
    VMW_INV U98 ( .A(A[26]), .Z(n398) );
    VMW_NAND2 U26 ( .A(n356), .B(A[11]), .Z(n357) );
    VMW_NAND2 U48 ( .A(n392), .B(B[24]), .Z(n391) );
    VMW_AO21 U9 ( .A(B[3]), .B(n330), .C(n326), .Z(n329) );
    VMW_NAND2 U12 ( .A(n334), .B(B[6]), .Z(n333) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n371), .C(n369), .D(n367), .Z(n370) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n400), .C(n396), .D(n391), .Z(n399) );
    VMW_INV U91 ( .A(A[28]), .Z(n405) );
    VMW_INV U74 ( .A(A[3]), .Z(n330) );
    VMW_INV U99 ( .A(B[23]), .Z(n394) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n354), .C(n357), .D(n355), .Z(n358) );
    VMW_NAND2 U40 ( .A(n380), .B(B[20]), .Z(n379) );
    VMW_INV U82 ( .A(A[15]), .Z(n371) );
    VMW_NAND2 U52 ( .A(n398), .B(B[26]), .Z(n397) );
    VMW_INV U67 ( .A(A[7]), .Z(n346) );
    VMW_INV U75 ( .A(B[25]), .Z(n400) );
    VMW_INV U90 ( .A(B[11]), .Z(n356) );
    VMW_NAND2 U20 ( .A(n348), .B(B[10]), .Z(n347) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n394), .C(n390), .D(n385), .Z(n393) );
    VMW_INV U69 ( .A(B[17]), .Z(n375) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n362), .C(n358), .D(n353), .Z(n361) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n386), .C(n389), .D(n387), .Z(n390) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n403), .C(n401), .D(n399), .Z(n402) );
    VMW_INV U72 ( .A(A[27]), .Z(n410) );
    VMW_INV U97 ( .A(B[13]), .Z(n362) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n412), .C(n409), .D(n404), .Z(n411) );
    VMW_INV U100 ( .A(A[6]), .Z(n334) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n339), .C(n337), .D(n335), .Z(n338) );
    VMW_INV U85 ( .A(A[24]), .Z(n392) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n343), .C(n338), .D(n333), .Z(n342) );
    VMW_NAND2 U22 ( .A(n350), .B(A[9]), .Z(n351) );
    VMW_NAND2 U32 ( .A(n366), .B(B[16]), .Z(n365) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n378), .C(n376), .D(n374), .Z(n377) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n407), .C(n402), .D(n397), .Z(n406) );
    VMW_INV U70 ( .A(A[17]), .Z(n378) );
    VMW_INV U95 ( .A(B[31]), .Z(n319) );
    VMW_NAND2 U30 ( .A(n362), .B(A[13]), .Z(n363) );
    VMW_INV U79 ( .A(A[10]), .Z(n348) );
    VMW_INV U87 ( .A(B[21]), .Z(n388) );
    VMW_OR2 U10 ( .A(B[4]), .B(n328), .Z(n331) );
    VMW_NAND2 U42 ( .A(n382), .B(A[19]), .Z(n383) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n388), .C(n384), .D(n379), .Z(n387) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n415), .C(n413), .D(n411), .Z(n414) );
    VMW_INV U65 ( .A(A[12]), .Z(n354) );
    VMW_INV U80 ( .A(B[9]), .Z(n350) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n330), .C(n331), .D(n329), .Z(n332) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n346), .C(n344), .D(n342), .Z(n345) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n356), .C(n352), .D(n347), .Z(n355) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n375), .C(n370), .D(n365), .Z(n374) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n410), .C(n408), .D(n406), .Z(n409) );
    VMW_INV U89 ( .A(A[14]), .Z(n360) );
    VMW_NAND2 U50 ( .A(n394), .B(A[23]), .Z(n395) );
    VMW_INV U77 ( .A(A[20]), .Z(n380) );
    VMW_INV U92 ( .A(A[5]), .Z(n339) );
    VMW_OR2 U58 ( .A(B[28]), .B(n405), .Z(n408) );
    VMW_NAND2 U36 ( .A(n373), .B(B[18]), .Z(n372) );
    VMW_INV U81 ( .A(B[29]), .Z(n412) );
    VMW_NOR2 U4 ( .A(n322), .B(B[1]), .Z(n321) );
    VMW_OR2 U18 ( .A(B[8]), .B(n341), .Z(n344) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n380), .C(n383), .D(n381), .Z(n384) );
    VMW_AO22 U64 ( .A(n414), .B(n416), .C(A[31]), .D(n319), .Z(n320) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n392), .C(n395), .D(n393), .Z(n396) );
    VMW_INV U76 ( .A(A[25]), .Z(n403) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n348), .C(n351), .D(n349), .Z(n352) );
    VMW_NAND2 U24 ( .A(n354), .B(B[12]), .Z(n353) );
    VMW_INV U88 ( .A(A[18]), .Z(n373) );
    VMW_INV U93 ( .A(B[5]), .Z(n336) );
    VMW_OR2 U38 ( .A(B[18]), .B(n373), .Z(n376) );
    VMW_NAND2 U44 ( .A(n386), .B(B[22]), .Z(n385) );
    VMW_NAND2 U56 ( .A(n405), .B(B[28]), .Z(n404) );
    VMW_INV U94 ( .A(A[1]), .Z(n322) );
    VMW_INV U71 ( .A(A[22]), .Z(n386) );
    VMW_NAND2 U63 ( .A(n415), .B(B[30]), .Z(n416) );
    VMW_INV U86 ( .A(A[8]), .Z(n341) );
    VMW_NAND2 U16 ( .A(n341), .B(B[8]), .Z(n340) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n360), .C(n363), .D(n361), .Z(n364) );
    VMW_INV U78 ( .A(B[19]), .Z(n382) );
endmodule


module BHeap_Node_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, Enable, 
    P_WR, P_In, P_Out, L_WR, L_In, L_Out, R_WR, R_In, R_Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
output [31:0] P_Out;
output [31:0] L_Out;
input  [31:0] R_In;
input  [31:0] P_In;
input  [31:0] L_In;
output [31:0] R_Out;
input  Clk, Reset, RD, WR, Enable;
output P_WR, L_WR, R_WR;
    wire n454, n100, n421, n433, n446, n428, n441, n434, n426, n448, n90, n453, 
        n435, n449, n98, n440, n452, n427, n420, n429, n447, n439, n432, n422, 
        n417, n430, n445, n442, n437, n425, n450, n419, n436, n443, n418, n451, 
        n92, n424, n423, n438, n444, n431;
    tri \P_Out[31] , \R_Out[25]1 , \R_Out[16]1 , \R_Out[24]1 , \R_Out[17]1 , 
        \P_Out[21]1 , \P_Out[12]1 , \P_Out[20]1 , \P_Out[13]1 , \P_Out[7]1 , 
        \R_Out[2]1 , \L_Out[20]1 , \L_Out[13]1 , \L_Out[6]1 , \R_Out[3]1 , 
        \R_Out[30]1 , \R_Out[29]1 , \P_Out[6]1 , \L_Out[7]1 , \R_Out[28]1 , 
        \L_Out[21]1 , \L_Out[12]1 , \P_Out[24]1 , \P_Out[17]1 , \P_Out[25]1 , 
        \P_Out[16]1 , \L_Out[30]1 , \R_Out[20]1 , \R_Out[13]1 , \L_Out[29]1 , 
        \L_Out[28]1 , \R_Out[21]1 , \R_Out[12]1 , \L_Out[3]1 , \P_Out[2]1 , 
        \L_Out[25]1 , \L_Out[16]1 , \P_Out[3]1 , \L_Out[2]1 , \L_Out[24]1 , 
        \L_Out[17]1 , \R_Out[7]1 , \P_Out[28]1 , \P_Out[30]1 , \P_Out[29]1 , 
        \R_Out[6]1 , \P_Out[26]1 , \P_Out[15]1 , \R_Out[9]1 , \R_Out[8]1 , 
        \P_Out[27]1 , \P_Out[14]1 , \L_Out[18]1 , \R_Out[22]1 , \R_Out[11]1 , 
        \P_Out[0]1 , \L_Out[27]1 , \L_Out[19]1 , \R_Out[23]1 , \R_Out[10]1 , 
        \L_Out[1]1 , \L_Out[14]1 , \L_Out[0]1 , \P_Out[1]1 , \L_Out[26]1 , 
        \L_Out[15]1 , \R_Out[5]1 , \P_Out[19]1 , \P_Out[18]1 , \L_Out[31] , 
        \P_Out[9]1 , \L_Out[8]1 , \R_Out[4]1 , \R_Out[27]1 , \R_Out[14]1 , 
        \P_Out[23]1 , \P_Out[10]1 , \P_Out[8]1 , \L_Out[9]1 , \R_Out[26]1 , 
        \R_Out[15]1 , \P_Out[22]1 , \P_Out[11]1 , \P_Out[5]1 , \R_Out[0]1 , 
        \R_Out[1]1 , \L_Out[22]1 , \L_Out[11]1 , \L_Out[4]1 , \R_Out[18]1 , 
        \R_Out[31] , \P_Out[4]1 , \L_Out[5]1 , \R_Out[19]1 , \L_Out[23]1 , 
        \L_Out[10]1 ;
    assign P_Out[31] = \P_Out[31] ;
    assign P_Out[30] = \P_Out[30]1 ;
    assign P_Out[29] = \P_Out[29]1 ;
    assign P_Out[28] = \P_Out[28]1 ;
    assign P_Out[27] = \P_Out[27]1 ;
    assign P_Out[26] = \P_Out[26]1 ;
    assign P_Out[25] = \P_Out[25]1 ;
    assign P_Out[24] = \P_Out[24]1 ;
    assign P_Out[23] = \P_Out[23]1 ;
    assign P_Out[22] = \P_Out[22]1 ;
    assign P_Out[21] = \P_Out[21]1 ;
    assign P_Out[20] = \P_Out[20]1 ;
    assign P_Out[19] = \P_Out[19]1 ;
    assign P_Out[18] = \P_Out[18]1 ;
    assign P_Out[17] = \P_Out[17]1 ;
    assign P_Out[16] = \P_Out[16]1 ;
    assign P_Out[15] = \P_Out[15]1 ;
    assign P_Out[14] = \P_Out[14]1 ;
    assign P_Out[13] = \P_Out[13]1 ;
    assign P_Out[12] = \P_Out[12]1 ;
    assign P_Out[11] = \P_Out[11]1 ;
    assign P_Out[10] = \P_Out[10]1 ;
    assign P_Out[9] = \P_Out[9]1 ;
    assign P_Out[8] = \P_Out[8]1 ;
    assign P_Out[7] = \P_Out[7]1 ;
    assign P_Out[6] = \P_Out[6]1 ;
    assign P_Out[5] = \P_Out[5]1 ;
    assign P_Out[4] = \P_Out[4]1 ;
    assign P_Out[3] = \P_Out[3]1 ;
    assign P_Out[2] = \P_Out[2]1 ;
    assign P_Out[1] = \P_Out[1]1 ;
    assign P_Out[0] = \P_Out[0]1 ;
    assign L_Out[31] = \L_Out[31] ;
    assign L_Out[30] = \L_Out[30]1 ;
    assign L_Out[29] = \L_Out[29]1 ;
    assign L_Out[28] = \L_Out[28]1 ;
    assign L_Out[27] = \L_Out[27]1 ;
    assign L_Out[26] = \L_Out[26]1 ;
    assign L_Out[25] = \L_Out[25]1 ;
    assign L_Out[24] = \L_Out[24]1 ;
    assign L_Out[23] = \L_Out[23]1 ;
    assign L_Out[22] = \L_Out[22]1 ;
    assign L_Out[21] = \L_Out[21]1 ;
    assign L_Out[20] = \L_Out[20]1 ;
    assign L_Out[19] = \L_Out[19]1 ;
    assign L_Out[18] = \L_Out[18]1 ;
    assign L_Out[17] = \L_Out[17]1 ;
    assign L_Out[16] = \L_Out[16]1 ;
    assign L_Out[15] = \L_Out[15]1 ;
    assign L_Out[14] = \L_Out[14]1 ;
    assign L_Out[13] = \L_Out[13]1 ;
    assign L_Out[12] = \L_Out[12]1 ;
    assign L_Out[11] = \L_Out[11]1 ;
    assign L_Out[10] = \L_Out[10]1 ;
    assign L_Out[9] = \L_Out[9]1 ;
    assign L_Out[8] = \L_Out[8]1 ;
    assign L_Out[7] = \L_Out[7]1 ;
    assign L_Out[6] = \L_Out[6]1 ;
    assign L_Out[5] = \L_Out[5]1 ;
    assign L_Out[4] = \L_Out[4]1 ;
    assign L_Out[3] = \L_Out[3]1 ;
    assign L_Out[2] = \L_Out[2]1 ;
    assign L_Out[1] = \L_Out[1]1 ;
    assign L_Out[0] = \L_Out[0]1 ;
    assign R_Out[31] = \R_Out[31] ;
    assign R_Out[30] = \R_Out[30]1 ;
    assign R_Out[29] = \R_Out[29]1 ;
    assign R_Out[28] = \R_Out[28]1 ;
    assign R_Out[27] = \R_Out[27]1 ;
    assign R_Out[26] = \R_Out[26]1 ;
    assign R_Out[25] = \R_Out[25]1 ;
    assign R_Out[24] = \R_Out[24]1 ;
    assign R_Out[23] = \R_Out[23]1 ;
    assign R_Out[22] = \R_Out[22]1 ;
    assign R_Out[21] = \R_Out[21]1 ;
    assign R_Out[20] = \R_Out[20]1 ;
    assign R_Out[19] = \R_Out[19]1 ;
    assign R_Out[18] = \R_Out[18]1 ;
    assign R_Out[17] = \R_Out[17]1 ;
    assign R_Out[16] = \R_Out[16]1 ;
    assign R_Out[15] = \R_Out[15]1 ;
    assign R_Out[14] = \R_Out[14]1 ;
    assign R_Out[13] = \R_Out[13]1 ;
    assign R_Out[12] = \R_Out[12]1 ;
    assign R_Out[11] = \R_Out[11]1 ;
    assign R_Out[10] = \R_Out[10]1 ;
    assign R_Out[9] = \R_Out[9]1 ;
    assign R_Out[8] = \R_Out[8]1 ;
    assign R_Out[7] = \R_Out[7]1 ;
    assign R_Out[6] = \R_Out[6]1 ;
    assign R_Out[5] = \R_Out[5]1 ;
    assign R_Out[4] = \R_Out[4]1 ;
    assign R_Out[3] = \R_Out[3]1 ;
    assign R_Out[2] = \R_Out[2]1 ;
    assign R_Out[1] = \R_Out[1]1 ;
    assign R_Out[0] = \R_Out[0]1 ;
    VMW_AO22 U54 ( .A(R_In[26]), .B(n417), .C(L_In[26]), .D(L_WR), .Z(n431) );
    VMW_AND3 U73 ( .A(n92), .B(Enable), .C(n90), .Z(L_WR) );
    VMW_BUFIZ U113 ( .A(P_In[3]), .E(L_WR), .Z(\L_Out[3]1 ) );
    VMW_BUFIZ U134 ( .A(P_In[22]), .E(R_WR), .Z(\R_Out[22]1 ) );
    VMW_AO22 U68 ( .A(R_In[13]), .B(n417), .C(L_In[13]), .D(L_WR), .Z(n426) );
    VMW_BUFIZ U96 ( .A(n421), .E(P_WR), .Z(\P_Out[17]1 ) );
    VMW_BUFIZ U108 ( .A(P_In[12]), .E(R_WR), .Z(\R_Out[12]1 ) );
    VMW_BUFIZ U141 ( .A(n444), .E(P_WR), .Z(\P_Out[3]1 ) );
    VMW_BUFIZ U166 ( .A(P_In[4]), .E(R_WR), .Z(\R_Out[4]1 ) );
    VMW_PULLDOWN U35 ( .Z(n451) );
    VMW_AO22 U41 ( .A(R_In[9]), .B(n417), .C(L_In[9]), .D(L_WR), .Z(n429) );
    VMW_AO22 U46 ( .A(R_In[4]), .B(n417), .C(L_In[4]), .D(L_WR), .Z(n433) );
    VMW_AO22 U61 ( .A(R_In[1]), .B(n417), .C(L_In[1]), .D(L_WR), .Z(n443) );
    VMW_BUFIZ U84 ( .A(P_In[24]), .E(L_WR), .Z(\L_Out[24]1 ) );
    VMW_BUFIZ U148 ( .A(P_In[13]), .E(R_WR), .Z(\R_Out[13]1 ) );
    VMW_BUFIZ U153 ( .A(n449), .E(P_WR), .Z(\P_Out[16]1 ) );
    VMW_BUFIZ U101 ( .A(n424), .E(P_WR), .Z(\P_Out[20]1 ) );
    VMW_BUFIZ U126 ( .A(n434), .E(P_WR), .Z(\P_Out[27]1 ) );
    VMW_AO22 U48 ( .A(R_In[31]), .B(n417), .C(L_In[31]), .D(L_WR), .Z(n440) );
    VMW_AO22 U66 ( .A(R_In[15]), .B(n417), .C(L_In[15]), .D(L_WR), .Z(n432) );
    VMW_BUFIZ U106 ( .A(P_In[28]), .E(R_WR), .Z(\R_Out[28]1 ) );
    VMW_BUFIZ U121 ( .A(n432), .E(P_WR), .Z(\P_Out[15]1 ) );
    VMW_BUFIZ U83 ( .A(P_In[15]), .E(L_WR), .Z(\L_Out[15]1 ) );
    VMW_BUFIZ U168 ( .A(P_In[9]), .E(R_WR), .Z(\R_Out[9]1 ) );
    VMW_BUFIZ U98 ( .A(P_In[16]), .E(R_WR), .Z(\R_Out[16]1 ) );
    VMW_BUFIZ U128 ( .A(n436), .E(P_WR), .Z(\P_Out[14]1 ) );
    VMW_BUFIZ U154 ( .A(P_In[24]), .E(R_WR), .Z(\R_Out[24]1 ) );
    VMW_AO22 U53 ( .A(R_In[27]), .B(n417), .C(L_In[27]), .D(L_WR), .Z(n434) );
    VMW_BUFIZ U91 ( .A(n420), .E(P_WR), .Z(\P_Out[6]1 ) );
    VMW_BUFIZ U146 ( .A(P_In[9]), .E(L_WR), .Z(\L_Out[9]1 ) );
    VMW_BUFIZ U161 ( .A(P_In[25]), .E(L_WR), .Z(\L_Out[25]1 ) );
    VMW_AND3 U74 ( .A(n98), .B(n100), .C(Enable), .Z(R_WR) );
    VMW_BUFIZ U114 ( .A(P_In[23]), .E(R_WR), .Z(\R_Out[23]1 ) );
    VMW_BUFIZ U133 ( .A(P_In[2]), .E(L_WR), .Z(\L_Out[2]1 ) );
    VMW_BUFIZ U99 ( .A(n422), .E(P_WR), .Z(\P_Out[29]1 ) );
    VMW_BUFIZ U155 ( .A(P_In[17]), .E(R_WR), .Z(\R_Out[17]1 ) );
    VMW_OR2 U40 ( .A(L_WR), .B(R_WR), .Z(P_WR) );
    VMW_BUFIZ U82 ( .A(P_In[26]), .E(L_WR), .Z(\L_Out[26]1 ) );
    VMW_BUFIZ U169 ( .A(P_In[23]), .E(L_WR), .Z(\L_Out[23]1 ) );
    VMW_AO22 U47 ( .A(R_In[3]), .B(n417), .C(L_In[3]), .D(L_WR), .Z(n444) );
    VMW_AO22 U49 ( .A(R_In[30]), .B(n417), .C(L_In[30]), .D(L_WR), .Z(n418) );
    VMW_AO22 U52 ( .A(R_In[28]), .B(n417), .C(L_In[28]), .D(L_WR), .Z(n441) );
    VMW_AO22 U67 ( .A(R_In[14]), .B(n417), .C(L_In[14]), .D(L_WR), .Z(n436) );
    VMW_BUFIZ U107 ( .A(P_In[21]), .E(R_WR), .Z(\R_Out[21]1 ) );
    VMW_BUFIZ U120 ( .A(n431), .E(P_WR), .Z(\P_Out[26]1 ) );
    VMW_INV U75 ( .A(L_WR), .Z(n417) );
    VMW_BUFIZ U115 ( .A(P_In[10]), .E(R_WR), .Z(\R_Out[10]1 ) );
    VMW_BUFIZ U132 ( .A(n439), .E(P_WR), .Z(\P_Out[8]1 ) );
    VMW_BUFIZ U90 ( .A(n419), .E(P_WR), .Z(\P_Out[24]1 ) );
    VMW_BUFIZ U129 ( .A(n437), .E(P_WR), .Z(\P_Out[5]1 ) );
    VMW_BUFIZ U147 ( .A(P_In[20]), .E(R_WR), .Z(\R_Out[20]1 ) );
    VMW_BUFIZ U160 ( .A(P_In[28]), .E(L_WR), .Z(\L_Out[28]1 ) );
    VMW_AO22 U55 ( .A(R_In[25]), .B(n417), .C(L_In[25]), .D(L_WR), .Z(n448) );
    VMW_AO22 U69 ( .A(R_In[12]), .B(n417), .C(L_In[12]), .D(L_WR), .Z(n446) );
    VMW_BUFIZ U109 ( .A(n426), .E(P_WR), .Z(\P_Out[13]1 ) );
    VMW_AO22 U72 ( .A(R_In[0]), .B(n417), .C(L_In[0]), .D(L_WR), .Z(n430) );
    VMW_BUFIZ U97 ( .A(P_In[25]), .E(R_WR), .Z(\R_Out[25]1 ) );
    VMW_BUFIZ U140 ( .A(n443), .E(P_WR), .Z(\P_Out[1]1 ) );
    VMW_BUFIZ U167 ( .A(P_In[19]), .E(L_WR), .Z(\L_Out[19]1 ) );
    VMW_BUFIZ U112 ( .A(n429), .E(P_WR), .Z(\P_Out[9]1 ) );
    VMW_BUFIZ U135 ( .A(P_In[11]), .E(R_WR), .Z(\R_Out[11]1 ) );
    VMW_AO22 U60 ( .A(R_In[20]), .B(n417), .C(L_In[20]), .D(L_WR), .Z(n424) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_1 gt_48_1 ( .A(L_In), .B(R_In), .LEQ(n452), 
        .TC(n452), .LT_LE(n100) );
    VMW_BUFIZ U100 ( .A(n423), .E(P_WR), .Z(\P_Out[22]1 ) );
    VMW_BUFIZ U127 ( .A(n435), .E(P_WR), .Z(\P_Out[23]1 ) );
    VMW_BUFIZ U85 ( .A(P_In[17]), .E(L_WR), .Z(\L_Out[17]1 ) );
    VMW_BUFIZ U149 ( .A(n446), .E(P_WR), .Z(\P_Out[12]1 ) );
    VMW_BUFIZ U152 ( .A(n448), .E(P_WR), .Z(\P_Out[25]1 ) );
    VMW_PULLUP U36 ( .Z(n450) );
    VMW_PULLDOWN U37 ( .Z(n452) );
    VMW_PULLDOWN U39 ( .Z(n454) );
    VMW_AO22 U57 ( .A(R_In[23]), .B(n417), .C(L_In[23]), .D(L_WR), .Z(n435) );
    VMW_BUFIZ U137 ( .A(n441), .E(P_WR), .Z(\P_Out[28]1 ) );
    VMW_AO22 U70 ( .A(R_In[11]), .B(n417), .C(L_In[11]), .D(L_WR), .Z(n428) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_2 gt_48 ( .A(P_In), .B(R_In), .LEQ(n453), 
        .TC(n453), .LT_LE(n98) );
    VMW_BUFIZ U110 ( .A(n427), .E(P_WR), .Z(\P_Out[18]1 ) );
    VMW_BUFIZ U159 ( .A(P_In[12]), .E(L_WR), .Z(\L_Out[12]1 ) );
    VMW_AO22 U42 ( .A(R_In[8]), .B(n417), .C(L_In[8]), .D(L_WR), .Z(n439) );
    VMW_AO22 U45 ( .A(R_In[5]), .B(n417), .C(L_In[5]), .D(L_WR), .Z(n437) );
    VMW_BUFIZ U79 ( .A(P_In[11]), .E(L_WR), .Z(\L_Out[11]1 ) );
    VMW_BUFIZ U95 ( .A(P_In[5]), .E(L_WR), .Z(\L_Out[5]1 ) );
    VMW_BUFIZ U119 ( .A(P_In[14]), .E(R_WR), .Z(\R_Out[14]1 ) );
    VMW_BUFIZ U142 ( .A(P_In[0]), .E(L_WR), .Z(\L_Out[0]1 ) );
    VMW_BUFIZ U165 ( .A(P_In[14]), .E(L_WR), .Z(\L_Out[14]1 ) );
    VMW_BUFIZ U87 ( .A(P_In[13]), .E(L_WR), .Z(\L_Out[13]1 ) );
    VMW_BUFIZ U150 ( .A(n447), .E(P_WR), .Z(\P_Out[7]1 ) );
    VMW_BUFIZ U125 ( .A(P_In[15]), .E(R_WR), .Z(\R_Out[15]1 ) );
    VMW_AO22 U62 ( .A(R_In[19]), .B(n417), .C(L_In[19]), .D(L_WR), .Z(n442) );
    VMW_AO22 U65 ( .A(R_In[16]), .B(n417), .C(L_In[16]), .D(L_WR), .Z(n449) );
    VMW_BUFIZ U102 ( .A(n425), .E(P_WR), .Z(\P_Out[2]1 ) );
    VMW_BUFIZ U105 ( .A(P_In[31]), .E(R_WR), .Z(\R_Out[31] ) );
    VMW_BUFIZ U80 ( .A(P_In[5]), .E(R_WR), .Z(\R_Out[5]1 ) );
    VMW_BUFIZ U122 ( .A(n433), .E(P_WR), .Z(\P_Out[4]1 ) );
    VMW_BUFIZ U157 ( .A(P_In[31]), .E(L_WR), .Z(\L_Out[31] ) );
    VMW_BUFIZ U170 ( .A(P_In[10]), .E(L_WR), .Z(\L_Out[10]1 ) );
    VMW_AO22 U50 ( .A(R_In[2]), .B(n417), .C(L_In[2]), .D(L_WR), .Z(n425) );
    VMW_AO22 U59 ( .A(R_In[21]), .B(n417), .C(L_In[21]), .D(L_WR), .Z(n445) );
    VMW_BUFIZ U139 ( .A(P_In[18]), .E(R_WR), .Z(\R_Out[18]1 ) );
    VMW_BUFIZ U77 ( .A(P_In[18]), .E(L_WR), .Z(\L_Out[18]1 ) );
    VMW_BUFIZ U89 ( .A(n418), .E(P_WR), .Z(\P_Out[30]1 ) );
    VMW_BUFIZ U92 ( .A(P_In[30]), .E(L_WR), .Z(\L_Out[30]1 ) );
    VMW_BUFIZ U145 ( .A(n445), .E(P_WR), .Z(\P_Out[21]1 ) );
    VMW_BUFIZ U162 ( .A(P_In[16]), .E(L_WR), .Z(\L_Out[16]1 ) );
    VMW_BUFIZ U117 ( .A(n430), .E(P_WR), .Z(\P_Out[0]1 ) );
    VMW_AO22 U58 ( .A(R_In[22]), .B(n417), .C(L_In[22]), .D(L_WR), .Z(n423) );
    VMW_BUFIZ U130 ( .A(P_In[6]), .E(L_WR), .Z(\L_Out[6]1 ) );
    VMW_BUFIZ U138 ( .A(n442), .E(P_WR), .Z(\P_Out[19]1 ) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_3 gt_47 ( .A(P_In), .B(L_In), .LEQ(n454), 
        .TC(n454), .LT_LE(n90) );
    VMW_BUFIZ U156 ( .A(P_In[2]), .E(R_WR), .Z(\R_Out[2]1 ) );
    VMW_BUFIZ U171 ( .A(P_In[0]), .E(R_WR), .Z(\R_Out[0]1 ) );
    VMW_PULLDOWN U38 ( .Z(n453) );
    VMW_AO22 U43 ( .A(R_In[7]), .B(n417), .C(L_In[7]), .D(L_WR), .Z(n447) );
    VMW_AO22 U64 ( .A(R_In[17]), .B(n417), .C(L_In[17]), .D(L_WR), .Z(n421) );
    VMW_BUFIZ U81 ( .A(P_In[1]), .E(R_WR), .Z(\R_Out[1]1 ) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_0 gte_47 ( .A(R_In), .B(L_In), .LEQ(n450), 
        .TC(n451), .LT_LE(n92) );
    VMW_BUFIZ U104 ( .A(P_In[1]), .E(L_WR), .Z(\L_Out[1]1 ) );
    VMW_AO22 U51 ( .A(R_In[29]), .B(n417), .C(L_In[29]), .D(L_WR), .Z(n422) );
    VMW_BUFIZ U76 ( .A(P_In[22]), .E(L_WR), .Z(\L_Out[22]1 ) );
    VMW_BUFIZ U116 ( .A(P_In[19]), .E(R_WR), .Z(\R_Out[19]1 ) );
    VMW_BUFIZ U123 ( .A(P_In[7]), .E(L_WR), .Z(\L_Out[7]1 ) );
    VMW_BUFIZ U88 ( .A(P_In[3]), .E(R_WR), .Z(\R_Out[3]1 ) );
    VMW_BUFIZ U93 ( .A(P_In[29]), .E(L_WR), .Z(\L_Out[29]1 ) );
    VMW_BUFIZ U131 ( .A(n438), .E(P_WR), .Z(\P_Out[10]1 ) );
    VMW_BUFIZ U143 ( .A(P_In[30]), .E(R_WR), .Z(\R_Out[30]1 ) );
    VMW_BUFIZ U144 ( .A(P_In[29]), .E(R_WR), .Z(\R_Out[29]1 ) );
    VMW_BUFIZ U163 ( .A(P_In[6]), .E(R_WR), .Z(\R_Out[6]1 ) );
    VMW_BUFIZ U158 ( .A(P_In[21]), .E(L_WR), .Z(\L_Out[21]1 ) );
    VMW_BUFIZ U164 ( .A(P_In[27]), .E(L_WR), .Z(\L_Out[27]1 ) );
    VMW_AO22 U44 ( .A(R_In[6]), .B(n417), .C(L_In[6]), .D(L_WR), .Z(n420) );
    VMW_AO22 U56 ( .A(R_In[24]), .B(n417), .C(L_In[24]), .D(L_WR), .Z(n419) );
    VMW_BUFIZ U94 ( .A(P_In[20]), .E(L_WR), .Z(\L_Out[20]1 ) );
    VMW_BUFIZ U136 ( .A(n440), .E(P_WR), .Z(\P_Out[31] ) );
    VMW_AO22 U71 ( .A(R_In[10]), .B(n417), .C(L_In[10]), .D(L_WR), .Z(n438) );
    VMW_BUFIZ U111 ( .A(n428), .E(P_WR), .Z(\P_Out[11]1 ) );
    VMW_BUFIZ U124 ( .A(P_In[26]), .E(R_WR), .Z(\R_Out[26]1 ) );
    VMW_AO22 U63 ( .A(R_In[18]), .B(n417), .C(L_In[18]), .D(L_WR), .Z(n427) );
    VMW_BUFIZ U78 ( .A(P_In[8]), .E(R_WR), .Z(\R_Out[8]1 ) );
    VMW_BUFIZ U86 ( .A(P_In[7]), .E(R_WR), .Z(\R_Out[7]1 ) );
    VMW_BUFIZ U103 ( .A(P_In[8]), .E(L_WR), .Z(\L_Out[8]1 ) );
    VMW_BUFIZ U118 ( .A(P_In[27]), .E(R_WR), .Z(\R_Out[27]1 ) );
    VMW_BUFIZ U151 ( .A(P_In[4]), .E(L_WR), .Z(\L_Out[4]1 ) );
endmodule


module BHeap_CtrlReg_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, In, 
    Out, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR, In;
output Out, Enable;
    wire n77, Out70;
    assign Enable = Out;
    VMW_NOR2 U12 ( .A(n77), .B(Reset), .Z(Out70) );
    VMW_INV U13 ( .A(In), .Z(n77) );
    VMW_FD Out_reg ( .D(Out70), .CP(Clk), .Q(Out) );
endmodule


module BHeap_Control_CWIDTH3_IDWIDTH1_WIDTH32_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, Go, Done );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR, Done;
output ScanEnable, Go;
    wire \Count[0] , n379, n362, n345, n387, n339, n395, n370, n357, n389, 
        n377, n350, n392, n380, n342, n365, \Count[2] , n359, n356, n393, n376, 
        n351, \ScanReg[15] , \ScanReg[26] , \ScanReg[2] , n388, \ScanReg[18] , 
        n358, n343, n364, n381, \ScanReg[11] , \ScanReg[6] , \ScanReg[22] , 
        n344, n386, \ScanReg[20] , \ScanReg[13] , \ScanReg[4] , n363, n378, 
        \ScanReg[29] , \ScanReg[30] , \ScanReg[17] , \ScanReg[24] , 
        \ScanReg[0] , n371, \ScanReg[9] , n338, n394, \ScanReg[16] , 
        \ScanReg[25] , Go259, \ScanReg[1] , \ScanReg[8] , n346, n361, 
        \ScanReg[7] , n384, \ScanReg[5] , n396, \ScanReg[21] , \ScanReg[12] , 
        n373, n354, n368, \ScanReg[28] , \ScanReg[31] , \ScanReg[19] , n348, 
        n374, n353, n391, \ScanReg[10] , n383, \ScanReg[23] , n341, n366, 
        \ScanReg[14] , \ScanReg[27] , \ScanReg[3] , n398, n390, n375, n352, 
        n349, n360, n340, n367, n382, n385, n347, \Count[1] , n369, n372, n355, 
        n397;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U68 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_AND2 U73 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_AO22 U96 ( .A(n344), .B(n343), .C(\Count[2] ), .D(n345), .Z(n396) );
    VMW_AND2 U113 ( .A(\ScanReg[21] ), .B(n346), .Z(n377) );
    VMW_NOR2 U134 ( .A(\Count[1] ), .B(\Count[0] ), .Z(n355) );
    VMW_FD \Count_reg[0]  ( .D(n398), .CP(Clk), .Q(\Count[0] ) );
    VMW_AND2 U108 ( .A(\ScanReg[20] ), .B(n346), .Z(n383) );
    VMW_OR2 U141 ( .A(Done), .B(n350), .Z(n343) );
    VMW_BUFIZ U166 ( .A(n373), .E(n368), .Z(\arr[16] ) );
    VMW_BUFIZ U183 ( .A(n390), .E(n368), .Z(\arr[15] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AND2 U66 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U84 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_OR2 U148 ( .A(Reset), .B(n356), .Z(n357) );
    VMW_INV U153 ( .A(\Count[0] ), .Z(n349) );
    VMW_BUFIZ U174 ( .A(n381), .E(n368), .Z(\arr[30] ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U101 ( .A(\ScanReg[15] ), .B(n346), .Z(n390) );
    VMW_AND2 U106 ( .A(\ScanReg[24] ), .B(n346), .Z(n385) );
    VMW_AND2 U121 ( .A(\ScanReg[4] ), .B(n346), .Z(n369) );
    VMW_AND2 U126 ( .A(\ScanReg[19] ), .B(n346), .Z(n363) );
    VMW_AND2 U74 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U83 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_BUFIZ U168 ( .A(n375), .E(n368), .Z(\arr[12] ) );
    VMW_AND2 U91 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_AND2 U98 ( .A(\ScanReg[11] ), .B(n346), .Z(n393) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_NOR3 U128 ( .A(DataIn[0]), .B(DataIn[2]), .C(DataIn[1]), .Z(n338) );
    VMW_INV U154 ( .A(n353), .Z(ScanEnable) );
    VMW_BUFIZ U173 ( .A(n380), .E(n368), .Z(\arr[13] ) );
    VMW_BUFIZ U184 ( .A(n391), .E(n368), .Z(\arr[18] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_OAI22 U146 ( .A(n362), .B(n339), .C(n350), .D(n360), .Z(n342) );
    VMW_BUFIZ U161 ( .A(n367), .E(n368), .Z(\arr[9] ) );
    VMW_AND2 U114 ( .A(\ScanReg[31] ), .B(n346), .Z(n376) );
    VMW_OAI21 U133 ( .A(RD), .B(WR), .C(n354), .Z(n353) );
    VMW_AND2 U99 ( .A(\ScanReg[22] ), .B(n346), .Z(n392) );
    VMW_FD \Count_reg[2]  ( .D(n396), .CP(Clk), .Q(\Count[2] ) );
    VMW_INV U155 ( .A(n355), .Z(n360) );
    VMW_BUFIZ U172 ( .A(n379), .E(n368), .Z(\arr[2] ) );
    VMW_AND2 U67 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U82 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_BUFIZ U169 ( .A(n376), .E(n368), .Z(\arr[31] ) );
    VMW_AND2 U107 ( .A(\ScanReg[3] ), .B(n346), .Z(n384) );
    VMW_AND2 U120 ( .A(\ScanReg[27] ), .B(n346), .Z(n370) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_AND2 U69 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U75 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AND2 U115 ( .A(\ScanReg[12] ), .B(n346), .Z(n375) );
    VMW_OR2 U132 ( .A(Reset), .B(n352), .Z(n339) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U90 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AND2 U109 ( .A(\ScanReg[29] ), .B(n346), .Z(n382) );
    VMW_XOR2 U129 ( .A(Addr[0]), .B(Id), .Z(n346) );
    VMW_XNOR2 U147 ( .A(Addr[0]), .B(ScanId), .Z(n354) );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_BUFIZ U160 ( .A(n366), .E(n368), .Z(\arr[10] ) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_BUFIZ U185 ( .A(n392), .E(n368), .Z(\arr[22] ) );
    VMW_BUFIZ U182 ( .A(n389), .E(n368), .Z(\arr[26] ) );
    VMW_AND2 U72 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_AND2 U97 ( .A(\ScanReg[8] ), .B(n346), .Z(n395) );
    VMW_OR3 U140 ( .A(n348), .B(n350), .C(n358), .Z(n340) );
    VMW_BUFIZ U167 ( .A(n374), .E(n368), .Z(\arr[6] ) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD Go_reg ( .D(Go259), .CP(Clk), .Q(Go) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_AND2 U85 ( .A(WR), .B(DataIn[9]), .Z(ScanOut[9]) );
    VMW_AND2 U100 ( .A(\ScanReg[18] ), .B(n346), .Z(n391) );
    VMW_AND2 U112 ( .A(\ScanReg[28] ), .B(n346), .Z(n378) );
    VMW_AO22 U135 ( .A(\Count[2] ), .B(n347), .C(\ScanReg[2] ), .D(n346), .Z(
        n379) );
    VMW_NOR3 U127 ( .A(\Count[2] ), .B(\Count[1] ), .C(n349), .Z(n348) );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_INV U149 ( .A(n346), .Z(n347) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_INV U152 ( .A(n352), .Z(n351) );
    VMW_BUFIZ U175 ( .A(n382), .E(n368), .Z(\arr[29] ) );
    VMW_OAI21 U62 ( .A(n338), .B(n339), .C(n340), .Z(Go259) );
    VMW_AND2 U70 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_AO22 U137 ( .A(\Count[0] ), .B(n347), .C(\ScanReg[0] ), .D(n346), .Z(
        n364) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AND2 U79 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_AO22 U95 ( .A(\Count[1] ), .B(n341), .C(n342), .D(n343), .Z(n397) );
    VMW_AND2 U110 ( .A(\ScanReg[30] ), .B(n346), .Z(n381) );
    VMW_BUFIZ U159 ( .A(n365), .E(n368), .Z(\arr[23] ) );
    VMW_AND2 U119 ( .A(\ScanReg[14] ), .B(n346), .Z(n371) );
    VMW_OR3 U142 ( .A(\Count[2] ), .B(n350), .C(n360), .Z(n359) );
    VMW_BUFIZ U165 ( .A(n372), .E(n368), .Z(\arr[25] ) );
    VMW_BUFIZ U180 ( .A(n387), .E(n368), .Z(\arr[7] ) );
    VMW_AND2 U87 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_INV U150 ( .A(DataIn[2]), .Z(n361) );
    VMW_BUFIZ U177 ( .A(n384), .E(n368), .Z(\arr[3] ) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO21 U125 ( .A(RD), .B(ScanEnable), .C(n347), .Z(n368) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U63 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U64 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U65 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U102 ( .A(\ScanReg[26] ), .B(n346), .Z(n389) );
    VMW_AND2 U105 ( .A(\ScanReg[17] ), .B(n346), .Z(n386) );
    VMW_AND2 U77 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AND2 U80 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U122 ( .A(\ScanReg[9] ), .B(n346), .Z(n367) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_AND2 U89 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_MUX2I U139 ( .A(n349), .B(n357), .S(n343), .Z(n398) );
    VMW_BUFIZ U157 ( .A(n363), .E(n368), .Z(\arr[19] ) );
    VMW_BUFIZ U170 ( .A(n377), .E(n368), .Z(\arr[21] ) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_BUFIZ U187 ( .A(n394), .E(n368), .Z(\arr[1] ) );
    VMW_AND2 U92 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_OAI21 U145 ( .A(n349), .B(n350), .C(n343), .Z(n341) );
    VMW_BUFIZ U162 ( .A(n369), .E(n368), .Z(\arr[4] ) );
    VMW_BUFIZ U179 ( .A(n386), .E(n368), .Z(\arr[17] ) );
    VMW_AND2 U117 ( .A(\ScanReg[16] ), .B(n346), .Z(n373) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AND2 U81 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_OR2 U130 ( .A(Reset), .B(n351), .Z(n350) );
    VMW_MUX2I U138 ( .A(DataIn[0]), .B(n349), .S(n352), .Z(n356) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_INV U156 ( .A(DataIn[1]), .Z(n362) );
    VMW_BUFIZ U171 ( .A(n378), .E(n368), .Z(\arr[28] ) );
    VMW_AND2 U104 ( .A(\ScanReg[7] ), .B(n346), .Z(n387) );
    VMW_AND2 U71 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U76 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AND2 U116 ( .A(\ScanReg[6] ), .B(n346), .Z(n374) );
    VMW_AND2 U123 ( .A(\ScanReg[10] ), .B(n346), .Z(n366) );
    VMW_AND2 U88 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_AND2 U93 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_NAND2 U131 ( .A(WR), .B(n347), .Z(n352) );
    VMW_BUFIZ U178 ( .A(n385), .E(n368), .Z(\arr[24] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_OAI21 U143 ( .A(n361), .B(n339), .C(n359), .Z(n344) );
    VMW_OAI21 U144 ( .A(n355), .B(n350), .C(n343), .Z(n345) );
    VMW_BUFIZ U163 ( .A(n370), .E(n368), .Z(\arr[27] ) );
    VMW_BUFIZ U181 ( .A(n388), .E(n368), .Z(\arr[5] ) );
    VMW_BUFIZ U186 ( .A(n393), .E(n368), .Z(\arr[11] ) );
    VMW_BUFIZ U158 ( .A(n364), .E(n368), .Z(\arr[0] ) );
    VMW_BUFIZ U164 ( .A(n371), .E(n368), .Z(\arr[14] ) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(\Count[1] ), .B(n347), .C(\ScanReg[1] ), .D(n346), .Z(
        n394) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AND2 U111 ( .A(\ScanReg[13] ), .B(n346), .Z(n380) );
    VMW_AND2 U124 ( .A(\ScanReg[23] ), .B(n346), .Z(n365) );
    VMW_AND2 U78 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_AND2 U86 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U103 ( .A(\ScanReg[5] ), .B(n346), .Z(n388) );
    VMW_BUFIZ U188 ( .A(n395), .E(n368), .Z(\arr[8] ) );
    VMW_FD \Count_reg[1]  ( .D(n397), .CP(Clk), .Q(\Count[1] ) );
    VMW_AND2 U118 ( .A(\ScanReg[25] ), .B(n346), .Z(n372) );
    VMW_INV U151 ( .A(Done), .Z(n358) );
    VMW_BUFIZ U176 ( .A(n383), .E(n368), .Z(\arr[20] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \wRegInTop_3_7[11] , \wRegOut_4_3[16] , \ScanLink0[13] , 
        \wRegInTop_1_0[15] , \ScanLink24[18] , \ScanLink50[8] , 
        \ScanLink51[31] , \ScanLink51[28] , \wRegInTop_5_19[16] , 
        \wRegInTop_1_0[26] , \wRegOut_3_1[3] , \wRegInTop_3_7[22] , 
        \wRegInTop_4_15[2] , \wRegOut_5_1[7] , \ScanLink29[3] , 
        \ScanLink1[19] , \ScanLink0[20] , \wRegInBot_3_2[31] , 
        \wRegInBot_3_2[28] , \wRegOut_4_3[25] , \wRegInTop_5_0[31] , 
        \wRegInTop_5_0[28] , \wRegOut_1_0[0] , \wRegEnBot_2_0[0] , 
        \wRegOut_3_2[0] , \wRegInTop_4_4[8] , \wRegInTop_5_19[25] , 
        \wRegInBot_2_0[7] , \wRegOut_3_0[20] , \ScanLink19[22] , 
        \wRegInTop_4_4[27] , \wRegOut_5_2[4] , \ScanLink9[6] , 
        \wRegOut_4_8[30] , \wRegOut_4_8[29] , \wRegOut_5_21[17] , 
        \ScanLink56[6] , \wRegOut_5_17[12] , \wRegInTop_5_12[29] , 
        \ScanLink55[5] , \wRegInBot_4_0[3] , \wRegInTop_4_1[5] , 
        \wRegInTop_5_12[30] , \wRegOut_5_17[21] , \wRegInTop_5_31[18] , 
        \ScanLink32[2] , \wRegOut_5_20[2] , \wRegOut_5_7[9] , 
        \wRegOut_5_21[24] , \ScanLink4[22] , \ScanLink4[11] , 
        \wRegInTop_2_1[1] , \wRegInTop_2_2[2] , \wRegInBot_2_3[4] , 
        \wRegOut_3_0[13] , \wRegInTop_4_2[6] , \ScanLink19[11] , 
        \wRegInTop_4_4[14] , \ScanLink31[1] , \wRegOut_5_7[19] , 
        \wRegOut_5_23[1] , \wRegInBot_4_3[0] , \wRegInBot_2_2[25] , 
        \wRegOut_5_3[31] , \wRegInTop_5_31[9] , \wRegOut_5_3[28] , 
        \wRegInBot_2_2[16] , \wRegOut_3_4[22] , \ScanLink15[7] , 
        \wRegOut_4_9[0] , \ScanLink16[4] , \wRegOut_5_13[10] , 
        \wRegOut_5_30[21] , \wRegOut_5_25[15] , \wRegInTop_4_0[25] , 
        \wRegInTop_5_16[18] , \wRegOut_3_4[11] , \wRegInTop_4_0[16] , 
        \wRegInTop_5_4[19] , \wRegOut_5_13[23] , \wRegOut_5_25[26] , 
        \wRegOut_5_30[12] , \wRegInTop_5_9[2] , \wRegInTop_3_3[13] , 
        \ScanLink13[9] , \wRegInTop_4_13[24] , \wRegInTop_5_13[1] , 
        \wRegInBot_4_13[23] , \wRegOut_5_8[17] , \wRegInTop_5_10[2] , 
        \wRegInBot_3_6[19] , \wRegOut_4_7[14] , \wRegInTop_4_13[17] , 
        \wRegInBot_4_13[10] , \wRegOut_5_8[24] , \wRegInTop_3_3[20] , 
        \wRegOut_4_7[27] , \wRegInBot_4_4[16] , \ScanLink20[30] , 
        \ScanLink20[29] , \wRegOut_5_12[30] , \ScanLink55[19] , 
        \wRegOut_5_31[18] , \wRegOut_5_12[29] , \wRegOut_5_2[11] , 
        \wRegInTop_5_17[12] , \wRegInTop_5_21[17] , \wRegInBot_1_0[24] , 
        \wRegInBot_3_0[8] , \wRegOut_3_5[31] , \ScanLink61[9] , 
        \wRegOut_3_5[28] , \wRegInBot_4_4[25] , \wRegOut_4_7[6] , 
        \ScanLink18[2] , \wRegOut_4_4[5] , \wRegEnTop_5_4[0] , 
        \wRegOut_5_2[22] , \wRegInTop_5_2[9] , \wRegInTop_5_21[24] , 
        \ScanLink21[23] , \wRegInTop_5_17[21] , \wRegInBot_1_0[17] , 
        \wRegOut_2_1[27] , \ScanLink5[28] , \wRegInBot_3_7[20] , 
        \ScanLink17[26] , \ScanLink54[13] , \wRegInBot_4_15[0] , 
        \ScanLink34[17] , \ScanLink62[16] , \ScanLink41[27] , 
        \wRegOut_5_19[16] , \ScanLink5[31] , \wRegInTop_3_2[19] , 
        \wRegInTop_5_5[20] , \wRegInBot_3_6[6] , \wRegInTop_3_7[0] , 
        \wRegInBot_3_7[13] , \wRegOut_5_19[25] , \ScanLink62[25] , 
        \ScanLink17[15] , \wRegOut_4_1[8] , \ScanLink34[24] , \ScanLink41[14] , 
        \wRegOut_5_12[0] , \ScanLink54[20] , \wRegOut_2_1[14] , 
        \wRegInTop_3_4[3] , \ScanLink21[10] , \wRegInTop_5_7[4] , 
        \wRegInBot_3_5[5] , \wRegInBot_4_12[30] , \wRegInBot_4_12[29] , 
        \wRegInTop_5_4[7] , \wRegOut_5_11[3] , \wRegInTop_5_5[13] , 
        \wRegInBot_3_3[22] , \wRegInTop_3_6[31] , \ScanLink27[5] , 
        \wRegOut_4_14[3] , \wRegInTop_5_1[22] , \wRegInTop_3_6[28] , 
        \ScanLink39[9] , \ScanLink13[24] , \wRegOut_4_13[24] , \ScanLink24[6] , 
        \ScanLink30[15] , \ScanLink45[25] , \ScanLink25[21] , \ScanLink50[11] , 
        \wRegInTop_2_2[27] , \wRegInTop_2_2[14] , \wRegInBot_3_3[11] , 
        \ScanLink13[17] , \ScanLink25[12] , \wRegInTop_5_1[11] , 
        \ScanLink40[2] , \ScanLink43[1] , \ScanLink50[22] , \wRegOut_4_13[17] , 
        \ScanLink30[26] , \ScanLink45[16] , \wRegOut_5_6[13] , 
        \wRegInTop_5_21[3] , \wRegInTop_5_25[15] , \wRegOut_3_1[19] , 
        \wRegInBot_4_0[14] , \wRegInTop_5_13[10] , \wRegInTop_5_30[21] , 
        \ScanLink22[8] , \wRegOut_5_30[8] , \wRegOut_4_9[10] , 
        \wRegInTop_5_22[0] , \wRegInTop_5_30[12] , \wRegOut_5_6[20] , 
        \wRegInTop_5_13[23] , \ScanLink58[0] , \wRegInTop_5_25[26] , 
        \wRegOut_0_0[6] , \wRegInBot_0_0[30] , \ScanLink4[3] , 
        \wRegInBot_0_0[29] , \wRegInBot_0_0[20] , \wRegOut_1_0[9] , 
        \wRegOut_2_1[5] , \ScanLink7[0] , \wRegInTop_3_2[10] , 
        \wRegInBot_4_0[27] , \ScanLink18[31] , \ScanLink18[28] , 
        \wRegOut_4_9[23] , \wRegOut_5_16[18] , \wRegOut_4_6[17] , 
        \ScanLink21[19] , \ScanLink54[29] , \wRegOut_5_12[9] , \ScanLink5[21] , 
        \ScanLink5[12] , \wRegOut_2_2[6] , \wRegInTop_3_7[9] , 
        \ScanLink54[30] , \wRegOut_4_1[1] , \wRegEnTop_3_1[0] , 
        \wRegInBot_4_12[20] , \wRegOut_5_9[14] , \wRegOut_4_2[2] , 
        \wRegInTop_4_12[27] , \wRegInTop_3_2[23] , \wRegInBot_4_15[9] , 
        \wRegInBot_3_7[30] , \wRegInBot_3_7[29] , \wRegOut_4_6[24] , 
        \wRegInTop_5_5[30] , \wRegInTop_5_5[29] , \wRegInBot_2_3[26] , 
        \wRegInBot_3_0[1] , \wRegInTop_3_1[7] , \wRegOut_3_5[21] , 
        \wRegInTop_4_1[26] , \wRegInTop_4_12[14] , \wRegInBot_4_12[13] , 
        \wRegOut_5_9[27] , \wRegInTop_5_1[3] , \wRegOut_5_14[7] , 
        \wRegOut_5_24[16] , \wRegOut_5_31[22] , \wRegOut_5_12[13] , 
        \wRegInTop_3_2[4] , \wRegInTop_5_2[0] , \wRegOut_5_17[4] , 
        \wRegInBot_3_3[2] , \wRegInTop_5_17[31] , \wRegInTop_5_17[28] , 
        \wRegInBot_2_3[15] , \wRegOut_3_5[12] , \wRegInBot_4_13[7] , 
        \wRegInTop_5_18[3] , \wRegOut_5_31[11] , \wRegOut_5_12[20] , 
        \ScanLink62[3] , \wRegOut_5_24[25] , \wRegInTop_4_1[15] , 
        \wRegEnTop_4_10[0] , \wRegInBot_4_10[4] , \wRegOut_5_2[18] , 
        \ScanLink61[0] , \wRegOut_5_6[30] , \wRegOut_5_6[29] , \ScanLink58[9] , 
        \wRegInBot_0_0[13] , \ScanLink7[9] , \ScanLink45[6] , 
        \wRegOut_5_16[11] , \wRegOut_3_1[23] , \ScanLink46[5] , 
        \wRegOut_5_20[14] , \ScanLink18[21] , \wRegInTop_4_5[24] , 
        \wRegEnTop_5_15[0] , \ScanLink21[2] , \ScanLink1[23] , \ScanLink1[10] , 
        \wRegOut_3_1[10] , \ScanLink18[12] , \wRegOut_4_12[4] , 
        \wRegOut_5_9[6] , \wRegInTop_5_30[28] , \wRegInTop_5_13[19] , 
        \wRegInTop_5_30[31] , \wRegInTop_4_5[17] , \ScanLink22[1] , 
        \wRegOut_4_11[7] , \wRegOut_5_20[27] , \wRegInTop_5_22[9] , 
        \wRegOut_5_30[1] , \wRegOut_4_9[19] , \wRegOut_5_16[22] , 
        \wRegInTop_5_1[18] , \ScanLink1[7] , \ScanLink2[4] , 
        \wRegInTop_5_18[15] , \wRegInTop_1_1[16] , \ScanLink43[8] , 
        \wRegInBot_3_3[18] , \wRegInTop_3_6[12] , \wRegOut_4_2[15] , 
        \wRegInTop_5_18[26] , \wRegInTop_5_27[4] , \wRegInTop_1_1[25] , 
        \wRegInTop_3_6[21] , \wRegOut_4_2[26] , \wRegInBot_4_8[2] , 
        \wRegInTop_4_9[4] , \wRegOut_5_28[3] , \ScanLink25[31] , 
        \ScanLink25[28] , \ScanLink39[0] , \ScanLink50[18] , 
        \wRegInTop_5_24[7] , \wRegInTop_2_1[8] , \wRegInTop_4_13[5] , 
        \wRegOut_5_7[0] , \wRegInTop_2_3[17] , \wRegOut_3_7[4] , 
        \wRegEnBot_4_5[0] , \wRegOut_5_17[28] , \wRegInBot_4_1[17] , 
        \ScanLink19[18] , \wRegOut_4_8[13] , \wRegOut_5_17[31] , 
        \wRegInTop_5_12[13] , \wRegOut_3_0[30] , \wRegOut_3_0[29] , 
        \wRegOut_3_4[7] , \wRegInBot_4_3[9] , \wRegInTop_4_10[6] , 
        \wRegOut_5_4[3] , \wRegOut_5_7[10] , \wRegInTop_5_24[16] , 
        \wRegInTop_5_31[22] , \ScanLink31[8] , \wRegInTop_5_31[0] , 
        \wRegOut_5_23[8] , \wRegInBot_4_1[24] , \wRegOut_4_8[20] , 
        \ScanLink0[30] , \wRegInTop_2_3[24] , \wRegOut_5_7[23] , 
        \wRegInTop_5_24[25] , \wRegInTop_5_12[20] , \wRegInTop_5_31[11] , 
        \wRegInBot_3_2[21] , \ScanLink12[27] , \ScanLink24[22] , 
        \ScanLink48[3] , \ScanLink31[16] , \ScanLink51[12] , \ScanLink34[5] , 
        \ScanLink44[26] , \wRegOut_5_26[5] , \wRegInBot_4_6[4] , 
        \wRegInTop_4_7[2] , \wRegOut_4_12[27] , \wRegInTop_5_29[2] , 
        \ScanLink0[29] , \wRegInTop_1_0[4] , \wRegInBot_1_1[2] , 
        \wRegOut_3_2[9] , \wRegInTop_4_4[1] , \wRegInTop_5_0[21] , 
        \wRegInBot_3_2[12] , \wRegInTop_3_7[18] , \wRegInBot_4_5[7] , 
        \ScanLink37[6] , \wRegOut_5_25[6] , \wRegOut_4_12[14] , 
        \ScanLink12[14] , \ScanLink31[25] , \ScanLink44[15] , \ScanLink24[11] , 
        \ScanLink50[1] , \ScanLink51[21] , \wRegInBot_1_1[27] , 
        \wRegOut_2_0[24] , \wRegInBot_4_13[19] , \wRegInTop_5_0[12] , 
        \ScanLink53[2] , \wEnable_1[0] , \wRegInTop_5_4[23] , 
        \wRegInTop_3_3[30] , \wRegInTop_3_3[29] , \wRegInBot_3_6[23] , 
        \ScanLink16[25] , \ScanLink35[14] , \wRegOut_5_18[15] , 
        \ScanLink40[24] , \ScanLink20[20] , \ScanLink63[15] , 
        \wRegOut_2_0[17] , \ScanLink55[10] , \ScanLink4[18] , 
        \wRegInTop_5_4[10] , \wRegInBot_1_1[14] , \ScanLink10[3] , 
        \ScanLink13[0] , \wRegInTop_5_13[8] , \ScanLink55[23] , 
        \wRegInTop_2_2[10] , \wRegOut_3_4[18] , \wRegInBot_3_6[10] , 
        \ScanLink16[16] , \ScanLink20[13] , \ScanLink35[27] , \ScanLink40[17] , 
        \ScanLink63[26] , \wRegOut_5_18[26] , \wRegInBot_4_5[15] , 
        \wRegOut_5_3[12] , \wRegInTop_5_20[14] , \wRegInTop_5_16[11] , 
        \wRegInBot_4_0[10] , \wRegInBot_4_5[26] , \wRegOut_4_9[9] , 
        \wRegOut_5_3[21] , \wRegInTop_5_16[22] , \wRegInTop_5_20[27] , 
        \wRegOut_5_13[19] , \wRegInTop_5_15[6] , \wRegInTop_5_16[5] , 
        \wRegOut_5_30[31] , \wRegOut_5_19[2] , \wRegOut_5_30[28] , 
        \wRegOut_4_9[14] , \wRegInTop_5_22[4] , \wRegInTop_5_13[14] , 
        \ScanLink7[4] , \wRegInBot_4_0[23] , \wRegOut_4_12[9] , 
        \wRegOut_5_6[17] , \wRegInTop_5_25[11] , \wRegInTop_5_30[25] , 
        \wRegInTop_5_21[7] , \wRegInTop_4_5[30] , \wRegInTop_4_5[29] , 
        \wRegOut_4_9[27] , \ScanLink46[8] , \wRegOut_5_20[19] , \ScanLink4[7] , 
        \wRegInTop_2_2[23] , \wRegOut_5_6[24] , \wRegInTop_5_25[22] , 
        \wRegInTop_5_13[27] , \wRegInTop_5_30[16] , \ScanLink58[4] , 
        \ScanLink0[17] , \ScanEnable[0] , \wRegOut_1_0[4] , 
        \wRegInBot_1_0[20] , \ScanLink2[9] , \wRegInTop_1_1[31] , 
        \ScanLink25[25] , \ScanLink30[11] , \ScanLink50[15] , 
        \wRegInTop_1_1[28] , \ScanLink13[20] , \ScanLink24[2] , 
        \ScanLink45[21] , \wRegInBot_3_3[26] , \wRegInBot_3_3[15] , 
        \wRegInTop_4_9[9] , \wRegOut_4_13[20] , \ScanLink27[1] , 
        \wRegInTop_5_1[26] , \wRegInTop_5_27[9] , \wRegOut_4_13[13] , 
        \wRegOut_4_14[7] , \ScanLink13[13] , \wRegOut_4_2[18] , 
        \ScanLink30[22] , \ScanLink45[12] , \ScanLink25[16] , \ScanLink40[6] , 
        \ScanLink50[26] , \ScanLink43[5] , \wRegInTop_5_18[18] , 
        \wRegOut_2_1[23] , \wRegInTop_4_12[19] , \wRegInTop_5_1[15] , 
        \wRegEnTop_5_10[0] , \wRegEnTop_4_15[0] , \wRegInTop_5_5[24] , 
        \wRegInBot_3_7[24] , \wRegOut_4_6[29] , \ScanLink17[22] , 
        \wRegOut_4_6[30] , \wRegOut_5_19[12] , \wRegInBot_4_15[4] , 
        \ScanLink34[13] , \ScanLink41[23] , \ScanLink21[27] , \ScanLink62[12] , 
        \wRegInBot_1_0[13] , \wRegOut_2_1[10] , \ScanLink54[17] , 
        \wRegOut_2_1[8] , \wRegInTop_3_4[7] , \wRegInTop_5_4[3] , 
        \wRegInTop_5_5[17] , \wRegOut_5_11[7] , \wRegOut_5_9[19] , 
        \wRegInBot_3_5[1] , \wRegInTop_5_7[0] , \ScanLink54[24] , 
        \wRegInBot_3_6[2] , \wRegInTop_3_7[4] , \ScanLink21[14] , 
        \wRegOut_5_12[4] , \ScanLink34[20] , \ScanLink41[10] , 
        \ScanLink62[21] , \ScanLink17[11] , \wRegInBot_3_7[17] , 
        \wRegOut_5_19[21] , \wRegInBot_4_10[9] , \wRegInBot_1_1[19] , 
        \wRegInBot_2_3[18] , \wRegInTop_5_21[13] , \wRegInTop_3_2[9] , 
        \wRegInTop_4_1[18] , \wRegInBot_4_4[12] , \wRegOut_5_2[15] , 
        \wRegInTop_5_17[16] , \ScanLink18[6] , \wRegInTop_5_17[25] , 
        \wRegOut_5_24[31] , \wRegOut_5_24[28] , \wRegOut_5_2[26] , 
        \wRegInTop_5_21[20] , \wRegOut_5_17[9] , \wRegInTop_3_3[17] , 
        \wRegEnTop_3_4[0] , \wRegOut_4_4[1] , \wRegInBot_4_4[21] , 
        \wRegOut_4_7[2] , \wRegOut_4_7[10] , \wRegOut_2_0[30] , 
        \wRegOut_2_0[29] , \ScanLink4[26] , \ScanLink4[15] , 
        \wRegInTop_4_13[20] , \wRegInBot_4_13[27] , \wRegOut_5_8[13] , 
        \wRegInTop_5_10[6] , \wRegInTop_5_9[6] , \wRegInTop_5_13[5] , 
        \wRegInTop_3_3[24] , \ScanLink16[31] , \ScanLink16[28] , 
        \ScanLink35[19] , \ScanLink40[30] , \ScanLink63[18] , \ScanLink40[29] , 
        \wRegOut_4_7[23] , \wRegOut_5_18[18] , \wRegOut_3_4[26] , 
        \wRegInTop_4_0[21] , \wRegInTop_4_13[13] , \wRegInBot_4_13[14] , 
        \wRegOut_5_8[20] , \ScanLink15[3] , \ScanLink16[0] , 
        \wRegOut_5_13[14] , \wRegOut_5_25[11] , \wRegOut_5_30[25] , 
        \wRegInTop_5_16[8] , \wRegInBot_2_0[3] , \wRegInTop_2_2[6] , 
        \wRegInBot_2_2[21] , \wRegInBot_2_2[12] , \wRegOut_3_4[15] , 
        \wRegInBot_4_5[18] , \wRegOut_4_9[4] , \wRegOut_5_13[27] , 
        \wRegOut_5_30[16] , \wRegOut_5_25[22] , \wEnable_4[0] , 
        \wRegInTop_4_0[12] , \wRegInTop_2_3[30] , \wRegInTop_2_3[29] , 
        \wRegInTop_5_20[19] , \wRegInTop_5_24[31] , \wRegInTop_5_24[28] , 
        \ScanLink9[2] , \wRegInBot_2_3[0] , \wRegOut_3_0[24] , 
        \wRegInBot_4_1[30] , \wRegOut_5_17[16] , \ScanLink55[1] , 
        \wRegOut_5_21[13] , \ScanLink56[2] , \wRegInBot_4_1[29] , 
        \ScanLink19[26] , \wRegInTop_4_4[23] , \wRegOut_3_0[17] , 
        \wRegInTop_4_2[2] , \wRegInBot_4_3[4] , \ScanLink19[15] , 
        \ScanLink31[5] , \wRegOut_5_23[5] , \wRegInTop_4_4[10] , 
        \wRegInTop_2_1[5] , \wRegInTop_4_13[8] , \wRegOut_3_7[9] , 
        \wRegInTop_4_1[1] , \ScanLink32[6] , \wRegOut_5_20[6] , 
        \wRegOut_5_21[20] , \wRegOut_5_17[25] , \wRegInBot_4_0[7] , 
        \wRegInTop_1_0[11] , \wRegInTop_1_0[9] , \wRegInTop_5_19[12] , 
        \ScanLink12[19] , \ScanLink31[31] , \ScanLink31[28] , \ScanLink44[18] , 
        \ScanLink0[24] , \wRegOut_3_2[4] , \wRegInTop_3_7[15] , 
        \wRegOut_4_3[12] , \wRegOut_4_12[19] , \wRegOut_5_2[0] , 
        \wRegInTop_5_19[21] , \wRegEnBot_4_0[0] , \wRegOut_4_3[21] , 
        \wRegInTop_1_0[22] , \wRegInTop_3_7[26] , \ScanLink29[7] , 
        \wRegInTop_4_15[6] , \wRegOut_5_1[3] , \wRegInBot_1_1[23] , 
        \wRegInBot_2_2[31] , \wRegInBot_2_2[28] , \wRegOut_3_1[7] , 
        \wRegInBot_4_6[9] , \wRegInTop_4_0[31] , \wRegInBot_4_5[22] , 
        \wRegInBot_4_5[11] , \ScanLink34[8] , \wRegOut_5_26[8] , 
        \wRegOut_5_3[16] , \wRegInTop_5_16[15] , \wRegInTop_5_20[10] , 
        \wRegInTop_4_0[28] , \ScanLink16[9] , \wRegInTop_5_16[1] , 
        \wRegOut_5_19[6] , \wRegOut_5_3[25] , \wRegInTop_5_15[2] , 
        \wRegOut_5_25[18] , \ScanLink20[24] , \wRegInTop_5_16[26] , 
        \wRegInTop_5_20[23] , \wRegInBot_1_1[10] , \wRegOut_2_0[20] , 
        \wRegInBot_3_6[27] , \ScanLink16[21] , \ScanLink55[14] , 
        \ScanLink35[10] , \ScanLink63[11] , \ScanLink40[20] , 
        \wRegOut_5_18[11] , \ScanLink10[7] , \wRegInBot_3_6[14] , 
        \wRegInTop_5_4[27] , \wRegOut_5_8[30] , \wRegOut_5_8[29] , 
        \wRegOut_5_18[22] , \ScanLink16[12] , \wRegOut_4_7[19] , 
        \ScanLink63[22] , \ScanLink35[23] , \ScanLink40[13] , \ScanLink55[27] , 
        \wRegOut_2_0[13] , \ScanLink13[4] , \ScanLink20[17] , 
        \wRegInTop_4_13[30] , \wRegInTop_4_13[29] , \wRegInTop_5_4[14] , 
        \wRegInTop_4_4[5] , \ScanLink37[2] , \wRegInTop_5_19[31] , 
        \wRegInTop_5_19[28] , \wRegOut_5_25[2] , \wRegInBot_4_5[3] , 
        \wRegInTop_5_0[25] , \wRegOut_5_2[9] , \wRegOut_0_0[2] , 
        \wRegInTop_1_0[18] , \wRegInTop_1_0[0] , \wRegInBot_1_1[6] , 
        \wRegInBot_3_2[25] , \wRegOut_4_3[31] , \wRegOut_4_3[28] , 
        \ScanLink12[23] , \wRegOut_4_12[23] , \wRegInTop_5_29[6] , 
        \wRegInBot_4_6[0] , \wRegInTop_4_7[6] , \ScanLink24[26] , 
        \ScanLink31[12] , \ScanLink34[1] , \ScanLink44[22] , \wRegOut_5_26[1] , 
        \wRegInTop_5_0[16] , \ScanLink51[16] , \ScanLink24[15] , 
        \ScanLink50[5] , \ScanLink51[25] , \ScanLink53[6] , 
        \wRegInTop_2_3[20] , \wRegInTop_2_3[13] , \wRegInBot_2_3[9] , 
        \wRegInBot_3_2[16] , \ScanLink12[10] , \wRegOut_4_12[10] , 
        \ScanLink31[21] , \ScanLink44[11] , \wRegOut_3_4[3] , 
        \wRegInTop_4_10[2] , \wRegOut_5_4[7] , \wRegOut_5_7[14] , 
        \wRegInTop_5_31[4] , \wRegInTop_5_24[12] , \wRegOut_3_7[0] , 
        \wRegInTop_4_1[8] , \wRegInBot_4_1[13] , \wRegInTop_5_12[17] , 
        \wRegInTop_5_31[26] , \wRegInTop_4_4[19] , \wRegOut_4_8[17] , 
        \wRegInTop_4_13[1] , \wRegOut_5_7[4] , \wRegOut_5_21[30] , 
        \wRegOut_5_21[29] , \wRegInTop_5_31[15] , \wRegOut_5_7[27] , 
        \wRegInTop_5_12[24] , \ScanLink48[7] , \ScanLink55[8] , 
        \wRegInTop_5_24[21] , \ScanLink1[27] , \ScanLink1[14] , \ScanLink1[3] , 
        \wRegInTop_3_6[16] , \wRegInBot_4_1[20] , \wRegOut_4_8[24] , 
        \wRegOut_4_2[11] , \ScanLink2[0] , \wRegInTop_1_1[12] , 
        \wRegInTop_5_18[11] , \wRegInTop_1_1[21] , \ScanLink13[30] , 
        \ScanLink30[18] , \ScanLink13[29] , \ScanLink45[28] , \ScanLink45[31] , 
        \wRegInTop_3_6[25] , \wRegInTop_5_24[3] , \wRegOut_4_2[22] , 
        \wRegOut_4_13[29] , \ScanLink39[4] , \wRegInBot_4_8[6] , 
        \wRegInTop_4_9[0] , \wRegOut_4_13[30] , \wRegOut_5_28[7] , 
        \wRegOut_3_1[27] , \ScanLink18[25] , \wRegInTop_4_5[20] , 
        \ScanLink27[8] , \wRegInTop_5_18[22] , \wRegInTop_5_27[0] , 
        \ScanLink46[1] , \wRegOut_5_16[15] , \wRegOut_5_20[10] , 
        \wRegInBot_0_0[26] , \wRegInBot_0_0[24] , \ScanLink45[2] , 
        \wRegInBot_0_0[17] , \wRegInTop_2_2[19] , \wRegOut_3_1[14] , 
        \wRegInBot_4_0[19] , \ScanLink22[5] , \wRegOut_4_11[3] , 
        \wRegOut_5_16[26] , \wRegOut_5_30[5] , \wRegOut_5_20[23] , 
        \ScanLink18[16] , \wRegInTop_4_5[13] , \wRegOut_5_9[2] , 
        \wRegInTop_5_25[18] , \ScanLink21[6] , \wRegOut_4_12[0] , 
        \ScanLink1[25] , \ScanLink1[16] , \wRegInBot_1_0[30] , 
        \wRegOut_2_1[19] , \wRegInBot_2_3[22] , \wRegInTop_5_21[30] , 
        \wRegInTop_5_21[29] , \wRegInBot_2_3[11] , \wRegInBot_3_0[5] , 
        \wRegInTop_3_1[3] , \wRegInTop_3_2[0] , \wRegInTop_5_18[7] , 
        \wRegInBot_3_3[6] , \wRegOut_4_4[8] , \wRegInTop_5_2[4] , 
        \wRegOut_5_17[0] , \wRegOut_5_12[17] , \wRegOut_3_5[25] , 
        \wRegInTop_5_1[7] , \wRegOut_5_14[3] , \wRegOut_5_31[26] , 
        \wRegOut_5_24[12] , \wRegInTop_4_1[22] , \wRegInBot_4_4[31] , 
        \wRegInBot_4_4[28] , \wRegInBot_4_10[0] , \ScanLink61[4] , 
        \wRegOut_3_5[16] , \wRegInTop_4_1[11] , \wRegInBot_4_13[3] , 
        \wRegOut_5_12[24] , \wRegOut_5_24[21] , \wRegOut_5_31[15] , 
        \ScanLink62[7] , \wRegOut_2_1[1] , \ScanLink5[16] , \wRegOut_2_2[2] , 
        \wRegInBot_3_5[8] , \wRegOut_4_2[6] , \wRegInTop_4_12[23] , 
        \wRegOut_4_1[5] , \ScanLink17[18] , \wRegInBot_4_12[24] , 
        \wRegOut_5_9[10] , \wRegEnTop_5_1[0] , \ScanLink34[29] , 
        \ScanLink41[19] , \ScanLink62[31] , \ScanLink62[28] , \ScanLink34[30] , 
        \ScanLink5[25] , \wRegInTop_3_2[14] , \wRegInTop_5_7[9] , 
        \wRegOut_4_6[13] , \wRegOut_5_19[28] , \wRegInTop_4_12[10] , 
        \wRegInBot_4_12[17] , \wRegOut_5_9[23] , \wRegOut_5_19[31] , 
        \wRegEnTop_5_29[0] , \wRegInTop_3_2[27] , \wRegOut_4_6[20] , 
        \wRegInBot_1_0[29] , \ScanLink1[1] , \ScanLink2[2] , 
        \wRegInTop_5_18[13] , \wRegInTop_1_1[10] , \ScanLink13[18] , 
        \ScanLink30[30] , \ScanLink30[29] , \ScanLink45[19] , 
        \wRegInTop_3_6[14] , \wRegOut_4_2[13] , \wRegOut_4_13[18] , 
        \wRegInTop_5_18[20] , \wRegInTop_5_27[2] , \wRegInTop_1_1[23] , 
        \wRegInTop_3_6[27] , \wRegOut_4_2[20] , \wRegInBot_4_8[4] , 
        \wRegInTop_4_9[2] , \wRegOut_5_28[5] , \ScanLink24[9] , 
        \ScanLink39[6] , \wRegInTop_5_24[1] , \wRegInTop_2_2[31] , 
        \wRegInTop_5_25[30] , \wRegInTop_5_25[29] , \wRegInTop_2_2[28] , 
        \wRegInBot_0_0[15] , \wRegOut_3_1[25] , \ScanLink45[0] , 
        \ScanLink46[3] , \wRegOut_5_16[17] , \wRegOut_5_20[12] , 
        \wRegInBot_4_0[31] , \wRegInBot_4_0[28] , \ScanLink18[27] , 
        \wRegInTop_4_5[22] , \ScanLink21[4] , \wRegInTop_1_0[30] , 
        \wRegInTop_1_0[29] , \wRegInBot_1_0[18] , \wRegOut_2_1[3] , 
        \wRegInBot_2_3[20] , \wRegInBot_3_0[7] , \wRegOut_3_1[16] , 
        \ScanLink18[14] , \wRegInTop_4_5[11] , \wRegOut_4_12[2] , 
        \wRegOut_5_9[0] , \wRegOut_3_5[27] , \wRegInTop_4_1[20] , 
        \ScanLink22[7] , \wRegOut_4_11[1] , \wRegOut_5_16[24] , 
        \wRegOut_5_20[21] , \wRegOut_5_30[7] , \wRegInTop_5_1[5] , 
        \wRegOut_5_14[1] , \wRegOut_5_24[10] , \wRegOut_5_12[15] , 
        \wRegInTop_3_1[1] , \wRegOut_4_7[9] , \wRegInTop_3_2[2] , 
        \wRegInBot_3_3[4] , \wRegInTop_5_2[6] , \wRegOut_5_31[24] , 
        \wRegOut_5_17[2] , \wRegInTop_5_18[5] , \wRegInBot_2_3[13] , 
        \wRegOut_3_5[14] , \wRegInBot_4_4[19] , \wRegInBot_4_13[1] , 
        \wRegOut_5_12[26] , \ScanLink62[5] , \wRegOut_5_31[17] , 
        \wRegOut_5_24[23] , \wRegEnTop_5_31[0] , \wRegInTop_4_1[13] , 
        \wRegInTop_5_21[18] , \wRegInTop_3_2[16] , \wRegOut_4_6[11] , 
        \wRegInBot_4_10[2] , \ScanLink61[6] , \wRegInBot_1_1[21] , 
        \wRegOut_2_0[22] , \wRegOut_2_1[31] , \ScanLink5[14] , 
        \wRegOut_2_2[0] , \wRegInBot_3_6[9] , \wRegOut_4_1[7] , 
        \wRegInBot_4_12[26] , \wRegInTop_5_4[8] , \wRegOut_5_9[12] , 
        \wRegEnBot_3_0[0] , \wRegOut_4_2[4] , \wRegInTop_4_12[21] , 
        \wRegInTop_3_2[25] , \ScanLink17[30] , \ScanLink41[28] , 
        \ScanLink17[29] , \ScanLink34[18] , \ScanLink41[31] , \ScanLink62[19] , 
        \wRegOut_4_6[22] , \wRegOut_5_19[19] , \wRegOut_2_1[28] , 
        \ScanLink5[27] , \wRegInBot_2_2[19] , \wRegInTop_4_12[12] , 
        \wRegInBot_4_12[15] , \wRegOut_5_9[21] , \ScanLink15[8] , 
        \wRegInTop_4_0[19] , \wRegInBot_4_5[13] , \wRegOut_5_3[14] , 
        \wRegInTop_5_16[17] , \wRegInTop_5_20[12] , \wRegOut_5_3[27] , 
        \wRegInTop_5_16[24] , \wRegOut_5_25[30] , \wRegOut_5_25[29] , 
        \wRegInTop_5_20[21] , \wRegInBot_4_5[20] , \wRegInTop_5_15[0] , 
        \wRegInTop_5_16[3] , \wRegOut_5_19[4] , \wRegInTop_4_13[18] , 
        \wRegInTop_5_4[25] , \wRegInBot_3_6[25] , \wRegOut_4_7[31] , 
        \wRegOut_4_7[28] , \wRegOut_5_18[13] , \ScanLink16[23] , 
        \ScanLink63[13] , \ScanLink35[12] , \ScanLink40[22] , \ScanLink55[16] , 
        \wRegInBot_1_1[12] , \wRegOut_2_0[11] , \ScanLink20[26] , 
        \ScanLink10[5] , \ScanLink13[6] , \wRegInTop_5_4[16] , 
        \wRegOut_5_8[18] , \ScanLink20[15] , \wRegInBot_3_6[16] , 
        \ScanLink16[10] , \ScanLink55[25] , \ScanLink35[21] , \ScanLink63[20] , 
        \ScanLink40[11] , \ScanLink24[24] , \wRegOut_5_18[20] , 
        \ScanLink51[14] , \wRegOut_5_1[8] , \ScanLink12[21] , 
        \wRegInBot_4_6[2] , \wRegInTop_4_7[4] , \ScanLink44[20] , 
        \wRegOut_5_26[3] , \wRegInBot_3_2[27] , \wRegOut_4_12[21] , 
        \ScanLink31[10] , \ScanLink34[3] , \wRegInTop_5_29[4] , 
        \wRegInTop_4_4[7] , \wRegInBot_4_5[1] , \wRegInTop_5_0[27] , 
        \ScanLink37[0] , \wRegOut_5_25[0] , \wRegOut_0_0[9] , \wRegOut_0_0[0] , 
        \wRegInTop_1_0[2] , \wRegInBot_3_2[14] , \ScanLink12[12] , 
        \wRegOut_4_3[19] , \wRegOut_4_12[12] , \ScanLink24[17] , 
        \ScanLink31[23] , \ScanLink44[13] , \ScanLink50[7] , 
        \wRegInTop_5_19[19] , \ScanLink51[27] , \wRegInBot_1_1[4] , 
        \ScanLink53[4] , \wRegInBot_2_0[8] , \wRegInTop_4_13[3] , 
        \wRegInTop_5_0[14] , \wRegInTop_2_3[11] , \wRegOut_3_7[2] , 
        \wRegOut_4_8[15] , \wRegOut_5_7[6] , \wRegInBot_4_1[11] , 
        \wRegEnTop_4_4[0] , \wRegInTop_5_31[24] , \wRegOut_3_4[1] , 
        \wRegInTop_4_10[0] , \wRegOut_5_7[16] , \wRegInTop_5_12[15] , 
        \wRegInTop_5_24[10] , \wRegInTop_5_31[6] , \wRegOut_5_4[5] , 
        \wRegInBot_4_1[22] , \wRegInTop_4_2[9] , \wRegInTop_4_4[31] , 
        \wRegInTop_4_4[28] , \wRegOut_4_8[26] , \wRegOut_5_21[18] , 
        \ScanLink56[9] , \wRegInBot_1_1[31] , \wRegInBot_1_1[28] , 
        \wRegOut_2_0[18] , \ScanLink4[17] , \wRegInTop_2_3[22] , 
        \wRegOut_5_7[25] , \wRegInTop_5_24[23] , \ScanLink9[9] , 
        \wRegInTop_5_12[26] , \ScanLink48[5] , \wRegInTop_5_31[17] , 
        \wRegInTop_5_9[4] , \ScanLink4[24] , \wRegInTop_3_3[15] , 
        \ScanLink16[19] , \wRegInTop_4_13[22] , \wRegInTop_5_13[7] , 
        \wRegInBot_4_13[25] , \ScanLink35[31] , \wRegOut_5_8[11] , 
        \ScanLink35[28] , \wRegInTop_5_10[4] , \ScanLink63[29] , 
        \ScanLink40[18] , \ScanLink63[30] , \wRegOut_4_7[12] , 
        \wRegOut_5_18[30] , \wRegInTop_4_13[11] , \wRegInBot_4_13[16] , 
        \wRegOut_5_18[29] , \wRegOut_5_8[22] , \wRegInTop_3_3[26] , 
        \wRegOut_4_7[21] , \wRegInBot_2_2[23] , \wRegOut_4_9[6] , 
        \wRegInBot_2_2[10] , \wRegOut_3_4[24] , \ScanLink15[1] , 
        \wRegInTop_5_15[9] , \wRegInTop_5_20[31] , \wRegInTop_5_20[28] , 
        \ScanLink16[2] , \wRegOut_5_13[16] , \wRegOut_5_30[27] , 
        \wCtrlOut_1[0] , \wRegInBot_4_5[30] , \wRegOut_5_25[13] , 
        \wRegInTop_4_0[23] , \wRegInBot_4_5[29] , \wRegEnTop_5_22[0] , 
        \wRegOut_3_0[26] , \wRegOut_3_4[17] , \wRegInTop_4_0[10] , 
        \ScanLink19[24] , \wRegOut_5_13[25] , \wRegOut_5_25[20] , 
        \wRegOut_5_30[14] , \wRegInTop_4_4[21] , \wRegOut_5_17[14] , 
        \wRegOut_5_21[11] , \ScanLink56[0] , \ScanLink55[3] , 
        \wRegInBot_2_0[1] , \wRegInTop_2_1[7] , \ScanLink9[0] , 
        \wRegInBot_4_0[5] , \ScanLink32[4] , \wRegOut_5_20[4] , 
        \wRegInTop_4_1[3] , \wRegOut_5_17[27] , \wRegInTop_2_2[4] , 
        \wRegInTop_2_3[18] , \wRegOut_3_0[15] , \wRegInBot_4_1[18] , 
        \wRegOut_5_21[22] , \ScanLink19[17] , \wRegInTop_4_4[12] , 
        \wRegInTop_5_24[19] , \wRegOut_3_4[8] , \wRegInTop_4_2[0] , 
        \wRegInBot_4_3[6] , \ScanLink31[7] , \wRegOut_5_23[7] , 
        \wRegInBot_2_3[2] , \wRegInTop_4_10[9] , \wRegOut_4_3[10] , 
        \ScanLink0[15] , \wRegInTop_1_0[13] , \wRegInTop_3_7[17] , 
        \wRegInTop_5_19[10] , \wRegInTop_1_0[20] , \wRegOut_3_1[5] , 
        \ScanLink44[30] , \ScanLink12[31] , \ScanLink12[28] , \ScanLink44[29] , 
        \wRegInTop_4_15[4] , \ScanLink31[19] , \wRegOut_5_1[1] , 
        \ScanLink0[26] , \wRegInTop_3_7[24] , \wRegOut_4_3[23] , 
        \wRegOut_4_12[31] , \ScanLink29[5] , \wRegOut_4_12[28] , 
        \wRegEnTop_2_1[0] , \wRegOut_3_2[6] , \wRegInBot_4_5[8] , 
        \wRegEnBot_4_15[0] , \ScanLink37[9] , \wRegOut_5_25[9] , 
        \wRegInTop_5_19[23] , \wRegInTop_2_2[21] , \wRegInTop_2_2[12] , 
        \wRegOut_5_2[2] , \wRegOut_5_6[15] , \wRegInTop_5_21[5] , 
        \wRegInTop_5_25[13] , \wRegOut_5_9[9] , \wRegInTop_5_13[16] , 
        \wRegInTop_5_30[27] , \wRegInBot_4_0[12] , \wRegInTop_4_5[18] , 
        \wRegOut_4_9[16] , \wRegOut_4_11[8] , \wRegInTop_5_13[25] , 
        \wRegOut_5_20[31] , \wRegOut_5_20[28] , \wRegInTop_5_22[6] , 
        \wRegOut_5_6[26] , \wRegInTop_5_25[20] , \ScanLink58[6] , 
        \wRegInTop_5_30[14] , \wRegOut_0_0[4] , \ScanLink1[8] , \ScanLink4[5] , 
        \ScanLink7[6] , \ScanLink45[9] , \wRegInBot_3_3[24] , 
        \wRegInBot_4_0[21] , \wRegOut_4_9[25] , \wRegOut_4_2[29] , 
        \ScanLink27[3] , \wRegInTop_5_18[29] , \wRegOut_4_13[22] , 
        \wRegOut_4_14[5] , \wRegInTop_5_1[24] , \wRegInTop_5_18[30] , 
        \ScanLink13[22] , \wRegOut_4_2[30] , \ScanLink24[0] , \ScanLink45[23] , 
        \ScanLink30[13] , \ScanLink25[27] , \ScanLink50[17] , 
        \wRegInTop_5_24[8] , \wRegInTop_5_1[17] , \ScanLink43[7] , 
        \wRegOut_1_0[6] , \wRegInBot_1_0[22] , \wRegInTop_1_1[19] , 
        \ScanLink13[11] , \ScanLink25[14] , \ScanLink40[4] , \ScanLink30[20] , 
        \ScanLink50[24] , \ScanLink45[10] , \wRegInBot_3_3[17] , 
        \wRegOut_4_13[11] , \ScanLink54[15] , \wRegInBot_1_0[11] , 
        \wRegOut_2_1[21] , \wRegInBot_3_7[26] , \ScanLink17[20] , 
        \ScanLink21[25] , \wRegInBot_4_15[6] , \ScanLink34[11] , 
        \ScanLink41[21] , \ScanLink62[10] , \wRegOut_5_19[10] , 
        \wRegInBot_3_6[0] , \wRegInBot_3_7[15] , \wRegInTop_5_5[26] , 
        \wRegOut_5_9[31] , \wRegOut_5_9[28] , \ScanLink17[13] , 
        \wRegOut_4_6[18] , \ScanLink34[22] , \wRegOut_5_19[23] , 
        \ScanLink41[12] , \wRegInTop_3_7[6] , \ScanLink21[16] , 
        \wRegInTop_5_7[2] , \ScanLink62[23] , \wRegOut_5_12[6] , 
        \wRegOut_2_1[12] , \wRegOut_2_2[9] , \wRegInTop_3_4[5] , 
        \wRegInBot_3_5[3] , \ScanLink54[26] , \wRegInTop_4_12[31] , 
        \wRegInTop_4_12[28] , \wRegInTop_5_4[1] , \wRegOut_5_11[5] , 
        \wRegInTop_5_5[15] , \wRegInBot_4_4[10] , \wRegInBot_4_13[8] , 
        \wRegOut_5_2[17] , \wRegInTop_5_17[14] , \wRegInTop_5_21[11] , 
        \wRegInTop_2_2[9] , \wRegInBot_2_3[30] , \wRegInTop_3_1[8] , 
        \wRegInTop_4_1[30] , \wRegInTop_4_1[29] , \wRegInBot_4_4[23] , 
        \wRegOut_4_7[0] , \wRegOut_4_4[3] , \wRegOut_5_14[8] , 
        \wRegOut_5_24[19] , \wRegInTop_5_21[22] , \wRegInBot_2_3[29] , 
        \wRegOut_5_2[24] , \wRegOut_3_4[5] , \ScanLink18[4] , 
        \wRegInTop_5_17[27] , \wRegInTop_2_3[26] , \wRegInTop_2_3[15] , 
        \wRegInTop_4_10[4] , \wRegInTop_5_31[2] , \wRegOut_5_4[1] , 
        \wRegOut_5_7[12] , \wRegInTop_5_24[14] , \wRegInTop_5_12[11] , 
        \wRegInTop_5_31[20] , \wRegOut_3_0[18] , \wRegInBot_4_1[15] , 
        \wRegOut_3_7[6] , \wRegInBot_4_0[8] , \wRegOut_4_8[11] , 
        \wRegEnBot_4_10[0] , \wRegInTop_4_13[7] , \ScanLink32[9] , 
        \wRegOut_5_20[9] , \wRegOut_5_7[2] , \wRegInTop_5_12[22] , 
        \wRegOut_5_7[21] , \ScanLink48[1] , \wRegInTop_5_24[27] , 
        \wRegInTop_5_31[13] , \ScanLink0[18] , \wRegOut_3_1[8] , 
        \wRegInBot_3_2[23] , \wRegInTop_3_7[30] , \wRegInTop_3_7[29] , 
        \wRegInBot_4_1[26] , \ScanLink19[30] , \wRegOut_4_8[22] , 
        \wRegOut_5_17[19] , \ScanLink19[29] , \wRegInTop_4_4[3] , 
        \wRegInBot_4_5[5] , \wRegInTop_5_0[23] , \ScanLink37[4] , 
        \wRegOut_5_25[4] , \ScanLink29[8] , \wRegOut_4_12[25] , 
        \wRegInTop_5_29[0] , \ScanLink31[14] , \ScanLink34[7] , 
        \ScanLink44[24] , \wRegOut_5_26[7] , \ScanLink12[25] , 
        \wRegInBot_4_6[6] , \wRegInTop_4_7[0] , \ScanLink24[20] , 
        \wRegInTop_4_15[9] , \ScanLink51[10] , \wRegInTop_1_0[6] , 
        \wRegInTop_5_0[10] , \wRegInBot_1_1[25] , \wRegInBot_1_1[0] , 
        \ScanLink53[0] , \wRegInBot_3_2[10] , \ScanLink12[16] , 
        \ScanLink24[13] , \ScanLink50[3] , \ScanLink31[27] , \ScanLink51[23] , 
        \ScanLink44[17] , \wRegOut_4_12[16] , \ScanLink55[12] , 
        \wRegInBot_1_1[16] , \wRegOut_2_0[26] , \ScanLink4[30] , 
        \wRegInBot_3_6[21] , \ScanLink16[27] , \ScanLink20[22] , 
        \ScanLink35[16] , \ScanLink40[26] , \ScanLink63[17] , 
        \wRegOut_5_18[17] , \wRegEnTop_5_27[0] , \ScanLink4[29] , 
        \ScanLink10[1] , \wRegInTop_3_3[18] , \wRegInTop_5_4[21] , 
        \wRegInBot_3_6[12] , \ScanLink16[14] , \ScanLink35[25] , 
        \wRegOut_5_18[24] , \ScanLink40[15] , \wRegInTop_5_10[9] , 
        \ScanLink63[24] , \ScanLink20[11] , \ScanLink13[2] , \ScanLink55[21] , 
        \wRegInBot_4_13[31] , \wRegInBot_0_0[22] , \wRegOut_2_0[15] , 
        \wRegInBot_4_13[28] , \wRegInTop_5_4[12] , \wCtrlOut_4[0] , 
        \wRegInTop_5_9[9] , \ScanLink4[8] , \wRegOut_2_1[7] , \ScanLink5[10] , 
        \wRegOut_3_4[30] , \wRegOut_3_4[29] , \wRegInBot_4_5[17] , 
        \wRegOut_5_13[31] , \wRegOut_5_13[28] , \wRegOut_5_30[19] , 
        \wRegOut_5_3[10] , \wRegInTop_5_16[13] , \wRegInTop_5_20[16] , 
        \wRegInBot_4_5[24] , \wRegOut_5_3[23] , \wRegInTop_5_15[4] , 
        \wRegInTop_5_16[7] , \wRegOut_5_19[0] , \wRegInTop_5_20[25] , 
        \wRegInTop_5_5[18] , \wRegInTop_5_16[20] , \wRegOut_2_2[4] , 
        \wRegInTop_3_4[8] , \wRegOut_4_2[0] , \wRegInTop_4_12[25] , 
        \wRegInBot_4_12[22] , \wRegOut_5_9[16] , \wRegOut_4_1[3] , 
        \wRegOut_5_11[8] , \ScanLink5[23] , \wRegInTop_3_2[12] , 
        \wRegInBot_3_7[18] , \wRegOut_4_6[15] , \wRegInTop_4_12[16] , 
        \wRegInBot_4_12[11] , \wRegOut_5_9[25] , \wRegInBot_2_3[24] , 
        \wRegInTop_3_2[21] , \wRegOut_4_6[26] , \ScanLink21[31] , 
        \ScanLink21[28] , \ScanLink54[18] , \wRegOut_5_2[29] , 
        \wRegInTop_5_18[1] , \wRegInBot_2_3[17] , \wRegInBot_3_0[3] , 
        \wRegInTop_3_2[6] , \wRegInBot_3_3[0] , \ScanLink18[9] , 
        \wRegOut_5_2[30] , \wRegInTop_5_2[2] , \wRegOut_5_17[6] , 
        \wRegOut_5_12[11] , \wRegOut_5_31[20] , \wRegInTop_3_1[5] , 
        \wRegOut_3_5[23] , \wRegInTop_5_1[1] , \wRegOut_5_14[5] , 
        \wRegOut_5_24[14] , \wRegInTop_4_1[24] , \wRegInBot_4_10[6] , 
        \ScanLink61[2] , \wRegInTop_5_17[19] , \wRegOut_3_1[21] , 
        \wRegOut_3_5[10] , \wRegInTop_4_1[17] , \ScanLink18[23] , 
        \wRegInBot_4_13[5] , \wRegOut_5_24[27] , \ScanLink62[1] , 
        \wRegOut_5_31[13] , \wRegOut_5_12[22] , \wRegInTop_4_5[26] , 
        \wRegOut_4_9[31] , \ScanLink46[7] , \wRegOut_5_20[16] , 
        \wRegOut_4_9[28] , \wRegOut_5_16[13] , \ScanLink45[4] , 
        \wRegInBot_0_0[18] , \wRegInBot_0_0[11] , \wRegOut_3_1[12] , 
        \ScanLink22[3] , \wRegOut_4_11[5] , \wRegInTop_5_13[31] , 
        \wRegInTop_5_30[19] , \wRegInTop_5_13[28] , \wRegOut_5_30[3] , 
        \wRegOut_5_16[20] , \wRegOut_5_20[25] , \ScanLink18[10] , 
        \wRegInTop_4_5[15] , \ScanLink21[0] , \wRegOut_5_6[18] , 
        \wRegOut_5_9[4] , \wRegOut_4_12[6] , \ScanLink1[31] , \ScanLink1[28] , 
        \ScanLink1[21] , \ScanLink1[12] , \ScanLink1[5] , \wRegInTop_3_6[10] , 
        \wRegOut_4_2[17] , \wRegInTop_5_21[8] , \ScanLink25[19] , 
        \ScanLink40[9] , \ScanLink50[29] , \ScanLink2[6] , \wRegInTop_1_1[14] , 
        \ScanLink50[30] , \wRegInTop_5_18[17] , \wRegInTop_1_1[27] , 
        \wRegInBot_3_3[30] , \wRegInTop_3_6[23] , \wRegInTop_5_24[5] , 
        \ScanLink39[2] , \wRegInBot_3_3[29] , \wRegOut_4_2[24] , 
        \wRegInBot_4_8[0] , \wRegInTop_5_1[29] , \wRegOut_5_28[1] , 
        \wRegInTop_4_9[6] , \wRegInTop_5_1[30] , \wRegOut_1_0[2] , 
        \wRegOut_4_14[8] , \wRegInTop_5_18[24] , \wRegInTop_5_27[6] , 
        \wRegInBot_1_0[26] , \wRegOut_2_1[25] , \wRegInBot_3_3[9] , 
        \wRegOut_3_5[19] , \wRegInBot_4_4[14] , \wRegOut_5_2[13] , 
        \wRegInTop_5_17[10] , \wRegInTop_5_21[15] , \ScanLink18[0] , 
        \ScanLink62[8] , \wRegOut_4_4[7] , \wRegOut_5_2[20] , 
        \wRegInTop_5_17[23] , \wRegInTop_5_18[8] , \wRegInTop_5_21[26] , 
        \wRegEnBot_3_5[0] , \wRegInTop_5_1[8] , \wRegOut_5_31[29] , 
        \wRegInBot_4_4[27] , \wRegOut_4_7[4] , \wRegOut_5_12[18] , 
        \wRegOut_5_31[30] , \wRegInBot_4_12[18] , \wRegInTop_5_5[22] , 
        \wRegInTop_3_2[31] , \wRegInTop_3_2[28] , \wRegInBot_3_7[22] , 
        \wRegOut_5_19[14] , \ScanLink17[24] , \ScanLink62[14] , 
        \wRegInBot_4_15[2] , \ScanLink34[15] , \ScanLink41[25] , 
        \ScanLink54[11] , \wRegInBot_1_0[15] , \wRegOut_2_1[16] , 
        \ScanLink5[19] , \ScanLink21[21] , \wRegInTop_3_4[1] , 
        \wRegInBot_3_5[7] , \wRegInTop_5_4[5] , \wRegInTop_5_5[11] , 
        \wRegOut_5_11[1] , \wRegOut_4_2[9] , \ScanLink21[12] , 
        \wRegInBot_3_3[20] , \ScanLink13[26] , \wRegInBot_3_6[4] , 
        \ScanLink17[17] , \wRegInTop_5_7[6] , \wRegOut_5_12[2] , 
        \ScanLink54[22] , \wRegInTop_3_7[2] , \wRegInBot_3_7[11] , 
        \ScanLink34[26] , \ScanLink62[27] , \ScanLink41[16] , \ScanLink25[23] , 
        \ScanLink50[13] , \wRegOut_5_19[27] , \ScanLink24[4] , 
        \ScanLink45[27] , \wRegOut_4_13[26] , \ScanLink30[17] , 
        \wRegInTop_2_2[16] , \wRegInBot_3_3[13] , \wRegInTop_3_6[19] , 
        \wRegInBot_4_8[9] , \wRegInTop_5_1[20] , \wRegOut_5_28[8] , 
        \ScanLink27[7] , \wRegOut_4_14[1] , \ScanLink13[15] , 
        \wRegOut_4_13[15] , \wRegInBot_4_0[16] , \ScanLink18[19] , 
        \wRegOut_4_9[12] , \ScanLink25[10] , \ScanLink30[24] , \ScanLink40[0] , 
        \ScanLink45[14] , \wRegInTop_5_1[13] , \ScanLink43[3] , 
        \ScanLink50[20] , \wRegOut_5_16[30] , \wRegInTop_5_22[2] , 
        \wRegOut_5_16[29] , \wRegInTop_5_30[23] , \ScanLink21[9] , 
        \wRegOut_5_6[11] , \wRegInTop_5_13[12] , \wRegInTop_5_21[1] , 
        \wRegInTop_5_25[17] , \ScanLink7[2] , \wRegOut_3_1[31] , 
        \wRegOut_3_1[28] , \wRegInBot_4_0[25] , \wRegOut_4_9[21] , 
        \ScanLink0[11] , \ScanLink4[1] , \wRegInTop_2_2[25] , 
        \wRegOut_5_6[22] , \wRegInTop_5_25[24] , \wRegInTop_5_0[19] , 
        \wRegInTop_5_13[21] , \ScanLink58[2] , \wRegInTop_5_30[10] , 
        \wRegInTop_1_0[17] , \wRegInBot_1_1[9] , \wRegInTop_5_19[14] , 
        \ScanLink53[9] , \wRegInTop_3_7[13] , \ScanLink0[22] , 
        \wRegOut_3_2[2] , \wRegInBot_3_2[19] , \wRegOut_4_3[14] , 
        \wRegOut_5_2[6] , \wRegEnTop_4_1[0] , \wRegInTop_5_19[27] , 
        \wRegInTop_3_7[20] , \wRegOut_4_3[27] , \wRegInTop_5_29[9] , 
        \ScanLink29[1] , \wRegInTop_1_0[24] , \ScanLink24[30] , 
        \wRegInTop_4_15[0] , \wRegOut_5_1[5] , \ScanLink24[29] , 
        \ScanLink51[19] , \wRegInBot_1_0[4] , \ScanLink2[24] , 
        \wRegInBot_2_0[5] , \wRegInTop_2_1[3] , \wRegInTop_2_2[0] , 
        \wRegOut_3_0[22] , \wRegOut_3_1[1] , \ScanLink9[4] , 
        \wRegInTop_4_7[9] , \wRegOut_5_7[31] , \wRegOut_5_7[28] , 
        \ScanLink48[8] , \wRegOut_5_17[10] , \ScanLink55[7] , 
        \wRegOut_5_21[15] , \ScanLink56[4] , \ScanLink19[20] , 
        \wRegInTop_4_4[25] , \wRegInBot_2_3[6] , \wRegOut_5_4[8] , 
        \wRegOut_3_0[11] , \wRegInTop_4_2[4] , \wRegInBot_4_3[2] , 
        \ScanLink31[3] , \wRegOut_5_23[3] , \ScanLink19[13] , 
        \wRegInTop_4_4[16] , \wRegInTop_5_12[18] , \wRegInTop_5_31[30] , 
        \wRegInTop_5_31[29] , \wRegOut_5_21[26] , \ScanLink4[20] , 
        \ScanLink4[13] , \wRegInBot_2_2[27] , \wRegOut_3_4[20] , 
        \wRegInTop_4_0[27] , \wRegInBot_4_0[1] , \wRegInTop_4_1[7] , 
        \wRegOut_4_8[18] , \ScanLink32[0] , \wRegOut_5_17[23] , 
        \wRegOut_5_20[0] , \wRegOut_5_19[9] , \ScanLink15[5] , \ScanLink16[6] , 
        \wRegOut_5_13[12] , \wRegOut_5_25[17] , \wRegOut_5_30[23] , 
        \wRegOut_4_9[2] , \wRegInTop_5_16[30] , \wRegInTop_5_16[29] , 
        \wRegInBot_2_2[14] , \wRegOut_3_4[13] , \wRegOut_5_13[21] , 
        \wRegOut_5_25[24] , \wRegOut_5_30[10] , \wRegInTop_4_0[14] , 
        \ScanLink10[8] , \wRegInTop_3_3[11] , \wRegOut_4_7[16] , 
        \wRegOut_5_3[19] , \ScanLink55[31] , \ScanLink20[18] , 
        \wRegInTop_4_13[26] , \wRegInBot_4_13[21] , \wRegOut_5_8[15] , 
        \wRegInTop_5_10[0] , \ScanLink55[28] , \wRegInTop_5_13[3] , 
        \wRegInTop_5_9[0] , \wRegInTop_3_3[22] , \wRegInBot_3_6[31] , 
        \wRegInBot_3_6[28] , \wRegOut_4_7[25] , \wRegInTop_5_4[31] , 
        \wRegInTop_5_4[28] , \wRegInTop_4_13[15] , \wRegInBot_4_13[12] , 
        \wRegOut_5_8[26] , \wRegInTop_4_15[11] , \wRegInBot_4_15[16] , 
        \wRegInTop_5_17[3] , \wRegOut_5_18[4] , \ScanLink2[17] , 
        \wRegInTop_3_5[26] , \ScanLink14[8] , \wRegOut_4_1[21] , 
        \wRegInBot_4_8[25] , \wRegInTop_5_14[0] , \wRegInTop_1_1[2] , 
        \wRegInTop_2_1[30] , \wRegOut_3_2[17] , \ScanLink10[19] , 
        \wRegInBot_4_8[16] , \wRegInTop_4_15[22] , \wRegInBot_4_15[25] , 
        \ScanLink33[28] , \ScanLink46[18] , \ScanLink11[5] , 
        \wRegInTop_3_5[15] , \wRegOut_4_1[12] , \ScanLink33[31] , 
        \wRegOut_4_10[19] , \wRegInTop_5_9[13] , \ScanLink12[6] , 
        \wRegInTop_4_6[10] , \ScanLink38[24] , \ScanLink58[20] , 
        \wRegOut_5_15[25] , \wRegOut_5_23[20] , \wRegInTop_2_1[29] , 
        \ScanLink9[31] , \wRegInTop_5_9[20] , \wRegInTop_5_26[31] , 
        \wRegInTop_5_26[28] , \ScanLink9[28] , \wRegOut_3_2[24] , 
        \wRegInBot_4_3[29] , \wRegInTop_4_6[23] , \ScanLink38[17] , 
        \wRegOut_5_15[16] , \wRegOut_5_23[13] , \wRegInBot_4_3[30] , 
        \ScanLink58[13] , \wRegOut_5_11[27] , \wRegOut_5_27[22] , 
        \ScanLink52[4] , \wRegOut_1_1[22] , \wRegOut_1_1[11] , 
        \wRegInBot_2_0[12] , \wRegOut_3_6[15] , \wRegInTop_4_2[12] , 
        \ScanLink49[16] , \wRegInBot_4_7[18] , \ScanLink29[12] , 
        \wRegInTop_5_22[19] , \wRegOut_3_6[26] , \ScanLink51[7] , 
        \wRegInTop_4_2[21] , \ScanLink29[21] , \ScanLink49[25] , 
        \wRegOut_5_11[14] , \wRegInBot_2_0[21] , \wRegInBot_4_4[1] , 
        \ScanLink36[0] , \wRegOut_5_24[0] , \wRegOut_5_27[11] , 
        \wRegInTop_4_5[7] , \wRegInTop_4_6[4] , \wRegInBot_4_7[2] , 
        \wRegOut_5_0[8] , \ScanLink35[3] , \wRegOut_5_27[3] , 
        \wRegInTop_5_28[4] , \wRegOut_2_2[30] , \ScanLink8[9] , 
        \wRegInTop_3_1[24] , \ScanLink14[31] , \ScanLink37[19] , 
        \ScanLink42[29] , \ScanLink14[28] , \ScanLink42[30] , \ScanLink61[18] , 
        \wRegOut_4_5[23] , \wRegOut_4_14[28] , \wRegOut_4_14[31] , 
        \ScanLink49[5] , \wRegOut_2_2[29] , \ScanLink6[26] , 
        \wRegInTop_3_1[17] , \wRegInTop_4_11[13] , \wRegInBot_4_11[14] , 
        \wRegInTop_5_29[26] , \ScanLink57[9] , \wRegOut_3_5[1] , 
        \wRegOut_4_5[10] , \wRegInTop_4_11[0] , \wRegInTop_5_30[6] , 
        \wRegOut_5_5[5] , \wRegInTop_4_3[9] , \ScanLink0[1] , 
        \wRegOut_1_0[31] , \wRegOut_1_0[28] , \wRegInBot_2_1[8] , 
        \wRegInTop_4_11[20] , \wRegInTop_4_12[3] , \ScanLink6[15] , 
        \wRegOut_3_6[2] , \wRegOut_5_6[6] , \wRegInTop_5_29[15] , 
        \wRegEnTop_4_5[0] , \wRegInBot_4_11[27] , \ScanLink25[9] , 
        \wRegOut_5_0[26] , \ScanLink38[6] , \wRegInTop_5_23[20] , 
        \wRegInTop_5_15[25] , \wRegInTop_5_25[1] , \wRegInTop_5_26[2] , 
        \wRegInBot_4_6[21] , \wRegInTop_4_8[2] , \wRegInBot_4_9[4] , 
        \wRegOut_5_29[5] , \ScanLink3[2] , \wRegInBot_2_1[18] , 
        \wRegOut_5_0[15] , \wRegInTop_5_15[16] , \wRegInTop_4_3[18] , 
        \wRegInTop_5_23[13] , \wRegInBot_4_6[12] , \ScanLink28[18] , 
        \wRegOut_5_26[31] , \wRegOut_5_26[28] , \wRegOut_2_3[23] , 
        \wRegOut_2_3[10] , \wRegInTop_5_7[17] , \wRegInBot_3_5[17] , 
        \ScanLink15[11] , \ScanLink23[7] , \wRegOut_4_10[1] , 
        \wRegOut_5_31[7] , \ScanLink20[4] , \ScanLink23[14] , 
        \wRegInTop_4_8[14] , \ScanLink36[20] , \ScanLink60[21] , 
        \wRegOut_4_13[2] , \ScanLink43[10] , \wRegOut_4_15[11] , 
        \wRegOut_5_8[0] , \ScanLink56[24] , \wRegInTop_4_10[19] , 
        \ScanLink47[3] , \wRegInBot_3_1[15] , \wRegInBot_3_5[24] , 
        \wRegOut_4_4[30] , \wRegInTop_5_7[24] , \ScanLink15[22] , 
        \wRegOut_4_4[29] , \ScanLink23[27] , \wRegOut_4_15[22] , 
        \ScanLink56[17] , \ScanLink60[12] , \wRegOut_4_0[18] , 
        \wRegInTop_4_8[27] , \ScanLink36[13] , \ScanLink43[23] , 
        \ScanLink44[0] , \wRegOut_4_11[13] , \wRegOut_5_29[26] , 
        \wRegOut_0_0[16] , \ScanLink11[13] , \wRegInBot_4_11[2] , 
        \ScanLink27[16] , \ScanLink52[26] , \ScanLink60[6] , 
        \wRegInBot_4_12[1] , \ScanLink32[22] , \ScanLink47[12] , 
        \ScanLink63[5] , \wRegInBot_3_2[4] , \ScanLink11[20] , 
        \wRegInTop_4_14[31] , \wRegInTop_4_14[28] , \wRegInTop_5_3[15] , 
        \wRegEnTop_5_30[0] , \wRegInTop_5_3[6] , \ScanLink27[25] , 
        \ScanLink32[11] , \ScanLink47[21] , \wRegOut_5_16[2] , 
        \ScanLink52[15] , \wRegInTop_3_3[2] , \wRegOut_5_29[15] , 
        \wRegOut_0_0[25] , \wRegInTop_3_0[1] , \wRegInBot_3_1[26] , 
        \wRegInTop_5_19[5] , \wRegInBot_3_1[7] , \wRegOut_4_11[20] , 
        \wRegInTop_5_0[5] , \wRegInTop_5_3[26] , \wRegOut_5_15[1] , 
        \wRegOut_4_6[9] , \wRegInBot_0_0[2] , \ScanLink0[8] , \wRegOut_2_0[3] , 
        \wRegInTop_2_0[23] , \ScanLink8[22] , \wRegInBot_4_2[23] , 
        \wRegInTop_4_7[30] , \wRegInTop_4_7[29] , \ScanLink59[19] , 
        \wRegOut_5_22[19] , \wRegInTop_2_0[10] , \wRegOut_2_3[0] , 
        \wRegOut_5_4[24] , \wRegInTop_5_11[27] , \wRegInTop_5_5[8] , 
        \wRegInTop_5_27[22] , \wRegEnBot_3_1[0] , \wRegInBot_4_2[10] , 
        \wRegOut_4_3[4] , \wRegOut_5_4[17] , \wRegInTop_5_27[11] , 
        \ScanLink8[11] , \wRegInTop_5_11[14] , \ScanLink5[5] , \ScanLink6[6] , 
        \wRegInBot_3_7[9] , \wRegOut_4_0[7] , \wRegInTop_5_8[19] , 
        \wRegInTop_4_10[10] , \ScanLink7[25] , \wRegInBot_4_10[17] , 
        \wRegInTop_5_28[25] , \wRegInTop_3_0[27] , \ScanLink59[6] , 
        \wRegOut_4_4[20] , \wRegOut_2_3[19] , \ScanLink7[16] , \ScanLink44[9] , 
        \wRegInTop_3_0[14] , \ScanLink15[18] , \wRegOut_4_10[8] , 
        \wRegInBot_4_10[24] , \wRegInTop_5_28[16] , \wRegInTop_4_10[23] , 
        \wRegInTop_5_23[6] , \wRegInTop_5_20[5] , \wRegOut_4_4[13] , 
        \ScanLink36[30] , \ScanLink36[29] , \ScanLink60[28] , \ScanLink43[19] , 
        \ScanLink60[31] , \wRegOut_4_15[18] , \wRegOut_5_8[9] , 
        \wRegOut_1_0[21] , \wRegOut_1_0[12] , \wRegInBot_2_1[11] , 
        \ScanLink41[4] , \wRegOut_3_7[16] , \ScanLink28[11] , 
        \wRegInTop_4_3[11] , \ScanLink42[7] , \ScanLink48[15] , 
        \wRegInBot_2_1[22] , \wRegOut_5_10[24] , \wRegInTop_5_23[30] , 
        \wRegOut_5_26[21] , \ScanLink25[0] , \wRegInTop_5_23[29] , 
        \ScanLink26[3] , \wRegOut_4_15[5] , \wRegInTop_5_25[8] , 
        \wRegOut_5_26[12] , \wRegInTop_2_0[19] , \wRegOut_2_3[9] , 
        \wRegInBot_3_4[3] , \wRegOut_3_7[25] , \wRegInTop_4_3[22] , 
        \wRegOut_5_10[17] , \ScanLink48[26] , \wRegInBot_4_6[31] , 
        \wRegInBot_4_6[28] , \ScanLink28[22] , \wRegInTop_3_5[5] , 
        \wRegInTop_5_5[1] , \wRegOut_5_10[5] , \wRegOut_5_22[23] , 
        \wRegOut_3_3[14] , \wRegInTop_4_7[13] , \ScanLink39[27] , 
        \wRegOut_5_14[26] , \ScanLink59[23] , \wRegInBot_4_2[19] , 
        \ScanLink8[18] , \wRegInTop_3_6[6] , \wRegInBot_3_7[0] , 
        \wRegInTop_5_8[10] , \wRegInTop_5_27[18] , \wRegInTop_5_6[2] , 
        \wRegOut_3_3[27] , \wRegOut_5_13[6] , \ScanLink59[10] , 
        \wRegInTop_4_7[20] , \ScanLink39[14] , \wRegOut_5_14[15] , 
        \wRegOut_5_22[10] , \ScanLink11[30] , \ScanLink11[29] , 
        \wRegOut_4_5[3] , \wRegInBot_4_9[26] , \wRegInBot_4_14[6] , 
        \wRegInTop_5_8[23] , \ScanLink47[31] , \ScanLink32[18] , 
        \ScanLink47[28] , \wRegInTop_3_4[25] , \wRegOut_4_0[22] , 
        \wRegOut_4_11[30] , \wRegOut_4_11[29] , \ScanLink19[4] , 
        \wRegOut_1_1[6] , \ScanLink3[27] , \wRegInTop_3_0[8] , 
        \wRegOut_4_6[0] , \wRegInBot_4_14[15] , \wRegInTop_3_4[16] , 
        \wRegInTop_4_14[12] , \wRegOut_5_15[8] , \wRegOut_4_0[11] , 
        \wRegInBot_4_9[15] , \wRegOut_0_0[12] , \wRegOut_1_1[18] , 
        \ScanLink3[14] , \wRegInBot_4_12[8] , \wRegInTop_4_14[21] , 
        \wRegInBot_4_14[26] , \wRegEnTop_2_0[0] , \wRegInTop_2_0[7] , 
        \wRegInTop_2_1[20] , \wRegOut_5_5[27] , \wRegInTop_5_26[21] , 
        \wRegInTop_5_10[24] , \wRegInTop_2_1[13] , \ScanLink9[21] , 
        \ScanLink9[12] , \wRegInBot_4_3[20] , \wRegInTop_5_9[30] , 
        \wRegInTop_5_9[29] , \wRegInTop_5_11[4] , \wRegInTop_5_10[17] , 
        \wRegInBot_2_2[2] , \wRegInTop_2_3[4] , \wRegInBot_3_0[25] , 
        \wRegInBot_3_0[16] , \ScanLink10[10] , \wRegInBot_4_3[13] , 
        \wRegInTop_4_6[19] , \wRegOut_5_5[14] , \wRegInTop_5_26[12] , 
        \wRegInTop_5_8[4] , \ScanLink58[30] , \ScanLink33[21] , 
        \wRegInTop_5_2[16] , \wRegInTop_5_12[7] , \wRegOut_5_23[29] , 
        \ScanLink58[29] , \wRegOut_5_23[30] , \ScanLink46[11] , 
        \wRegOut_4_10[10] , \ScanLink26[15] , \ScanLink53[25] , 
        \wRegOut_5_28[25] , \ScanLink17[2] , \wRegInTop_4_15[18] , 
        \wRegEnTop_5_23[0] , \wCtrlOut_0[0] , \wRegOut_4_8[6] , 
        \wRegInTop_5_2[25] , \ScanLink10[23] , \ScanLink14[1] , 
        \wRegOut_4_1[31] , \wRegOut_4_1[28] , \wRegOut_4_10[23] , 
        \ScanLink26[26] , \wRegInTop_5_14[9] , \wRegOut_5_28[16] , 
        \ScanLink53[16] , \ScanLink33[12] , \ScanLink46[22] , 
        \wRegInBot_3_4[14] , \wRegOut_4_5[19] , \wRegOut_4_14[12] , 
        \wRegOut_3_5[8] , \wRegInBot_4_2[6] , \wRegInTop_4_3[0] , 
        \ScanLink22[17] , \wRegOut_5_22[7] , \wRegInTop_4_9[17] , 
        \ScanLink30[7] , \ScanLink37[23] , \ScanLink57[27] , 
        \wRegInTop_4_11[9] , \ScanLink42[13] , \ScanLink14[12] , 
        \wRegInTop_4_0[3] , \wRegInBot_4_1[5] , \ScanLink33[4] , 
        \ScanLink61[22] , \wRegOut_5_21[4] , \wRegInBot_2_1[1] , 
        \wRegInTop_4_11[29] , \wRegOut_2_2[20] , \wRegOut_2_2[13] , 
        \wRegInTop_4_11[30] , \ScanLink8[0] , \ScanLink14[21] , 
        \wRegInTop_4_9[24] , \ScanLink37[10] , \wRegInTop_5_6[14] , 
        \ScanLink42[20] , \ScanLink54[3] , \ScanLink61[11] , \ScanLink22[24] , 
        \ScanLink57[14] , \wRegInBot_3_4[27] , \wRegOut_4_14[21] , 
        \wRegInTop_5_6[27] , \wRegOut_3_3[6] , \wRegInTop_4_2[31] , 
        \wRegInTop_4_2[28] , \ScanLink57[0] , \wRegInBot_4_4[8] , 
        \wRegInBot_4_7[22] , \ScanLink29[31] , \ScanLink29[28] , 
        \wRegEnBot_4_14[0] , \ScanLink36[9] , \wRegOut_5_24[9] , 
        \wRegOut_5_27[18] , \wRegInBot_2_0[31] , \wRegOut_3_0[5] , 
        \wRegOut_5_3[2] , \ScanLink28[5] , \wRegInTop_4_14[4] , 
        \wRegOut_5_0[1] , \wRegInTop_5_14[26] , \wRegInBot_2_0[28] , 
        \wRegInTop_5_22[23] , \wRegOut_5_1[25] , \ScanLink3[19] , 
        \wRegOut_2_0[7] , \wRegInTop_2_0[27] , \wRegInBot_4_7[11] , 
        \wRegOut_5_1[16] , \wRegInTop_5_22[10] , \wRegOut_5_4[20] , 
        \wRegInTop_5_14[15] , \wRegInTop_5_27[26] , \wRegInTop_5_11[23] , 
        \ScanLink8[26] , \ScanLink8[15] , \wRegOut_4_0[3] , 
        \wRegInBot_4_2[27] , \wRegOut_5_14[18] , \ScanLink39[19] , 
        \wRegInTop_2_0[14] , \wRegInTop_5_11[10] , \wRegOut_2_3[4] , 
        \wRegOut_3_3[19] , \wRegOut_5_4[13] , \wRegInTop_5_27[15] , 
        \wRegInTop_3_5[8] , \wRegInBot_4_2[14] , \wRegOut_4_3[0] , 
        \wRegInTop_5_3[11] , \wRegOut_5_10[8] , \ScanLink63[1] , 
        \ScanLink11[17] , \wRegInBot_4_12[5] , \ScanLink32[26] , 
        \ScanLink47[16] , \wRegInBot_4_9[18] , \wRegInBot_4_11[6] , 
        \ScanLink27[12] , \ScanLink52[22] , \ScanLink60[2] , 
        \wRegOut_5_29[22] , \wRegOut_0_0[21] , \wRegInBot_3_1[11] , 
        \wRegOut_4_11[17] , \wRegInTop_3_0[5] , \wRegInBot_3_1[3] , 
        \wRegInBot_4_14[18] , \wRegInBot_3_1[22] , \wRegInTop_5_0[1] , 
        \wRegInTop_5_3[22] , \wRegOut_5_15[5] , \wRegInTop_5_19[1] , 
        \ScanLink19[9] , \wRegOut_4_11[24] , \wRegOut_5_29[11] , 
        \ScanLink0[5] , \ScanLink3[6] , \ScanLink5[8] , \wRegOut_2_3[14] , 
        \wRegInTop_3_0[19] , \wRegInBot_3_2[0] , \wRegInTop_3_4[31] , 
        \wRegInTop_3_4[28] , \wRegInTop_3_3[6] , \ScanLink11[24] , 
        \ScanLink27[21] , \ScanLink52[11] , \ScanLink32[15] , \ScanLink47[25] , 
        \wRegOut_5_16[6] , \wRegInTop_5_3[2] , \wRegInBot_3_5[13] , 
        \wRegOut_4_15[15] , \ScanLink15[15] , \ScanLink20[0] , 
        \ScanLink23[10] , \wRegOut_5_8[4] , \wRegOut_4_13[6] , 
        \wRegInTop_4_8[10] , \ScanLink36[24] , \ScanLink56[20] , 
        \ScanLink43[14] , \wRegInTop_5_20[8] , \ScanLink23[3] , 
        \wRegInBot_4_10[30] , \ScanLink60[25] , \wRegOut_4_10[5] , 
        \wRegOut_5_31[3] , \wRegInBot_4_10[29] , \wRegInTop_4_8[23] , 
        \ScanLink36[17] , \wRegInTop_5_7[13] , \ScanLink43[27] , 
        \ScanLink44[4] , \ScanLink60[16] , \wRegOut_2_3[27] , \ScanLink7[31] , 
        \wRegInBot_3_5[20] , \ScanLink15[26] , \ScanLink23[23] , 
        \ScanLink56[13] , \wRegOut_4_15[26] , \wRegInTop_5_7[20] , 
        \ScanLink7[28] , \wRegOut_3_7[31] , \wRegOut_3_7[28] , 
        \wRegInBot_4_6[25] , \wRegInTop_4_8[6] , \wRegInBot_4_9[0] , 
        \ScanLink47[7] , \wRegInTop_5_28[31] , \wRegInTop_5_28[28] , 
        \wRegOut_5_29[1] , \wRegOut_4_15[8] , \wRegOut_5_0[22] , 
        \ScanLink38[2] , \wRegInTop_5_15[21] , \wRegInTop_5_25[5] , 
        \wRegInTop_5_26[6] , \wRegInTop_5_23[24] , \wRegInBot_4_6[16] , 
        \wRegOut_5_10[30] , \wRegOut_5_10[29] , \wRegOut_5_0[11] , 
        \ScanLink48[18] , \wRegInTop_5_23[17] , \ScanLink41[9] , 
        \wRegInTop_5_15[12] , \ScanLink6[22] , \wRegInTop_4_11[17] , 
        \wRegInBot_4_11[10] , \wRegInTop_5_29[22] , \ScanLink6[11] , 
        \wRegInTop_3_1[20] , \ScanLink49[1] , \wRegOut_4_5[27] , 
        \ScanLink22[30] , \ScanLink22[29] , \wRegInTop_4_9[30] , 
        \wRegInTop_4_9[29] , \ScanLink57[19] , \wRegOut_3_6[6] , 
        \wRegInBot_4_1[8] , \wRegEnBot_4_11[0] , \wRegInTop_5_6[19] , 
        \wRegInBot_4_11[23] , \wRegInTop_4_11[24] , \wRegInTop_4_12[7] , 
        \ScanLink33[9] , \wRegOut_5_21[9] , \wRegInTop_5_29[11] , 
        \wRegOut_5_6[2] , \wRegOut_0_0[31] , \wRegOut_0_0[28] , 
        \wRegInBot_1_0[9] , \wRegInBot_1_0[0] , \wRegOut_1_1[15] , 
        \wRegInTop_1_1[6] , \wRegInBot_2_0[16] , \wRegInTop_2_3[9] , 
        \wRegOut_3_5[5] , \wRegInTop_4_11[4] , \wRegInTop_5_30[2] , 
        \wRegInTop_3_1[13] , \wRegInBot_3_4[19] , \wRegOut_4_5[14] , 
        \wRegOut_5_5[1] , \ScanLink51[3] , \wRegOut_3_6[11] , \ScanLink29[16] , 
        \wRegInTop_5_14[18] , \wRegInTop_4_2[16] , \ScanLink49[12] , 
        \ScanLink52[0] , \ScanLink2[20] , \wRegOut_1_1[26] , 
        \wRegInBot_2_0[25] , \ScanLink28[8] , \wRegOut_5_11[23] , 
        \wRegOut_5_27[26] , \wRegInTop_5_28[0] , \wRegOut_3_0[8] , 
        \wRegOut_5_1[31] , \wRegOut_5_1[28] , \ScanLink35[7] , 
        \wRegOut_5_27[7] , \wRegInBot_4_4[5] , \wRegInTop_4_6[0] , 
        \wRegInBot_4_7[6] , \wRegInTop_4_14[9] , \wRegInTop_4_5[3] , 
        \ScanLink36[4] , \wRegOut_5_24[4] , \wRegOut_5_27[15] , 
        \wRegInBot_3_0[31] , \wRegOut_3_2[20] , \wRegOut_3_2[13] , 
        \ScanLink12[2] , \wRegOut_3_6[22] , \wRegInTop_4_2[25] , 
        \wRegOut_5_11[10] , \ScanLink49[21] , \ScanLink29[25] , 
        \wRegOut_5_23[24] , \wRegInTop_4_6[14] , \ScanLink38[20] , 
        \wRegOut_5_15[21] , \wCtrlOut_5[0] , \wRegInTop_5_8[9] , 
        \ScanLink58[24] , \ScanLink11[1] , \wRegOut_5_5[19] , 
        \wRegInTop_5_9[17] , \wRegInTop_5_11[9] , \ScanLink58[17] , 
        \wRegInTop_4_6[27] , \ScanLink38[13] , \wRegInBot_4_8[21] , 
        \wRegInTop_5_9[24] , \wRegOut_5_15[12] , \wRegOut_5_23[17] , 
        \wRegInTop_5_10[30] , \wRegInTop_5_10[29] , \wRegEnTop_5_26[0] , 
        \wRegInTop_5_14[4] , \wRegInBot_3_0[28] , \wRegInTop_3_5[22] , 
        \wRegOut_4_1[25] , \ScanLink2[13] , \wRegInTop_3_5[11] , 
        \wRegInTop_4_15[15] , \wRegInBot_4_15[12] , \wRegInTop_5_2[31] , 
        \wRegInTop_5_2[28] , \wRegOut_5_18[0] , \wRegInTop_5_17[7] , 
        \wRegOut_5_28[31] , \wRegOut_5_28[28] , \wRegOut_4_1[16] , 
        \wRegInBot_4_8[12] , \ScanLink26[18] , \ScanLink53[28] , 
        \wRegInTop_4_15[26] , \ScanLink53[31] , \wRegInBot_4_15[21] , 
        \wRegOut_3_0[1] , \ScanLink28[1] , \wRegOut_5_1[21] , 
        \wRegInTop_5_28[9] , \wRegInTop_5_22[27] , \wRegInTop_4_14[0] , 
        \wRegInTop_5_14[22] , \wRegOut_5_0[5] , \wRegOut_3_3[2] , 
        \wRegInTop_4_6[9] , \wRegOut_5_3[6] , \wRegOut_5_11[19] , 
        \wRegOut_3_6[18] , \wRegEnTop_4_0[0] , \wRegInBot_4_7[26] , 
        \wRegOut_5_1[12] , \wRegInTop_5_14[11] , \ScanLink49[31] , 
        \ScanLink49[28] , \wRegInTop_5_22[14] , \wRegInBot_4_7[15] , 
        \ScanLink52[9] , \ScanLink2[30] , \ScanLink2[29] , \wRegInTop_2_0[3] , 
        \wRegOut_2_2[17] , \ScanLink6[18] , \wRegInTop_5_6[10] , 
        \wRegInBot_2_1[5] , \wRegOut_2_2[24] , \wRegInBot_2_2[6] , 
        \wRegInTop_2_3[0] , \wRegInTop_4_0[7] , \wRegInBot_4_1[1] , 
        \ScanLink33[0] , \wRegInTop_5_29[18] , \wRegOut_5_21[0] , 
        \ScanLink14[16] , \wRegOut_5_5[8] , \wRegInBot_3_4[10] , 
        \wRegInBot_4_2[2] , \ScanLink22[13] , \wRegInTop_4_9[13] , 
        \ScanLink37[27] , \ScanLink61[26] , \ScanLink42[17] , 
        \wRegOut_5_22[3] , \ScanLink30[3] , \ScanLink57[23] , 
        \wRegInTop_4_3[4] , \wRegOut_4_14[16] , \wRegInBot_4_11[19] , 
        \ScanLink57[4] , \wRegInBot_3_0[21] , \wRegInBot_3_0[12] , 
        \ScanLink8[4] , \wRegInTop_3_1[30] , \wRegInBot_3_4[23] , 
        \wRegInTop_5_6[23] , \wRegOut_4_14[25] , \wRegInTop_3_1[29] , 
        \ScanLink49[8] , \ScanLink14[25] , \ScanLink22[20] , \ScanLink57[10] , 
        \ScanLink61[15] , \wRegInTop_4_9[20] , \ScanLink37[14] , 
        \ScanLink42[24] , \ScanLink54[7] , \wRegOut_4_10[14] , 
        \ScanLink10[27] , \ScanLink10[14] , \wRegInTop_3_5[18] , 
        \wRegOut_5_28[21] , \ScanLink26[11] , \ScanLink53[21] , 
        \wRegInBot_4_15[31] , \wRegInBot_4_15[28] , \ScanLink33[25] , 
        \ScanLink46[15] , \wRegInTop_5_2[12] , \ScanLink14[5] , 
        \wRegOut_4_8[2] , \wRegInBot_4_8[31] , \ScanLink33[16] , 
        \ScanLink46[26] , \wRegInBot_4_8[28] , \ScanLink26[22] , 
        \ScanLink53[12] , \wRegOut_5_28[12] , \wRegOut_4_10[27] , 
        \wRegInTop_5_2[21] , \wRegOut_5_18[9] , \wRegInTop_2_1[24] , 
        \ScanLink9[25] , \wRegOut_3_2[30] , \ScanLink17[6] , \wRegOut_3_2[29] , 
        \wRegInBot_4_3[24] , \wRegInTop_2_1[17] , \wRegInBot_4_3[17] , 
        \wRegOut_5_5[23] , \wRegInTop_5_10[20] , \wRegInTop_5_8[0] , 
        \wRegInTop_5_12[3] , \wRegOut_5_15[31] , \wRegInTop_5_26[25] , 
        \wRegOut_5_15[28] , \wRegOut_5_5[10] , \ScanLink38[30] , 
        \ScanLink38[29] , \wRegInTop_5_26[16] , \ScanLink9[16] , 
        \wRegInTop_5_10[13] , \ScanLink11[8] , \wRegInTop_4_14[16] , 
        \wRegInTop_5_0[8] , \wRegInTop_5_11[0] , \ScanLink3[23] , 
        \wRegEnBot_3_4[0] , \wRegOut_4_6[4] , \wRegInBot_4_14[11] , 
        \ScanLink3[10] , \wRegInBot_3_2[9] , \wRegInTop_3_4[21] , 
        \ScanLink19[0] , \wRegOut_5_29[18] , \wRegOut_4_0[26] , 
        \wRegInTop_5_19[8] , \wRegOut_4_5[7] , \wRegInBot_4_9[22] , 
        \ScanLink27[31] , \ScanLink27[28] , \ScanLink52[18] , 
        \wRegInBot_4_14[22] , \wRegInTop_5_3[18] , \ScanLink63[8] , 
        \wRegInBot_0_0[6] , \wRegOut_1_1[2] , \wRegInBot_4_9[11] , 
        \wRegInTop_4_14[25] , \wRegInBot_3_1[18] , \wRegOut_4_0[15] , 
        \wRegOut_3_3[10] , \wRegInTop_3_4[12] , \wRegInTop_3_6[2] , 
        \wRegInBot_3_7[4] , \wRegInTop_5_6[6] , \wRegOut_5_13[2] , 
        \wRegInTop_5_8[14] , \wRegInTop_5_11[19] , \wRegInBot_3_4[7] , 
        \wRegInTop_4_7[17] , \ScanLink39[23] , \ScanLink59[27] , 
        \wRegInTop_5_5[5] , \wRegOut_5_10[1] , \wRegOut_5_14[22] , 
        \wRegOut_5_22[27] , \wRegInTop_3_5[1] , \wRegOut_4_3[9] , 
        \wRegInBot_4_14[2] , \wRegOut_5_4[30] , \wRegOut_5_4[29] , 
        \wRegInTop_5_8[27] , \wRegOut_5_22[14] , \wRegOut_1_0[16] , 
        \wRegOut_3_3[23] , \wRegInTop_4_7[24] , \ScanLink39[10] , 
        \wRegOut_5_14[11] , \wRegOut_5_10[20] , \wRegOut_5_26[25] , 
        \ScanLink59[14] , \ScanLink42[3] , \wRegInTop_4_3[15] , 
        \ScanLink48[11] , \wRegOut_1_0[25] , \wRegInBot_2_1[15] , 
        \wRegOut_3_7[12] , \ScanLink28[15] , \wRegOut_5_0[18] , 
        \wRegOut_3_7[21] , \ScanLink41[0] , \wRegInTop_4_3[26] , 
        \ScanLink28[26] , \ScanLink48[22] , \wRegOut_5_29[8] , 
        \wRegInBot_4_9[9] , \wRegOut_5_10[13] , \wRegOut_1_1[0] , 
        \ScanLink3[21] , \wRegInBot_2_1[26] , \ScanLink25[4] , \ScanLink26[7] , 
        \wRegOut_4_15[1] , \wRegOut_5_26[16] , \ScanLink5[1] , 
        \wRegInTop_5_15[31] , \wRegInTop_5_15[28] , \ScanLink6[2] , 
        \ScanLink7[21] , \wRegInTop_3_0[23] , \wRegInBot_3_5[30] , 
        \wRegInBot_3_5[29] , \wRegOut_4_4[24] , \ScanLink59[2] , 
        \wRegInTop_4_10[14] , \wRegInBot_4_10[13] , \wRegInTop_5_7[30] , 
        \wRegInTop_5_7[29] , \wRegInTop_5_28[21] , \ScanLink7[12] , 
        \wRegInTop_3_0[10] , \wRegOut_4_4[17] , \ScanLink20[9] , 
        \ScanLink23[19] , \wRegInTop_4_8[19] , \wRegInTop_5_20[1] , 
        \ScanLink56[30] , \wRegInTop_4_10[27] , \wRegInTop_5_23[2] , 
        \ScanLink56[29] , \wRegInBot_4_10[20] , \wRegInTop_5_28[12] , 
        \wRegInBot_3_1[30] , \wRegInBot_3_1[29] , \wRegOut_4_5[5] , 
        \wRegInBot_4_9[20] , \wRegInTop_5_3[9] , \wRegOut_4_0[24] , 
        \wRegInTop_3_4[23] , \ScanLink19[2] , \wRegInBot_3_1[8] , 
        \wRegOut_4_6[6] , \wRegInBot_4_14[13] , \wRegInTop_5_3[30] , 
        \wRegInTop_5_3[29] , \wRegInTop_3_4[10] , \wRegInTop_4_14[14] , 
        \wRegEnTop_5_5[0] , \wRegOut_5_29[29] , \wRegOut_4_0[17] , 
        \wRegOut_5_29[30] , \wRegInBot_4_9[13] , \ScanLink52[30] , 
        \ScanLink27[19] , \ScanLink52[29] , \wRegInTop_4_14[27] , 
        \ScanLink60[9] , \wRegOut_0_0[19] , \wRegInBot_0_0[4] , 
        \ScanLink3[12] , \wRegInBot_4_14[20] , \wRegOut_3_3[21] , 
        \wRegOut_3_3[12] , \wRegInBot_3_4[5] , \wRegInTop_3_5[3] , 
        \wRegOut_5_22[25] , \wRegInTop_4_7[15] , \wRegInTop_5_5[7] , 
        \wRegOut_5_14[20] , \wRegOut_5_10[3] , \ScanLink39[21] , 
        \wRegInTop_3_6[0] , \wRegOut_5_4[18] , \ScanLink59[25] , 
        \wRegInBot_3_7[6] , \wRegOut_4_0[8] , \wRegInTop_5_6[4] , 
        \wRegInTop_5_8[16] , \wRegOut_5_13[0] , \wRegInTop_4_7[26] , 
        \ScanLink59[16] , \ScanLink39[12] , \wRegOut_5_14[13] , 
        \wRegOut_5_22[16] , \wRegOut_1_0[27] , \wRegOut_1_0[14] , 
        \wRegInBot_2_1[17] , \wRegInBot_4_14[0] , \wRegInTop_5_8[25] , 
        \ScanLink41[2] , \wRegInTop_5_11[31] , \wRegInTop_5_11[28] , 
        \wRegOut_3_7[10] , \wRegInTop_5_15[19] , \wRegInTop_4_3[17] , 
        \ScanLink28[17] , \ScanLink48[13] , \wRegOut_5_10[22] , 
        \wRegInBot_2_1[24] , \wRegOut_5_0[30] , \ScanLink38[9] , 
        \ScanLink42[1] , \wRegOut_5_26[27] , \ScanLink25[6] , 
        \wRegOut_5_0[29] , \ScanLink26[5] , \wRegOut_4_15[3] , 
        \wRegOut_5_26[14] , \wRegOut_5_10[11] , \wRegEnBot_2_1[0] , 
        \ScanLink5[3] , \ScanLink6[0] , \wRegOut_3_7[23] , \wRegInTop_4_3[24] , 
        \ScanLink48[20] , \ScanLink28[24] , \ScanLink7[23] , 
        \wRegInTop_4_10[16] , \wRegInBot_4_10[11] , \wRegInTop_5_28[23] , 
        \wRegInTop_3_0[21] , \ScanLink59[0] , \wRegOut_4_4[26] , 
        \wRegInTop_4_8[28] , \ScanLink7[10] , \ScanLink23[31] , 
        \wRegInTop_4_8[31] , \ScanLink23[28] , \ScanLink56[18] , 
        \wRegInTop_3_0[12] , \wRegInBot_3_5[18] , \wRegOut_4_4[15] , 
        \ScanLink23[8] , \wRegInTop_5_7[18] , \wRegInTop_5_28[10] , 
        \wRegInTop_4_10[25] , \wRegInBot_4_10[22] , \wRegOut_5_31[8] , 
        \wRegInTop_5_20[3] , \wRegInTop_5_23[0] , \wRegOut_3_3[0] , 
        \wRegOut_3_6[30] , \wRegOut_3_6[29] , \wRegInBot_4_7[24] , 
        \wRegInTop_4_5[8] , \wRegOut_5_3[4] , \wRegOut_3_0[3] , 
        \wRegInTop_3_1[18] , \wRegInBot_3_4[12] , \wRegInBot_4_7[17] , 
        \ScanLink28[3] , \wRegInTop_4_14[2] , \wRegOut_5_0[7] , 
        \wRegOut_5_1[23] , \wRegInTop_5_14[20] , \wRegOut_5_11[31] , 
        \wRegInTop_5_22[25] , \wRegOut_5_11[28] , \wRegOut_5_1[10] , 
        \ScanLink49[19] , \wRegInTop_5_14[13] , \wRegInTop_5_22[16] , 
        \ScanLink51[8] , \wRegOut_4_14[14] , \ScanLink2[18] , 
        \wRegInTop_2_0[1] , \wRegInBot_2_1[7] , \wRegInBot_2_2[4] , 
        \wRegInBot_4_2[0] , \wRegInTop_4_3[6] , \ScanLink22[11] , 
        \ScanLink57[21] , \ScanLink30[1] , \wRegOut_5_22[1] , 
        \wRegInTop_2_3[2] , \ScanLink14[14] , \ScanLink61[24] , 
        \wRegInTop_5_30[9] , \wRegInTop_4_0[5] , \wRegInTop_4_9[11] , 
        \ScanLink42[15] , \ScanLink37[25] , \wRegInBot_4_1[3] , 
        \wRegInBot_4_11[28] , \wRegInBot_4_11[31] , \ScanLink33[2] , 
        \wRegOut_5_6[9] , \wRegOut_5_21[2] , \wRegOut_2_2[26] , 
        \wRegOut_2_2[15] , \ScanLink6[29] , \ScanLink8[6] , \ScanLink14[27] , 
        \wRegInTop_5_6[12] , \ScanLink22[22] , \wRegInTop_4_9[22] , 
        \ScanLink61[17] , \ScanLink37[16] , \ScanLink42[26] , \ScanLink54[5] , 
        \ScanLink57[12] , \wRegInBot_3_4[21] , \wRegOut_4_14[27] , 
        \wRegInTop_5_6[21] , \ScanLink6[30] , \wRegInTop_5_2[10] , 
        \ScanLink57[6] , \wRegInTop_5_29[30] , \wRegInTop_5_29[29] , 
        \wRegInTop_2_1[26] , \wRegInBot_3_0[23] , \wRegInBot_3_0[10] , 
        \ScanLink10[16] , \wRegInBot_4_8[19] , \ScanLink26[13] , 
        \ScanLink33[27] , \ScanLink46[17] , \ScanLink53[23] , 
        \wRegOut_5_28[23] , \ScanLink17[4] , \wRegOut_4_10[16] , 
        \wRegInBot_4_15[19] , \wRegOut_4_10[25] , \wRegInTop_5_2[23] , 
        \ScanLink10[25] , \wRegInTop_3_5[30] , \wRegOut_4_8[0] , 
        \wRegInTop_3_5[29] , \wRegOut_5_28[10] , \ScanLink26[20] , 
        \ScanLink53[10] , \ScanLink14[7] , \ScanLink33[14] , \wRegOut_5_5[21] , 
        \ScanLink46[24] , \wRegInTop_5_26[27] , \wRegInTop_2_1[15] , 
        \ScanLink9[27] , \wRegInTop_5_10[22] , \ScanLink9[14] , 
        \wRegInBot_4_3[26] , \wRegOut_5_15[19] , \ScanLink38[18] , 
        \wRegInTop_5_11[2] , \ScanLink6[20] , \wRegInTop_3_1[22] , 
        \wRegOut_3_2[18] , \wRegOut_5_5[12] , \wRegInTop_5_10[11] , 
        \wRegInTop_5_26[14] , \wRegInBot_3_4[31] , \ScanLink12[9] , 
        \wRegInBot_4_3[15] , \wRegInTop_5_8[2] , \wRegInTop_5_12[1] , 
        \wRegInBot_3_4[28] , \wRegOut_4_5[25] , \ScanLink49[3] , 
        \wRegInTop_3_1[11] , \wRegInTop_4_11[15] , \wRegInBot_4_11[12] , 
        \wRegInTop_5_6[31] , \wRegInTop_5_6[28] , \wRegInTop_5_29[20] , 
        \wRegOut_4_5[16] , \wRegInTop_4_9[18] , \wRegInTop_4_11[6] , 
        \wRegOut_5_5[3] , \wRegInTop_5_30[0] , \ScanLink57[28] , 
        \wRegInBot_1_0[2] , \wRegInTop_2_0[8] , \wRegOut_3_5[7] , 
        \wRegInBot_4_2[9] , \ScanLink22[18] , \wRegOut_5_22[8] , 
        \ScanLink30[8] , \ScanLink57[31] , \wRegInTop_4_11[26] , 
        \wRegOut_5_6[0] , \ScanLink6[13] , \wRegOut_3_6[4] , 
        \wRegInTop_4_12[5] , \wRegEnBot_4_4[0] , \wRegInBot_4_11[21] , 
        \wRegInTop_5_29[13] , \wRegOut_5_27[24] , \wRegOut_1_1[17] , 
        \wRegInTop_1_1[4] , \ScanLink52[2] , \wRegInBot_2_0[14] , 
        \wRegOut_3_6[13] , \wRegInTop_4_2[14] , \wRegOut_5_11[21] , 
        \ScanLink49[10] , \ScanLink29[14] , \wRegOut_5_1[19] , 
        \wRegOut_3_6[20] , \ScanLink29[27] , \ScanLink51[1] , \ScanLink2[22] , 
        \wRegOut_1_1[24] , \wRegInTop_4_2[27] , \ScanLink49[23] , 
        \wRegInBot_2_0[27] , \wRegOut_3_3[9] , \wRegInTop_4_5[1] , 
        \wRegOut_5_11[12] , \wRegInBot_4_4[7] , \wRegInTop_4_6[2] , 
        \ScanLink35[5] , \ScanLink36[6] , \wRegOut_5_24[6] , 
        \wRegOut_5_27[17] , \wRegOut_5_27[5] , \wRegInBot_4_7[4] , 
        \wRegOut_3_2[22] , \wRegOut_3_2[11] , \ScanLink11[3] , 
        \wRegInTop_5_14[30] , \wRegInTop_5_28[2] , \wRegInTop_5_14[29] , 
        \wRegInTop_5_9[15] , \wRegInTop_5_10[18] , \ScanLink58[26] , 
        \ScanLink12[0] , \wRegInTop_4_6[16] , \ScanLink38[22] , 
        \wRegInTop_4_6[25] , \wRegOut_5_5[31] , \wRegOut_5_5[28] , 
        \wRegInTop_5_12[8] , \wRegOut_5_15[23] , \wRegOut_5_23[26] , 
        \wRegInTop_5_9[26] , \wRegOut_5_15[10] , \wRegOut_5_23[15] , 
        \wEnable_0[0] , \ScanLink38[11] , \ScanLink58[15] , 
        \wRegInTop_4_15[17] , \wRegInBot_4_15[10] , \wRegInTop_5_17[5] , 
        \wRegOut_5_18[2] , \ScanLink2[11] , \wRegInTop_3_5[20] , 
        \wRegOut_5_28[19] , \wRegOut_4_1[27] , \wRegOut_4_8[9] , 
        \wRegInBot_4_8[23] , \ScanLink26[30] , \ScanLink26[29] , 
        \ScanLink53[19] , \wRegInTop_5_14[6] , \wRegOut_2_0[5] , 
        \wRegInTop_2_0[25] , \wRegInBot_3_0[19] , \wRegOut_4_1[14] , 
        \wRegInBot_4_8[10] , \wRegInTop_4_15[24] , \wRegInBot_4_15[23] , 
        \wRegInTop_5_2[19] , \ScanLink8[24] , \wRegOut_3_3[31] , 
        \wRegOut_3_3[28] , \wRegInTop_3_5[13] , \wRegInBot_4_2[25] , 
        \wRegInBot_4_14[9] , \wRegInTop_5_11[21] , \wRegInTop_2_0[16] , 
        \wRegOut_2_3[6] , \wRegOut_5_4[22] , \wRegInTop_5_27[24] , 
        \wRegEnTop_3_0[0] , \wRegOut_5_14[30] , \wRegOut_5_14[29] , 
        \wRegInBot_4_2[16] , \wRegOut_4_3[2] , \wRegOut_5_4[11] , 
        \ScanLink39[31] , \ScanLink39[28] , \wRegInTop_5_27[17] , 
        \wRegInTop_5_11[12] , \wRegOut_5_13[9] , \ScanLink8[17] , 
        \wRegInBot_3_1[13] , \wRegInTop_3_6[9] , \wRegOut_4_0[1] , 
        \wRegOut_4_11[15] , \wRegOut_5_29[20] , \wRegOut_0_0[10] , 
        \wRegOut_1_1[9] , \wRegInTop_3_4[19] , \wRegInBot_4_11[4] , 
        \ScanLink52[20] , \ScanLink27[10] , \ScanLink60[0] , \ScanLink11[15] , 
        \ScanLink32[24] , \ScanLink47[14] , \wRegInBot_4_12[7] , 
        \wRegInBot_3_2[2] , \wRegInTop_3_3[4] , \ScanLink11[26] , 
        \wRegEnTop_4_11[0] , \wRegInBot_4_14[30] , \ScanLink63[3] , 
        \wRegInBot_4_14[29] , \ScanLink32[17] , \wRegInTop_5_3[13] , 
        \ScanLink47[27] , \wRegOut_5_16[4] , \wRegInTop_5_3[0] , 
        \wRegInBot_4_9[29] , \wRegInBot_4_9[30] , \ScanLink27[23] , 
        \ScanLink52[13] , \wRegOut_5_29[13] , \wRegOut_0_0[23] , 
        \ScanLink3[31] , \wRegInBot_3_1[20] , \wRegOut_4_11[26] , 
        \wRegInTop_5_3[20] , \wRegInTop_5_19[3] , \ScanLink3[28] , 
        \wRegInTop_5_0[3] , \wRegOut_5_15[7] , \wRegInBot_0_0[0] , 
        \ScanLink0[7] , \ScanLink6[9] , \wRegOut_2_3[16] , \wRegInTop_3_0[7] , 
        \wRegInBot_3_1[1] , \wRegInTop_5_7[11] , \ScanLink7[19] , 
        \wRegInBot_3_5[11] , \ScanLink15[17] , \ScanLink23[1] , 
        \wRegInTop_5_23[9] , \wRegInTop_4_8[12] , \wRegOut_4_10[7] , 
        \wRegInTop_5_28[19] , \ScanLink43[16] , \wRegOut_5_31[1] , 
        \ScanLink36[26] , \ScanLink60[27] , \ScanLink20[2] , \ScanLink23[12] , 
        \wRegOut_4_13[4] , \ScanLink56[22] , \wRegOut_5_8[6] , 
        \wRegInBot_4_10[18] , \wRegOut_4_15[17] , \wRegOut_2_3[25] , 
        \ScanLink47[5] , \wRegInTop_3_0[31] , \wRegInTop_3_0[28] , 
        \wRegInBot_3_5[22] , \wRegOut_4_15[24] , \wRegInTop_5_7[22] , 
        \wRegEnTop_5_14[0] , \ScanLink59[9] , \ScanLink15[24] , 
        \ScanLink23[21] , \wRegInTop_4_8[21] , \ScanLink56[11] , 
        \ScanLink36[15] , \ScanLink43[25] , \ScanLink44[6] , 
        \wRegInBot_4_6[27] , \wRegOut_5_0[20] , \wRegInTop_5_23[26] , 
        \ScanLink60[14] , \ScanLink38[0] , \wRegInTop_5_15[23] , 
        \wRegOut_5_10[18] , \wRegInTop_5_25[7] , \wRegInTop_5_26[4] , 
        \wRegInTop_4_8[4] , \ScanLink48[29] , \wRegOut_5_29[3] , 
        \wRegInBot_4_9[2] , \ScanLink48[30] , \wRegOut_1_0[23] , 
        \wRegOut_1_0[10] , \wRegOut_1_1[30] , \ScanLink3[4] , 
        \wRegOut_3_7[19] , \wRegOut_5_0[13] , \wRegInTop_5_15[10] , 
        \wRegInTop_5_23[15] , \wRegInBot_4_6[14] , \wRegInTop_2_0[5] , 
        \wRegInTop_2_1[22] , \ScanLink9[23] , \wRegInBot_4_3[22] , 
        \wRegInTop_4_6[31] , \wRegInTop_4_6[28] , \ScanLink42[8] , 
        \wRegOut_5_23[18] , \ScanLink58[18] , \wRegInTop_5_10[26] , 
        \wRegInTop_2_1[11] , \wRegInBot_4_3[11] , \wRegOut_5_5[25] , 
        \wRegInTop_5_26[23] , \wRegInTop_5_12[5] , \wRegOut_5_5[16] , 
        \wRegInTop_5_8[6] , \wRegInTop_5_26[10] , \wRegInTop_5_10[15] , 
        \wRegInBot_2_1[3] , \wRegOut_2_2[11] , \wRegInBot_3_0[27] , 
        \wRegInBot_3_0[14] , \ScanLink9[10] , \wRegOut_4_1[19] , 
        \wRegInTop_5_9[18] , \wRegInTop_5_11[6] , \ScanLink10[21] , 
        \ScanLink10[12] , \wRegOut_4_10[12] , \ScanLink26[17] , 
        \ScanLink53[27] , \wRegOut_5_28[27] , \ScanLink33[23] , 
        \ScanLink46[13] , \ScanLink14[3] , \wRegInTop_4_15[30] , 
        \wRegInTop_4_15[29] , \ScanLink33[10] , \wRegInTop_5_2[14] , 
        \ScanLink46[20] , \wRegOut_4_10[21] , \ScanLink26[24] , 
        \ScanLink53[14] , \wRegOut_5_28[14] , \ScanLink17[0] , 
        \wRegOut_4_8[4] , \wRegInTop_5_2[27] , \wRegInTop_5_6[16] , 
        \wRegInTop_5_17[8] , \wRegOut_2_2[22] , \wRegInBot_2_2[0] , 
        \wRegOut_3_6[9] , \wRegInTop_4_0[1] , \wRegInTop_4_12[8] , 
        \ScanLink33[6] , \wRegOut_5_21[6] , \wRegInBot_4_1[7] , 
        \wRegInTop_4_9[15] , \ScanLink42[11] , \ScanLink37[21] , 
        \wRegInTop_2_3[6] , \ScanLink14[10] , \ScanLink61[20] , 
        \wRegInBot_3_4[16] , \wRegInBot_4_2[4] , \wRegInTop_4_3[2] , 
        \ScanLink22[15] , \ScanLink57[25] , \ScanLink30[5] , \wRegOut_5_22[5] , 
        \wRegInTop_4_11[18] , \wRegOut_4_14[10] , \ScanLink57[2] , 
        \wRegOut_3_0[7] , \ScanLink8[2] , \wRegInBot_3_4[25] , 
        \wRegOut_4_14[23] , \wRegInTop_5_6[25] , \wRegOut_4_5[31] , 
        \wRegOut_4_5[28] , \ScanLink14[23] , \ScanLink22[26] , 
        \wRegInTop_4_9[26] , \ScanLink57[16] , \ScanLink37[12] , 
        \ScanLink42[22] , \ScanLink54[1] , \wRegInBot_4_7[9] , \ScanLink28[7] , 
        \wRegOut_5_1[27] , \wRegInTop_5_22[21] , \ScanLink61[13] , 
        \wRegInTop_5_14[24] , \wRegInTop_4_14[6] , \wRegOut_5_0[3] , 
        \wRegOut_5_3[0] , \ScanLink35[8] , \wRegOut_5_27[8] , 
        \wRegOut_1_1[29] , \wRegInTop_1_1[9] , \wRegInBot_2_0[19] , 
        \wRegOut_3_3[4] , \wRegEnBot_4_1[0] , \wRegInBot_4_7[20] , 
        \wRegOut_5_1[14] , \wRegInTop_5_14[17] , \wRegInTop_5_22[12] , 
        \wRegInTop_4_2[19] , \wRegInBot_4_7[13] , \ScanLink29[19] , 
        \wRegOut_5_27[30] , \wRegOut_5_27[29] , \ScanLink5[7] , \ScanLink6[4] , 
        \wRegOut_2_3[31] , \wRegOut_2_3[28] , \ScanLink7[27] , 
        \wRegInTop_3_0[25] , \ScanLink15[30] , \ScanLink15[29] , 
        \ScanLink43[31] , \ScanLink60[19] , \wRegOut_4_4[22] , 
        \wRegOut_4_15[30] , \ScanLink36[18] , \ScanLink43[28] , 
        \wRegOut_4_15[29] , \ScanLink59[4] , \wRegInBot_4_10[15] , 
        \ScanLink47[8] , \wRegInTop_5_28[27] , \ScanLink7[14] , 
        \wRegInTop_3_0[16] , \wRegInTop_4_10[12] , \wRegOut_4_4[11] , 
        \wRegInTop_4_10[21] , \wRegOut_4_13[9] , \wRegInTop_5_20[7] , 
        \wRegInBot_4_10[26] , \wRegInTop_5_23[4] , \wRegInTop_5_28[14] , 
        \wRegOut_5_26[23] , \ScanLink3[9] , \ScanLink42[5] , 
        \wRegInBot_2_1[13] , \wRegOut_3_7[14] , \wRegInTop_4_3[13] , 
        \wRegOut_5_10[26] , \ScanLink48[17] , \ScanLink28[13] , 
        \wRegInBot_4_6[19] , \wRegEnTop_5_11[0] , \wRegOut_3_7[27] , 
        \ScanLink28[20] , \ScanLink41[6] , \wRegInTop_5_23[18] , 
        \wRegInTop_4_3[20] , \wRegInTop_4_8[9] , \ScanLink48[24] , 
        \wRegOut_2_0[8] , \wRegInBot_2_1[20] , \ScanLink25[2] , 
        \ScanLink26[1] , \wRegOut_4_15[7] , \wRegOut_5_10[15] , 
        \wRegInTop_5_26[9] , \wRegOut_5_26[10] , \wRegInTop_2_0[31] , 
        \wRegInTop_2_0[28] , \wRegOut_3_3[16] , \wRegInTop_3_6[4] , 
        \wRegInTop_5_6[0] , \wRegInTop_5_8[12] , \wRegOut_5_13[4] , 
        \wRegInBot_3_7[2] , \ScanLink59[21] , \wRegInBot_3_4[1] , 
        \wRegInTop_3_5[7] , \wRegInTop_4_7[11] , \wRegInTop_5_5[3] , 
        \ScanLink39[25] , \wRegOut_5_10[7] , \wRegOut_5_14[24] , 
        \wRegOut_5_22[21] , \ScanLink8[30] , \ScanLink8[29] , 
        \wRegInBot_4_14[4] , \wRegInTop_5_27[30] , \wRegInTop_5_27[29] , 
        \wRegInTop_5_8[21] , \wRegOut_5_22[12] , \ScanLink3[25] , 
        \wRegOut_3_3[25] , \wRegInBot_4_2[31] , \wRegInTop_4_7[22] , 
        \wRegEnTop_4_14[0] , \wRegOut_5_14[17] , \ScanLink39[16] , 
        \wRegInBot_4_2[28] , \ScanLink59[12] , \wRegEnTop_3_5[0] , 
        \wRegInTop_4_14[10] , \wRegInBot_4_14[17] , \wRegOut_4_6[2] , 
        \ScanLink3[16] , \wRegInTop_3_3[9] , \wRegInTop_3_4[27] , 
        \ScanLink19[6] , \wRegOut_4_0[20] , \wRegOut_5_16[9] , 
        \wRegOut_4_5[1] , \wRegInBot_4_9[24] , \wRegInTop_4_14[23] , 
        \wRegInBot_4_14[24] , \wRegOut_1_1[4] , \ScanLink11[18] , 
        \wRegInBot_4_9[17] , \wRegInBot_4_11[9] , \ScanLink32[30] , 
        \wRegOut_4_0[13] , \wRegOut_4_11[18] , \ScanLink32[29] , 
        \ScanLink47[19] , \wRegInTop_3_4[14] , \ScanLink0[3] , 
        \wRegOut_1_0[19] , \wRegInBot_2_1[30] , \wRegInBot_2_1[29] , 
        \wRegInTop_4_3[30] , \wRegInTop_4_8[0] , \wRegInTop_4_3[29] , 
        \wRegInBot_4_9[6] , \wRegInBot_4_6[23] , \ScanLink28[30] , 
        \ScanLink28[29] , \wRegOut_5_29[7] , \ScanLink26[8] , 
        \wRegOut_5_26[19] , \ScanLink38[4] , \wRegInTop_5_25[3] , 
        \wRegInTop_5_26[0] , \wRegInTop_5_15[27] , \wRegOut_5_0[24] , 
        \wRegInTop_5_23[22] , \ScanLink3[0] , \wRegInBot_4_6[10] , 
        \wRegOut_5_0[17] , \wRegInTop_5_15[14] , \wRegInTop_5_23[11] , 
        \wRegOut_2_3[21] , \wRegOut_2_3[12] , \wRegInBot_3_5[15] , 
        \wRegOut_4_4[18] , \ScanLink15[13] , \ScanLink20[6] , \ScanLink23[16] , 
        \wRegOut_4_15[13] , \wRegOut_5_8[2] , \ScanLink56[26] , 
        \wRegOut_4_13[0] , \ScanLink60[23] , \ScanLink23[5] , 
        \wRegInTop_4_8[16] , \ScanLink43[12] , \ScanLink36[22] , 
        \wRegOut_4_10[3] , \wRegInTop_4_10[31] , \wRegOut_5_31[5] , 
        \wRegInTop_4_10[28] , \wRegInBot_3_5[26] , \ScanLink15[20] , 
        \wRegInTop_5_7[15] , \ScanLink23[25] , \wRegInTop_4_8[25] , 
        \ScanLink60[10] , \ScanLink36[11] , \ScanLink43[21] , \ScanLink44[2] , 
        \wRegOut_4_15[20] , \ScanLink56[15] , \wRegInTop_5_7[26] , 
        \wRegInTop_5_3[17] , \ScanLink47[1] , \wRegOut_0_0[14] , 
        \ScanLink11[11] , \wRegInBot_4_12[3] , \ScanLink63[7] , 
        \wRegInBot_4_11[0] , \ScanLink32[20] , \ScanLink47[10] , 
        \ScanLink52[24] , \ScanLink27[14] , \ScanLink60[4] , 
        \wRegOut_5_29[24] , \wRegOut_0_0[27] , \wRegInTop_3_0[3] , 
        \wRegInBot_3_1[17] , \wRegOut_4_11[11] , \wRegInBot_3_1[5] , 
        \wRegInBot_3_1[24] , \wRegOut_4_0[30] , \wRegInTop_4_14[19] , 
        \wRegOut_5_15[3] , \wRegInTop_5_0[7] , \wRegInTop_5_3[24] , 
        \wRegOut_4_11[22] , \wRegOut_4_0[29] , \wRegInTop_5_19[7] , 
        \wRegOut_5_29[17] , \wRegInBot_0_0[9] , \wRegInTop_2_0[21] , 
        \wRegInBot_3_2[6] , \wRegInTop_3_3[0] , \ScanLink27[27] , 
        \ScanLink52[17] , \ScanLink11[22] , \wRegOut_4_5[8] , \ScanLink32[13] , 
        \wRegInTop_5_3[4] , \wRegOut_5_4[26] , \ScanLink47[23] , 
        \wRegOut_5_16[0] , \wRegInTop_5_27[20] , \ScanLink8[20] , 
        \wRegInTop_5_11[25] , \wRegInTop_5_8[31] , \wRegInTop_5_8[28] , 
        \wRegEnTop_5_28[0] , \wRegInBot_1_0[6] , \ScanLink2[26] , 
        \wRegOut_2_0[1] , \wRegOut_4_0[5] , \wRegInBot_4_2[21] , 
        \wRegInTop_2_0[12] , \ScanLink8[13] , \wRegInTop_5_6[9] , 
        \wRegOut_2_3[2] , \wRegInBot_3_4[8] , \wRegInBot_4_2[12] , 
        \wRegInTop_4_7[18] , \wRegOut_5_4[15] , \wRegInTop_5_11[16] , 
        \wRegInTop_5_27[13] , \ScanLink59[28] , \wRegOut_4_3[6] , 
        \wRegOut_5_22[31] , \ScanLink59[31] , \wRegOut_5_22[28] , 
        \ScanLink10[31] , \wRegInBot_4_8[27] , \wRegEnTop_5_0[0] , 
        \wRegInTop_5_14[2] , \ScanLink10[28] , \ScanLink33[19] , 
        \ScanLink46[29] , \wRegInTop_3_5[24] , \wRegOut_4_1[23] , 
        \ScanLink46[30] , \wRegOut_4_10[31] , \wRegOut_4_10[28] , 
        \ScanLink2[15] , \wRegInTop_3_5[17] , \ScanLink17[9] , 
        \wRegInTop_4_15[13] , \wRegInBot_4_15[14] , \wRegOut_5_18[6] , 
        \wRegInTop_5_17[1] , \wRegOut_4_1[10] , \wRegInBot_4_8[14] , 
        \wRegInTop_4_15[20] , \wRegInBot_4_15[27] , \wRegOut_1_1[13] , 
        \wRegInBot_2_0[10] , \wRegInTop_2_1[18] , \wRegOut_3_2[15] , 
        \ScanLink12[4] , \wRegOut_5_15[27] , \wRegOut_5_23[22] , 
        \wRegInTop_4_6[12] , \ScanLink38[26] , \wRegInBot_4_3[18] , 
        \ScanLink58[22] , \ScanLink9[19] , \ScanLink11[7] , 
        \wRegInTop_5_9[11] , \wRegInTop_5_26[19] , \wRegOut_3_2[26] , 
        \wRegInTop_4_6[21] , \ScanLink58[11] , \ScanLink38[15] , 
        \wRegInTop_5_9[22] , \wRegOut_5_15[14] , \wRegOut_5_23[11] , 
        \ScanLink51[5] , \wRegOut_3_6[17] , \wRegInTop_4_2[10] , 
        \ScanLink29[10] , \ScanLink49[14] , \wRegOut_5_11[25] , 
        \wRegOut_1_1[20] , \wRegInTop_1_1[0] , \ScanLink52[6] , 
        \wRegInBot_2_0[23] , \wRegInTop_5_22[28] , \wRegOut_5_27[20] , 
        \wRegInBot_4_4[3] , \wRegInTop_4_5[5] , \wRegInTop_4_6[6] , 
        \wRegInTop_5_22[31] , \wRegInTop_5_28[6] , \wRegInBot_4_7[0] , 
        \ScanLink35[1] , \ScanLink36[2] , \wRegOut_5_24[2] , 
        \wRegOut_5_27[13] , \wRegOut_5_27[1] , \wRegOut_5_3[9] , 
        \wRegOut_5_11[16] , \wRegOut_2_2[18] , \ScanLink6[24] , 
        \wRegOut_3_6[24] , \wRegInTop_4_2[23] , \wRegInBot_4_7[29] , 
        \ScanLink49[27] , \wRegInBot_4_7[30] , \ScanLink29[23] , 
        \wRegInTop_4_11[11] , \wRegInBot_4_11[16] , \wRegInTop_5_29[24] , 
        \wRegInTop_3_1[26] , \ScanLink49[7] , \wRegOut_4_5[21] , 
        \ScanLink54[8] , \ScanLink6[17] , \wRegOut_3_5[3] , \wRegOut_3_6[0] , 
        \wRegInTop_4_0[8] , \wRegInTop_5_29[17] , \wRegInBot_4_11[25] , 
        \wRegInTop_4_11[22] , \wRegInTop_4_12[1] , \wRegOut_5_6[4] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[11] , \wRegOut_1_1[31] , 
        \wRegOut_1_1[28] , \wRegInTop_2_1[23] , \wRegInBot_2_2[9] , 
        \ScanLink37[28] , \ScanLink42[18] , \ScanLink61[30] , 
        \wRegInBot_3_0[26] , \wRegInBot_3_0[15] , \wRegInTop_3_1[15] , 
        \ScanLink14[19] , \wRegInTop_4_11[2] , \wRegOut_5_5[7] , 
        \ScanLink61[29] , \ScanLink37[31] , \wRegInTop_5_30[4] , 
        \wRegOut_4_5[12] , \wRegOut_4_14[19] , \wRegInTop_4_15[31] , 
        \wRegInTop_4_15[28] , \wRegInTop_5_2[15] , \wRegEnTop_5_20[0] , 
        \wRegOut_5_28[26] , \ScanLink10[20] , \ScanLink10[13] , 
        \wRegOut_4_1[18] , \wRegOut_4_10[13] , \ScanLink17[1] , 
        \ScanLink26[16] , \ScanLink33[22] , \ScanLink46[12] , \ScanLink53[26] , 
        \wRegInTop_5_2[26] , \wRegEnTop_5_8[0] , \wRegInTop_5_17[9] , 
        \ScanLink26[25] , \ScanLink53[15] , \ScanLink14[2] , \ScanLink33[11] , 
        \wCtrlOut_3[0] , \ScanLink46[21] , \wRegOut_4_10[20] , \ScanLink9[22] , 
        \wRegOut_4_8[5] , \wRegOut_5_28[15] , \wRegOut_5_5[24] , 
        \wRegInTop_5_26[22] , \wRegInTop_2_1[10] , \wRegInBot_4_3[23] , 
        \wRegInTop_5_10[27] , \ScanLink58[19] , \wRegInTop_4_6[30] , 
        \wRegInTop_4_6[29] , \wRegOut_5_23[19] , \ScanLink9[11] , 
        \wRegOut_5_5[17] , \wRegInTop_5_10[14] , \wRegInTop_5_9[19] , 
        \wRegInTop_5_26[11] , \wRegInTop_5_11[7] , \wRegOut_3_3[5] , 
        \wRegInBot_4_3[10] , \wRegInTop_5_12[4] , \wRegInTop_5_8[7] , 
        \wRegOut_5_3[1] , \wRegInTop_1_1[8] , \wRegEnTop_2_3[0] , 
        \wRegOut_3_0[6] , \wRegInBot_4_7[21] , \ScanLink28[6] , 
        \wRegOut_5_1[26] , \wRegInTop_5_14[25] , \ScanLink35[9] , 
        \wRegInTop_5_22[20] , \wRegOut_5_27[9] , \wRegInBot_4_7[8] , 
        \wRegInTop_4_14[7] , \wRegOut_5_0[2] , \wRegInTop_4_2[18] , 
        \wRegInBot_4_7[12] , \ScanLink29[18] , \ScanLink3[8] , 
        \wRegInTop_2_0[4] , \wRegInBot_2_0[18] , \wRegOut_5_27[31] , 
        \wRegOut_5_27[28] , \wRegInBot_2_1[2] , \wRegOut_2_2[10] , 
        \wRegInBot_2_2[1] , \wRegInBot_4_2[5] , \wRegInTop_4_3[3] , 
        \ScanLink22[14] , \ScanLink30[4] , \wRegOut_5_1[15] , 
        \wRegInTop_5_14[16] , \wRegInTop_5_22[13] , \ScanLink57[24] , 
        \wRegOut_5_22[4] , \ScanLink61[21] , \wRegInTop_2_3[7] , 
        \ScanLink14[11] , \wRegInBot_3_4[17] , \wRegInTop_4_9[14] , 
        \ScanLink37[20] , \ScanLink42[10] , \wRegOut_4_14[11] , 
        \wRegOut_3_6[8] , \wRegInTop_4_0[0] , \wRegInTop_5_6[17] , 
        \wRegInBot_4_1[6] , \ScanLink33[7] , \wRegOut_5_21[7] , 
        \wRegInTop_4_12[9] , \wRegInBot_2_1[12] , \wRegOut_2_2[23] , 
        \ScanLink8[3] , \wRegInBot_3_4[24] , \wRegOut_4_5[30] , 
        \wRegOut_4_5[29] , \wRegOut_4_14[22] , \ScanLink14[22] , 
        \ScanLink22[27] , \wRegInTop_4_9[27] , \ScanLink37[13] , 
        \ScanLink61[12] , \ScanLink42[23] , \ScanLink54[0] , 
        \wRegInTop_4_11[19] , \ScanLink57[17] , \ScanLink57[3] , 
        \wRegInTop_5_6[24] , \wRegInTop_5_23[19] , \ScanLink41[7] , 
        \wRegOut_5_10[27] , \wRegInBot_2_1[21] , \wRegOut_3_7[15] , 
        \wRegInBot_4_6[18] , \ScanLink42[4] , \wRegOut_5_26[22] , 
        \wRegInTop_4_3[12] , \ScanLink28[12] , \ScanLink48[16] , 
        \ScanLink25[3] , \wRegOut_3_7[26] , \wRegInTop_4_3[21] , 
        \wRegInTop_4_8[8] , \ScanLink48[25] , \ScanLink26[0] , 
        \ScanLink28[21] , \wRegOut_4_15[6] , \wRegOut_5_26[11] , 
        \wRegOut_5_10[14] , \wRegInTop_5_26[8] , \wRegOut_1_1[5] , 
        \ScanLink3[24] , \ScanLink5[6] , \ScanLink6[5] , \wRegOut_2_3[30] , 
        \wRegOut_2_3[29] , \ScanLink7[26] , \ScanLink15[31] , 
        \wRegInTop_4_10[13] , \wRegInBot_4_10[14] , \ScanLink47[9] , 
        \wRegInTop_5_28[26] , \ScanLink15[28] , \ScanLink36[19] , 
        \ScanLink43[29] , \ScanLink7[15] , \wRegInTop_3_0[24] , 
        \ScanLink43[30] , \ScanLink60[18] , \wRegOut_4_4[23] , \ScanLink59[5] , 
        \wRegInTop_4_10[20] , \wRegInBot_4_10[27] , \wRegOut_4_15[31] , 
        \wRegOut_4_15[28] , \wRegInTop_5_28[15] , \wRegInTop_5_23[5] , 
        \wRegInTop_3_0[17] , \wRegOut_4_4[10] , \wRegInTop_3_3[8] , 
        \wRegInTop_3_4[26] , \wRegOut_4_0[21] , \wRegOut_4_13[8] , 
        \wRegInTop_5_20[6] , \ScanLink19[7] , \wRegOut_4_5[0] , 
        \wRegOut_4_6[3] , \wRegInBot_4_9[25] , \wRegInBot_4_14[16] , 
        \wRegOut_5_16[8] , \wRegInTop_4_14[11] , \ScanLink47[18] , 
        \ScanLink11[19] , \ScanLink32[31] , \ScanLink32[28] , 
        \wRegInTop_3_4[15] , \wRegInBot_4_9[16] , \wRegInBot_4_11[8] , 
        \ScanLink3[17] , \wRegOut_4_0[12] , \wRegOut_4_11[19] , 
        \wRegInTop_4_14[22] , \wRegInBot_0_0[8] , \wRegInBot_0_0[1] , 
        \wRegOut_2_0[9] , \wRegOut_3_3[17] , \wRegInTop_4_7[10] , 
        \wRegInBot_4_14[25] , \ScanLink39[24] , \wRegInBot_3_4[0] , 
        \wRegInTop_3_5[6] , \wRegOut_5_22[20] , \ScanLink59[20] , 
        \wRegInTop_3_6[5] , \wRegInTop_5_5[2] , \wRegOut_5_14[25] , 
        \wRegOut_5_10[6] , \wRegInBot_3_7[3] , \wRegInTop_5_8[13] , 
        \wRegOut_5_13[5] , \wRegInTop_5_6[1] , \wRegOut_5_14[16] , 
        \ScanLink0[2] , \wRegInTop_2_0[30] , \wRegOut_3_3[24] , 
        \wRegOut_5_22[13] , \wRegInBot_4_2[30] , \wRegInBot_4_2[29] , 
        \wRegInTop_4_7[23] , \ScanLink39[17] , \ScanLink59[13] , 
        \wRegInTop_5_27[31] , \wRegInTop_5_27[28] , \wRegInTop_2_0[29] , 
        \wRegInBot_2_1[31] , \wRegOut_2_3[20] , \wRegOut_2_3[13] , 
        \ScanLink8[31] , \ScanLink8[28] , \ScanLink23[4] , \wRegOut_4_10[2] , 
        \wRegInTop_4_10[30] , \wRegInTop_4_10[29] , \wRegInBot_4_14[5] , 
        \wRegInTop_5_8[20] , \wRegOut_5_31[4] , \wRegInTop_5_7[14] , 
        \wRegInBot_3_5[14] , \wRegEnBot_4_9[0] , \wRegOut_5_8[3] , 
        \ScanLink15[12] , \wRegOut_4_4[19] , \wRegInTop_4_8[17] , 
        \wRegOut_4_15[12] , \ScanLink36[23] , \ScanLink43[13] , 
        \ScanLink60[22] , \ScanLink20[7] , \ScanLink56[27] , \ScanLink23[17] , 
        \wRegOut_4_13[1] , \wRegInBot_3_5[27] , \ScanLink15[21] , 
        \ScanLink23[24] , \wRegInTop_5_7[27] , \ScanLink47[0] , 
        \wRegInTop_4_8[24] , \ScanLink36[10] , \ScanLink56[14] , 
        \ScanLink43[20] , \ScanLink44[3] , \wRegOut_4_15[21] , 
        \ScanLink60[11] , \wRegInTop_5_25[2] , \wRegInBot_2_1[28] , 
        \wRegOut_5_0[25] , \wRegInTop_5_23[23] , \wRegInTop_4_3[31] , 
        \wRegInTop_4_3[28] , \wRegInBot_4_6[22] , \ScanLink28[31] , 
        \ScanLink38[5] , \wRegInTop_5_15[26] , \ScanLink28[28] , 
        \wRegOut_5_29[6] , \wRegInTop_4_8[1] , \wRegInBot_4_9[7] , 
        \ScanLink26[9] , \wRegInTop_5_26[1] , \wRegOut_5_0[16] , 
        \wRegInTop_5_15[15] , \wRegOut_5_26[18] , \wRegInTop_5_23[10] , 
        \wRegOut_1_0[18] , \ScanLink3[1] , \wRegInBot_4_6[11] , 
        \wRegOut_2_0[0] , \wRegInTop_2_0[20] , \wRegInBot_4_2[20] , 
        \wRegInTop_5_11[24] , \wRegOut_2_3[3] , \ScanLink8[21] , 
        \wRegOut_5_4[27] , \wRegInTop_5_27[21] , \wRegInTop_5_8[30] , 
        \wRegInTop_5_8[29] , \wRegInBot_4_2[13] , \wRegInTop_4_7[19] , 
        \ScanLink59[30] , \ScanLink59[29] , \wRegInBot_3_4[9] , 
        \wRegOut_5_22[30] , \wRegOut_5_22[29] , \wRegOut_4_3[7] , 
        \wRegInTop_2_0[13] , \ScanLink8[12] , \wRegEnBot_3_2[0] , 
        \wRegInTop_5_6[8] , \wRegOut_4_0[4] , \wRegOut_5_4[14] , 
        \wRegInTop_5_27[12] , \wRegInTop_5_11[17] , \wRegInBot_3_1[16] , 
        \ScanLink11[10] , \wRegInBot_4_11[1] , \ScanLink27[15] , 
        \ScanLink52[25] , \ScanLink60[5] , \ScanLink32[21] , \ScanLink47[11] , 
        \wRegOut_4_11[10] , \wRegOut_0_0[15] , \wRegInBot_4_12[2] , 
        \wRegInTop_5_3[16] , \wRegOut_5_29[25] , \ScanLink63[6] , 
        \wRegOut_0_0[26] , \wRegInBot_3_1[25] , \wRegOut_4_0[28] , 
        \wRegOut_4_11[23] , \wRegOut_5_29[16] , \wRegInBot_3_2[7] , 
        \wRegInTop_3_3[1] , \ScanLink11[23] , \wRegOut_4_0[31] , 
        \wRegInTop_5_19[6] , \ScanLink32[12] , \ScanLink47[22] , 
        \wRegOut_5_16[1] , \wRegInTop_5_3[5] , \wRegOut_4_5[9] , 
        \ScanLink27[26] , \wRegInTop_4_14[18] , \wRegInTop_5_0[6] , 
        \ScanLink52[16] , \wRegOut_5_15[2] , \wRegEnBot_1_0[0] , 
        \ScanLink2[27] , \wRegInTop_2_1[19] , \wRegInTop_3_0[2] , 
        \wRegInBot_3_1[4] , \wRegInTop_5_3[25] , \wRegInTop_5_26[18] , 
        \ScanLink9[18] , \wRegOut_3_2[27] , \wRegOut_3_2[14] , \ScanLink11[6] , 
        \ScanLink12[5] , \wRegInTop_5_9[10] , \wRegInBot_4_3[19] , 
        \wRegOut_5_15[26] , \wRegOut_5_23[23] , \ScanLink58[23] , 
        \wRegInTop_4_6[20] , \wRegInTop_4_6[13] , \ScanLink38[27] , 
        \ScanLink38[14] , \wRegInTop_5_9[23] , \ScanLink58[10] , 
        \wRegOut_5_15[15] , \wRegOut_5_23[10] , \wRegOut_5_18[7] , 
        \ScanLink2[14] , \ScanLink10[30] , \ScanLink10[29] , \ScanLink17[8] , 
        \wRegInTop_4_15[12] , \wRegInBot_4_15[15] , \wRegInTop_5_17[0] , 
        \ScanLink46[31] , \wRegInTop_3_5[25] , \wRegInBot_4_8[26] , 
        \ScanLink33[18] , \wRegInTop_5_14[3] , \ScanLink46[28] , 
        \wRegOut_4_1[22] , \wRegOut_4_10[30] , \wRegOut_4_10[29] , 
        \wRegInTop_4_15[21] , \wRegInBot_4_15[26] , \wRegInTop_3_1[27] , 
        \wRegInTop_3_5[16] , \wRegOut_4_1[11] , \wRegOut_4_5[20] , 
        \wRegInBot_4_8[15] , \wRegInBot_4_11[17] , \ScanLink49[6] , 
        \ScanLink54[9] , \wRegInTop_5_29[25] , \wRegInBot_2_2[8] , 
        \ScanLink6[25] , \wRegInTop_4_11[10] , \wRegEnTop_5_19[0] , 
        \wRegOut_5_5[6] , \ScanLink61[28] , \ScanLink14[18] , \ScanLink37[30] , 
        \wRegInTop_4_11[3] , \ScanLink37[29] , \ScanLink42[19] , 
        \ScanLink61[31] , \wRegInTop_5_30[5] , \wRegOut_0_0[18] , 
        \wRegInBot_0_0[5] , \wRegInBot_1_0[7] , \wRegOut_2_2[19] , 
        \wRegInTop_3_1[14] , \wRegOut_3_5[2] , \wRegEnTop_4_6[0] , 
        \wRegOut_4_5[13] , \wRegOut_4_14[18] , \ScanLink6[16] , 
        \wRegOut_3_6[16] , \wRegOut_3_6[1] , \wRegInTop_4_0[9] , 
        \wRegInTop_4_11[23] , \wRegOut_5_6[5] , \wRegInTop_4_12[0] , 
        \wRegInTop_4_2[11] , \wRegInBot_4_11[24] , \ScanLink49[15] , 
        \wRegInTop_5_29[16] , \ScanLink29[11] , \wRegOut_5_27[21] , 
        \wRegOut_1_1[21] , \wRegOut_1_1[12] , \wRegInTop_1_1[1] , 
        \wRegInBot_2_0[11] , \wRegOut_5_11[24] , \ScanLink52[7] , 
        \ScanLink51[4] , \wRegInBot_2_0[22] , \wRegOut_3_6[25] , 
        \wRegInBot_4_4[2] , \wRegInTop_4_5[4] , \wRegOut_5_3[8] , 
        \wRegOut_5_11[17] , \wRegInBot_4_7[31] , \ScanLink29[22] , 
        \ScanLink36[3] , \wRegOut_5_24[3] , \wRegOut_5_27[12] , 
        \wRegInTop_4_2[22] , \wRegInBot_4_7[28] , \ScanLink49[26] , 
        \wRegInTop_5_22[30] , \wRegOut_3_3[20] , \wRegOut_3_3[13] , 
        \wRegInBot_3_4[4] , \wRegInTop_3_5[2] , \wRegInTop_3_6[1] , 
        \wRegInTop_4_6[7] , \ScanLink35[0] , \wRegInTop_5_22[29] , 
        \wRegInTop_5_28[7] , \wRegOut_5_27[0] , \wRegInBot_4_7[1] , 
        \wRegOut_5_4[19] , \wRegInTop_5_6[5] , \wRegInTop_5_8[17] , 
        \wRegOut_5_13[1] , \wRegInBot_3_7[7] , \wRegOut_4_0[9] , 
        \wRegInTop_5_5[6] , \wRegOut_5_10[2] , \wRegOut_5_14[21] , 
        \wRegOut_5_22[24] , \ScanLink59[24] , \wRegInTop_4_7[27] , 
        \wRegInTop_4_7[14] , \ScanLink39[20] , \wRegInBot_4_14[1] , 
        \wRegInTop_5_8[24] , \ScanLink39[13] , \wRegInTop_5_11[30] , 
        \wRegInTop_5_11[29] , \ScanLink59[17] , \ScanLink3[20] , 
        \wRegInTop_5_3[31] , \wRegInTop_5_3[28] , \wRegOut_5_14[12] , 
        \wRegOut_5_22[17] , \wRegInBot_3_1[31] , \wRegInBot_3_1[9] , 
        \wRegInTop_4_14[15] , \wRegInBot_4_14[12] , \wRegInTop_3_4[22] , 
        \wRegEnBot_3_7[0] , \wRegOut_4_5[4] , \wRegOut_4_6[7] , 
        \wRegInTop_5_3[8] , \wRegInBot_4_9[21] , \ScanLink19[3] , 
        \wRegInBot_3_1[28] , \wRegOut_4_0[25] , \wRegInBot_4_14[21] , 
        \wRegInTop_4_14[26] , \wRegOut_1_0[26] , \wRegOut_1_0[15] , 
        \wRegOut_1_1[1] , \ScanLink3[13] , \wRegInTop_3_4[11] , 
        \wRegOut_4_0[16] , \wRegOut_5_29[31] , \wRegInBot_4_9[12] , 
        \ScanLink27[18] , \ScanLink52[28] , \wRegOut_5_29[28] , 
        \ScanLink60[8] , \ScanLink52[31] , \ScanLink5[2] , \wRegInTop_3_0[20] , 
        \wRegOut_4_4[27] , \ScanLink23[30] , \ScanLink23[29] , \ScanLink59[1] , 
        \ScanLink56[19] , \wRegInTop_4_8[30] , \ScanLink6[1] , 
        \wRegInTop_4_8[29] , \wRegInBot_4_10[10] , \wRegInTop_5_28[22] , 
        \ScanLink7[22] , \wRegInTop_4_10[17] , \ScanLink7[11] , 
        \wRegInTop_3_0[13] , \wRegInTop_5_20[2] , \wRegInBot_3_5[19] , 
        \wRegOut_4_4[14] , \wRegInTop_5_7[19] , \wRegOut_3_7[11] , 
        \wRegInTop_4_3[16] , \ScanLink23[9] , \wRegInTop_4_10[24] , 
        \wRegInBot_4_10[23] , \wRegInTop_5_23[1] , \wRegInTop_5_28[11] , 
        \wRegOut_5_31[9] , \ScanLink48[12] , \ScanLink28[16] , 
        \wRegOut_5_26[26] , \wRegInBot_2_1[16] , \ScanLink41[3] , 
        \wRegOut_5_10[23] , \ScanLink42[0] , \wRegInTop_5_15[18] , 
        \wRegInTop_2_0[0] , \wRegInBot_2_1[25] , \wRegOut_3_7[22] , 
        \ScanLink26[4] , \wRegOut_5_10[10] , \ScanLink28[25] , 
        \wRegOut_4_15[2] , \wRegOut_5_26[15] , \wRegInTop_4_3[25] , 
        \wRegOut_5_0[28] , \ScanLink48[21] , \wRegInBot_2_1[6] , 
        \ScanLink25[7] , \wRegOut_5_0[31] , \ScanLink38[8] , \wRegOut_5_6[8] , 
        \wRegOut_2_2[14] , \wRegInTop_4_0[4] , \wRegInBot_4_11[30] , 
        \ScanLink33[3] , \wRegOut_5_21[3] , \wRegInBot_4_1[2] , 
        \wRegInBot_4_11[29] , \wRegInTop_5_6[13] , \wRegInBot_2_2[5] , 
        \wRegInTop_3_1[19] , \wRegInBot_3_4[13] , \wRegInTop_4_9[10] , 
        \wRegOut_4_14[15] , \ScanLink37[24] , \ScanLink42[14] , 
        \ScanLink61[25] , \wRegInTop_2_3[3] , \ScanLink14[15] , 
        \wRegInBot_4_2[1] , \wRegInTop_4_3[7] , \wRegInTop_5_30[8] , 
        \wRegInBot_1_0[3] , \ScanLink2[19] , \wRegInTop_2_1[27] , 
        \wRegOut_2_2[27] , \ScanLink6[31] , \ScanLink22[10] , \ScanLink30[0] , 
        \ScanLink57[20] , \wRegOut_5_22[0] , \ScanLink6[28] , \wRegOut_3_0[2] , 
        \ScanLink8[7] , \wRegInBot_3_4[20] , \ScanLink14[26] , 
        \ScanLink22[23] , \wRegInTop_5_6[20] , \ScanLink57[7] , 
        \wRegInTop_5_29[31] , \wRegInTop_5_29[28] , \wRegInTop_4_9[23] , 
        \ScanLink37[17] , \ScanLink57[13] , \ScanLink42[27] , \ScanLink54[4] , 
        \wRegOut_4_14[26] , \ScanLink61[16] , \wRegEnTop_4_3[0] , 
        \wRegInTop_4_14[3] , \wRegOut_5_0[6] , \wRegOut_3_3[1] , 
        \wRegOut_3_6[31] , \wRegOut_3_6[28] , \ScanLink28[2] , 
        \wRegOut_5_1[22] , \wRegInTop_5_22[24] , \wRegInTop_5_14[21] , 
        \wRegInBot_4_7[25] , \wRegInTop_4_5[9] , \wRegOut_5_3[5] , 
        \wRegInBot_4_3[27] , \wRegInBot_4_7[16] , \wRegOut_5_1[11] , 
        \wRegInTop_5_14[12] , \wRegInTop_5_22[17] , \wRegOut_5_11[30] , 
        \wRegOut_5_11[29] , \ScanLink51[9] , \ScanLink49[18] , 
        \ScanLink38[19] , \wRegOut_5_15[18] , \wRegInTop_5_10[23] , 
        \wRegInTop_2_1[14] , \ScanLink9[26] , \wRegOut_5_5[20] , 
        \wRegInTop_5_26[26] , \ScanLink9[15] , \wRegOut_3_2[19] , 
        \wRegInBot_4_3[14] , \ScanLink12[8] , \wRegInTop_5_8[3] , 
        \wRegInTop_5_12[0] , \wRegOut_5_5[13] , \wRegInTop_5_11[3] , 
        \wRegInTop_5_26[15] , \wRegInTop_5_10[10] , \wRegInBot_3_0[11] , 
        \ScanLink10[17] , \wRegInBot_4_8[18] , \ScanLink26[12] , 
        \ScanLink53[22] , \ScanLink33[26] , \ScanLink46[16] , 
        \wRegOut_4_10[17] , \wRegOut_5_28[22] , \wRegOut_1_1[16] , 
        \wRegInBot_2_0[15] , \wRegInBot_3_0[22] , \wRegInTop_3_5[31] , 
        \wRegInTop_3_5[28] , \wRegInTop_5_2[11] , \wRegOut_5_28[11] , 
        \wRegOut_4_10[24] , \ScanLink10[24] , \ScanLink14[6] , 
        \wRegOut_4_8[1] , \ScanLink33[15] , \ScanLink46[25] , \ScanLink17[5] , 
        \ScanLink26[21] , \ScanLink53[11] , \wRegInBot_4_15[18] , 
        \wRegInTop_5_2[22] , \wRegOut_5_1[18] , \wRegOut_5_11[20] , 
        \ScanLink51[0] , \wRegOut_1_1[25] , \wRegInTop_1_1[5] , 
        \wRegInBot_2_0[26] , \wRegOut_3_6[12] , \ScanLink52[3] , 
        \wRegOut_5_27[25] , \wRegInTop_4_2[15] , \ScanLink29[15] , 
        \ScanLink49[11] , \wRegInTop_4_6[3] , \wRegInBot_4_7[5] , 
        \ScanLink35[4] , \wRegOut_5_27[4] , \wRegInTop_5_14[31] , 
        \wRegInTop_5_14[28] , \wRegOut_3_3[8] , \wRegOut_3_6[21] , 
        \wRegInTop_4_2[26] , \wRegInTop_5_28[3] , \ScanLink49[22] , 
        \wRegInBot_4_4[6] , \wRegInTop_4_5[0] , \ScanLink29[26] , 
        \ScanLink36[7] , \wRegOut_5_24[7] , \wRegOut_5_27[16] , 
        \wRegOut_5_11[13] , \wRegInTop_2_0[9] , \ScanLink6[21] , 
        \wRegInTop_5_6[30] , \wRegInTop_5_6[29] , \wRegInTop_3_1[23] , 
        \wRegInTop_4_11[14] , \wRegInBot_4_11[13] , \wRegInTop_5_29[21] , 
        \wRegInBot_3_4[30] , \wRegInBot_3_4[29] , \wRegOut_4_5[24] , 
        \ScanLink49[2] , \wRegOut_3_6[5] , \wRegInBot_4_11[20] , 
        \wRegInTop_5_29[12] , \wRegInTop_4_11[27] , \wRegOut_5_6[1] , 
        \wRegInTop_4_12[4] , \ScanLink6[12] , \wRegInTop_3_1[10] , 
        \wRegOut_4_5[17] , \wRegOut_3_5[6] , \wRegEnBot_4_12[0] , 
        \ScanLink57[30] , \wRegInBot_4_2[8] , \ScanLink57[29] , 
        \wRegOut_0_0[11] , \ScanLink2[23] , \wRegInTop_3_5[21] , 
        \wRegOut_4_1[26] , \ScanLink22[19] , \ScanLink30[9] , 
        \wRegOut_5_22[9] , \wRegInTop_4_9[19] , \wRegInTop_4_11[7] , 
        \wRegOut_5_5[2] , \wRegInTop_5_30[1] , \wRegOut_4_8[8] , 
        \wRegInBot_4_8[22] , \ScanLink26[31] , \wRegOut_5_28[18] , 
        \wRegInTop_5_14[7] , \ScanLink26[28] , \wRegInTop_4_15[16] , 
        \wRegInBot_4_15[11] , \ScanLink53[18] , \wRegInTop_5_17[4] , 
        \ScanLink2[10] , \wRegInBot_3_0[18] , \wRegInTop_3_5[12] , 
        \wRegInBot_4_8[11] , \wRegOut_5_18[3] , \wRegOut_4_1[15] , 
        \wRegInTop_5_2[18] , \wRegOut_3_2[23] , \wRegOut_3_2[10] , 
        \wRegInTop_4_6[17] , \wRegInTop_4_15[25] , \wRegInBot_4_15[22] , 
        \ScanLink38[23] , \ScanLink11[2] , \ScanLink12[1] , 
        \wRegInTop_5_12[9] , \wRegOut_5_23[27] , \ScanLink58[27] , 
        \wRegOut_5_15[22] , \wRegInTop_5_9[14] , \wRegInTop_5_10[19] , 
        \wRegOut_5_15[11] , \wRegOut_5_23[14] , \wRegInTop_4_6[24] , 
        \ScanLink38[10] , \ScanLink58[14] , \wRegInBot_4_14[28] , 
        \wRegOut_5_5[30] , \wRegEnTop_5_25[0] , \wRegOut_5_5[29] , 
        \wRegInTop_5_9[27] , \wRegInBot_4_12[6] , \wRegInBot_4_14[31] , 
        \ScanLink63[2] , \wRegInTop_5_3[12] , \wRegOut_0_0[22] , 
        \wRegOut_1_1[8] , \wRegInBot_3_1[12] , \wRegInTop_3_4[18] , 
        \wRegOut_5_29[21] , \ScanLink11[14] , \wRegOut_4_11[14] , 
        \ScanLink47[15] , \ScanLink3[30] , \ScanLink3[29] , 
        \wRegInBot_4_11[5] , \ScanLink32[25] , \ScanLink27[11] , 
        \ScanLink52[21] , \ScanLink60[1] , \wRegInTop_3_0[6] , 
        \wRegInTop_5_3[21] , \wRegInBot_3_1[0] , \wRegInBot_3_1[21] , 
        \wRegInBot_3_2[3] , \wRegInTop_3_3[5] , \wRegInBot_4_9[31] , 
        \ScanLink27[22] , \wRegInTop_5_0[2] , \wRegOut_5_15[6] , 
        \ScanLink52[12] , \ScanLink11[27] , \wRegInBot_4_9[28] , 
        \wRegOut_4_11[27] , \ScanLink32[16] , \wRegInTop_5_3[1] , 
        \ScanLink47[26] , \wRegOut_5_16[5] , \wRegInTop_5_19[2] , 
        \ScanLink0[6] , \ScanLink3[5] , \wRegOut_2_0[4] , \wRegInTop_2_0[24] , 
        \ScanLink8[25] , \wRegOut_5_29[12] , \wRegInBot_4_14[8] , 
        \wRegOut_5_4[23] , \wRegInTop_5_27[25] , \wRegInTop_2_0[17] , 
        \wRegOut_3_3[30] , \wRegInTop_5_11[20] , \wRegOut_3_3[29] , 
        \wRegInBot_4_2[24] , \wRegInTop_3_6[8] , \wRegOut_5_4[10] , 
        \wRegInTop_5_11[13] , \wRegInTop_5_27[16] , \wRegOut_4_0[0] , 
        \wRegOut_2_3[7] , \ScanLink8[16] , \wRegOut_4_3[3] , \wRegOut_5_13[8] , 
        \wRegOut_5_14[31] , \wRegOut_5_14[28] , \wRegOut_3_7[18] , 
        \wRegInBot_4_2[17] , \ScanLink39[30] , \ScanLink39[29] , 
        \wRegInBot_4_6[26] , \wRegInTop_4_8[5] , \wRegOut_5_10[19] , 
        \wRegInTop_5_26[5] , \wRegInBot_4_9[3] , \ScanLink48[31] , 
        \ScanLink48[28] , \wRegOut_5_29[2] , \wRegInBot_4_6[15] , 
        \wRegOut_5_0[21] , \ScanLink38[1] , \wRegInTop_5_15[22] , 
        \wRegInTop_5_23[27] , \wRegInTop_5_25[6] , \ScanLink42[9] , 
        \ScanLink6[8] , \wRegOut_2_3[17] , \wRegInBot_3_5[10] , 
        \ScanLink15[16] , \ScanLink20[3] , \wRegOut_5_0[12] , 
        \wRegInTop_5_15[11] , \wRegInTop_5_23[14] , \ScanLink56[23] , 
        \ScanLink23[13] , \wRegOut_4_13[5] , \ScanLink60[26] , 
        \wRegInTop_4_8[13] , \ScanLink36[27] , \ScanLink43[17] , 
        \wRegOut_4_15[16] , \wRegOut_5_8[7] , \ScanLink7[18] , 
        \wRegInTop_3_0[30] , \ScanLink23[0] , \wRegOut_4_10[6] , 
        \wRegInTop_5_7[10] , \wRegOut_5_31[0] , \wRegInTop_5_23[8] , 
        \wRegInTop_5_28[18] , \wRegInTop_3_0[29] , \wRegInBot_3_5[23] , 
        \wRegOut_4_15[25] , \ScanLink59[8] , \ScanLink15[25] , 
        \ScanLink23[20] , \wRegInTop_4_8[20] , \ScanLink36[14] , 
        \ScanLink60[15] , \ScanLink43[24] , \ScanLink44[7] , \ScanLink47[4] , 
        \ScanLink56[10] , \wRegOut_2_3[24] , \wRegInBot_4_10[19] , 
        \wRegInTop_5_7[23] , \wRegInBot_3_1[10] , \ScanLink11[16] , 
        \wRegInBot_4_9[19] , \wRegInBot_4_11[7] , \ScanLink27[13] , 
        \ScanLink60[3] , \ScanLink52[23] , \wRegOut_4_11[16] , 
        \wRegEnTop_4_12[0] , \ScanLink32[27] , \ScanLink47[17] , 
        \wRegOut_0_0[13] , \ScanLink3[18] , \wRegOut_5_29[23] , 
        \wRegInBot_4_12[4] , \wRegInTop_5_3[10] , \ScanLink63[0] , 
        \wRegInTop_3_4[30] , \wRegOut_0_0[20] , \wRegInTop_3_0[4] , 
        \wRegInBot_3_1[23] , \wRegInTop_3_4[29] , \ScanLink19[8] , 
        \wRegOut_5_29[10] , \wRegInTop_5_19[0] , \wRegInBot_3_1[2] , 
        \wRegInBot_3_2[1] , \ScanLink11[25] , \wRegOut_4_11[25] , 
        \wRegInTop_5_3[3] , \ScanLink27[20] , \ScanLink32[14] , 
        \ScanLink47[24] , \wRegOut_5_16[7] , \ScanLink52[10] , 
        \wRegInTop_3_3[7] , \wRegInTop_5_0[0] , \wRegOut_5_15[4] , 
        \wRegInBot_4_14[19] , \ScanLink0[4] , \wRegOut_2_0[6] , 
        \wRegInTop_2_0[26] , \wRegInBot_4_2[26] , \wRegInTop_5_3[23] , 
        \ScanLink39[18] , \wRegOut_5_14[19] , \wRegOut_2_3[5] , 
        \ScanLink8[27] , \wRegOut_5_4[21] , \wRegInTop_5_11[22] , 
        \wRegInTop_5_27[27] , \wRegOut_3_3[18] , \wRegInBot_4_2[15] , 
        \wRegOut_5_10[9] , \ScanLink8[14] , \wRegInTop_3_5[9] , 
        \wRegOut_4_3[1] , \wRegInTop_2_0[15] , \wRegEnTop_3_3[0] , 
        \wRegOut_4_0[2] , \wRegOut_5_4[12] , \wRegInTop_5_27[14] , 
        \wRegOut_3_7[30] , \wRegOut_5_0[23] , \wRegInTop_5_11[11] , 
        \wRegInTop_5_25[4] , \ScanLink38[3] , \wRegInTop_5_23[25] , 
        \wRegInTop_5_15[20] , \wRegOut_3_7[29] , \wRegInBot_4_6[24] , 
        \wRegInTop_4_8[7] , \wRegInBot_4_9[1] , \wRegOut_4_15[9] , 
        \wRegInTop_5_26[7] , \wRegOut_5_29[0] , \wRegOut_5_0[10] , 
        \wRegInTop_5_15[13] , \wRegInTop_5_23[16] , \wRegInBot_1_0[1] , 
        \wRegInTop_1_1[7] , \ScanLink3[7] , \ScanLink41[8] , 
        \wRegOut_5_10[31] , \wRegOut_5_10[28] , \ScanLink5[9] , 
        \wRegOut_2_3[26] , \wRegOut_2_3[15] , \wRegInBot_4_6[17] , 
        \ScanLink48[19] , \ScanLink23[2] , \wRegOut_4_10[4] , 
        \wRegInBot_4_10[28] , \wRegOut_5_31[2] , \wRegInBot_4_10[31] , 
        \wRegInTop_5_7[12] , \wRegInTop_3_0[18] , \wRegEnTop_4_8[0] , 
        \wRegOut_5_8[5] , \wRegInBot_3_5[12] , \wRegOut_4_15[14] , 
        \ScanLink15[14] , \ScanLink20[1] , \wRegInTop_4_8[11] , 
        \wRegInTop_5_20[9] , \ScanLink60[24] , \ScanLink36[25] , 
        \ScanLink43[15] , \ScanLink23[11] , \wRegOut_4_13[7] , 
        \ScanLink56[21] , \ScanLink7[30] , \ScanLink7[29] , \ScanLink15[27] , 
        \ScanLink23[22] , \wRegInTop_5_7[21] , \ScanLink47[6] , 
        \wRegInTop_5_28[30] , \wRegInTop_5_28[29] , \ScanLink56[12] , 
        \ScanLink60[17] , \wRegInBot_3_5[21] , \wRegInTop_4_8[22] , 
        \ScanLink43[26] , \ScanLink44[5] , \ScanLink36[16] , \wRegOut_3_6[10] , 
        \wRegInTop_4_2[17] , \wRegOut_4_15[27] , \wRegEnTop_5_17[0] , 
        \ScanLink49[13] , \ScanLink29[17] , \wRegOut_5_11[22] , 
        \wRegOut_5_27[27] , \ScanLink52[1] , \wRegOut_1_1[27] , 
        \wRegOut_1_1[14] , \wRegInBot_2_0[17] , \wRegInTop_5_14[19] , 
        \ScanLink51[2] , \wRegOut_5_11[11] , \wRegEnTop_1_1[0] , 
        \wRegInBot_2_0[24] , \wRegOut_3_6[23] , \wRegInBot_4_4[4] , 
        \ScanLink36[5] , \wRegOut_5_24[5] , \wRegOut_5_27[14] , 
        \wRegInTop_4_5[2] , \wRegInTop_4_2[24] , \ScanLink29[24] , 
        \ScanLink49[20] , \wRegOut_5_1[30] , \wRegOut_5_1[29] , 
        \wRegInTop_5_28[1] , \wRegOut_3_0[9] , \wRegInBot_4_7[7] , 
        \ScanLink28[9] , \wRegInTop_4_14[8] , \wRegInTop_3_1[21] , 
        \wRegOut_4_5[26] , \wRegInTop_4_6[1] , \ScanLink35[6] , 
        \wRegOut_5_27[6] , \ScanLink22[31] , \ScanLink49[0] , \ScanLink22[28] , 
        \ScanLink57[18] , \wRegInTop_4_9[31] , \wRegInTop_4_9[28] , 
        \wRegInTop_4_11[16] , \wRegInBot_4_11[11] , \wRegInTop_5_29[23] , 
        \ScanLink6[23] , \wRegInTop_2_3[8] , \wRegOut_3_5[4] , 
        \wRegInTop_4_11[5] , \wRegInTop_5_30[3] , \wRegOut_5_5[0] , 
        \wRegEnBot_4_7[0] , \wRegInBot_1_0[8] , \ScanLink2[21] , 
        \ScanLink6[10] , \wRegInTop_3_1[12] , \wRegInBot_3_4[18] , 
        \wRegOut_4_5[15] , \wRegInTop_5_6[18] , \wRegOut_3_6[7] , 
        \wRegInTop_4_11[25] , \wRegInTop_4_12[6] , \wRegOut_5_6[3] , 
        \ScanLink33[8] , \wRegOut_5_21[8] , \wRegInTop_5_29[10] , 
        \wRegInBot_4_1[9] , \wRegInBot_4_11[22] , \wRegInTop_5_2[30] , 
        \wRegInTop_5_2[29] , \wRegOut_5_18[1] , \ScanLink2[12] , 
        \wRegInBot_3_0[30] , \wRegInBot_3_0[29] , \wRegInTop_3_5[23] , 
        \wRegInBot_4_8[20] , \wRegInTop_4_15[14] , \wRegInBot_4_15[13] , 
        \wRegInTop_5_17[6] , \wRegInTop_5_14[5] , \wRegOut_4_1[24] , 
        \wRegInTop_4_15[27] , \wRegInBot_4_15[20] , \wRegInTop_2_0[2] , 
        \wRegOut_2_2[16] , \wRegInBot_2_2[7] , \wRegInTop_2_3[1] , 
        \wRegOut_3_2[21] , \wRegOut_3_2[12] , \ScanLink11[0] , 
        \wRegInTop_3_5[10] , \wRegOut_4_1[17] , \wRegInBot_4_8[13] , 
        \wRegOut_5_28[30] , \wRegOut_5_28[29] , \ScanLink26[19] , 
        \ScanLink53[30] , \wRegOut_5_5[18] , \ScanLink53[29] , \ScanLink12[3] , 
        \wRegInTop_5_9[16] , \wRegInTop_5_11[8] , \wRegOut_5_15[20] , 
        \wRegInTop_5_8[8] , \wRegOut_5_23[25] , \wRegInTop_4_6[26] , 
        \wRegInTop_4_6[15] , \ScanLink58[25] , \ScanLink38[21] , 
        \wRegInTop_5_9[25] , \wRegInTop_5_10[31] , \wRegInTop_5_10[28] , 
        \wEnable_3[0] , \ScanLink38[12] , \wRegInBot_4_2[3] , 
        \wRegOut_5_15[13] , \wRegOut_5_23[16] , \ScanLink58[16] , 
        \wRegInTop_4_3[5] , \ScanLink22[12] , \ScanLink30[2] , 
        \wRegOut_5_22[2] , \wRegInTop_4_9[12] , \ScanLink57[22] , 
        \ScanLink37[26] , \ScanLink42[16] , \ScanLink14[17] , \ScanLink61[27] , 
        \ScanLink6[19] , \wRegInBot_3_4[11] , \wRegOut_4_14[17] , 
        \wRegOut_5_5[9] , \wRegInTop_4_0[6] , \wRegInBot_4_1[0] , 
        \ScanLink33[1] , \wRegInTop_5_6[11] , \wRegOut_5_21[1] , 
        \wRegInTop_5_29[19] , \wRegInBot_2_1[4] , \wRegOut_2_2[25] , 
        \ScanLink8[5] , \wRegInTop_3_1[31] , \wRegInTop_3_1[28] , 
        \ScanLink49[9] , \wRegInBot_3_4[22] , \ScanLink14[24] , 
        \wRegInTop_4_9[21] , \wRegOut_4_14[24] , \ScanLink42[25] , 
        \ScanLink54[6] , \ScanLink37[15] , \ScanLink61[14] , \ScanLink22[21] , 
        \ScanLink57[11] , \wRegInBot_4_11[18] , \ScanLink57[5] , 
        \wRegInTop_5_6[22] , \wRegEnBot_2_2[0] , \wRegOut_3_0[0] , 
        \wRegOut_3_3[3] , \wRegInBot_4_7[27] , \wRegOut_5_3[7] , 
        \wRegOut_5_11[18] , \ScanLink49[30] , \ScanLink49[29] , 
        \ScanLink28[0] , \wRegInTop_5_14[23] , \wRegOut_5_1[20] , 
        \wRegInTop_5_22[26] , \wRegInTop_5_28[8] , \wRegInTop_4_6[8] , 
        \wRegInTop_4_14[1] , \wRegOut_5_0[4] , \wRegOut_3_6[19] , 
        \wRegInBot_4_7[14] , \ScanLink52[8] , \ScanLink2[31] , 
        \wRegInTop_2_1[25] , \ScanLink9[24] , \wRegOut_5_1[13] , 
        \wRegInTop_5_22[15] , \wRegInTop_5_14[10] , \wRegOut_5_5[22] , 
        \wRegInTop_5_26[24] , \wRegInTop_5_10[21] , \wRegInTop_2_1[16] , 
        \wRegOut_3_2[31] , \wRegOut_3_2[28] , \wRegInBot_4_3[25] , 
        \wRegInTop_5_10[12] , \wRegInBot_3_0[13] , \ScanLink9[17] , 
        \ScanLink11[9] , \wRegOut_5_5[11] , \wRegInTop_5_26[17] , 
        \wRegInTop_5_11[1] , \wRegInTop_3_5[19] , \wRegInBot_4_3[16] , 
        \ScanLink38[31] , \ScanLink38[28] , \wRegInTop_5_12[2] , 
        \wRegOut_5_15[30] , \wRegOut_5_15[29] , \wRegInTop_5_8[1] , 
        \wRegInBot_4_15[30] , \wRegInBot_4_15[29] , \wRegInTop_5_2[13] , 
        \wRegOut_4_10[15] , \wRegOut_5_28[20] , \ScanLink10[15] , 
        \ScanLink33[24] , \ScanLink46[14] , \ScanLink26[10] , \ScanLink53[20] , 
        \ScanLink2[28] , \wRegInBot_3_0[20] , \ScanLink10[26] , 
        \ScanLink14[4] , \ScanLink17[7] , \wRegInTop_5_2[20] , 
        \wRegOut_5_18[8] , \wRegInBot_4_8[30] , \wRegInBot_4_8[29] , 
        \ScanLink26[23] , \ScanLink53[13] , \ScanLink46[27] , \ScanLink33[17] , 
        \wRegOut_4_8[3] , \wRegOut_3_3[11] , \wRegInTop_4_7[16] , 
        \wRegOut_4_10[26] , \wRegOut_5_28[13] , \ScanLink39[22] , 
        \ScanLink59[26] , \wRegInBot_3_4[6] , \wRegOut_4_3[8] , 
        \wRegInTop_3_5[0] , \wRegInTop_3_6[3] , \wRegInBot_3_7[5] , 
        \wRegInTop_5_5[4] , \wRegOut_5_10[0] , \wRegOut_5_22[26] , 
        \wRegInTop_5_8[15] , \wRegOut_5_14[23] , \wRegInTop_5_6[7] , 
        \wRegOut_5_13[3] , \wRegOut_0_0[30] , \wRegInBot_0_0[7] , 
        \wRegInTop_5_11[18] , \wRegOut_5_14[10] , \wRegInBot_3_2[8] , 
        \wRegOut_3_3[22] , \wRegOut_5_22[15] , \ScanLink59[15] , 
        \wRegInTop_3_4[20] , \wRegOut_4_0[27] , \wRegInTop_4_7[25] , 
        \wRegInBot_4_14[3] , \wRegOut_5_4[31] , \wRegOut_5_4[28] , 
        \ScanLink39[11] , \wRegInTop_5_8[26] , \wRegInTop_5_19[9] , 
        \ScanLink19[1] , \ScanLink27[29] , \ScanLink52[19] , 
        \wRegOut_5_29[19] , \wRegOut_4_5[6] , \wRegOut_4_6[5] , 
        \wRegInBot_4_9[23] , \ScanLink27[30] , \wRegEnTop_5_6[0] , 
        \wRegOut_0_0[29] , \wRegInBot_4_14[10] , \wRegOut_1_1[3] , 
        \ScanLink3[22] , \wRegInTop_4_14[17] , \wRegInTop_5_0[9] , 
        \ScanLink3[11] , \wRegInBot_3_1[19] , \wRegInTop_3_4[13] , 
        \wRegInBot_4_9[10] , \wRegOut_4_0[14] , \wRegInTop_5_3[19] , 
        \wRegEnBot_0_0[0] , \wRegInTop_4_14[24] , \wRegInBot_4_14[23] , 
        \wRegOut_1_0[24] , \wRegOut_1_0[17] , \wRegInBot_2_1[14] , 
        \ScanLink5[0] , \ScanLink6[3] , \ScanLink7[20] , \wRegInTop_5_7[31] , 
        \wRegInTop_5_7[28] , \ScanLink63[9] , \wRegInTop_4_10[15] , 
        \wRegInBot_4_10[12] , \wRegInTop_5_28[20] , \ScanLink7[13] , 
        \wRegInTop_3_0[22] , \wRegInBot_3_5[31] , \ScanLink59[3] , 
        \wRegInBot_3_5[28] , \wRegOut_4_4[25] , \wRegInTop_4_10[26] , 
        \wRegInBot_4_10[21] , \wRegInTop_5_23[3] , \wRegInTop_5_28[13] , 
        \wRegInTop_3_0[11] , \wRegOut_4_4[16] , \ScanLink20[8] , 
        \ScanLink23[18] , \wRegInTop_4_8[18] , \wRegInTop_5_20[0] , 
        \ScanLink56[31] , \ScanLink56[28] , \wRegOut_5_0[19] , \ScanLink41[1] , 
        \ScanLink42[2] , \wRegInBot_2_1[27] , \wRegOut_3_7[13] , 
        \ScanLink28[14] , \wRegOut_5_10[21] , \wRegOut_5_26[24] , 
        \wRegInTop_4_3[14] , \ScanLink25[5] , \ScanLink48[10] , 
        \wRegInTop_5_15[30] , \wRegInTop_5_15[29] , \wRegOut_3_7[20] , 
        \wRegInTop_4_3[27] , \wRegInBot_4_9[8] , \ScanLink48[23] , 
        \wRegOut_5_29[9] , \ScanLink28[27] , \ScanLink26[6] , 
        \wRegOut_4_15[0] , \wRegOut_5_26[17] , \ScanLink2[25] , 
        \wRegInTop_2_1[31] , \wRegInTop_2_1[28] , \wRegOut_3_2[25] , 
        \wRegOut_3_2[16] , \wRegInTop_4_6[11] , \wRegOut_5_10[12] , 
        \ScanLink38[25] , \ScanLink58[21] , \ScanLink11[4] , \ScanLink12[7] , 
        \wRegOut_5_23[21] , \wRegInTop_5_9[12] , \wRegOut_5_15[24] , 
        \wRegInBot_4_3[31] , \wRegOut_5_15[17] , \wRegOut_5_23[12] , 
        \ScanLink58[12] , \wRegInBot_4_3[28] , \wRegInTop_4_6[22] , 
        \ScanLink38[16] , \wRegInTop_5_26[30] , \wRegInTop_5_26[29] , 
        \ScanLink9[30] , \ScanLink9[29] , \wRegInTop_3_5[27] , 
        \wRegOut_4_1[20] , \wRegInTop_5_9[21] , \ScanLink14[9] , 
        \wRegInBot_4_8[24] , \wRegInTop_5_14[1] , \wRegInTop_4_15[10] , 
        \wRegInBot_4_15[17] , \wRegInTop_5_17[2] , \ScanLink2[16] , 
        \ScanLink10[18] , \wRegOut_5_18[5] , \wRegInTop_3_5[14] , 
        \wRegInBot_4_8[17] , \ScanLink33[30] , \ScanLink33[29] , 
        \ScanLink46[19] , \wRegOut_4_1[13] , \wRegOut_4_10[18] , 
        \wRegInBot_2_1[9] , \wRegOut_2_2[31] , \wRegOut_2_2[28] , 
        \wRegInTop_4_15[23] , \wRegInBot_4_15[24] , \ScanLink6[27] , 
        \ScanLink8[8] , \ScanLink14[30] , \ScanLink14[29] , 
        \wRegInTop_4_11[12] , \ScanLink57[8] , \wRegInBot_4_11[15] , 
        \ScanLink42[31] , \wRegInTop_5_29[27] , \ScanLink61[19] , 
        \ScanLink37[18] , \ScanLink42[28] , \wRegInTop_3_1[25] , 
        \wRegOut_3_6[3] , \wRegOut_4_5[22] , \wRegOut_4_14[30] , 
        \ScanLink49[4] , \wRegOut_4_14[29] , \wRegInBot_4_11[26] , 
        \wRegInTop_4_12[2] , \wRegInTop_5_29[14] , \wRegOut_5_6[7] , 
        \ScanLink6[14] , \wRegInTop_4_11[21] , \wRegInTop_3_1[16] , 
        \wRegOut_4_5[11] , \wRegOut_0_0[17] , \ScanLink0[0] , 
        \wRegOut_1_0[30] , \wRegInBot_1_0[5] , \wRegOut_1_1[10] , 
        \wRegInTop_1_1[3] , \wRegInBot_2_0[13] , \wRegOut_3_5[0] , 
        \wRegInTop_4_3[8] , \wRegInTop_4_11[1] , \wRegInTop_5_30[7] , 
        \wRegOut_5_5[4] , \ScanLink51[6] , \wRegInTop_5_22[18] , 
        \ScanLink52[5] , \wRegOut_1_1[23] , \wRegInBot_2_0[20] , 
        \wRegOut_3_6[14] , \wRegInBot_4_7[19] , \ScanLink29[13] , 
        \wRegOut_5_11[26] , \wRegOut_5_27[23] , \wRegInTop_4_2[13] , 
        \wRegInTop_4_6[5] , \wRegInBot_4_7[3] , \ScanLink35[2] , 
        \ScanLink49[17] , \wRegOut_5_27[2] , \wRegOut_5_0[9] , 
        \wRegInTop_5_28[5] , \wRegOut_3_6[27] , \wRegInTop_4_2[20] , 
        \ScanLink49[24] , \ScanLink29[20] , \wRegInBot_4_4[0] , 
        \wRegInTop_4_5[6] , \ScanLink36[1] , \wRegOut_5_24[1] , 
        \wRegOut_5_27[10] , \wRegOut_2_3[22] , \wRegOut_2_3[11] , 
        \wRegInBot_3_5[16] , \ScanLink15[10] , \ScanLink20[5] , 
        \wRegOut_5_11[15] , \ScanLink23[15] , \wRegInTop_4_8[15] , 
        \wRegOut_4_13[3] , \ScanLink56[25] , \ScanLink36[21] , 
        \ScanLink43[11] , \wRegOut_4_15[10] , \ScanLink60[20] , 
        \wRegOut_5_8[1] , \wRegInBot_3_5[25] , \wRegOut_4_4[28] , 
        \ScanLink23[6] , \wRegOut_4_10[0] , \wRegInTop_5_7[16] , 
        \wRegOut_5_31[6] , \ScanLink15[23] , \wRegOut_4_4[31] , 
        \wRegOut_4_15[23] , \wRegInTop_4_8[26] , \ScanLink43[22] , 
        \ScanLink44[1] , \ScanLink36[12] , \ScanLink60[13] , \ScanLink23[26] , 
        \ScanLink56[16] , \wRegInTop_4_10[18] , \wRegInTop_5_7[25] , 
        \ScanLink47[2] , \wRegInTop_5_26[3] , \wRegOut_1_0[29] , 
        \ScanLink3[3] , \wRegInTop_4_3[19] , \wRegInBot_4_6[20] , 
        \wRegInTop_4_8[3] , \wRegInBot_4_9[5] , \wRegOut_5_29[4] , 
        \wRegInBot_4_6[13] , \ScanLink25[8] , \wRegOut_5_0[27] , 
        \ScanLink38[7] , \wRegInTop_5_15[24] , \wRegInTop_5_23[21] , 
        \wRegInTop_5_25[0] , \ScanLink28[19] , \wRegOut_5_26[30] , 
        \wRegOut_5_26[29] , \wRegOut_2_0[2] , \wRegInTop_2_0[22] , 
        \wRegInBot_2_1[19] , \wRegInTop_5_23[12] , \ScanLink8[23] , 
        \wRegOut_5_0[14] , \wRegInTop_5_15[17] , \wRegOut_5_4[25] , 
        \wRegInTop_5_27[23] , \wRegInTop_5_11[26] , \wRegInTop_2_0[11] , 
        \wRegInBot_4_2[22] , \wRegInTop_4_7[31] , \wRegInTop_4_7[28] , 
        \ScanLink59[18] , \wRegInTop_5_11[15] , \wRegOut_5_22[18] , 
        \ScanLink8[10] , \wRegInBot_3_7[8] , \wRegOut_5_4[16] , 
        \wRegInTop_5_27[10] , \wRegOut_4_0[6] , \wRegEnTop_5_3[0] , 
        \wRegInTop_5_8[18] , \wRegOut_2_3[1] , \wRegOut_4_3[5] , 
        \wRegInTop_5_5[9] , \wRegInBot_4_2[11] , \wRegInTop_4_14[30] , 
        \wRegInTop_4_14[29] , \ScanLink63[4] , \wRegInBot_4_12[0] , 
        \wRegInTop_5_3[14] , \wRegOut_0_0[24] , \wRegInBot_3_1[14] , 
        \wRegOut_4_11[12] , \wRegOut_5_29[27] , \ScanLink11[12] , 
        \wRegOut_4_0[19] , \ScanLink32[23] , \ScanLink47[13] , 
        \wRegInBot_4_11[3] , \ScanLink27[17] , \ScanLink60[7] , 
        \wRegInTop_5_3[27] , \ScanLink52[27] , \wRegInTop_3_0[0] , 
        \wRegInBot_3_1[6] , \wRegOut_4_6[8] , \wRegInBot_3_1[27] , 
        \wRegInBot_3_2[5] , \wRegInTop_5_0[4] , \wRegOut_5_15[0] , 
        \wRegInTop_3_3[3] , \ScanLink11[21] , \ScanLink27[24] , 
        \ScanLink52[14] , \ScanLink32[10] , \ScanLink47[20] , 
        \wRegOut_5_16[3] , \wRegInTop_5_3[7] , \wRegInTop_5_19[4] , 
        \wRegOut_4_11[21] , \ScanLink0[9] , \wRegOut_1_0[13] , 
        \wRegOut_3_7[17] , \wRegInTop_4_3[10] , \wRegOut_5_29[14] , 
        \ScanLink48[14] , \ScanLink28[10] , \wRegOut_5_10[25] , 
        \wRegOut_5_26[20] , \ScanLink42[6] , \ScanLink41[5] , 
        \wRegOut_1_0[20] , \wRegInBot_2_1[10] , \wRegEnTop_5_12[0] , 
        \wRegOut_5_10[16] , \ScanLink3[26] , \wRegInBot_2_1[23] , 
        \wRegOut_3_7[24] , \ScanLink26[2] , \wRegOut_4_15[4] , 
        \wRegOut_5_26[13] , \wRegInTop_4_3[23] , \wRegInBot_4_6[30] , 
        \wRegInBot_4_6[29] , \ScanLink28[23] , \ScanLink48[27] , 
        \wRegInTop_5_23[28] , \ScanLink5[4] , \wRegInTop_3_0[26] , 
        \wRegOut_4_4[21] , \ScanLink25[1] , \wRegInTop_5_23[31] , 
        \wRegInTop_5_25[9] , \ScanLink44[8] , \ScanLink59[7] , \ScanLink6[7] , 
        \wRegInTop_4_10[11] , \wRegInBot_4_10[16] , \wRegInTop_5_28[24] , 
        \wRegOut_2_3[18] , \ScanLink7[24] , \ScanLink7[17] , 
        \wRegInTop_3_0[15] , \ScanLink15[19] , \ScanLink36[28] , 
        \ScanLink43[18] , \ScanLink60[30] , \ScanLink36[31] , 
        \wRegInTop_5_20[4] , \ScanLink60[29] , \wRegOut_4_4[12] , 
        \wRegOut_5_8[8] , \wRegOut_4_15[19] , \wRegOut_4_10[9] , 
        \wRegInTop_4_10[22] , \wRegInTop_5_23[7] , \wRegInBot_4_10[25] , 
        \wRegInTop_5_28[17] , \wRegInTop_3_0[9] , \wRegOut_4_6[1] , 
        \wRegInTop_4_14[13] , \wRegOut_5_15[9] , \ScanLink11[31] , 
        \wRegInBot_4_14[14] , \ScanLink32[19] , \ScanLink47[29] , 
        \ScanLink11[28] , \ScanLink47[30] , \wRegInTop_3_4[24] , 
        \wRegEnTop_3_6[0] , \wRegOut_4_5[2] , \wRegInBot_4_9[27] , 
        \wRegOut_4_0[23] , \ScanLink19[5] , \wRegOut_4_11[28] , 
        \wRegOut_4_11[31] , \wRegInBot_4_12[9] , \wRegInBot_4_14[27] , 
        \wRegOut_0_0[5] , \wRegInBot_0_0[3] , \wRegOut_1_1[7] , 
        \ScanLink3[15] , \wRegInTop_4_14[20] , \wRegInTop_3_4[17] , 
        \wRegOut_4_0[10] , \wRegInBot_4_9[14] , \wRegInTop_2_0[18] , 
        \wRegInTop_5_27[19] , \wRegOut_2_3[8] , \ScanLink8[19] , 
        \wRegOut_5_13[7] , \wRegInTop_3_6[7] , \wRegInBot_3_7[1] , 
        \wRegInTop_5_6[3] , \wRegInTop_5_5[0] , \wRegInTop_5_8[11] , 
        \wRegOut_5_14[27] , \wRegOut_3_3[26] , \wRegOut_3_3[15] , 
        \wRegInBot_3_4[2] , \wRegOut_5_10[4] , \wRegOut_5_22[22] , 
        \wRegInTop_3_5[4] , \wRegInBot_4_2[18] , \wRegInTop_4_7[21] , 
        \wRegInTop_4_7[12] , \ScanLink59[22] , \wRegInBot_4_14[7] , 
        \ScanLink39[26] , \wRegInTop_5_8[22] , \ScanLink39[15] , 
        \ScanLink59[11] , \ScanLink0[19] , \wRegOut_1_1[19] , 
        \wRegInBot_2_0[30] , \wRegInBot_2_0[29] , \wRegInTop_2_1[21] , 
        \wRegInBot_3_0[24] , \wRegInBot_3_0[17] , \ScanLink10[11] , 
        \ScanLink26[14] , \wRegOut_5_14[14] , \wRegOut_5_22[11] , 
        \ScanLink53[24] , \wRegOut_4_10[11] , \ScanLink33[20] , 
        \ScanLink46[10] , \wRegOut_4_1[30] , \wRegInTop_5_2[17] , 
        \wRegOut_5_28[24] , \wRegOut_5_28[17] , \wRegOut_4_1[29] , 
        \wRegOut_4_8[7] , \ScanLink10[22] , \wRegOut_4_10[22] , 
        \ScanLink14[0] , \ScanLink46[23] , \ScanLink17[3] , \ScanLink26[27] , 
        \ScanLink33[13] , \ScanLink53[17] , \wRegInTop_5_14[8] , 
        \wRegInBot_4_3[21] , \wRegInTop_4_15[19] , \wRegInTop_5_2[24] , 
        \wRegInTop_2_1[12] , \ScanLink9[20] , \wRegOut_5_5[26] , 
        \wRegInTop_5_10[25] , \wRegInTop_5_9[31] , \wRegInTop_5_9[28] , 
        \wRegInTop_5_26[20] , \ScanLink9[13] , \wRegInBot_4_3[12] , 
        \wRegInTop_5_8[5] , \ScanLink58[28] , \ScanLink58[31] , 
        \wRegInTop_4_6[18] , \wRegInTop_5_12[6] , \wRegOut_5_23[31] , 
        \wRegOut_5_23[28] , \wRegOut_5_5[15] , \wRegInTop_5_11[5] , 
        \wRegInTop_5_26[13] , \wRegOut_3_0[4] , \wRegEnBot_4_2[0] , 
        \wRegInTop_4_14[5] , \wRegInTop_5_10[16] , \wRegOut_5_0[0] , 
        \wRegOut_5_1[24] , \wRegInTop_5_22[22] , \wRegOut_3_3[7] , 
        \wRegInTop_4_2[30] , \wRegInBot_4_7[23] , \ScanLink28[4] , 
        \ScanLink29[29] , \wRegInTop_5_14[27] , \ScanLink29[30] , 
        \wRegInTop_4_2[29] , \wRegOut_5_3[3] , \wRegInBot_4_4[9] , 
        \wRegOut_5_1[17] , \ScanLink36[8] , \wRegInTop_5_14[14] , 
        \wRegOut_5_24[8] , \wRegOut_5_27[19] , \wRegInTop_5_22[11] , 
        \wRegInTop_2_0[6] , \wRegInBot_4_7[10] , \wRegInTop_4_11[31] , 
        \wRegInBot_2_1[0] , \wRegOut_2_2[21] , \wRegOut_2_2[12] , 
        \wRegInTop_4_0[2] , \wRegInBot_4_1[4] , \wRegInTop_4_11[28] , 
        \ScanLink33[5] , \wRegOut_5_21[5] , \wRegInTop_5_6[15] , 
        \wRegInBot_2_2[3] , \wRegInTop_2_3[5] , \wRegInBot_3_4[15] , 
        \wRegOut_4_14[13] , \wRegOut_4_5[18] , \ScanLink14[13] , 
        \wRegInTop_4_11[8] , \ScanLink61[23] , \wRegOut_3_5[9] , 
        \wRegInBot_4_2[7] , \ScanLink22[16] , \wRegInTop_4_9[16] , 
        \ScanLink30[6] , \ScanLink37[22] , \ScanLink42[12] , \wRegOut_5_22[6] , 
        \ScanLink57[26] , \wRegInTop_4_3[1] , \ScanLink8[1] , 
        \wRegInBot_3_4[26] , \ScanLink14[20] , \ScanLink22[25] , 
        \wRegInTop_5_6[26] , \ScanLink57[15] , \ScanLink57[1] , 
        \ScanLink61[10] , \wRegInTop_4_9[25] , \ScanLink42[21] , 
        \ScanLink54[2] , \ScanLink37[11] , \wRegOut_4_14[20] , 
        \wRegOut_3_1[9] , \wRegInBot_3_2[22] , \wRegOut_4_12[24] , 
        \wRegInTop_5_29[1] , \wRegInTop_3_7[31] , \wRegInTop_3_7[28] , 
        \ScanLink29[9] , \wRegInBot_4_6[7] , \ScanLink24[21] , 
        \ScanLink51[11] , \wRegInTop_4_15[8] , \wRegInBot_3_2[11] , 
        \ScanLink12[24] , \wRegInTop_4_7[1] , \ScanLink12[17] , 
        \wRegInTop_4_4[2] , \wRegInBot_4_5[4] , \ScanLink31[15] , 
        \ScanLink34[6] , \ScanLink44[25] , \wRegOut_5_26[6] , \ScanLink37[5] , 
        \wRegOut_5_25[5] , \wRegInTop_5_0[22] , \ScanLink24[12] , 
        \ScanLink31[26] , \ScanLink44[16] , \ScanLink50[2] , \ScanLink51[22] , 
        \wRegOut_4_12[17] , \wRegInTop_5_0[11] , \wRegEnTop_1_0[0] , 
        \wRegInTop_1_0[7] , \ScanLink53[1] , \wRegInBot_1_1[1] , 
        \wRegInTop_2_2[8] , \wRegOut_3_0[19] , \wRegOut_3_7[7] , 
        \wRegInBot_4_1[14] , \wRegOut_4_8[10] , \wRegInTop_4_13[6] , 
        \ScanLink32[8] , \wRegOut_5_7[3] , \wRegOut_5_20[8] , 
        \wRegInBot_4_0[9] , \wRegInTop_4_10[5] , \wRegInTop_5_31[3] , 
        \wRegInTop_2_3[14] , \wRegOut_3_4[4] , \wRegEnBot_4_6[0] , 
        \wRegOut_5_4[0] , \wRegInTop_5_31[21] , \wRegOut_4_8[23] , 
        \wRegOut_5_7[13] , \wRegInTop_5_12[10] , \wRegOut_5_17[18] , 
        \wRegInTop_5_24[15] , \wRegInTop_2_3[27] , \wRegInBot_4_1[27] , 
        \ScanLink19[31] , \ScanLink19[28] , \wRegOut_5_7[20] , \ScanLink48[0] , 
        \wRegInTop_5_24[26] , \wRegInTop_5_12[23] , \wRegInTop_5_31[12] , 
        \wRegInBot_1_1[24] , \wRegOut_2_0[27] , \wRegOut_3_4[31] , 
        \wRegInBot_4_5[16] , \wRegOut_5_3[11] , \wRegOut_5_13[30] , 
        \wRegInTop_5_16[12] , \wRegInTop_5_20[17] , \wRegOut_5_13[29] , 
        \wRegOut_5_30[18] , \wRegOut_5_3[22] , \wRegInTop_5_15[5] , 
        \wRegInTop_5_16[21] , \wRegOut_5_19[1] , \wRegInTop_5_20[24] , 
        \wRegOut_3_4[28] , \wRegInBot_4_5[25] , \wRegInTop_5_4[20] , 
        \wRegInTop_5_16[6] , \ScanLink4[31] , \ScanLink4[28] , 
        \ScanLink16[26] , \ScanLink63[16] , \ScanLink35[17] , \ScanLink40[27] , 
        \ScanLink55[13] , \wEnable_2[0] , \ScanLink13[3] , \wRegInBot_3_6[20] , 
        \ScanLink20[23] , \wRegOut_5_18[16] , \wRegInBot_4_13[29] , 
        \wRegInBot_0_0[23] , \ScanLink1[20] , \ScanLink1[13] , \ScanLink2[7] , 
        \wRegInBot_1_1[17] , \wRegOut_2_0[14] , \wRegInBot_4_13[30] , 
        \wRegInTop_5_9[8] , \wRegInTop_3_3[19] , \wRegInBot_3_6[13] , 
        \wRegInTop_5_4[13] , \wRegOut_5_18[25] , \ScanLink20[10] , 
        \wRegOut_2_1[6] , \wRegInBot_2_3[25] , \wRegInBot_3_0[2] , 
        \ScanLink10[0] , \ScanLink16[15] , \wRegInTop_5_10[8] , 
        \ScanLink55[20] , \wRegInTop_5_1[0] , \ScanLink35[24] , 
        \ScanLink63[25] , \ScanLink40[14] , \wRegOut_5_14[4] , 
        \wRegOut_5_24[15] , \wRegInTop_3_1[4] , \wRegOut_5_12[10] , 
        \wRegOut_3_5[22] , \wRegInTop_4_1[25] , \wRegOut_5_31[21] , 
        \ScanLink18[8] , \wRegOut_5_2[31] , \wRegInTop_5_18[0] , 
        \wRegInBot_2_3[16] , \wRegInTop_3_2[7] , \wRegInBot_3_3[1] , 
        \wRegOut_5_2[28] , \wRegInTop_5_2[3] , \wRegOut_5_17[7] , 
        \wRegOut_3_5[11] , \wRegInTop_4_1[16] , \wRegInBot_4_10[7] , 
        \wRegInBot_4_13[4] , \wRegOut_5_12[23] , \ScanLink62[0] , 
        \wRegOut_5_24[26] , \wRegOut_5_31[12] , \ScanLink61[3] , 
        \wRegEnTop_4_13[0] , \wRegInTop_5_17[18] , \ScanLink5[22] , 
        \ScanLink5[11] , \wRegEnTop_3_2[0] , \wRegOut_4_1[2] , 
        \wRegInTop_3_2[13] , \wRegInBot_3_7[19] , \wRegOut_4_6[14] , 
        \wRegOut_2_2[5] , \wRegInBot_4_12[23] , \wRegInTop_5_5[19] , 
        \wRegOut_5_11[9] , \wRegOut_5_9[17] , \wRegInTop_3_2[20] , 
        \wRegInTop_3_4[9] , \wRegOut_4_2[1] , \wRegInTop_4_12[24] , 
        \ScanLink21[30] , \wRegOut_4_6[27] , \ScanLink21[29] , 
        \ScanLink54[19] , \wRegInTop_4_12[17] , \wRegInBot_4_12[10] , 
        \wRegOut_5_9[24] , \wRegInTop_5_18[16] , \ScanLink1[4] , 
        \wRegInTop_1_1[15] , \wRegInTop_3_6[11] , \wRegOut_4_2[16] , 
        \ScanLink50[31] , \ScanLink25[18] , \ScanLink40[8] , \ScanLink50[28] , 
        \wRegInTop_1_1[26] , \wRegInBot_4_8[1] , \wRegInTop_4_9[7] , 
        \wRegOut_4_14[9] , \wRegInTop_5_1[31] , \wRegInTop_5_1[28] , 
        \wRegOut_5_28[0] , \wRegInTop_5_18[25] , \wRegInTop_5_27[7] , 
        \wRegInTop_5_24[4] , \wRegInBot_3_3[31] , \wRegInBot_3_3[28] , 
        \wRegOut_4_2[25] , \wRegInTop_3_6[22] , \ScanLink39[3] , 
        \wRegInBot_0_0[19] , \wRegInBot_0_0[10] , \ScanLink4[9] , 
        \wRegOut_3_1[20] , \wRegInTop_5_13[30] , \wRegInTop_5_13[29] , 
        \ScanLink45[5] , \wRegEnTop_5_16[0] , \wRegInTop_5_30[18] , 
        \ScanLink18[22] , \wRegInTop_4_5[27] , \wRegOut_4_9[30] , 
        \wRegOut_4_9[29] , \wRegOut_5_16[12] , \wRegOut_5_6[19] , 
        \wRegOut_5_9[5] , \ScanLink46[6] , \wRegOut_5_20[17] , 
        \wRegInTop_5_21[9] , \wRegOut_1_0[3] , \wRegInBot_1_0[27] , 
        \wRegOut_3_1[13] , \ScanLink18[11] , \wRegInTop_4_5[14] , 
        \ScanLink21[1] , \wRegOut_4_12[7] , \ScanLink22[2] , 
        \wRegOut_5_16[21] , \wRegOut_5_20[24] , \wRegOut_4_11[4] , 
        \wRegOut_5_30[2] , \wRegEnTop_4_9[0] , \wRegInTop_3_2[30] , 
        \wRegInTop_3_2[29] , \wRegInBot_3_7[23] , \wRegOut_5_19[15] , 
        \ScanLink54[10] , \wRegInBot_1_0[14] , \wRegOut_2_1[24] , 
        \ScanLink17[25] , \ScanLink21[20] , \wRegInBot_4_15[3] , 
        \ScanLink41[24] , \ScanLink34[14] , \ScanLink62[15] , 
        \wRegInBot_4_12[19] , \wRegInBot_3_6[5] , \ScanLink34[27] , 
        \wRegInTop_5_5[23] , \ScanLink41[17] , \wRegInTop_3_7[3] , 
        \ScanLink17[16] , \ScanLink21[13] , \wRegInTop_5_7[7] , 
        \ScanLink62[26] , \wRegOut_5_12[3] , \wRegOut_2_1[17] , 
        \ScanLink5[18] , \wRegInBot_3_7[10] , \ScanLink54[23] , 
        \wRegInTop_5_5[10] , \wRegOut_5_19[26] , \wRegInTop_3_4[0] , 
        \wRegInBot_3_5[6] , \wRegOut_4_2[8] , \wRegOut_3_5[18] , 
        \wRegInTop_5_4[4] , \wRegOut_5_11[0] , \wRegInBot_4_4[15] , 
        \ScanLink62[9] , \wRegInTop_2_2[17] , \wRegInBot_3_3[8] , 
        \ScanLink18[1] , \wRegInBot_4_4[26] , \wRegOut_4_7[5] , 
        \wRegOut_5_2[12] , \wRegInTop_5_17[11] , \wRegInTop_5_21[14] , 
        \wRegInTop_5_1[9] , \wRegOut_5_12[19] , \wRegOut_5_31[31] , 
        \wRegOut_5_31[28] , \wRegOut_5_2[21] , \wRegInTop_5_18[9] , 
        \wRegInTop_5_21[27] , \wRegInTop_5_17[22] , \wRegOut_4_4[6] , 
        \wRegOut_5_6[10] , \wRegEnTop_5_7[0] , \wRegInTop_5_25[16] , 
        \wRegInTop_5_13[13] , \wRegInTop_5_30[22] , \ScanLink4[0] , 
        \wRegInBot_4_0[17] , \ScanLink21[8] , \wRegOut_4_9[13] , 
        \wRegInTop_5_21[0] , \wRegOut_5_16[31] , \wRegOut_5_16[28] , 
        \wRegInTop_5_22[3] , \ScanLink18[18] , \ScanLink1[30] , 
        \wRegInTop_2_2[24] , \wRegInTop_5_13[20] , \ScanLink58[3] , 
        \ScanLink7[3] , \wRegOut_3_1[30] , \wRegOut_3_1[29] , 
        \wRegInBot_4_0[24] , \wRegOut_5_6[23] , \wRegInTop_5_25[25] , 
        \wRegInTop_5_30[11] , \wRegInBot_4_8[8] , \wRegOut_4_9[20] , 
        \wRegInTop_5_1[21] , \wRegOut_5_28[9] , \ScanLink1[29] , 
        \wRegInTop_1_0[16] , \wRegInBot_2_0[4] , \wRegInTop_2_1[2] , 
        \wRegOut_3_0[23] , \wRegInBot_3_3[21] , \ScanLink13[27] , 
        \ScanLink24[5] , \ScanLink27[6] , \wRegOut_4_14[0] , \ScanLink30[16] , 
        \ScanLink45[26] , \ScanLink25[22] , \ScanLink50[12] , 
        \wRegOut_4_13[27] , \wRegInBot_3_3[12] , \wRegInTop_5_1[12] , 
        \ScanLink43[2] , \ScanLink13[14] , \wRegInTop_3_6[18] , 
        \wRegOut_4_13[14] , \ScanLink25[11] , \ScanLink30[25] , 
        \ScanLink40[1] , \ScanLink50[21] , \ScanLink45[15] , \ScanLink19[21] , 
        \wRegOut_5_17[11] , \wRegOut_5_21[14] , \ScanLink56[5] , 
        \wRegInTop_4_4[24] , \wRegOut_3_0[10] , \ScanLink9[5] , 
        \ScanLink48[9] , \wRegOut_5_7[30] , \wRegOut_5_7[29] , \ScanLink55[6] , 
        \wRegInBot_4_0[0] , \ScanLink19[12] , \wRegInTop_4_4[17] , 
        \ScanLink32[1] , \wRegOut_5_20[1] , \wRegInTop_4_1[6] , 
        \wRegOut_4_8[19] , \wRegOut_5_17[22] , \wRegInTop_2_2[1] , 
        \wRegInTop_4_2[5] , \wRegInBot_4_3[3] , \wRegOut_5_21[27] , 
        \ScanLink31[2] , \wRegOut_5_23[2] , \wRegInBot_2_3[7] , 
        \wRegOut_5_4[9] , \wRegInTop_5_12[19] , \wRegInTop_5_31[28] , 
        \wRegInTop_5_31[31] , \wRegInBot_3_2[18] , \wRegOut_4_3[15] , 
        \ScanLink0[10] , \wRegInTop_3_7[12] , \wRegInBot_1_1[8] , 
        \wRegInTop_5_0[18] , \ScanLink53[8] , \wRegInTop_5_19[15] , 
        \wRegInBot_0_0[27] , \ScanLink0[23] , \wRegInTop_1_0[25] , 
        \wRegOut_3_1[0] , \wRegInTop_3_7[21] , \ScanLink29[0] , 
        \wRegOut_4_3[26] , \wRegInTop_5_29[8] , \wRegEnBot_2_3[0] , 
        \wRegInTop_4_7[8] , \ScanLink24[28] , \ScanLink51[18] , 
        \wRegInTop_4_15[1] , \wRegOut_3_2[3] , \ScanLink24[31] , 
        \wRegOut_5_1[4] , \wRegOut_5_2[7] , \wRegInTop_5_19[26] , 
        \ScanLink4[21] , \ScanLink4[12] , \wRegInTop_4_13[27] , 
        \wRegInTop_5_13[2] , \wRegInBot_4_13[20] , \wRegOut_5_8[14] , 
        \ScanLink10[9] , \wRegInTop_3_3[10] , \wRegInTop_5_9[1] , 
        \ScanLink20[19] , \wRegOut_4_7[17] , \wRegInTop_5_10[1] , 
        \ScanLink55[30] , \ScanLink55[29] , \wRegInTop_2_2[30] , 
        \wRegInTop_2_2[29] , \wRegInBot_2_2[26] , \wRegInTop_3_3[23] , 
        \wRegInBot_3_6[30] , \wRegInTop_4_13[14] , \wRegInBot_4_13[13] , 
        \wRegInTop_5_4[30] , \wRegInTop_5_4[29] , \wRegOut_5_8[27] , 
        \wRegInBot_3_6[29] , \wRegOut_4_7[24] , \ScanLink15[4] , 
        \wRegOut_4_9[3] , \wRegInBot_2_2[15] , \wRegOut_3_4[21] , 
        \wRegInTop_5_16[31] , \wRegInTop_5_16[28] , \wRegInTop_4_0[26] , 
        \wRegOut_5_19[8] , \ScanLink16[7] , \wRegOut_5_13[13] , 
        \wRegOut_5_30[22] , \wRegOut_5_25[16] , \wRegOut_5_3[18] , 
        \wRegOut_3_1[24] , \wRegOut_3_4[12] , \wRegInTop_4_0[15] , 
        \wRegOut_5_13[20] , \wRegOut_5_25[25] , \wRegOut_5_30[11] , 
        \wRegInBot_4_0[30] , \ScanLink18[26] , \ScanLink46[2] , 
        \wRegOut_5_20[13] , \wRegOut_5_16[16] , \wRegInTop_4_5[23] , 
        \wRegInBot_4_0[29] , \ScanLink45[1] , \wRegInTop_5_25[31] , 
        \wRegInTop_5_25[28] , \wRegInBot_0_0[14] , \wRegOut_3_1[17] , 
        \ScanLink18[15] , \wRegInTop_4_5[10] , \ScanLink22[6] , 
        \wRegOut_4_11[0] , \wRegOut_5_30[6] , \wRegOut_4_12[3] , 
        \wRegOut_5_16[25] , \wRegOut_5_20[20] , \ScanLink1[24] , 
        \ScanLink1[17] , \ScanLink1[0] , \ScanLink21[5] , \wRegOut_5_9[1] , 
        \wRegInTop_1_1[11] , \ScanLink13[19] , \ScanLink30[31] , 
        \wRegInTop_3_6[15] , \wRegOut_4_2[12] , \wRegOut_4_13[19] , 
        \ScanLink30[28] , \ScanLink45[18] , \ScanLink2[3] , 
        \wRegInTop_1_1[22] , \wRegInTop_3_6[26] , \ScanLink39[7] , 
        \wRegInTop_5_18[12] , \wRegOut_4_2[21] , \wRegInBot_4_8[5] , 
        \ScanLink24[8] , \wRegInTop_5_18[21] , \wRegInTop_5_24[0] , 
        \wRegInTop_5_27[3] , \wRegOut_5_28[4] , \wRegInTop_4_9[3] , 
        \wRegInBot_1_0[19] , \ScanLink5[15] , \wRegOut_2_2[1] , 
        \wRegOut_4_2[5] , \wRegInTop_4_12[20] , \wRegInBot_4_12[27] , 
        \wRegOut_5_9[13] , \wRegInTop_5_4[9] , \wRegInTop_3_2[17] , 
        \wRegInBot_3_6[8] , \wRegOut_4_6[10] , \wRegOut_4_1[6] , 
        \wRegInBot_1_1[20] , \wRegOut_2_1[30] , \wRegOut_2_1[29] , 
        \wRegOut_2_1[2] , \wRegEnTop_5_2[0] , \ScanLink5[26] , 
        \wRegInBot_2_3[21] , \wRegInTop_3_2[24] , \ScanLink17[31] , 
        \ScanLink17[28] , \wRegInTop_4_12[13] , \wRegInBot_4_12[14] , 
        \wRegOut_5_9[20] , \ScanLink41[30] , \ScanLink62[18] , 
        \ScanLink41[29] , \wRegOut_4_6[23] , \ScanLink34[19] , 
        \wRegOut_5_19[18] , \wRegInTop_3_2[3] , \wRegInBot_3_3[5] , 
        \wRegInTop_5_2[7] , \wRegOut_5_17[3] , \wRegInTop_5_18[4] , 
        \wRegInBot_2_3[12] , \wRegInBot_3_0[6] , \wRegOut_3_5[26] , 
        \wRegInTop_4_1[21] , \wRegOut_4_7[8] , \wRegOut_5_31[25] , 
        \wRegInTop_3_1[0] , \wRegOut_5_12[14] , \wRegInTop_5_1[4] , 
        \wRegOut_5_14[0] , \wRegOut_5_24[11] , \wRegOut_3_5[15] , 
        \wRegInTop_4_1[12] , \wRegInBot_4_10[3] , \wRegInTop_5_21[19] , 
        \ScanLink61[7] , \wRegInBot_4_13[0] , \wRegOut_5_24[22] , 
        \ScanLink62[4] , \wRegOut_5_12[27] , \wRegOut_5_31[16] , 
        \wRegInBot_3_6[24] , \wRegInBot_4_4[18] , \wRegOut_5_18[12] , 
        \wRegOut_4_7[30] , \wRegOut_4_7[29] , \ScanLink55[17] , 
        \wRegInBot_1_1[13] , \wRegOut_2_0[23] , \ScanLink16[22] , 
        \ScanLink20[27] , \ScanLink35[13] , \ScanLink40[23] , \ScanLink63[12] , 
        \wRegInTop_4_13[19] , \ScanLink16[11] , \ScanLink35[20] , 
        \wRegInTop_5_4[24] , \ScanLink40[10] , \ScanLink20[14] , 
        \ScanLink63[21] , \wRegOut_2_0[10] , \ScanLink10[4] , 
        \wRegInBot_3_6[17] , \ScanLink55[24] , \wRegInTop_5_4[17] , 
        \wRegOut_5_18[21] , \ScanLink13[7] , \wRegOut_0_0[1] , 
        \wRegInBot_2_0[9] , \wRegInBot_2_2[18] , \wRegInTop_4_0[18] , 
        \wRegOut_5_8[19] , \wRegInBot_4_5[12] , \wRegOut_5_3[15] , 
        \wRegInTop_5_16[16] , \wRegOut_5_25[31] , \wRegOut_5_25[28] , 
        \wRegInTop_5_20[13] , \wRegInTop_2_3[10] , \ScanLink15[9] , 
        \wRegInBot_4_5[21] , \wRegInTop_5_16[2] , \wRegOut_5_3[26] , 
        \wRegOut_5_19[5] , \wRegInTop_5_20[20] , \wRegInTop_5_15[1] , 
        \wRegInTop_5_16[25] , \wRegOut_5_7[17] , \wRegInTop_5_24[11] , 
        \wRegInTop_5_12[14] , \wRegInTop_5_31[25] , \wRegOut_3_4[0] , 
        \wRegOut_3_7[3] , \wRegInTop_4_2[8] , \wRegOut_4_8[14] , 
        \wRegInTop_4_10[1] , \wRegInTop_5_31[7] , \wRegOut_5_4[4] , 
        \wRegInTop_4_13[2] , \wRegOut_5_7[7] , \wRegInBot_4_1[10] , 
        \wRegInTop_1_0[31] , \wRegInTop_2_3[23] , \ScanLink9[8] , 
        \wRegInTop_5_12[27] , \ScanLink48[4] , \wRegInBot_4_1[23] , 
        \wRegInTop_4_4[30] , \wRegInTop_4_4[29] , \wRegOut_5_7[24] , 
        \wRegInTop_5_24[22] , \wRegInTop_5_31[16] , \wRegInTop_4_4[6] , 
        \wRegInBot_4_5[0] , \wRegOut_4_8[27] , \wRegOut_5_21[19] , 
        \ScanLink56[8] , \wRegInTop_5_0[26] , \ScanLink34[2] , \ScanLink37[1] , 
        \wRegOut_5_25[1] , \wRegOut_5_26[2] , \wRegInTop_1_0[28] , 
        \wRegInBot_4_6[3] , \ScanLink31[11] , \ScanLink44[21] , 
        \wRegInTop_1_0[3] , \wRegInBot_3_2[26] , \ScanLink12[20] , 
        \wRegInTop_4_7[5] , \ScanLink24[25] , \wRegOut_5_1[9] , 
        \ScanLink51[15] , \wRegOut_4_12[20] , \wRegInTop_5_29[5] , 
        \ScanLink53[5] , \wRegInBot_1_1[5] , \wRegInBot_3_2[15] , 
        \wRegOut_4_3[18] , \wRegInTop_5_0[15] , \wRegInTop_5_19[18] , 
        \wRegOut_4_12[13] , \ScanLink0[14] , \wRegInBot_1_1[30] , 
        \wRegOut_2_0[19] , \ScanLink4[16] , \wRegInBot_2_2[22] , 
        \wRegOut_3_4[25] , \ScanLink12[13] , \ScanLink24[16] , 
        \ScanLink31[22] , \ScanLink50[6] , \ScanLink51[26] , \ScanLink44[12] , 
        \wRegInTop_4_0[22] , \ScanLink16[3] , \wRegOut_5_25[12] , 
        \wRegOut_5_13[17] , \wRegOut_5_30[26] , \wRegInBot_4_5[28] , 
        \wRegInBot_4_5[31] , \wRegOut_4_9[7] , \wRegInTop_5_20[29] , 
        \wRegInTop_5_20[30] , \wRegInBot_2_2[11] , \wRegOut_3_4[16] , 
        \ScanLink15[0] , \wRegInTop_5_15[8] , \wRegInTop_4_0[11] , 
        \wRegOut_5_13[24] , \wRegOut_5_25[21] , \wRegOut_5_30[15] , 
        \wRegInTop_3_3[14] , \ScanLink16[18] , \ScanLink35[30] , 
        \ScanLink35[29] , \ScanLink40[19] , \ScanLink63[31] , 
        \wRegInTop_5_10[5] , \wRegOut_4_7[13] , \ScanLink63[28] , 
        \wRegOut_5_18[31] , \wRegOut_5_18[28] , \wRegInTop_5_9[5] , 
        \wRegInTop_3_3[27] , \wRegInTop_4_13[23] , \wRegInBot_4_13[24] , 
        \wRegOut_5_8[10] , \wRegInTop_5_13[6] , \wRegOut_4_7[20] , 
        \wRegInBot_1_1[29] , \ScanLink4[25] , \wRegInTop_4_13[10] , 
        \wRegInBot_4_13[17] , \wRegOut_5_8[23] , \wRegInTop_5_19[11] , 
        \wRegInTop_3_7[16] , \ScanLink0[27] , \wRegInTop_1_0[12] , 
        \wRegOut_4_3[11] , \wRegInTop_1_0[21] , \wRegOut_3_1[4] , 
        \wRegOut_3_2[7] , \wRegOut_5_2[3] , \ScanLink12[30] , 
        \wRegInBot_4_5[9] , \wRegInTop_4_15[5] , \ScanLink37[8] , 
        \wRegInTop_5_19[22] , \wRegOut_5_25[8] , \wRegOut_5_1[0] , 
        \ScanLink44[28] , \ScanLink31[18] , \wRegEnBot_4_3[0] , 
        \ScanLink44[31] , \ScanLink12[29] , \wRegInTop_3_7[25] , 
        \wRegOut_4_3[22] , \wRegOut_4_12[30] , \wRegOut_4_12[29] , 
        \ScanLink29[4] , \wRegOut_0_0[8] , \ScanLink1[9] , \wRegInTop_1_1[18] , 
        \wRegInBot_2_0[0] , \wRegInTop_2_1[6] , \wRegInTop_2_2[5] , 
        \wRegInTop_2_3[19] , \wRegOut_3_0[27] , \ScanLink9[1] , 
        \ScanLink55[2] , \ScanLink19[25] , \wRegInTop_4_4[20] , 
        \wRegOut_5_17[15] , \wRegOut_5_21[10] , \ScanLink56[1] , 
        \wRegInTop_4_10[8] , \wRegInTop_5_24[18] , \wRegInBot_2_3[3] , 
        \wRegOut_3_4[9] , \wRegInBot_4_3[7] , \ScanLink31[6] , 
        \wRegOut_5_23[6] , \wRegInTop_4_2[1] , \wRegOut_5_21[23] , 
        \wRegOut_3_0[14] , \wRegInBot_4_0[4] , \wRegInTop_4_1[2] , 
        \ScanLink19[16] , \wRegInTop_4_4[13] , \ScanLink32[5] , 
        \wRegOut_5_17[26] , \wRegOut_5_20[5] , \wRegInBot_3_3[25] , 
        \wRegInBot_4_1[19] , \wRegOut_4_2[31] , \wRegOut_4_13[23] , 
        \ScanLink13[23] , \wRegOut_4_2[28] , \ScanLink25[26] , 
        \ScanLink50[16] , \wRegInTop_5_24[9] , \ScanLink13[10] , 
        \ScanLink24[1] , \ScanLink27[2] , \wRegOut_4_14[4] , \ScanLink30[12] , 
        \ScanLink45[22] , \wRegInTop_5_1[25] , \wRegInTop_5_18[31] , 
        \wRegInTop_5_18[28] , \ScanLink25[15] , \ScanLink30[21] , 
        \ScanLink45[11] , \ScanLink40[5] , \ScanLink50[25] , \ScanLink4[4] , 
        \wRegInTop_2_2[20] , \wRegInTop_2_2[13] , \wRegInBot_3_3[16] , 
        \wRegInBot_4_0[13] , \wRegInTop_4_5[19] , \wRegOut_4_13[10] , 
        \wRegInTop_5_1[16] , \wRegEnTop_5_13[0] , \ScanLink43[6] , 
        \wRegOut_4_9[17] , \wRegOut_4_11[9] , \wRegOut_5_20[30] , 
        \wRegInTop_5_22[7] , \wRegOut_5_20[29] , \wRegInTop_5_21[4] , 
        \wRegInTop_5_30[26] , \ScanLink7[7] , \wRegOut_4_9[24] , 
        \wRegOut_5_6[14] , \wRegOut_5_9[8] , \wRegInTop_5_13[17] , 
        \wRegInTop_5_25[12] , \wRegInBot_4_0[20] , \wRegOut_5_6[27] , 
        \wRegInTop_5_25[21] , \ScanLink58[7] , \wRegInTop_5_13[24] , 
        \wRegInTop_5_30[15] , \ScanLink45[8] , \wRegOut_1_0[7] , 
        \wRegOut_5_2[16] , \wRegInTop_5_17[15] , \wRegInTop_5_21[10] , 
        \wRegInBot_1_0[23] , \wRegOut_2_1[20] , \wRegInBot_2_3[31] , 
        \wRegInBot_2_3[28] , \wRegEnTop_3_7[0] , \wRegOut_4_4[2] , 
        \wRegInBot_4_4[11] , \wRegInBot_4_13[9] , \ScanLink18[5] , 
        \wRegInTop_5_17[26] , \wRegOut_5_2[25] , \wRegInTop_3_1[9] , 
        \wRegInTop_4_1[31] , \wRegInTop_5_21[23] , \wRegInTop_4_1[28] , 
        \wRegInBot_4_4[22] , \wRegOut_4_7[1] , \wRegOut_5_14[9] , 
        \wRegOut_5_24[18] , \wRegInTop_5_5[27] , \ScanLink17[21] , 
        \wRegOut_5_9[30] , \wRegOut_5_9[29] , \ScanLink62[11] , 
        \wRegInBot_4_15[7] , \ScanLink41[20] , \ScanLink34[10] , 
        \ScanLink54[14] , \wRegInBot_1_0[10] , \wRegOut_2_1[13] , 
        \wRegOut_2_2[8] , \wRegInBot_3_7[27] , \ScanLink21[24] , 
        \wRegOut_5_19[11] , \wRegInTop_5_4[0] , \wRegInTop_3_4[4] , 
        \wRegInBot_3_5[2] , \wRegInTop_4_12[30] , \wRegOut_5_11[4] , 
        \wRegInTop_4_12[29] , \wRegInBot_3_7[14] , \wRegOut_4_6[19] , 
        \wRegInTop_5_5[14] , \ScanLink21[17] , \wRegOut_5_19[22] , 
        \ScanLink2[8] , \wRegInTop_1_1[30] , \wRegInTop_1_1[29] , 
        \ScanLink13[21] , \wRegInBot_3_6[1] , \wRegInTop_5_7[3] , 
        \wRegOut_5_12[7] , \ScanLink54[27] , \wRegInTop_3_7[7] , 
        \ScanLink17[12] , \wRegInTop_4_9[8] , \wRegInTop_5_1[27] , 
        \ScanLink34[23] , \ScanLink62[22] , \ScanLink41[13] , \ScanLink27[0] , 
        \wRegOut_4_14[6] , \wRegInTop_5_27[8] , \ScanLink24[3] , 
        \ScanLink30[10] , \ScanLink45[20] , \wRegInBot_3_3[27] , 
        \ScanLink25[24] , \ScanLink50[14] , \wRegOut_4_13[21] , \ScanLink4[6] , 
        \wRegInTop_2_2[11] , \wRegInBot_3_3[14] , \wRegOut_4_2[19] , 
        \wRegOut_4_13[12] , \wRegInTop_5_1[14] , \ScanLink43[4] , 
        \wRegInTop_5_18[19] , \ScanLink13[12] , \ScanLink25[17] , 
        \ScanLink50[27] , \ScanLink40[7] , \ScanLink30[23] , \ScanLink45[13] , 
        \wRegOut_5_6[16] , \wRegInTop_5_25[10] , \wRegInBot_4_0[11] , 
        \wRegOut_4_9[15] , \wRegOut_4_12[8] , \wRegInTop_5_13[15] , 
        \wRegInTop_5_30[24] , \wRegInTop_5_21[6] , \wRegInTop_5_22[5] , 
        \wRegOut_1_0[5] , \wRegInTop_2_2[22] , \ScanLink58[5] , 
        \wRegInTop_5_30[17] , \ScanLink7[5] , \wRegInBot_4_0[22] , 
        \wRegInTop_4_5[31] , \wRegOut_5_6[25] , \wRegInTop_5_13[26] , 
        \wRegInTop_5_25[23] , \wRegInTop_4_5[28] , \wRegInTop_4_1[19] , 
        \wRegOut_4_9[26] , \ScanLink46[9] , \wRegOut_5_20[18] , 
        \wRegInBot_4_4[13] , \wRegOut_5_24[30] , \wRegOut_5_24[29] , 
        \wRegInTop_1_0[10] , \wRegInBot_1_0[21] , \wRegInBot_2_3[19] , 
        \wRegInBot_4_10[8] , \wRegOut_5_2[14] , \wRegInTop_5_17[17] , 
        \wRegInTop_3_2[8] , \ScanLink18[7] , \wRegInBot_4_4[20] , 
        \wRegOut_4_7[3] , \wRegInTop_5_21[12] , \wRegOut_5_2[27] , 
        \wRegInTop_5_21[21] , \wRegInTop_5_17[24] , \wRegInBot_3_7[25] , 
        \wRegOut_4_4[0] , \wRegOut_4_6[31] , \wRegOut_5_17[8] , 
        \ScanLink21[26] , \wRegOut_4_6[28] , \wRegOut_5_19[13] , 
        \wRegInBot_1_0[12] , \wRegOut_2_1[22] , \ScanLink17[23] , 
        \ScanLink54[16] , \wRegInTop_4_12[18] , \wRegInBot_4_15[5] , 
        \ScanLink62[13] , \ScanLink34[12] , \ScanLink41[22] , 
        \wRegInBot_3_6[3] , \wRegInTop_3_7[5] , \wRegInTop_5_5[25] , 
        \ScanLink62[20] , \ScanLink17[10] , \ScanLink34[21] , \ScanLink41[11] , 
        \wRegOut_5_12[5] , \ScanLink54[25] , \wRegInBot_1_1[18] , 
        \ScanLink4[14] , \wRegOut_2_1[11] , \wRegOut_2_1[9] , \ScanLink21[15] , 
        \wRegInBot_3_7[16] , \wRegInTop_5_7[1] , \wRegOut_5_19[20] , 
        \wRegInTop_5_5[16] , \wRegInBot_2_2[20] , \wRegInTop_3_4[6] , 
        \wRegInBot_3_5[0] , \ScanLink15[2] , \wRegInTop_5_4[2] , 
        \wRegOut_5_9[18] , \wRegOut_5_11[6] , \wCtrlOut_2[0] , 
        \wRegInBot_2_2[13] , \wRegOut_3_4[27] , \wRegOut_4_9[5] , 
        \wRegInTop_4_0[20] , \ScanLink16[1] , \wRegEnTop_5_9[0] , 
        \wRegOut_5_13[15] , \wRegInTop_5_16[9] , \wRegOut_5_25[10] , 
        \wRegOut_5_30[24] , \wRegInTop_5_20[18] , \wRegOut_3_4[14] , 
        \wRegInTop_4_0[13] , \wRegOut_5_13[26] , \wRegOut_5_25[23] , 
        \wRegOut_5_30[17] , \wRegInBot_4_5[19] , \wRegInTop_4_13[21] , 
        \wRegEnTop_5_21[0] , \wRegInBot_4_13[26] , \wRegInTop_5_13[4] , 
        \wRegOut_5_8[12] , \wRegInTop_3_3[16] , \wRegInTop_5_9[7] , 
        \wRegOut_4_7[11] , \wRegInTop_5_10[7] , \wRegOut_2_0[31] , 
        \wRegOut_2_0[28] , \ScanLink4[27] , \wRegInTop_3_3[25] , 
        \ScanLink16[30] , \wRegInTop_4_13[12] , \wRegInBot_4_13[15] , 
        \wRegOut_5_8[21] , \ScanLink35[18] , \ScanLink16[29] , 
        \ScanLink40[28] , \wRegOut_4_7[22] , \ScanLink40[31] , 
        \ScanLink63[19] , \wRegOut_5_18[19] , \ScanLink31[29] , 
        \ScanLink44[19] , \ScanLink12[18] , \wRegInTop_3_7[14] , 
        \wRegOut_4_3[13] , \ScanLink31[30] , \wRegOut_4_12[18] , 
        \ScanLink0[16] , \wRegInTop_1_0[8] , \wRegInTop_3_7[27] , 
        \ScanLink29[6] , \wRegInTop_5_19[13] , \wRegOut_0_0[3] , 
        \ScanLink0[25] , \wRegInTop_1_0[23] , \wRegOut_3_1[6] , 
        \wRegOut_4_3[20] , \ScanLink34[9] , \wRegOut_5_26[9] , 
        \wRegInBot_4_6[8] , \wRegEnTop_2_2[0] , \wRegInTop_4_15[7] , 
        \wRegOut_5_1[2] , \wRegOut_3_2[5] , \wRegInTop_5_19[20] , 
        \wRegOut_5_2[1] , \wRegEnBot_1_1[0] , \wRegInBot_1_1[22] , 
        \wRegOut_2_0[21] , \wRegInBot_2_0[2] , \wRegInTop_2_3[31] , 
        \wRegOut_3_0[25] , \wRegInBot_4_1[28] , \ScanLink19[27] , 
        \wRegInTop_4_4[22] , \wRegOut_5_17[17] , \wRegOut_5_21[12] , 
        \ScanLink56[3] , \ScanLink9[3] , \wRegInBot_4_1[31] , 
        \wRegInTop_2_3[28] , \wRegOut_3_0[16] , \ScanLink55[0] , 
        \wRegInTop_5_24[30] , \wRegInTop_5_24[29] , \wRegOut_3_7[8] , 
        \wRegInBot_4_0[6] , \wRegInTop_4_1[0] , \ScanLink19[14] , 
        \wRegInTop_4_4[11] , \wRegOut_5_17[24] , \ScanLink32[7] , 
        \wRegOut_5_20[7] , \wRegOut_5_21[21] , \wRegInTop_2_1[4] , 
        \wRegInTop_2_2[7] , \wRegInBot_2_3[1] , \wRegInTop_4_2[3] , 
        \wRegInTop_4_13[9] , \ScanLink31[4] , \wRegOut_5_23[4] , 
        \wRegInBot_4_3[5] , \wRegInTop_5_4[26] , \ScanLink16[20] , 
        \ScanLink35[11] , \wRegOut_5_8[31] , \wRegOut_5_8[28] , 
        \ScanLink40[21] , \ScanLink20[25] , \ScanLink63[10] , 
        \wRegInBot_1_1[11] , \wRegOut_2_0[12] , \ScanLink13[5] , 
        \wRegInBot_3_6[26] , \ScanLink55[15] , \wRegOut_5_18[10] , 
        \wRegInTop_4_13[31] , \wRegInTop_4_13[28] , \wRegInBot_3_6[15] , 
        \wRegOut_4_7[18] , \wRegInTop_5_4[15] , \wRegOut_5_18[23] , 
        \ScanLink55[26] , \wRegInBot_2_2[30] , \ScanLink10[6] , 
        \ScanLink20[16] , \ScanLink16[13] , \ScanLink35[22] , \ScanLink40[12] , 
        \ScanLink63[23] , \wRegInBot_4_5[10] , \wRegOut_5_3[17] , 
        \wRegInTop_5_20[11] , \wRegInTop_5_16[14] , \wRegInTop_5_15[3] , 
        \wRegInTop_5_16[27] , \wRegInTop_5_20[22] , \wRegInBot_2_2[29] , 
        \wRegInTop_2_3[12] , \wRegInBot_2_3[8] , \wRegOut_3_7[1] , 
        \wRegInTop_4_0[30] , \wRegInTop_4_0[29] , \wRegOut_5_3[24] , 
        \wRegOut_5_19[7] , \ScanLink16[8] , \wRegInBot_4_5[23] , 
        \wRegOut_5_25[19] , \wRegInTop_4_1[9] , \wRegInBot_4_1[12] , 
        \wRegInTop_4_4[18] , \wRegInTop_5_16[0] , \wRegInTop_4_13[0] , 
        \wRegOut_5_7[5] , \wRegOut_5_21[31] , \wRegOut_5_21[28] , 
        \wRegOut_4_8[16] , \wRegOut_5_4[6] , \wRegOut_3_4[2] , 
        \wRegEnTop_4_7[0] , \wRegInTop_4_10[3] , \wRegInTop_5_31[5] , 
        \wRegInTop_5_12[16] , \wRegOut_4_8[25] , \wRegOut_5_7[15] , 
        \wRegInTop_5_24[13] , \wRegInTop_5_31[27] , \wRegInTop_2_3[21] , 
        \wRegInBot_4_1[21] , \wRegEnTop_5_18[0] , \wRegOut_5_7[26] , 
        \wRegInTop_5_24[20] , \wRegInTop_5_12[25] , \ScanLink48[6] , 
        \wRegInTop_5_31[14] , \wRegInBot_3_2[24] , \ScanLink55[9] , 
        \wRegOut_4_3[30] , \wRegOut_4_3[29] , \wRegOut_4_12[22] , 
        \wRegInTop_5_29[7] , \wRegInBot_0_0[25] , \wRegInTop_1_0[19] , 
        \ScanLink12[22] , \ScanLink24[27] , \ScanLink31[13] , \ScanLink51[17] , 
        \ScanLink34[0] , \ScanLink44[23] , \wRegOut_5_26[0] , 
        \wRegInTop_4_4[4] , \wRegInBot_4_6[1] , \wRegInTop_4_7[7] , 
        \wRegOut_5_2[8] , \wRegInBot_4_5[2] , \wRegInTop_5_19[29] , 
        \ScanLink31[20] , \wRegInTop_5_0[24] , \ScanLink37[3] , 
        \wRegInTop_5_19[30] , \wRegOut_5_25[3] , \ScanLink44[10] , 
        \wRegInTop_1_0[1] , \wRegInBot_1_1[7] , \wRegInBot_3_2[17] , 
        \ScanLink12[11] , \ScanLink24[14] , \ScanLink51[24] , 
        \wRegOut_4_12[11] , \ScanLink50[4] , \wRegInTop_5_0[17] , 
        \ScanLink53[7] , \ScanLink45[3] , \wRegInBot_0_0[16] , 
        \wRegInTop_2_2[18] , \wRegOut_3_1[26] , \ScanLink18[24] , 
        \wRegInTop_4_5[21] , \ScanLink46[0] , \wRegOut_5_16[14] , 
        \wRegOut_5_20[11] , \wRegOut_5_9[3] , \wRegInTop_5_25[19] , 
        \ScanLink1[26] , \ScanLink1[15] , \ScanLink2[1] , \wRegOut_3_1[15] , 
        \ScanLink18[17] , \ScanLink21[7] , \wRegOut_4_12[1] , \ScanLink22[4] , 
        \wRegOut_5_20[22] , \wRegOut_4_11[2] , \wRegOut_5_16[27] , 
        \wRegOut_5_30[4] , \wRegInTop_4_5[12] , \wRegInBot_4_0[18] , 
        \wRegEnBot_4_8[0] , \wRegInTop_5_18[10] , \ScanLink1[2] , 
        \wRegInTop_1_1[13] , \wRegInTop_3_6[17] , \wRegOut_4_2[10] , 
        \ScanLink0[12] , \wRegInBot_1_0[31] , \wRegInBot_1_0[28] , 
        \wRegInTop_1_1[20] , \ScanLink13[28] , \wRegInBot_4_8[7] , 
        \wRegInTop_4_9[1] , \wRegOut_5_28[6] , \ScanLink27[9] , 
        \wRegInTop_5_27[1] , \wRegInTop_5_18[23] , \wRegInTop_5_24[2] , 
        \wRegOut_2_1[18] , \wRegOut_2_1[0] , \ScanLink13[31] , 
        \ScanLink30[19] , \ScanLink45[30] , \wRegInTop_3_6[24] , 
        \wRegOut_4_2[23] , \wRegOut_4_13[31] , \ScanLink45[29] , 
        \wRegOut_4_13[28] , \ScanLink39[5] , \wRegInTop_3_2[15] , 
        \wRegEnBot_3_3[0] , \wRegOut_4_1[4] , \wRegInTop_5_7[8] , 
        \ScanLink62[29] , \ScanLink17[19] , \ScanLink34[31] , 
        \wRegOut_4_6[12] , \ScanLink34[28] , \ScanLink41[18] , 
        \ScanLink62[30] , \wRegOut_5_19[30] , \wRegOut_5_19[29] , 
        \ScanLink5[17] , \wRegOut_2_2[3] , \wRegInTop_3_2[26] , 
        \wRegInBot_3_5[9] , \wRegInTop_4_12[22] , \wRegInBot_4_12[25] , 
        \wRegOut_5_9[11] , \wRegOut_4_2[7] , \wRegOut_4_6[21] , 
        \wRegInBot_2_0[6] , \ScanLink5[24] , \wRegInTop_4_12[11] , 
        \wRegInBot_4_12[16] , \wRegOut_5_9[22] , \wRegInTop_2_2[3] , 
        \wRegInBot_2_3[23] , \wRegInBot_3_0[4] , \wRegInTop_3_1[2] , 
        \wRegInTop_5_1[6] , \wRegOut_5_14[2] , \wRegOut_5_24[13] , 
        \wRegOut_5_31[27] , \wRegOut_3_5[24] , \wRegInTop_4_1[23] , 
        \wRegOut_5_12[16] , \wRegInBot_4_4[30] , \wRegInBot_4_4[29] , 
        \wRegInBot_2_3[10] , \wRegInTop_3_2[1] , \wRegInTop_5_2[5] , 
        \wRegOut_5_17[1] , \wRegInTop_5_18[6] , \wRegInTop_5_21[31] , 
        \wRegInTop_5_21[28] , \wRegInBot_3_3[7] , \wRegOut_4_4[9] , 
        \wRegOut_3_5[17] , \wRegInTop_4_1[10] , \wRegInBot_4_10[1] , 
        \wRegInBot_4_13[2] , \wRegOut_5_12[25] , \ScanLink62[6] , 
        \wRegOut_5_31[14] , \wRegOut_5_24[20] , \ScanLink61[5] , 
        \wRegInBot_2_3[5] , \wRegOut_3_0[21] , \ScanLink9[7] , 
        \wRegInTop_5_12[31] , \ScanLink55[4] , \wRegInTop_5_31[19] , 
        \wRegInTop_5_12[28] , \ScanLink19[23] , \wRegInTop_4_4[26] , 
        \wRegOut_4_8[31] , \wRegOut_4_8[28] , \wRegOut_5_7[18] , 
        \wRegOut_5_17[13] , \wRegOut_5_21[16] , \ScanLink56[7] , 
        \wRegInTop_5_31[8] , \wRegInTop_4_2[7] , \wRegInBot_4_3[1] , 
        \ScanLink31[0] , \wRegOut_5_23[0] , \wRegInTop_2_1[0] , 
        \wRegOut_5_7[8] , \wRegOut_3_0[12] , \wRegInBot_4_0[2] , 
        \wRegInTop_4_1[4] , \ScanLink32[3] , \wRegOut_5_21[25] , 
        \wRegOut_5_17[20] , \wRegOut_5_20[3] , \ScanLink19[10] , 
        \wRegInTop_4_4[15] , \wRegInTop_5_19[17] , \ScanLink0[21] , 
        \wRegInTop_1_0[14] , \wRegInTop_3_7[10] , \wRegOut_4_3[17] , 
        \ScanLink24[19] , \ScanLink51[29] , \ScanLink50[9] , \ScanLink51[30] , 
        \wRegInTop_1_0[27] , \wRegOut_3_1[2] , \wRegOut_3_2[1] , 
        \wRegInTop_4_4[9] , \wRegInTop_5_0[30] , \wRegInTop_5_0[29] , 
        \wRegOut_5_2[5] , \wRegInTop_5_19[24] , \wRegEnTop_4_2[0] , 
        \wRegInTop_4_15[3] , \wRegOut_5_1[6] , \wRegInBot_3_2[30] , 
        \wRegInBot_3_2[29] , \wRegOut_4_3[24] , \wRegInBot_0_0[31] , 
        \wRegInBot_0_0[28] , \wRegOut_1_0[1] , \wRegInBot_1_0[25] , 
        \ScanLink4[23] , \ScanLink4[10] , \wRegInTop_3_3[12] , 
        \wRegInBot_3_6[18] , \wRegInTop_3_7[23] , \ScanLink29[2] , 
        \wRegOut_4_7[15] , \wRegInTop_5_10[3] , \wRegInTop_3_3[21] , 
        \ScanLink13[8] , \wRegInBot_4_13[22] , \wRegInTop_5_4[18] , 
        \wRegInTop_5_9[3] , \wRegOut_5_8[16] , \wRegInTop_4_13[25] , 
        \wRegInTop_5_13[0] , \ScanLink20[31] , \ScanLink20[28] , 
        \wRegOut_4_7[26] , \ScanLink55[18] , \wRegInTop_4_13[16] , 
        \wRegInBot_4_13[11] , \wRegOut_5_8[25] , \wRegOut_2_1[26] , 
        \ScanLink5[30] , \wRegInBot_2_2[24] , \wRegOut_3_4[23] , 
        \wRegInTop_4_0[24] , \ScanLink16[5] , \wRegOut_5_25[14] , 
        \wRegOut_5_13[11] , \wRegOut_5_30[20] , \wRegInBot_2_2[17] , 
        \wRegOut_3_4[10] , \ScanLink15[6] , \wRegOut_4_9[1] , 
        \wRegOut_5_3[29] , \wRegOut_5_3[30] , \wRegInTop_4_0[17] , 
        \wRegOut_5_13[22] , \wRegOut_5_30[13] , \wRegOut_5_25[27] , 
        \wRegInTop_5_5[21] , \wRegInTop_5_16[19] , \ScanLink5[29] , 
        \ScanLink17[27] , \wRegInBot_4_15[1] , \ScanLink34[16] , 
        \ScanLink41[26] , \ScanLink21[22] , \ScanLink62[17] , 
        \wRegInBot_1_0[16] , \wRegOut_2_1[15] , \wRegInTop_3_4[2] , 
        \wRegInBot_3_7[21] , \ScanLink54[12] , \wRegInBot_4_12[31] , 
        \wRegOut_5_19[17] , \wRegInBot_4_12[28] , \wRegOut_5_11[2] , 
        \wRegInTop_5_4[6] , \wRegInBot_3_5[4] , \wRegInTop_3_2[18] , 
        \wRegInBot_3_7[12] , \wRegInTop_5_5[12] , \wRegOut_5_19[24] , 
        \wRegInTop_5_7[5] , \ScanLink54[21] , \wRegInBot_3_6[7] , 
        \wRegInTop_3_7[1] , \ScanLink21[11] , \wRegOut_5_12[1] , 
        \ScanLink34[25] , \ScanLink41[15] , \ScanLink62[24] , \wRegOut_4_1[9] , 
        \ScanLink17[14] , \wRegOut_5_2[10] , \wRegInTop_5_21[16] , 
        \wRegInTop_5_17[13] , \ScanLink61[8] , \wRegInTop_2_2[26] , 
        \wRegInTop_2_2[15] , \wRegInBot_3_0[9] , \wRegOut_3_5[30] , 
        \wRegOut_3_5[29] , \wRegEnBot_3_6[0] , \wRegInBot_4_4[17] , 
        \wRegOut_5_12[31] , \wRegOut_5_12[28] , \wRegOut_5_31[19] , 
        \wRegInTop_5_2[8] , \ScanLink18[3] , \wRegOut_4_4[4] , 
        \wRegInTop_5_17[20] , \wRegInBot_4_4[24] , \wRegOut_5_2[23] , 
        \wRegInTop_5_21[25] , \wRegOut_3_1[18] , \wRegOut_4_7[7] , 
        \wRegInBot_4_0[15] , \ScanLink22[9] , \wRegOut_4_9[11] , 
        \wRegInTop_5_22[1] , \wRegInTop_5_13[11] , \wRegInTop_5_21[2] , 
        \wRegOut_5_30[9] , \ScanLink7[1] , \wRegOut_4_9[22] , 
        \wRegOut_5_6[12] , \wRegInTop_5_25[14] , \wRegInTop_5_30[20] , 
        \wRegOut_5_16[19] , \wRegInBot_4_0[26] , \ScanLink18[30] , 
        \ScanLink18[29] , \wRegOut_5_6[21] , \wRegInTop_5_25[27] , 
        \wRegInTop_5_13[22] , \ScanLink58[1] , \wRegInTop_5_30[13] , 
        \ScanLink4[2] , \wRegOut_0_0[7] , \wRegInBot_0_0[21] , \ScanLink1[22] , 
        \ScanLink1[18] , \wRegInBot_3_3[23] , \wRegInBot_3_3[10] , 
        \ScanLink13[25] , \wRegInTop_3_6[30] , \wRegInTop_3_6[29] , 
        \wRegOut_4_13[25] , \ScanLink39[8] , \ScanLink24[7] , \ScanLink25[20] , 
        \ScanLink30[14] , \ScanLink50[10] , \ScanLink45[24] , \ScanLink13[16] , 
        \ScanLink27[4] , \wRegOut_4_14[2] , \ScanLink30[27] , 
        \wRegInTop_5_1[23] , \ScanLink45[17] , \ScanLink25[13] , 
        \ScanLink50[23] , \wRegOut_4_13[16] , \ScanLink40[3] , 
        \wRegInTop_5_1[10] , \ScanLink1[11] , \ScanLink1[6] , \wRegOut_1_0[8] , 
        \wRegInBot_2_3[27] , \wRegInTop_3_2[5] , \ScanLink43[0] , 
        \wRegInBot_3_3[3] , \wRegInTop_5_2[1] , \wRegOut_5_17[5] , 
        \wRegInBot_2_3[14] , \wRegInBot_3_0[0] , \wRegInTop_3_1[6] , 
        \wRegOut_3_5[20] , \wRegInTop_5_17[30] , \wRegInTop_5_17[29] , 
        \wRegInTop_5_18[2] , \wRegInTop_4_1[27] , \wRegInTop_5_1[2] , 
        \wRegOut_5_12[12] , \wRegOut_5_14[6] , \wRegOut_5_31[23] , 
        \wRegOut_5_24[17] , \wRegOut_5_2[19] , \wRegOut_2_1[4] , 
        \ScanLink5[13] , \wRegOut_2_2[7] , \wRegOut_3_5[13] , 
        \wRegInTop_4_1[14] , \wRegInBot_4_10[5] , \wRegInBot_4_13[6] , 
        \wRegOut_5_12[21] , \wRegOut_5_24[24] , \ScanLink61[1] , 
        \ScanLink62[2] , \wRegOut_5_31[10] , \wRegOut_4_2[3] , 
        \wRegInTop_4_12[26] , \wRegInBot_4_12[21] , \wRegOut_5_9[15] , 
        \wRegInTop_3_2[11] , \wRegInTop_3_7[8] , \wRegOut_4_6[16] , 
        \wRegOut_4_1[0] , \ScanLink54[31] , \ScanLink5[20] , \ScanLink21[18] , 
        \ScanLink54[28] , \wRegOut_5_12[8] , \wRegInTop_3_2[22] , 
        \wRegInBot_3_7[31] , \wRegInBot_3_7[28] , \wRegInTop_4_12[15] , 
        \wRegInBot_4_12[12] , \wRegInTop_5_5[31] , \wRegInTop_5_5[28] , 
        \wRegOut_5_9[26] , \wRegInBot_4_15[8] , \wRegOut_4_6[25] , 
        \wRegInTop_1_1[17] , \wRegInBot_3_3[19] , \wRegOut_4_2[14] , 
        \wRegInTop_3_6[13] , \ScanLink2[5] , \wRegInTop_5_1[19] , 
        \ScanLink43[9] , \wRegInTop_1_1[24] , \wRegInTop_3_6[20] , 
        \ScanLink39[1] , \wRegInTop_5_18[14] , \wRegOut_4_2[27] , 
        \wRegInBot_4_8[3] , \wRegInTop_4_9[5] , \ScanLink25[30] , 
        \ScanLink25[29] , \wRegInTop_5_24[6] , \wRegInTop_5_18[27] , 
        \ScanLink50[19] , \wRegInTop_5_27[5] , \wRegOut_5_28[2] , 
        \ScanLink7[8] , \ScanLink46[4] , \wRegOut_5_20[15] , \wRegOut_3_1[22] , 
        \ScanLink18[20] , \wRegInTop_4_5[25] , \wRegOut_5_16[10] , 
        \wRegOut_5_6[31] , \ScanLink58[8] , \wRegOut_5_6[28] , \ScanLink45[7] , 
        \wRegInBot_0_0[12] , \wRegOut_3_1[11] , \ScanLink18[13] , 
        \wRegInTop_4_5[16] , \ScanLink22[0] , \wRegOut_4_9[18] , 
        \wRegOut_5_16[23] , \wRegOut_4_11[6] , \wRegOut_4_12[5] , 
        \wRegOut_5_20[26] , \wRegOut_5_30[0] , \wRegInTop_5_22[8] , 
        \ScanLink0[31] , \ScanLink0[28] , \ScanLink21[3] , \wRegInTop_5_0[20] , 
        \wRegOut_5_9[7] , \wRegInTop_5_13[18] , \wRegInTop_5_30[30] , 
        \wRegInTop_5_30[29] , \wRegInTop_1_0[5] , \wRegInBot_1_1[3] , 
        \wRegOut_3_2[8] , \wRegInTop_4_4[0] , \ScanLink37[7] , 
        \wRegOut_5_25[7] , \wRegInBot_4_5[6] , \wRegInBot_3_2[20] , 
        \ScanLink12[26] , \wRegInBot_4_6[5] , \wRegInTop_4_7[3] , 
        \ScanLink24[23] , \ScanLink31[17] , \ScanLink34[4] , \ScanLink44[27] , 
        \wRegOut_5_26[4] , \ScanLink51[13] , \wRegOut_4_12[26] , 
        \wRegInTop_5_29[3] , \ScanLink53[3] , \wRegInTop_2_1[9] , 
        \wRegInTop_2_3[16] , \wRegInBot_3_2[13] , \wRegOut_4_12[15] , 
        \wRegInTop_5_0[13] , \ScanLink12[15] , \wRegInTop_3_7[19] , 
        \ScanLink24[10] , \ScanLink51[20] , \ScanLink50[0] , 
        \wRegEnBot_4_13[0] , \ScanLink31[24] , \ScanLink44[14] , 
        \wRegOut_5_7[11] , \wRegInTop_5_24[17] , \wRegOut_3_4[6] , 
        \wRegInTop_5_12[12] , \wRegInTop_5_31[23] , \wRegOut_3_7[5] , 
        \wRegInBot_4_3[8] , \wRegInTop_4_10[7] , \ScanLink31[9] , 
        \wRegOut_5_23[9] , \wRegOut_5_4[2] , \wRegOut_5_17[30] , 
        \wRegInTop_5_31[1] , \wRegOut_5_17[29] , \wRegOut_4_8[12] , 
        \wRegOut_5_7[1] , \wRegInBot_4_1[16] , \wRegInTop_4_13[4] , 
        \ScanLink19[19] , \wRegInBot_1_1[26] , \wRegInTop_2_3[25] , 
        \ScanLink48[2] , \wRegInTop_5_31[10] , \wRegOut_3_0[31] , 
        \wRegOut_5_7[22] , \wRegInTop_5_12[21] , \wRegInTop_5_24[24] , 
        \wRegOut_3_0[28] , \wRegInBot_4_1[25] , \wRegInTop_3_3[31] , 
        \wRegOut_3_4[19] , \wRegOut_4_8[21] , \wRegInBot_3_6[22] , 
        \wRegInBot_4_5[27] , \wRegInBot_4_5[14] , \wRegOut_5_3[13] , 
        \wRegInTop_5_16[10] , \wRegOut_5_13[18] , \wRegInTop_5_16[4] , 
        \wRegInTop_5_20[15] , \wRegOut_5_30[29] , \wRegOut_5_30[30] , 
        \wRegOut_4_9[8] , \wRegOut_5_3[20] , \wRegOut_5_19[3] , 
        \wRegInTop_5_15[7] , \wRegInTop_5_16[23] , \wRegInTop_5_20[26] , 
        \wRegOut_5_18[14] , \wRegInTop_3_3[28] , \ScanLink20[21] , 
        \wRegInBot_1_1[15] , \wRegOut_2_0[25] , \ScanLink16[24] , 
        \ScanLink55[11] , \wRegInBot_4_13[18] , \ScanLink35[15] , 
        \ScanLink63[14] , \ScanLink40[25] , \ScanLink16[17] , 
        \wRegInTop_5_4[22] , \wRegEnTop_5_24[0] , \ScanLink63[27] , 
        \ScanLink35[26] , \ScanLink40[16] , \ScanLink55[22] , 
        \wRegOut_2_0[16] , \ScanLink10[2] , \ScanLink20[12] , 
        \wRegInBot_3_6[11] , \wRegOut_5_18[27] , \wRegInTop_5_4[11] , 
        \ScanLink4[19] , \wRegInTop_5_13[9] , \ScanLink13[1] ;
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink13[31] , \ScanLink13[30] , \ScanLink13[29] , 
        \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , \ScanLink13[25] , 
        \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , \ScanLink13[21] , 
        \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , \ScanLink13[17] , 
        \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , \ScanLink13[13] , 
        \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , \ScanLink13[9] , 
        \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , \ScanLink13[5] , 
        \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , \ScanLink13[1] , 
        \ScanLink13[0] }), .ScanOut({\ScanLink12[31] , \ScanLink12[30] , 
        \ScanLink12[29] , \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , 
        \ScanLink12[25] , \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , 
        \ScanLink12[21] , \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , 
        \ScanLink12[17] , \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , 
        \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , 
        \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , 
        \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , 
        \ScanLink12[1] , \ScanLink12[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_5[31] , \wRegOut_3_5[30] , \wRegOut_3_5[29] , 
        \wRegOut_3_5[28] , \wRegOut_3_5[27] , \wRegOut_3_5[26] , 
        \wRegOut_3_5[25] , \wRegOut_3_5[24] , \wRegOut_3_5[23] , 
        \wRegOut_3_5[22] , \wRegOut_3_5[21] , \wRegOut_3_5[20] , 
        \wRegOut_3_5[19] , \wRegOut_3_5[18] , \wRegOut_3_5[17] , 
        \wRegOut_3_5[16] , \wRegOut_3_5[15] , \wRegOut_3_5[14] , 
        \wRegOut_3_5[13] , \wRegOut_3_5[12] , \wRegOut_3_5[11] , 
        \wRegOut_3_5[10] , \wRegOut_3_5[9] , \wRegOut_3_5[8] , 
        \wRegOut_3_5[7] , \wRegOut_3_5[6] , \wRegOut_3_5[5] , \wRegOut_3_5[4] , 
        \wRegOut_3_5[3] , \wRegOut_3_5[2] , \wRegOut_3_5[1] , \wRegOut_3_5[0] 
        }), .Enable1(\wRegEnTop_3_5[0] ), .Enable2(\wRegEnBot_3_5[0] ), .In1({
        \wRegInTop_3_5[31] , \wRegInTop_3_5[30] , \wRegInTop_3_5[29] , 
        \wRegInTop_3_5[28] , \wRegInTop_3_5[27] , \wRegInTop_3_5[26] , 
        \wRegInTop_3_5[25] , \wRegInTop_3_5[24] , \wRegInTop_3_5[23] , 
        \wRegInTop_3_5[22] , \wRegInTop_3_5[21] , \wRegInTop_3_5[20] , 
        \wRegInTop_3_5[19] , \wRegInTop_3_5[18] , \wRegInTop_3_5[17] , 
        \wRegInTop_3_5[16] , \wRegInTop_3_5[15] , \wRegInTop_3_5[14] , 
        \wRegInTop_3_5[13] , \wRegInTop_3_5[12] , \wRegInTop_3_5[11] , 
        \wRegInTop_3_5[10] , \wRegInTop_3_5[9] , \wRegInTop_3_5[8] , 
        \wRegInTop_3_5[7] , \wRegInTop_3_5[6] , \wRegInTop_3_5[5] , 
        \wRegInTop_3_5[4] , \wRegInTop_3_5[3] , \wRegInTop_3_5[2] , 
        \wRegInTop_3_5[1] , \wRegInTop_3_5[0] }), .In2({\wRegInBot_3_5[31] , 
        \wRegInBot_3_5[30] , \wRegInBot_3_5[29] , \wRegInBot_3_5[28] , 
        \wRegInBot_3_5[27] , \wRegInBot_3_5[26] , \wRegInBot_3_5[25] , 
        \wRegInBot_3_5[24] , \wRegInBot_3_5[23] , \wRegInBot_3_5[22] , 
        \wRegInBot_3_5[21] , \wRegInBot_3_5[20] , \wRegInBot_3_5[19] , 
        \wRegInBot_3_5[18] , \wRegInBot_3_5[17] , \wRegInBot_3_5[16] , 
        \wRegInBot_3_5[15] , \wRegInBot_3_5[14] , \wRegInBot_3_5[13] , 
        \wRegInBot_3_5[12] , \wRegInBot_3_5[11] , \wRegInBot_3_5[10] , 
        \wRegInBot_3_5[9] , \wRegInBot_3_5[8] , \wRegInBot_3_5[7] , 
        \wRegInBot_3_5[6] , \wRegInBot_3_5[5] , \wRegInBot_3_5[4] , 
        \wRegInBot_3_5[3] , \wRegInBot_3_5[2] , \wRegInBot_3_5[1] , 
        \wRegInBot_3_5[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_26 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink58[31] , \ScanLink58[30] , \ScanLink58[29] , 
        \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , \ScanLink58[25] , 
        \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , \ScanLink58[21] , 
        \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , \ScanLink58[17] , 
        \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , \ScanLink58[13] , 
        \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , \ScanLink58[9] , 
        \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , \ScanLink58[5] , 
        \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , \ScanLink58[1] , 
        \ScanLink58[0] }), .ScanOut({\ScanLink57[31] , \ScanLink57[30] , 
        \ScanLink57[29] , \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , 
        \ScanLink57[25] , \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , 
        \ScanLink57[21] , \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , 
        \ScanLink57[17] , \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , 
        \ScanLink57[13] , \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , 
        \ScanLink57[9] , \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , 
        \ScanLink57[5] , \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , 
        \ScanLink57[1] , \ScanLink57[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_26[31] , \wRegOut_5_26[30] , 
        \wRegOut_5_26[29] , \wRegOut_5_26[28] , \wRegOut_5_26[27] , 
        \wRegOut_5_26[26] , \wRegOut_5_26[25] , \wRegOut_5_26[24] , 
        \wRegOut_5_26[23] , \wRegOut_5_26[22] , \wRegOut_5_26[21] , 
        \wRegOut_5_26[20] , \wRegOut_5_26[19] , \wRegOut_5_26[18] , 
        \wRegOut_5_26[17] , \wRegOut_5_26[16] , \wRegOut_5_26[15] , 
        \wRegOut_5_26[14] , \wRegOut_5_26[13] , \wRegOut_5_26[12] , 
        \wRegOut_5_26[11] , \wRegOut_5_26[10] , \wRegOut_5_26[9] , 
        \wRegOut_5_26[8] , \wRegOut_5_26[7] , \wRegOut_5_26[6] , 
        \wRegOut_5_26[5] , \wRegOut_5_26[4] , \wRegOut_5_26[3] , 
        \wRegOut_5_26[2] , \wRegOut_5_26[1] , \wRegOut_5_26[0] }), .Enable1(
        \wRegEnTop_5_26[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_26[31] , 
        \wRegInTop_5_26[30] , \wRegInTop_5_26[29] , \wRegInTop_5_26[28] , 
        \wRegInTop_5_26[27] , \wRegInTop_5_26[26] , \wRegInTop_5_26[25] , 
        \wRegInTop_5_26[24] , \wRegInTop_5_26[23] , \wRegInTop_5_26[22] , 
        \wRegInTop_5_26[21] , \wRegInTop_5_26[20] , \wRegInTop_5_26[19] , 
        \wRegInTop_5_26[18] , \wRegInTop_5_26[17] , \wRegInTop_5_26[16] , 
        \wRegInTop_5_26[15] , \wRegInTop_5_26[14] , \wRegInTop_5_26[13] , 
        \wRegInTop_5_26[12] , \wRegInTop_5_26[11] , \wRegInTop_5_26[10] , 
        \wRegInTop_5_26[9] , \wRegInTop_5_26[8] , \wRegInTop_5_26[7] , 
        \wRegInTop_5_26[6] , \wRegInTop_5_26[5] , \wRegInTop_5_26[4] , 
        \wRegInTop_5_26[3] , \wRegInTop_5_26[2] , \wRegInTop_5_26[1] , 
        \wRegInTop_5_26[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_7[0] ), .P_In({\wRegOut_3_7[31] , 
        \wRegOut_3_7[30] , \wRegOut_3_7[29] , \wRegOut_3_7[28] , 
        \wRegOut_3_7[27] , \wRegOut_3_7[26] , \wRegOut_3_7[25] , 
        \wRegOut_3_7[24] , \wRegOut_3_7[23] , \wRegOut_3_7[22] , 
        \wRegOut_3_7[21] , \wRegOut_3_7[20] , \wRegOut_3_7[19] , 
        \wRegOut_3_7[18] , \wRegOut_3_7[17] , \wRegOut_3_7[16] , 
        \wRegOut_3_7[15] , \wRegOut_3_7[14] , \wRegOut_3_7[13] , 
        \wRegOut_3_7[12] , \wRegOut_3_7[11] , \wRegOut_3_7[10] , 
        \wRegOut_3_7[9] , \wRegOut_3_7[8] , \wRegOut_3_7[7] , \wRegOut_3_7[6] , 
        \wRegOut_3_7[5] , \wRegOut_3_7[4] , \wRegOut_3_7[3] , \wRegOut_3_7[2] , 
        \wRegOut_3_7[1] , \wRegOut_3_7[0] }), .P_Out({\wRegInBot_3_7[31] , 
        \wRegInBot_3_7[30] , \wRegInBot_3_7[29] , \wRegInBot_3_7[28] , 
        \wRegInBot_3_7[27] , \wRegInBot_3_7[26] , \wRegInBot_3_7[25] , 
        \wRegInBot_3_7[24] , \wRegInBot_3_7[23] , \wRegInBot_3_7[22] , 
        \wRegInBot_3_7[21] , \wRegInBot_3_7[20] , \wRegInBot_3_7[19] , 
        \wRegInBot_3_7[18] , \wRegInBot_3_7[17] , \wRegInBot_3_7[16] , 
        \wRegInBot_3_7[15] , \wRegInBot_3_7[14] , \wRegInBot_3_7[13] , 
        \wRegInBot_3_7[12] , \wRegInBot_3_7[11] , \wRegInBot_3_7[10] , 
        \wRegInBot_3_7[9] , \wRegInBot_3_7[8] , \wRegInBot_3_7[7] , 
        \wRegInBot_3_7[6] , \wRegInBot_3_7[5] , \wRegInBot_3_7[4] , 
        \wRegInBot_3_7[3] , \wRegInBot_3_7[2] , \wRegInBot_3_7[1] , 
        \wRegInBot_3_7[0] }), .L_WR(\wRegEnTop_4_14[0] ), .L_In({
        \wRegOut_4_14[31] , \wRegOut_4_14[30] , \wRegOut_4_14[29] , 
        \wRegOut_4_14[28] , \wRegOut_4_14[27] , \wRegOut_4_14[26] , 
        \wRegOut_4_14[25] , \wRegOut_4_14[24] , \wRegOut_4_14[23] , 
        \wRegOut_4_14[22] , \wRegOut_4_14[21] , \wRegOut_4_14[20] , 
        \wRegOut_4_14[19] , \wRegOut_4_14[18] , \wRegOut_4_14[17] , 
        \wRegOut_4_14[16] , \wRegOut_4_14[15] , \wRegOut_4_14[14] , 
        \wRegOut_4_14[13] , \wRegOut_4_14[12] , \wRegOut_4_14[11] , 
        \wRegOut_4_14[10] , \wRegOut_4_14[9] , \wRegOut_4_14[8] , 
        \wRegOut_4_14[7] , \wRegOut_4_14[6] , \wRegOut_4_14[5] , 
        \wRegOut_4_14[4] , \wRegOut_4_14[3] , \wRegOut_4_14[2] , 
        \wRegOut_4_14[1] , \wRegOut_4_14[0] }), .L_Out({\wRegInTop_4_14[31] , 
        \wRegInTop_4_14[30] , \wRegInTop_4_14[29] , \wRegInTop_4_14[28] , 
        \wRegInTop_4_14[27] , \wRegInTop_4_14[26] , \wRegInTop_4_14[25] , 
        \wRegInTop_4_14[24] , \wRegInTop_4_14[23] , \wRegInTop_4_14[22] , 
        \wRegInTop_4_14[21] , \wRegInTop_4_14[20] , \wRegInTop_4_14[19] , 
        \wRegInTop_4_14[18] , \wRegInTop_4_14[17] , \wRegInTop_4_14[16] , 
        \wRegInTop_4_14[15] , \wRegInTop_4_14[14] , \wRegInTop_4_14[13] , 
        \wRegInTop_4_14[12] , \wRegInTop_4_14[11] , \wRegInTop_4_14[10] , 
        \wRegInTop_4_14[9] , \wRegInTop_4_14[8] , \wRegInTop_4_14[7] , 
        \wRegInTop_4_14[6] , \wRegInTop_4_14[5] , \wRegInTop_4_14[4] , 
        \wRegInTop_4_14[3] , \wRegInTop_4_14[2] , \wRegInTop_4_14[1] , 
        \wRegInTop_4_14[0] }), .R_WR(\wRegEnTop_4_15[0] ), .R_In({
        \wRegOut_4_15[31] , \wRegOut_4_15[30] , \wRegOut_4_15[29] , 
        \wRegOut_4_15[28] , \wRegOut_4_15[27] , \wRegOut_4_15[26] , 
        \wRegOut_4_15[25] , \wRegOut_4_15[24] , \wRegOut_4_15[23] , 
        \wRegOut_4_15[22] , \wRegOut_4_15[21] , \wRegOut_4_15[20] , 
        \wRegOut_4_15[19] , \wRegOut_4_15[18] , \wRegOut_4_15[17] , 
        \wRegOut_4_15[16] , \wRegOut_4_15[15] , \wRegOut_4_15[14] , 
        \wRegOut_4_15[13] , \wRegOut_4_15[12] , \wRegOut_4_15[11] , 
        \wRegOut_4_15[10] , \wRegOut_4_15[9] , \wRegOut_4_15[8] , 
        \wRegOut_4_15[7] , \wRegOut_4_15[6] , \wRegOut_4_15[5] , 
        \wRegOut_4_15[4] , \wRegOut_4_15[3] , \wRegOut_4_15[2] , 
        \wRegOut_4_15[1] , \wRegOut_4_15[0] }), .R_Out({\wRegInTop_4_15[31] , 
        \wRegInTop_4_15[30] , \wRegInTop_4_15[29] , \wRegInTop_4_15[28] , 
        \wRegInTop_4_15[27] , \wRegInTop_4_15[26] , \wRegInTop_4_15[25] , 
        \wRegInTop_4_15[24] , \wRegInTop_4_15[23] , \wRegInTop_4_15[22] , 
        \wRegInTop_4_15[21] , \wRegInTop_4_15[20] , \wRegInTop_4_15[19] , 
        \wRegInTop_4_15[18] , \wRegInTop_4_15[17] , \wRegInTop_4_15[16] , 
        \wRegInTop_4_15[15] , \wRegInTop_4_15[14] , \wRegInTop_4_15[13] , 
        \wRegInTop_4_15[12] , \wRegInTop_4_15[11] , \wRegInTop_4_15[10] , 
        \wRegInTop_4_15[9] , \wRegInTop_4_15[8] , \wRegInTop_4_15[7] , 
        \wRegInTop_4_15[6] , \wRegInTop_4_15[5] , \wRegInTop_4_15[4] , 
        \wRegInTop_4_15[3] , \wRegInTop_4_15[2] , \wRegInTop_4_15[1] , 
        \wRegInTop_4_15[0] }) );
    BHeap_Node_WIDTH32 BHN_4_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_14[0] ), .P_In({\wRegOut_4_14[31] , 
        \wRegOut_4_14[30] , \wRegOut_4_14[29] , \wRegOut_4_14[28] , 
        \wRegOut_4_14[27] , \wRegOut_4_14[26] , \wRegOut_4_14[25] , 
        \wRegOut_4_14[24] , \wRegOut_4_14[23] , \wRegOut_4_14[22] , 
        \wRegOut_4_14[21] , \wRegOut_4_14[20] , \wRegOut_4_14[19] , 
        \wRegOut_4_14[18] , \wRegOut_4_14[17] , \wRegOut_4_14[16] , 
        \wRegOut_4_14[15] , \wRegOut_4_14[14] , \wRegOut_4_14[13] , 
        \wRegOut_4_14[12] , \wRegOut_4_14[11] , \wRegOut_4_14[10] , 
        \wRegOut_4_14[9] , \wRegOut_4_14[8] , \wRegOut_4_14[7] , 
        \wRegOut_4_14[6] , \wRegOut_4_14[5] , \wRegOut_4_14[4] , 
        \wRegOut_4_14[3] , \wRegOut_4_14[2] , \wRegOut_4_14[1] , 
        \wRegOut_4_14[0] }), .P_Out({\wRegInBot_4_14[31] , 
        \wRegInBot_4_14[30] , \wRegInBot_4_14[29] , \wRegInBot_4_14[28] , 
        \wRegInBot_4_14[27] , \wRegInBot_4_14[26] , \wRegInBot_4_14[25] , 
        \wRegInBot_4_14[24] , \wRegInBot_4_14[23] , \wRegInBot_4_14[22] , 
        \wRegInBot_4_14[21] , \wRegInBot_4_14[20] , \wRegInBot_4_14[19] , 
        \wRegInBot_4_14[18] , \wRegInBot_4_14[17] , \wRegInBot_4_14[16] , 
        \wRegInBot_4_14[15] , \wRegInBot_4_14[14] , \wRegInBot_4_14[13] , 
        \wRegInBot_4_14[12] , \wRegInBot_4_14[11] , \wRegInBot_4_14[10] , 
        \wRegInBot_4_14[9] , \wRegInBot_4_14[8] , \wRegInBot_4_14[7] , 
        \wRegInBot_4_14[6] , \wRegInBot_4_14[5] , \wRegInBot_4_14[4] , 
        \wRegInBot_4_14[3] , \wRegInBot_4_14[2] , \wRegInBot_4_14[1] , 
        \wRegInBot_4_14[0] }), .L_WR(\wRegEnTop_5_28[0] ), .L_In({
        \wRegOut_5_28[31] , \wRegOut_5_28[30] , \wRegOut_5_28[29] , 
        \wRegOut_5_28[28] , \wRegOut_5_28[27] , \wRegOut_5_28[26] , 
        \wRegOut_5_28[25] , \wRegOut_5_28[24] , \wRegOut_5_28[23] , 
        \wRegOut_5_28[22] , \wRegOut_5_28[21] , \wRegOut_5_28[20] , 
        \wRegOut_5_28[19] , \wRegOut_5_28[18] , \wRegOut_5_28[17] , 
        \wRegOut_5_28[16] , \wRegOut_5_28[15] , \wRegOut_5_28[14] , 
        \wRegOut_5_28[13] , \wRegOut_5_28[12] , \wRegOut_5_28[11] , 
        \wRegOut_5_28[10] , \wRegOut_5_28[9] , \wRegOut_5_28[8] , 
        \wRegOut_5_28[7] , \wRegOut_5_28[6] , \wRegOut_5_28[5] , 
        \wRegOut_5_28[4] , \wRegOut_5_28[3] , \wRegOut_5_28[2] , 
        \wRegOut_5_28[1] , \wRegOut_5_28[0] }), .L_Out({\wRegInTop_5_28[31] , 
        \wRegInTop_5_28[30] , \wRegInTop_5_28[29] , \wRegInTop_5_28[28] , 
        \wRegInTop_5_28[27] , \wRegInTop_5_28[26] , \wRegInTop_5_28[25] , 
        \wRegInTop_5_28[24] , \wRegInTop_5_28[23] , \wRegInTop_5_28[22] , 
        \wRegInTop_5_28[21] , \wRegInTop_5_28[20] , \wRegInTop_5_28[19] , 
        \wRegInTop_5_28[18] , \wRegInTop_5_28[17] , \wRegInTop_5_28[16] , 
        \wRegInTop_5_28[15] , \wRegInTop_5_28[14] , \wRegInTop_5_28[13] , 
        \wRegInTop_5_28[12] , \wRegInTop_5_28[11] , \wRegInTop_5_28[10] , 
        \wRegInTop_5_28[9] , \wRegInTop_5_28[8] , \wRegInTop_5_28[7] , 
        \wRegInTop_5_28[6] , \wRegInTop_5_28[5] , \wRegInTop_5_28[4] , 
        \wRegInTop_5_28[3] , \wRegInTop_5_28[2] , \wRegInTop_5_28[1] , 
        \wRegInTop_5_28[0] }), .R_WR(\wRegEnTop_5_29[0] ), .R_In({
        \wRegOut_5_29[31] , \wRegOut_5_29[30] , \wRegOut_5_29[29] , 
        \wRegOut_5_29[28] , \wRegOut_5_29[27] , \wRegOut_5_29[26] , 
        \wRegOut_5_29[25] , \wRegOut_5_29[24] , \wRegOut_5_29[23] , 
        \wRegOut_5_29[22] , \wRegOut_5_29[21] , \wRegOut_5_29[20] , 
        \wRegOut_5_29[19] , \wRegOut_5_29[18] , \wRegOut_5_29[17] , 
        \wRegOut_5_29[16] , \wRegOut_5_29[15] , \wRegOut_5_29[14] , 
        \wRegOut_5_29[13] , \wRegOut_5_29[12] , \wRegOut_5_29[11] , 
        \wRegOut_5_29[10] , \wRegOut_5_29[9] , \wRegOut_5_29[8] , 
        \wRegOut_5_29[7] , \wRegOut_5_29[6] , \wRegOut_5_29[5] , 
        \wRegOut_5_29[4] , \wRegOut_5_29[3] , \wRegOut_5_29[2] , 
        \wRegOut_5_29[1] , \wRegOut_5_29[0] }), .R_Out({\wRegInTop_5_29[31] , 
        \wRegInTop_5_29[30] , \wRegInTop_5_29[29] , \wRegInTop_5_29[28] , 
        \wRegInTop_5_29[27] , \wRegInTop_5_29[26] , \wRegInTop_5_29[25] , 
        \wRegInTop_5_29[24] , \wRegInTop_5_29[23] , \wRegInTop_5_29[22] , 
        \wRegInTop_5_29[21] , \wRegInTop_5_29[20] , \wRegInTop_5_29[19] , 
        \wRegInTop_5_29[18] , \wRegInTop_5_29[17] , \wRegInTop_5_29[16] , 
        \wRegInTop_5_29[15] , \wRegInTop_5_29[14] , \wRegInTop_5_29[13] , 
        \wRegInTop_5_29[12] , \wRegInTop_5_29[11] , \wRegInTop_5_29[10] , 
        \wRegInTop_5_29[9] , \wRegInTop_5_29[8] , \wRegInTop_5_29[7] , 
        \wRegInTop_5_29[6] , \wRegInTop_5_29[5] , \wRegInTop_5_29[4] , 
        \wRegInTop_5_29[3] , \wRegInTop_5_29[2] , \wRegInTop_5_29[1] , 
        \wRegInTop_5_29[0] }) );
    BHeap_CtrlReg_WIDTH32 BHCR_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_4[0] ), 
        .Out(\wCtrlOut_3[0] ), .Enable(\wEnable_3[0] ) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_0_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink1[31] , \ScanLink1[30] , \ScanLink1[29] , 
        \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , \ScanLink1[25] , 
        \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , \ScanLink1[21] , 
        \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , \ScanLink1[17] , 
        \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , \ScanLink1[13] , 
        \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , \ScanLink1[9] , 
        \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , \ScanLink1[5] , 
        \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , \ScanLink1[1] , 
        \ScanLink1[0] }), .ScanOut({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_0_0[31] , \wRegOut_0_0[30] , \wRegOut_0_0[29] , 
        \wRegOut_0_0[28] , \wRegOut_0_0[27] , \wRegOut_0_0[26] , 
        \wRegOut_0_0[25] , \wRegOut_0_0[24] , \wRegOut_0_0[23] , 
        \wRegOut_0_0[22] , \wRegOut_0_0[21] , \wRegOut_0_0[20] , 
        \wRegOut_0_0[19] , \wRegOut_0_0[18] , \wRegOut_0_0[17] , 
        \wRegOut_0_0[16] , \wRegOut_0_0[15] , \wRegOut_0_0[14] , 
        \wRegOut_0_0[13] , \wRegOut_0_0[12] , \wRegOut_0_0[11] , 
        \wRegOut_0_0[10] , \wRegOut_0_0[9] , \wRegOut_0_0[8] , 
        \wRegOut_0_0[7] , \wRegOut_0_0[6] , \wRegOut_0_0[5] , \wRegOut_0_0[4] , 
        \wRegOut_0_0[3] , \wRegOut_0_0[2] , \wRegOut_0_0[1] , \wRegOut_0_0[0] 
        }), .Enable1(1'b0), .Enable2(\wRegEnBot_0_0[0] ), .In1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .In2({\wRegInBot_0_0[31] , 
        \wRegInBot_0_0[30] , \wRegInBot_0_0[29] , \wRegInBot_0_0[28] , 
        \wRegInBot_0_0[27] , \wRegInBot_0_0[26] , \wRegInBot_0_0[25] , 
        \wRegInBot_0_0[24] , \wRegInBot_0_0[23] , \wRegInBot_0_0[22] , 
        \wRegInBot_0_0[21] , \wRegInBot_0_0[20] , \wRegInBot_0_0[19] , 
        \wRegInBot_0_0[18] , \wRegInBot_0_0[17] , \wRegInBot_0_0[16] , 
        \wRegInBot_0_0[15] , \wRegInBot_0_0[14] , \wRegInBot_0_0[13] , 
        \wRegInBot_0_0[12] , \wRegInBot_0_0[11] , \wRegInBot_0_0[10] , 
        \wRegInBot_0_0[9] , \wRegInBot_0_0[8] , \wRegInBot_0_0[7] , 
        \wRegInBot_0_0[6] , \wRegInBot_0_0[5] , \wRegInBot_0_0[4] , 
        \wRegInBot_0_0[3] , \wRegInBot_0_0[2] , \wRegInBot_0_0[1] , 
        \wRegInBot_0_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_1_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink2[31] , \ScanLink2[30] , \ScanLink2[29] , 
        \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , \ScanLink2[25] , 
        \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , \ScanLink2[21] , 
        \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , \ScanLink2[17] , 
        \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , \ScanLink2[13] , 
        \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , \ScanLink2[9] , 
        \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , \ScanLink2[5] , 
        \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , \ScanLink2[1] , 
        \ScanLink2[0] }), .ScanOut({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_1_0[31] , \wRegOut_1_0[30] , \wRegOut_1_0[29] , 
        \wRegOut_1_0[28] , \wRegOut_1_0[27] , \wRegOut_1_0[26] , 
        \wRegOut_1_0[25] , \wRegOut_1_0[24] , \wRegOut_1_0[23] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[21] , \wRegOut_1_0[20] , 
        \wRegOut_1_0[19] , \wRegOut_1_0[18] , \wRegOut_1_0[17] , 
        \wRegOut_1_0[16] , \wRegOut_1_0[15] , \wRegOut_1_0[14] , 
        \wRegOut_1_0[13] , \wRegOut_1_0[12] , \wRegOut_1_0[11] , 
        \wRegOut_1_0[10] , \wRegOut_1_0[9] , \wRegOut_1_0[8] , 
        \wRegOut_1_0[7] , \wRegOut_1_0[6] , \wRegOut_1_0[5] , \wRegOut_1_0[4] , 
        \wRegOut_1_0[3] , \wRegOut_1_0[2] , \wRegOut_1_0[1] , \wRegOut_1_0[0] 
        }), .Enable1(\wRegEnTop_1_0[0] ), .Enable2(\wRegEnBot_1_0[0] ), .In1({
        \wRegInTop_1_0[31] , \wRegInTop_1_0[30] , \wRegInTop_1_0[29] , 
        \wRegInTop_1_0[28] , \wRegInTop_1_0[27] , \wRegInTop_1_0[26] , 
        \wRegInTop_1_0[25] , \wRegInTop_1_0[24] , \wRegInTop_1_0[23] , 
        \wRegInTop_1_0[22] , \wRegInTop_1_0[21] , \wRegInTop_1_0[20] , 
        \wRegInTop_1_0[19] , \wRegInTop_1_0[18] , \wRegInTop_1_0[17] , 
        \wRegInTop_1_0[16] , \wRegInTop_1_0[15] , \wRegInTop_1_0[14] , 
        \wRegInTop_1_0[13] , \wRegInTop_1_0[12] , \wRegInTop_1_0[11] , 
        \wRegInTop_1_0[10] , \wRegInTop_1_0[9] , \wRegInTop_1_0[8] , 
        \wRegInTop_1_0[7] , \wRegInTop_1_0[6] , \wRegInTop_1_0[5] , 
        \wRegInTop_1_0[4] , \wRegInTop_1_0[3] , \wRegInTop_1_0[2] , 
        \wRegInTop_1_0[1] , \wRegInTop_1_0[0] }), .In2({\wRegInBot_1_0[31] , 
        \wRegInBot_1_0[30] , \wRegInBot_1_0[29] , \wRegInBot_1_0[28] , 
        \wRegInBot_1_0[27] , \wRegInBot_1_0[26] , \wRegInBot_1_0[25] , 
        \wRegInBot_1_0[24] , \wRegInBot_1_0[23] , \wRegInBot_1_0[22] , 
        \wRegInBot_1_0[21] , \wRegInBot_1_0[20] , \wRegInBot_1_0[19] , 
        \wRegInBot_1_0[18] , \wRegInBot_1_0[17] , \wRegInBot_1_0[16] , 
        \wRegInBot_1_0[15] , \wRegInBot_1_0[14] , \wRegInBot_1_0[13] , 
        \wRegInBot_1_0[12] , \wRegInBot_1_0[11] , \wRegInBot_1_0[10] , 
        \wRegInBot_1_0[9] , \wRegInBot_1_0[8] , \wRegInBot_1_0[7] , 
        \wRegInBot_1_0[6] , \wRegInBot_1_0[5] , \wRegInBot_1_0[4] , 
        \wRegInBot_1_0[3] , \wRegInBot_1_0[2] , \wRegInBot_1_0[1] , 
        \wRegInBot_1_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink22[31] , \ScanLink22[30] , \ScanLink22[29] , 
        \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , \ScanLink22[25] , 
        \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , \ScanLink22[21] , 
        \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , \ScanLink22[17] , 
        \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , \ScanLink22[13] , 
        \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , \ScanLink22[9] , 
        \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , \ScanLink22[5] , 
        \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , \ScanLink22[1] , 
        \ScanLink22[0] }), .ScanOut({\ScanLink21[31] , \ScanLink21[30] , 
        \ScanLink21[29] , \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , 
        \ScanLink21[25] , \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , 
        \ScanLink21[21] , \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , 
        \ScanLink21[17] , \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , 
        \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , 
        \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , 
        \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , 
        \ScanLink21[1] , \ScanLink21[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_6[31] , \wRegOut_4_6[30] , \wRegOut_4_6[29] , 
        \wRegOut_4_6[28] , \wRegOut_4_6[27] , \wRegOut_4_6[26] , 
        \wRegOut_4_6[25] , \wRegOut_4_6[24] , \wRegOut_4_6[23] , 
        \wRegOut_4_6[22] , \wRegOut_4_6[21] , \wRegOut_4_6[20] , 
        \wRegOut_4_6[19] , \wRegOut_4_6[18] , \wRegOut_4_6[17] , 
        \wRegOut_4_6[16] , \wRegOut_4_6[15] , \wRegOut_4_6[14] , 
        \wRegOut_4_6[13] , \wRegOut_4_6[12] , \wRegOut_4_6[11] , 
        \wRegOut_4_6[10] , \wRegOut_4_6[9] , \wRegOut_4_6[8] , 
        \wRegOut_4_6[7] , \wRegOut_4_6[6] , \wRegOut_4_6[5] , \wRegOut_4_6[4] , 
        \wRegOut_4_6[3] , \wRegOut_4_6[2] , \wRegOut_4_6[1] , \wRegOut_4_6[0] 
        }), .Enable1(\wRegEnTop_4_6[0] ), .Enable2(\wRegEnBot_4_6[0] ), .In1({
        \wRegInTop_4_6[31] , \wRegInTop_4_6[30] , \wRegInTop_4_6[29] , 
        \wRegInTop_4_6[28] , \wRegInTop_4_6[27] , \wRegInTop_4_6[26] , 
        \wRegInTop_4_6[25] , \wRegInTop_4_6[24] , \wRegInTop_4_6[23] , 
        \wRegInTop_4_6[22] , \wRegInTop_4_6[21] , \wRegInTop_4_6[20] , 
        \wRegInTop_4_6[19] , \wRegInTop_4_6[18] , \wRegInTop_4_6[17] , 
        \wRegInTop_4_6[16] , \wRegInTop_4_6[15] , \wRegInTop_4_6[14] , 
        \wRegInTop_4_6[13] , \wRegInTop_4_6[12] , \wRegInTop_4_6[11] , 
        \wRegInTop_4_6[10] , \wRegInTop_4_6[9] , \wRegInTop_4_6[8] , 
        \wRegInTop_4_6[7] , \wRegInTop_4_6[6] , \wRegInTop_4_6[5] , 
        \wRegInTop_4_6[4] , \wRegInTop_4_6[3] , \wRegInTop_4_6[2] , 
        \wRegInTop_4_6[1] , \wRegInTop_4_6[0] }), .In2({\wRegInBot_4_6[31] , 
        \wRegInBot_4_6[30] , \wRegInBot_4_6[29] , \wRegInBot_4_6[28] , 
        \wRegInBot_4_6[27] , \wRegInBot_4_6[26] , \wRegInBot_4_6[25] , 
        \wRegInBot_4_6[24] , \wRegInBot_4_6[23] , \wRegInBot_4_6[22] , 
        \wRegInBot_4_6[21] , \wRegInBot_4_6[20] , \wRegInBot_4_6[19] , 
        \wRegInBot_4_6[18] , \wRegInBot_4_6[17] , \wRegInBot_4_6[16] , 
        \wRegInBot_4_6[15] , \wRegInBot_4_6[14] , \wRegInBot_4_6[13] , 
        \wRegInBot_4_6[12] , \wRegInBot_4_6[11] , \wRegInBot_4_6[10] , 
        \wRegInBot_4_6[9] , \wRegInBot_4_6[8] , \wRegInBot_4_6[7] , 
        \wRegInBot_4_6[6] , \wRegInBot_4_6[5] , \wRegInBot_4_6[4] , 
        \wRegInBot_4_6[3] , \wRegInBot_4_6[2] , \wRegInBot_4_6[1] , 
        \wRegInBot_4_6[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink28[31] , \ScanLink28[30] , \ScanLink28[29] , 
        \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , \ScanLink28[25] , 
        \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , \ScanLink28[21] , 
        \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , \ScanLink28[17] , 
        \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , \ScanLink28[13] , 
        \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , \ScanLink28[9] , 
        \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , \ScanLink28[5] , 
        \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , \ScanLink28[1] , 
        \ScanLink28[0] }), .ScanOut({\ScanLink27[31] , \ScanLink27[30] , 
        \ScanLink27[29] , \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , 
        \ScanLink27[25] , \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , 
        \ScanLink27[21] , \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , 
        \ScanLink27[17] , \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , 
        \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , 
        \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , 
        \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , 
        \ScanLink27[1] , \ScanLink27[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_12[31] , \wRegOut_4_12[30] , 
        \wRegOut_4_12[29] , \wRegOut_4_12[28] , \wRegOut_4_12[27] , 
        \wRegOut_4_12[26] , \wRegOut_4_12[25] , \wRegOut_4_12[24] , 
        \wRegOut_4_12[23] , \wRegOut_4_12[22] , \wRegOut_4_12[21] , 
        \wRegOut_4_12[20] , \wRegOut_4_12[19] , \wRegOut_4_12[18] , 
        \wRegOut_4_12[17] , \wRegOut_4_12[16] , \wRegOut_4_12[15] , 
        \wRegOut_4_12[14] , \wRegOut_4_12[13] , \wRegOut_4_12[12] , 
        \wRegOut_4_12[11] , \wRegOut_4_12[10] , \wRegOut_4_12[9] , 
        \wRegOut_4_12[8] , \wRegOut_4_12[7] , \wRegOut_4_12[6] , 
        \wRegOut_4_12[5] , \wRegOut_4_12[4] , \wRegOut_4_12[3] , 
        \wRegOut_4_12[2] , \wRegOut_4_12[1] , \wRegOut_4_12[0] }), .Enable1(
        \wRegEnTop_4_12[0] ), .Enable2(\wRegEnBot_4_12[0] ), .In1({
        \wRegInTop_4_12[31] , \wRegInTop_4_12[30] , \wRegInTop_4_12[29] , 
        \wRegInTop_4_12[28] , \wRegInTop_4_12[27] , \wRegInTop_4_12[26] , 
        \wRegInTop_4_12[25] , \wRegInTop_4_12[24] , \wRegInTop_4_12[23] , 
        \wRegInTop_4_12[22] , \wRegInTop_4_12[21] , \wRegInTop_4_12[20] , 
        \wRegInTop_4_12[19] , \wRegInTop_4_12[18] , \wRegInTop_4_12[17] , 
        \wRegInTop_4_12[16] , \wRegInTop_4_12[15] , \wRegInTop_4_12[14] , 
        \wRegInTop_4_12[13] , \wRegInTop_4_12[12] , \wRegInTop_4_12[11] , 
        \wRegInTop_4_12[10] , \wRegInTop_4_12[9] , \wRegInTop_4_12[8] , 
        \wRegInTop_4_12[7] , \wRegInTop_4_12[6] , \wRegInTop_4_12[5] , 
        \wRegInTop_4_12[4] , \wRegInTop_4_12[3] , \wRegInTop_4_12[2] , 
        \wRegInTop_4_12[1] , \wRegInTop_4_12[0] }), .In2({\wRegInBot_4_12[31] , 
        \wRegInBot_4_12[30] , \wRegInBot_4_12[29] , \wRegInBot_4_12[28] , 
        \wRegInBot_4_12[27] , \wRegInBot_4_12[26] , \wRegInBot_4_12[25] , 
        \wRegInBot_4_12[24] , \wRegInBot_4_12[23] , \wRegInBot_4_12[22] , 
        \wRegInBot_4_12[21] , \wRegInBot_4_12[20] , \wRegInBot_4_12[19] , 
        \wRegInBot_4_12[18] , \wRegInBot_4_12[17] , \wRegInBot_4_12[16] , 
        \wRegInBot_4_12[15] , \wRegInBot_4_12[14] , \wRegInBot_4_12[13] , 
        \wRegInBot_4_12[12] , \wRegInBot_4_12[11] , \wRegInBot_4_12[10] , 
        \wRegInBot_4_12[9] , \wRegInBot_4_12[8] , \wRegInBot_4_12[7] , 
        \wRegInBot_4_12[6] , \wRegInBot_4_12[5] , \wRegInBot_4_12[4] , 
        \wRegInBot_4_12[3] , \wRegInBot_4_12[2] , \wRegInBot_4_12[1] , 
        \wRegInBot_4_12[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink38[31] , \ScanLink38[30] , \ScanLink38[29] , 
        \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , \ScanLink38[25] , 
        \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , \ScanLink38[21] , 
        \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , \ScanLink38[17] , 
        \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , \ScanLink38[13] , 
        \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , \ScanLink38[9] , 
        \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , \ScanLink38[5] , 
        \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , \ScanLink38[1] , 
        \ScanLink38[0] }), .ScanOut({\ScanLink37[31] , \ScanLink37[30] , 
        \ScanLink37[29] , \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , 
        \ScanLink37[25] , \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , 
        \ScanLink37[21] , \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , 
        \ScanLink37[17] , \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , 
        \ScanLink37[13] , \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , 
        \ScanLink37[9] , \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , 
        \ScanLink37[5] , \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , 
        \ScanLink37[1] , \ScanLink37[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_6[31] , \wRegOut_5_6[30] , \wRegOut_5_6[29] , 
        \wRegOut_5_6[28] , \wRegOut_5_6[27] , \wRegOut_5_6[26] , 
        \wRegOut_5_6[25] , \wRegOut_5_6[24] , \wRegOut_5_6[23] , 
        \wRegOut_5_6[22] , \wRegOut_5_6[21] , \wRegOut_5_6[20] , 
        \wRegOut_5_6[19] , \wRegOut_5_6[18] , \wRegOut_5_6[17] , 
        \wRegOut_5_6[16] , \wRegOut_5_6[15] , \wRegOut_5_6[14] , 
        \wRegOut_5_6[13] , \wRegOut_5_6[12] , \wRegOut_5_6[11] , 
        \wRegOut_5_6[10] , \wRegOut_5_6[9] , \wRegOut_5_6[8] , 
        \wRegOut_5_6[7] , \wRegOut_5_6[6] , \wRegOut_5_6[5] , \wRegOut_5_6[4] , 
        \wRegOut_5_6[3] , \wRegOut_5_6[2] , \wRegOut_5_6[1] , \wRegOut_5_6[0] 
        }), .Enable1(\wRegEnTop_5_6[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_6[31] , \wRegInTop_5_6[30] , \wRegInTop_5_6[29] , 
        \wRegInTop_5_6[28] , \wRegInTop_5_6[27] , \wRegInTop_5_6[26] , 
        \wRegInTop_5_6[25] , \wRegInTop_5_6[24] , \wRegInTop_5_6[23] , 
        \wRegInTop_5_6[22] , \wRegInTop_5_6[21] , \wRegInTop_5_6[20] , 
        \wRegInTop_5_6[19] , \wRegInTop_5_6[18] , \wRegInTop_5_6[17] , 
        \wRegInTop_5_6[16] , \wRegInTop_5_6[15] , \wRegInTop_5_6[14] , 
        \wRegInTop_5_6[13] , \wRegInTop_5_6[12] , \wRegInTop_5_6[11] , 
        \wRegInTop_5_6[10] , \wRegInTop_5_6[9] , \wRegInTop_5_6[8] , 
        \wRegInTop_5_6[7] , \wRegInTop_5_6[6] , \wRegInTop_5_6[5] , 
        \wRegInTop_5_6[4] , \wRegInTop_5_6[3] , \wRegInTop_5_6[2] , 
        \wRegInTop_5_6[1] , \wRegInTop_5_6[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_4[0] ), .P_In({\wRegOut_4_4[31] , 
        \wRegOut_4_4[30] , \wRegOut_4_4[29] , \wRegOut_4_4[28] , 
        \wRegOut_4_4[27] , \wRegOut_4_4[26] , \wRegOut_4_4[25] , 
        \wRegOut_4_4[24] , \wRegOut_4_4[23] , \wRegOut_4_4[22] , 
        \wRegOut_4_4[21] , \wRegOut_4_4[20] , \wRegOut_4_4[19] , 
        \wRegOut_4_4[18] , \wRegOut_4_4[17] , \wRegOut_4_4[16] , 
        \wRegOut_4_4[15] , \wRegOut_4_4[14] , \wRegOut_4_4[13] , 
        \wRegOut_4_4[12] , \wRegOut_4_4[11] , \wRegOut_4_4[10] , 
        \wRegOut_4_4[9] , \wRegOut_4_4[8] , \wRegOut_4_4[7] , \wRegOut_4_4[6] , 
        \wRegOut_4_4[5] , \wRegOut_4_4[4] , \wRegOut_4_4[3] , \wRegOut_4_4[2] , 
        \wRegOut_4_4[1] , \wRegOut_4_4[0] }), .P_Out({\wRegInBot_4_4[31] , 
        \wRegInBot_4_4[30] , \wRegInBot_4_4[29] , \wRegInBot_4_4[28] , 
        \wRegInBot_4_4[27] , \wRegInBot_4_4[26] , \wRegInBot_4_4[25] , 
        \wRegInBot_4_4[24] , \wRegInBot_4_4[23] , \wRegInBot_4_4[22] , 
        \wRegInBot_4_4[21] , \wRegInBot_4_4[20] , \wRegInBot_4_4[19] , 
        \wRegInBot_4_4[18] , \wRegInBot_4_4[17] , \wRegInBot_4_4[16] , 
        \wRegInBot_4_4[15] , \wRegInBot_4_4[14] , \wRegInBot_4_4[13] , 
        \wRegInBot_4_4[12] , \wRegInBot_4_4[11] , \wRegInBot_4_4[10] , 
        \wRegInBot_4_4[9] , \wRegInBot_4_4[8] , \wRegInBot_4_4[7] , 
        \wRegInBot_4_4[6] , \wRegInBot_4_4[5] , \wRegInBot_4_4[4] , 
        \wRegInBot_4_4[3] , \wRegInBot_4_4[2] , \wRegInBot_4_4[1] , 
        \wRegInBot_4_4[0] }), .L_WR(\wRegEnTop_5_8[0] ), .L_In({
        \wRegOut_5_8[31] , \wRegOut_5_8[30] , \wRegOut_5_8[29] , 
        \wRegOut_5_8[28] , \wRegOut_5_8[27] , \wRegOut_5_8[26] , 
        \wRegOut_5_8[25] , \wRegOut_5_8[24] , \wRegOut_5_8[23] , 
        \wRegOut_5_8[22] , \wRegOut_5_8[21] , \wRegOut_5_8[20] , 
        \wRegOut_5_8[19] , \wRegOut_5_8[18] , \wRegOut_5_8[17] , 
        \wRegOut_5_8[16] , \wRegOut_5_8[15] , \wRegOut_5_8[14] , 
        \wRegOut_5_8[13] , \wRegOut_5_8[12] , \wRegOut_5_8[11] , 
        \wRegOut_5_8[10] , \wRegOut_5_8[9] , \wRegOut_5_8[8] , 
        \wRegOut_5_8[7] , \wRegOut_5_8[6] , \wRegOut_5_8[5] , \wRegOut_5_8[4] , 
        \wRegOut_5_8[3] , \wRegOut_5_8[2] , \wRegOut_5_8[1] , \wRegOut_5_8[0] 
        }), .L_Out({\wRegInTop_5_8[31] , \wRegInTop_5_8[30] , 
        \wRegInTop_5_8[29] , \wRegInTop_5_8[28] , \wRegInTop_5_8[27] , 
        \wRegInTop_5_8[26] , \wRegInTop_5_8[25] , \wRegInTop_5_8[24] , 
        \wRegInTop_5_8[23] , \wRegInTop_5_8[22] , \wRegInTop_5_8[21] , 
        \wRegInTop_5_8[20] , \wRegInTop_5_8[19] , \wRegInTop_5_8[18] , 
        \wRegInTop_5_8[17] , \wRegInTop_5_8[16] , \wRegInTop_5_8[15] , 
        \wRegInTop_5_8[14] , \wRegInTop_5_8[13] , \wRegInTop_5_8[12] , 
        \wRegInTop_5_8[11] , \wRegInTop_5_8[10] , \wRegInTop_5_8[9] , 
        \wRegInTop_5_8[8] , \wRegInTop_5_8[7] , \wRegInTop_5_8[6] , 
        \wRegInTop_5_8[5] , \wRegInTop_5_8[4] , \wRegInTop_5_8[3] , 
        \wRegInTop_5_8[2] , \wRegInTop_5_8[1] , \wRegInTop_5_8[0] }), .R_WR(
        \wRegEnTop_5_9[0] ), .R_In({\wRegOut_5_9[31] , \wRegOut_5_9[30] , 
        \wRegOut_5_9[29] , \wRegOut_5_9[28] , \wRegOut_5_9[27] , 
        \wRegOut_5_9[26] , \wRegOut_5_9[25] , \wRegOut_5_9[24] , 
        \wRegOut_5_9[23] , \wRegOut_5_9[22] , \wRegOut_5_9[21] , 
        \wRegOut_5_9[20] , \wRegOut_5_9[19] , \wRegOut_5_9[18] , 
        \wRegOut_5_9[17] , \wRegOut_5_9[16] , \wRegOut_5_9[15] , 
        \wRegOut_5_9[14] , \wRegOut_5_9[13] , \wRegOut_5_9[12] , 
        \wRegOut_5_9[11] , \wRegOut_5_9[10] , \wRegOut_5_9[9] , 
        \wRegOut_5_9[8] , \wRegOut_5_9[7] , \wRegOut_5_9[6] , \wRegOut_5_9[5] , 
        \wRegOut_5_9[4] , \wRegOut_5_9[3] , \wRegOut_5_9[2] , \wRegOut_5_9[1] , 
        \wRegOut_5_9[0] }), .R_Out({\wRegInTop_5_9[31] , \wRegInTop_5_9[30] , 
        \wRegInTop_5_9[29] , \wRegInTop_5_9[28] , \wRegInTop_5_9[27] , 
        \wRegInTop_5_9[26] , \wRegInTop_5_9[25] , \wRegInTop_5_9[24] , 
        \wRegInTop_5_9[23] , \wRegInTop_5_9[22] , \wRegInTop_5_9[21] , 
        \wRegInTop_5_9[20] , \wRegInTop_5_9[19] , \wRegInTop_5_9[18] , 
        \wRegInTop_5_9[17] , \wRegInTop_5_9[16] , \wRegInTop_5_9[15] , 
        \wRegInTop_5_9[14] , \wRegInTop_5_9[13] , \wRegInTop_5_9[12] , 
        \wRegInTop_5_9[11] , \wRegInTop_5_9[10] , \wRegInTop_5_9[9] , 
        \wRegInTop_5_9[8] , \wRegInTop_5_9[7] , \wRegInTop_5_9[6] , 
        \wRegInTop_5_9[5] , \wRegInTop_5_9[4] , \wRegInTop_5_9[3] , 
        \wRegInTop_5_9[2] , \wRegInTop_5_9[1] , \wRegInTop_5_9[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink45[31] , \ScanLink45[30] , \ScanLink45[29] , 
        \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , \ScanLink45[25] , 
        \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , \ScanLink45[21] , 
        \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , \ScanLink45[17] , 
        \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , \ScanLink45[13] , 
        \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , \ScanLink45[9] , 
        \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , \ScanLink45[5] , 
        \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , \ScanLink45[1] , 
        \ScanLink45[0] }), .ScanOut({\ScanLink44[31] , \ScanLink44[30] , 
        \ScanLink44[29] , \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , 
        \ScanLink44[25] , \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , 
        \ScanLink44[21] , \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , 
        \ScanLink44[17] , \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , 
        \ScanLink44[13] , \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , 
        \ScanLink44[9] , \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , 
        \ScanLink44[5] , \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , 
        \ScanLink44[1] , \ScanLink44[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_13[31] , \wRegOut_5_13[30] , 
        \wRegOut_5_13[29] , \wRegOut_5_13[28] , \wRegOut_5_13[27] , 
        \wRegOut_5_13[26] , \wRegOut_5_13[25] , \wRegOut_5_13[24] , 
        \wRegOut_5_13[23] , \wRegOut_5_13[22] , \wRegOut_5_13[21] , 
        \wRegOut_5_13[20] , \wRegOut_5_13[19] , \wRegOut_5_13[18] , 
        \wRegOut_5_13[17] , \wRegOut_5_13[16] , \wRegOut_5_13[15] , 
        \wRegOut_5_13[14] , \wRegOut_5_13[13] , \wRegOut_5_13[12] , 
        \wRegOut_5_13[11] , \wRegOut_5_13[10] , \wRegOut_5_13[9] , 
        \wRegOut_5_13[8] , \wRegOut_5_13[7] , \wRegOut_5_13[6] , 
        \wRegOut_5_13[5] , \wRegOut_5_13[4] , \wRegOut_5_13[3] , 
        \wRegOut_5_13[2] , \wRegOut_5_13[1] , \wRegOut_5_13[0] }), .Enable1(
        \wRegEnTop_5_13[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_13[31] , 
        \wRegInTop_5_13[30] , \wRegInTop_5_13[29] , \wRegInTop_5_13[28] , 
        \wRegInTop_5_13[27] , \wRegInTop_5_13[26] , \wRegInTop_5_13[25] , 
        \wRegInTop_5_13[24] , \wRegInTop_5_13[23] , \wRegInTop_5_13[22] , 
        \wRegInTop_5_13[21] , \wRegInTop_5_13[20] , \wRegInTop_5_13[19] , 
        \wRegInTop_5_13[18] , \wRegInTop_5_13[17] , \wRegInTop_5_13[16] , 
        \wRegInTop_5_13[15] , \wRegInTop_5_13[14] , \wRegInTop_5_13[13] , 
        \wRegInTop_5_13[12] , \wRegInTop_5_13[11] , \wRegInTop_5_13[10] , 
        \wRegInTop_5_13[9] , \wRegInTop_5_13[8] , \wRegInTop_5_13[7] , 
        \wRegInTop_5_13[6] , \wRegInTop_5_13[5] , \wRegInTop_5_13[4] , 
        \wRegInTop_5_13[3] , \wRegInTop_5_13[2] , \wRegInTop_5_13[1] , 
        \wRegInTop_5_13[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_1_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink3[31] , \ScanLink3[30] , \ScanLink3[29] , 
        \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , \ScanLink3[25] , 
        \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , \ScanLink3[21] , 
        \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , \ScanLink3[17] , 
        \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , \ScanLink3[13] , 
        \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , \ScanLink3[9] , 
        \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , \ScanLink3[5] , 
        \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , \ScanLink3[1] , 
        \ScanLink3[0] }), .ScanOut({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_1_1[31] , \wRegOut_1_1[30] , \wRegOut_1_1[29] , 
        \wRegOut_1_1[28] , \wRegOut_1_1[27] , \wRegOut_1_1[26] , 
        \wRegOut_1_1[25] , \wRegOut_1_1[24] , \wRegOut_1_1[23] , 
        \wRegOut_1_1[22] , \wRegOut_1_1[21] , \wRegOut_1_1[20] , 
        \wRegOut_1_1[19] , \wRegOut_1_1[18] , \wRegOut_1_1[17] , 
        \wRegOut_1_1[16] , \wRegOut_1_1[15] , \wRegOut_1_1[14] , 
        \wRegOut_1_1[13] , \wRegOut_1_1[12] , \wRegOut_1_1[11] , 
        \wRegOut_1_1[10] , \wRegOut_1_1[9] , \wRegOut_1_1[8] , 
        \wRegOut_1_1[7] , \wRegOut_1_1[6] , \wRegOut_1_1[5] , \wRegOut_1_1[4] , 
        \wRegOut_1_1[3] , \wRegOut_1_1[2] , \wRegOut_1_1[1] , \wRegOut_1_1[0] 
        }), .Enable1(\wRegEnTop_1_1[0] ), .Enable2(\wRegEnBot_1_1[0] ), .In1({
        \wRegInTop_1_1[31] , \wRegInTop_1_1[30] , \wRegInTop_1_1[29] , 
        \wRegInTop_1_1[28] , \wRegInTop_1_1[27] , \wRegInTop_1_1[26] , 
        \wRegInTop_1_1[25] , \wRegInTop_1_1[24] , \wRegInTop_1_1[23] , 
        \wRegInTop_1_1[22] , \wRegInTop_1_1[21] , \wRegInTop_1_1[20] , 
        \wRegInTop_1_1[19] , \wRegInTop_1_1[18] , \wRegInTop_1_1[17] , 
        \wRegInTop_1_1[16] , \wRegInTop_1_1[15] , \wRegInTop_1_1[14] , 
        \wRegInTop_1_1[13] , \wRegInTop_1_1[12] , \wRegInTop_1_1[11] , 
        \wRegInTop_1_1[10] , \wRegInTop_1_1[9] , \wRegInTop_1_1[8] , 
        \wRegInTop_1_1[7] , \wRegInTop_1_1[6] , \wRegInTop_1_1[5] , 
        \wRegInTop_1_1[4] , \wRegInTop_1_1[3] , \wRegInTop_1_1[2] , 
        \wRegInTop_1_1[1] , \wRegInTop_1_1[0] }), .In2({\wRegInBot_1_1[31] , 
        \wRegInBot_1_1[30] , \wRegInBot_1_1[29] , \wRegInBot_1_1[28] , 
        \wRegInBot_1_1[27] , \wRegInBot_1_1[26] , \wRegInBot_1_1[25] , 
        \wRegInBot_1_1[24] , \wRegInBot_1_1[23] , \wRegInBot_1_1[22] , 
        \wRegInBot_1_1[21] , \wRegInBot_1_1[20] , \wRegInBot_1_1[19] , 
        \wRegInBot_1_1[18] , \wRegInBot_1_1[17] , \wRegInBot_1_1[16] , 
        \wRegInBot_1_1[15] , \wRegInBot_1_1[14] , \wRegInBot_1_1[13] , 
        \wRegInBot_1_1[12] , \wRegInBot_1_1[11] , \wRegInBot_1_1[10] , 
        \wRegInBot_1_1[9] , \wRegInBot_1_1[8] , \wRegInBot_1_1[7] , 
        \wRegInBot_1_1[6] , \wRegInBot_1_1[5] , \wRegInBot_1_1[4] , 
        \wRegInBot_1_1[3] , \wRegInBot_1_1[2] , \wRegInBot_1_1[1] , 
        \wRegInBot_1_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_2_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink6[31] , \ScanLink6[30] , \ScanLink6[29] , 
        \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , \ScanLink6[25] , 
        \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , \ScanLink6[21] , 
        \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , \ScanLink6[17] , 
        \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , \ScanLink6[13] , 
        \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , \ScanLink6[9] , 
        \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , \ScanLink6[5] , 
        \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , \ScanLink6[1] , 
        \ScanLink6[0] }), .ScanOut({\ScanLink5[31] , \ScanLink5[30] , 
        \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , 
        \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , 
        \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , 
        \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , 
        \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , 
        \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_2_2[31] , \wRegOut_2_2[30] , \wRegOut_2_2[29] , 
        \wRegOut_2_2[28] , \wRegOut_2_2[27] , \wRegOut_2_2[26] , 
        \wRegOut_2_2[25] , \wRegOut_2_2[24] , \wRegOut_2_2[23] , 
        \wRegOut_2_2[22] , \wRegOut_2_2[21] , \wRegOut_2_2[20] , 
        \wRegOut_2_2[19] , \wRegOut_2_2[18] , \wRegOut_2_2[17] , 
        \wRegOut_2_2[16] , \wRegOut_2_2[15] , \wRegOut_2_2[14] , 
        \wRegOut_2_2[13] , \wRegOut_2_2[12] , \wRegOut_2_2[11] , 
        \wRegOut_2_2[10] , \wRegOut_2_2[9] , \wRegOut_2_2[8] , 
        \wRegOut_2_2[7] , \wRegOut_2_2[6] , \wRegOut_2_2[5] , \wRegOut_2_2[4] , 
        \wRegOut_2_2[3] , \wRegOut_2_2[2] , \wRegOut_2_2[1] , \wRegOut_2_2[0] 
        }), .Enable1(\wRegEnTop_2_2[0] ), .Enable2(\wRegEnBot_2_2[0] ), .In1({
        \wRegInTop_2_2[31] , \wRegInTop_2_2[30] , \wRegInTop_2_2[29] , 
        \wRegInTop_2_2[28] , \wRegInTop_2_2[27] , \wRegInTop_2_2[26] , 
        \wRegInTop_2_2[25] , \wRegInTop_2_2[24] , \wRegInTop_2_2[23] , 
        \wRegInTop_2_2[22] , \wRegInTop_2_2[21] , \wRegInTop_2_2[20] , 
        \wRegInTop_2_2[19] , \wRegInTop_2_2[18] , \wRegInTop_2_2[17] , 
        \wRegInTop_2_2[16] , \wRegInTop_2_2[15] , \wRegInTop_2_2[14] , 
        \wRegInTop_2_2[13] , \wRegInTop_2_2[12] , \wRegInTop_2_2[11] , 
        \wRegInTop_2_2[10] , \wRegInTop_2_2[9] , \wRegInTop_2_2[8] , 
        \wRegInTop_2_2[7] , \wRegInTop_2_2[6] , \wRegInTop_2_2[5] , 
        \wRegInTop_2_2[4] , \wRegInTop_2_2[3] , \wRegInTop_2_2[2] , 
        \wRegInTop_2_2[1] , \wRegInTop_2_2[0] }), .In2({\wRegInBot_2_2[31] , 
        \wRegInBot_2_2[30] , \wRegInBot_2_2[29] , \wRegInBot_2_2[28] , 
        \wRegInBot_2_2[27] , \wRegInBot_2_2[26] , \wRegInBot_2_2[25] , 
        \wRegInBot_2_2[24] , \wRegInBot_2_2[23] , \wRegInBot_2_2[22] , 
        \wRegInBot_2_2[21] , \wRegInBot_2_2[20] , \wRegInBot_2_2[19] , 
        \wRegInBot_2_2[18] , \wRegInBot_2_2[17] , \wRegInBot_2_2[16] , 
        \wRegInBot_2_2[15] , \wRegInBot_2_2[14] , \wRegInBot_2_2[13] , 
        \wRegInBot_2_2[12] , \wRegInBot_2_2[11] , \wRegInBot_2_2[10] , 
        \wRegInBot_2_2[9] , \wRegInBot_2_2[8] , \wRegInBot_2_2[7] , 
        \wRegInBot_2_2[6] , \wRegInBot_2_2[5] , \wRegInBot_2_2[4] , 
        \wRegInBot_2_2[3] , \wRegInBot_2_2[2] , \wRegInBot_2_2[1] , 
        \wRegInBot_2_2[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink10[31] , \ScanLink10[30] , \ScanLink10[29] , 
        \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , \ScanLink10[25] , 
        \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , \ScanLink10[21] , 
        \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , \ScanLink10[17] , 
        \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , \ScanLink10[13] , 
        \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , \ScanLink10[9] , 
        \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , \ScanLink10[5] , 
        \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , \ScanLink10[1] , 
        \ScanLink10[0] }), .ScanOut({\ScanLink9[31] , \ScanLink9[30] , 
        \ScanLink9[29] , \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , 
        \ScanLink9[25] , \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , 
        \ScanLink9[21] , \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , 
        \ScanLink9[17] , \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , 
        \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , 
        \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , 
        \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , 
        \ScanLink9[1] , \ScanLink9[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_2[31] , \wRegOut_3_2[30] , \wRegOut_3_2[29] , 
        \wRegOut_3_2[28] , \wRegOut_3_2[27] , \wRegOut_3_2[26] , 
        \wRegOut_3_2[25] , \wRegOut_3_2[24] , \wRegOut_3_2[23] , 
        \wRegOut_3_2[22] , \wRegOut_3_2[21] , \wRegOut_3_2[20] , 
        \wRegOut_3_2[19] , \wRegOut_3_2[18] , \wRegOut_3_2[17] , 
        \wRegOut_3_2[16] , \wRegOut_3_2[15] , \wRegOut_3_2[14] , 
        \wRegOut_3_2[13] , \wRegOut_3_2[12] , \wRegOut_3_2[11] , 
        \wRegOut_3_2[10] , \wRegOut_3_2[9] , \wRegOut_3_2[8] , 
        \wRegOut_3_2[7] , \wRegOut_3_2[6] , \wRegOut_3_2[5] , \wRegOut_3_2[4] , 
        \wRegOut_3_2[3] , \wRegOut_3_2[2] , \wRegOut_3_2[1] , \wRegOut_3_2[0] 
        }), .Enable1(\wRegEnTop_3_2[0] ), .Enable2(\wRegEnBot_3_2[0] ), .In1({
        \wRegInTop_3_2[31] , \wRegInTop_3_2[30] , \wRegInTop_3_2[29] , 
        \wRegInTop_3_2[28] , \wRegInTop_3_2[27] , \wRegInTop_3_2[26] , 
        \wRegInTop_3_2[25] , \wRegInTop_3_2[24] , \wRegInTop_3_2[23] , 
        \wRegInTop_3_2[22] , \wRegInTop_3_2[21] , \wRegInTop_3_2[20] , 
        \wRegInTop_3_2[19] , \wRegInTop_3_2[18] , \wRegInTop_3_2[17] , 
        \wRegInTop_3_2[16] , \wRegInTop_3_2[15] , \wRegInTop_3_2[14] , 
        \wRegInTop_3_2[13] , \wRegInTop_3_2[12] , \wRegInTop_3_2[11] , 
        \wRegInTop_3_2[10] , \wRegInTop_3_2[9] , \wRegInTop_3_2[8] , 
        \wRegInTop_3_2[7] , \wRegInTop_3_2[6] , \wRegInTop_3_2[5] , 
        \wRegInTop_3_2[4] , \wRegInTop_3_2[3] , \wRegInTop_3_2[2] , 
        \wRegInTop_3_2[1] , \wRegInTop_3_2[0] }), .In2({\wRegInBot_3_2[31] , 
        \wRegInBot_3_2[30] , \wRegInBot_3_2[29] , \wRegInBot_3_2[28] , 
        \wRegInBot_3_2[27] , \wRegInBot_3_2[26] , \wRegInBot_3_2[25] , 
        \wRegInBot_3_2[24] , \wRegInBot_3_2[23] , \wRegInBot_3_2[22] , 
        \wRegInBot_3_2[21] , \wRegInBot_3_2[20] , \wRegInBot_3_2[19] , 
        \wRegInBot_3_2[18] , \wRegInBot_3_2[17] , \wRegInBot_3_2[16] , 
        \wRegInBot_3_2[15] , \wRegInBot_3_2[14] , \wRegInBot_3_2[13] , 
        \wRegInBot_3_2[12] , \wRegInBot_3_2[11] , \wRegInBot_3_2[10] , 
        \wRegInBot_3_2[9] , \wRegInBot_3_2[8] , \wRegInBot_3_2[7] , 
        \wRegInBot_3_2[6] , \wRegInBot_3_2[5] , \wRegInBot_3_2[4] , 
        \wRegInBot_3_2[3] , \wRegInBot_3_2[2] , \wRegInBot_3_2[1] , 
        \wRegInBot_3_2[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink17[31] , \ScanLink17[30] , \ScanLink17[29] , 
        \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , \ScanLink17[25] , 
        \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , \ScanLink17[21] , 
        \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , \ScanLink17[17] , 
        \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , \ScanLink17[13] , 
        \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , \ScanLink17[9] , 
        \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , \ScanLink17[5] , 
        \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , \ScanLink17[1] , 
        \ScanLink17[0] }), .ScanOut({\ScanLink16[31] , \ScanLink16[30] , 
        \ScanLink16[29] , \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , 
        \ScanLink16[25] , \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , 
        \ScanLink16[21] , \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , 
        \ScanLink16[17] , \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , 
        \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , 
        \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , 
        \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , 
        \ScanLink16[1] , \ScanLink16[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_1[31] , \wRegOut_4_1[30] , \wRegOut_4_1[29] , 
        \wRegOut_4_1[28] , \wRegOut_4_1[27] , \wRegOut_4_1[26] , 
        \wRegOut_4_1[25] , \wRegOut_4_1[24] , \wRegOut_4_1[23] , 
        \wRegOut_4_1[22] , \wRegOut_4_1[21] , \wRegOut_4_1[20] , 
        \wRegOut_4_1[19] , \wRegOut_4_1[18] , \wRegOut_4_1[17] , 
        \wRegOut_4_1[16] , \wRegOut_4_1[15] , \wRegOut_4_1[14] , 
        \wRegOut_4_1[13] , \wRegOut_4_1[12] , \wRegOut_4_1[11] , 
        \wRegOut_4_1[10] , \wRegOut_4_1[9] , \wRegOut_4_1[8] , 
        \wRegOut_4_1[7] , \wRegOut_4_1[6] , \wRegOut_4_1[5] , \wRegOut_4_1[4] , 
        \wRegOut_4_1[3] , \wRegOut_4_1[2] , \wRegOut_4_1[1] , \wRegOut_4_1[0] 
        }), .Enable1(\wRegEnTop_4_1[0] ), .Enable2(\wRegEnBot_4_1[0] ), .In1({
        \wRegInTop_4_1[31] , \wRegInTop_4_1[30] , \wRegInTop_4_1[29] , 
        \wRegInTop_4_1[28] , \wRegInTop_4_1[27] , \wRegInTop_4_1[26] , 
        \wRegInTop_4_1[25] , \wRegInTop_4_1[24] , \wRegInTop_4_1[23] , 
        \wRegInTop_4_1[22] , \wRegInTop_4_1[21] , \wRegInTop_4_1[20] , 
        \wRegInTop_4_1[19] , \wRegInTop_4_1[18] , \wRegInTop_4_1[17] , 
        \wRegInTop_4_1[16] , \wRegInTop_4_1[15] , \wRegInTop_4_1[14] , 
        \wRegInTop_4_1[13] , \wRegInTop_4_1[12] , \wRegInTop_4_1[11] , 
        \wRegInTop_4_1[10] , \wRegInTop_4_1[9] , \wRegInTop_4_1[8] , 
        \wRegInTop_4_1[7] , \wRegInTop_4_1[6] , \wRegInTop_4_1[5] , 
        \wRegInTop_4_1[4] , \wRegInTop_4_1[3] , \wRegInTop_4_1[2] , 
        \wRegInTop_4_1[1] , \wRegInTop_4_1[0] }), .In2({\wRegInBot_4_1[31] , 
        \wRegInBot_4_1[30] , \wRegInBot_4_1[29] , \wRegInBot_4_1[28] , 
        \wRegInBot_4_1[27] , \wRegInBot_4_1[26] , \wRegInBot_4_1[25] , 
        \wRegInBot_4_1[24] , \wRegInBot_4_1[23] , \wRegInBot_4_1[22] , 
        \wRegInBot_4_1[21] , \wRegInBot_4_1[20] , \wRegInBot_4_1[19] , 
        \wRegInBot_4_1[18] , \wRegInBot_4_1[17] , \wRegInBot_4_1[16] , 
        \wRegInBot_4_1[15] , \wRegInBot_4_1[14] , \wRegInBot_4_1[13] , 
        \wRegInBot_4_1[12] , \wRegInBot_4_1[11] , \wRegInBot_4_1[10] , 
        \wRegInBot_4_1[9] , \wRegInBot_4_1[8] , \wRegInBot_4_1[7] , 
        \wRegInBot_4_1[6] , \wRegInBot_4_1[5] , \wRegInBot_4_1[4] , 
        \wRegInBot_4_1[3] , \wRegInBot_4_1[2] , \wRegInBot_4_1[1] , 
        \wRegInBot_4_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink46[31] , \ScanLink46[30] , \ScanLink46[29] , 
        \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , \ScanLink46[25] , 
        \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , \ScanLink46[21] , 
        \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , \ScanLink46[17] , 
        \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , \ScanLink46[13] , 
        \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , \ScanLink46[9] , 
        \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , \ScanLink46[5] , 
        \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , \ScanLink46[1] , 
        \ScanLink46[0] }), .ScanOut({\ScanLink45[31] , \ScanLink45[30] , 
        \ScanLink45[29] , \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , 
        \ScanLink45[25] , \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , 
        \ScanLink45[21] , \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , 
        \ScanLink45[17] , \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , 
        \ScanLink45[13] , \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , 
        \ScanLink45[9] , \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , 
        \ScanLink45[5] , \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , 
        \ScanLink45[1] , \ScanLink45[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_14[31] , \wRegOut_5_14[30] , 
        \wRegOut_5_14[29] , \wRegOut_5_14[28] , \wRegOut_5_14[27] , 
        \wRegOut_5_14[26] , \wRegOut_5_14[25] , \wRegOut_5_14[24] , 
        \wRegOut_5_14[23] , \wRegOut_5_14[22] , \wRegOut_5_14[21] , 
        \wRegOut_5_14[20] , \wRegOut_5_14[19] , \wRegOut_5_14[18] , 
        \wRegOut_5_14[17] , \wRegOut_5_14[16] , \wRegOut_5_14[15] , 
        \wRegOut_5_14[14] , \wRegOut_5_14[13] , \wRegOut_5_14[12] , 
        \wRegOut_5_14[11] , \wRegOut_5_14[10] , \wRegOut_5_14[9] , 
        \wRegOut_5_14[8] , \wRegOut_5_14[7] , \wRegOut_5_14[6] , 
        \wRegOut_5_14[5] , \wRegOut_5_14[4] , \wRegOut_5_14[3] , 
        \wRegOut_5_14[2] , \wRegOut_5_14[1] , \wRegOut_5_14[0] }), .Enable1(
        \wRegEnTop_5_14[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_14[31] , 
        \wRegInTop_5_14[30] , \wRegInTop_5_14[29] , \wRegInTop_5_14[28] , 
        \wRegInTop_5_14[27] , \wRegInTop_5_14[26] , \wRegInTop_5_14[25] , 
        \wRegInTop_5_14[24] , \wRegInTop_5_14[23] , \wRegInTop_5_14[22] , 
        \wRegInTop_5_14[21] , \wRegInTop_5_14[20] , \wRegInTop_5_14[19] , 
        \wRegInTop_5_14[18] , \wRegInTop_5_14[17] , \wRegInTop_5_14[16] , 
        \wRegInTop_5_14[15] , \wRegInTop_5_14[14] , \wRegInTop_5_14[13] , 
        \wRegInTop_5_14[12] , \wRegInTop_5_14[11] , \wRegInTop_5_14[10] , 
        \wRegInTop_5_14[9] , \wRegInTop_5_14[8] , \wRegInTop_5_14[7] , 
        \wRegInTop_5_14[6] , \wRegInTop_5_14[5] , \wRegInTop_5_14[4] , 
        \wRegInTop_5_14[3] , \wRegInTop_5_14[2] , \wRegInTop_5_14[1] , 
        \wRegInTop_5_14[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink31[31] , \ScanLink31[30] , \ScanLink31[29] , 
        \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , \ScanLink31[25] , 
        \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , \ScanLink31[21] , 
        \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , \ScanLink31[17] , 
        \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , \ScanLink31[13] , 
        \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , \ScanLink31[9] , 
        \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , \ScanLink31[5] , 
        \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , \ScanLink31[1] , 
        \ScanLink31[0] }), .ScanOut({\ScanLink30[31] , \ScanLink30[30] , 
        \ScanLink30[29] , \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , 
        \ScanLink30[25] , \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , 
        \ScanLink30[21] , \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , 
        \ScanLink30[17] , \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , 
        \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , 
        \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , 
        \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , 
        \ScanLink30[1] , \ScanLink30[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_15[31] , \wRegOut_4_15[30] , 
        \wRegOut_4_15[29] , \wRegOut_4_15[28] , \wRegOut_4_15[27] , 
        \wRegOut_4_15[26] , \wRegOut_4_15[25] , \wRegOut_4_15[24] , 
        \wRegOut_4_15[23] , \wRegOut_4_15[22] , \wRegOut_4_15[21] , 
        \wRegOut_4_15[20] , \wRegOut_4_15[19] , \wRegOut_4_15[18] , 
        \wRegOut_4_15[17] , \wRegOut_4_15[16] , \wRegOut_4_15[15] , 
        \wRegOut_4_15[14] , \wRegOut_4_15[13] , \wRegOut_4_15[12] , 
        \wRegOut_4_15[11] , \wRegOut_4_15[10] , \wRegOut_4_15[9] , 
        \wRegOut_4_15[8] , \wRegOut_4_15[7] , \wRegOut_4_15[6] , 
        \wRegOut_4_15[5] , \wRegOut_4_15[4] , \wRegOut_4_15[3] , 
        \wRegOut_4_15[2] , \wRegOut_4_15[1] , \wRegOut_4_15[0] }), .Enable1(
        \wRegEnTop_4_15[0] ), .Enable2(\wRegEnBot_4_15[0] ), .In1({
        \wRegInTop_4_15[31] , \wRegInTop_4_15[30] , \wRegInTop_4_15[29] , 
        \wRegInTop_4_15[28] , \wRegInTop_4_15[27] , \wRegInTop_4_15[26] , 
        \wRegInTop_4_15[25] , \wRegInTop_4_15[24] , \wRegInTop_4_15[23] , 
        \wRegInTop_4_15[22] , \wRegInTop_4_15[21] , \wRegInTop_4_15[20] , 
        \wRegInTop_4_15[19] , \wRegInTop_4_15[18] , \wRegInTop_4_15[17] , 
        \wRegInTop_4_15[16] , \wRegInTop_4_15[15] , \wRegInTop_4_15[14] , 
        \wRegInTop_4_15[13] , \wRegInTop_4_15[12] , \wRegInTop_4_15[11] , 
        \wRegInTop_4_15[10] , \wRegInTop_4_15[9] , \wRegInTop_4_15[8] , 
        \wRegInTop_4_15[7] , \wRegInTop_4_15[6] , \wRegInTop_4_15[5] , 
        \wRegInTop_4_15[4] , \wRegInTop_4_15[3] , \wRegInTop_4_15[2] , 
        \wRegInTop_4_15[1] , \wRegInTop_4_15[0] }), .In2({\wRegInBot_4_15[31] , 
        \wRegInBot_4_15[30] , \wRegInBot_4_15[29] , \wRegInBot_4_15[28] , 
        \wRegInBot_4_15[27] , \wRegInBot_4_15[26] , \wRegInBot_4_15[25] , 
        \wRegInBot_4_15[24] , \wRegInBot_4_15[23] , \wRegInBot_4_15[22] , 
        \wRegInBot_4_15[21] , \wRegInBot_4_15[20] , \wRegInBot_4_15[19] , 
        \wRegInBot_4_15[18] , \wRegInBot_4_15[17] , \wRegInBot_4_15[16] , 
        \wRegInBot_4_15[15] , \wRegInBot_4_15[14] , \wRegInBot_4_15[13] , 
        \wRegInBot_4_15[12] , \wRegInBot_4_15[11] , \wRegInBot_4_15[10] , 
        \wRegInBot_4_15[9] , \wRegInBot_4_15[8] , \wRegInBot_4_15[7] , 
        \wRegInBot_4_15[6] , \wRegInBot_4_15[5] , \wRegInBot_4_15[4] , 
        \wRegInBot_4_15[3] , \wRegInBot_4_15[2] , \wRegInBot_4_15[1] , 
        \wRegInBot_4_15[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink33[31] , \ScanLink33[30] , \ScanLink33[29] , 
        \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , \ScanLink33[25] , 
        \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , \ScanLink33[21] , 
        \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , \ScanLink33[17] , 
        \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , \ScanLink33[13] , 
        \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , \ScanLink33[9] , 
        \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , \ScanLink33[5] , 
        \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , \ScanLink33[1] , 
        \ScanLink33[0] }), .ScanOut({\ScanLink32[31] , \ScanLink32[30] , 
        \ScanLink32[29] , \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , 
        \ScanLink32[25] , \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , 
        \ScanLink32[21] , \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , 
        \ScanLink32[17] , \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , 
        \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , 
        \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , 
        \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , 
        \ScanLink32[1] , \ScanLink32[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_1[31] , \wRegOut_5_1[30] , \wRegOut_5_1[29] , 
        \wRegOut_5_1[28] , \wRegOut_5_1[27] , \wRegOut_5_1[26] , 
        \wRegOut_5_1[25] , \wRegOut_5_1[24] , \wRegOut_5_1[23] , 
        \wRegOut_5_1[22] , \wRegOut_5_1[21] , \wRegOut_5_1[20] , 
        \wRegOut_5_1[19] , \wRegOut_5_1[18] , \wRegOut_5_1[17] , 
        \wRegOut_5_1[16] , \wRegOut_5_1[15] , \wRegOut_5_1[14] , 
        \wRegOut_5_1[13] , \wRegOut_5_1[12] , \wRegOut_5_1[11] , 
        \wRegOut_5_1[10] , \wRegOut_5_1[9] , \wRegOut_5_1[8] , 
        \wRegOut_5_1[7] , \wRegOut_5_1[6] , \wRegOut_5_1[5] , \wRegOut_5_1[4] , 
        \wRegOut_5_1[3] , \wRegOut_5_1[2] , \wRegOut_5_1[1] , \wRegOut_5_1[0] 
        }), .Enable1(\wRegEnTop_5_1[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_1[31] , \wRegInTop_5_1[30] , \wRegInTop_5_1[29] , 
        \wRegInTop_5_1[28] , \wRegInTop_5_1[27] , \wRegInTop_5_1[26] , 
        \wRegInTop_5_1[25] , \wRegInTop_5_1[24] , \wRegInTop_5_1[23] , 
        \wRegInTop_5_1[22] , \wRegInTop_5_1[21] , \wRegInTop_5_1[20] , 
        \wRegInTop_5_1[19] , \wRegInTop_5_1[18] , \wRegInTop_5_1[17] , 
        \wRegInTop_5_1[16] , \wRegInTop_5_1[15] , \wRegInTop_5_1[14] , 
        \wRegInTop_5_1[13] , \wRegInTop_5_1[12] , \wRegInTop_5_1[11] , 
        \wRegInTop_5_1[10] , \wRegInTop_5_1[9] , \wRegInTop_5_1[8] , 
        \wRegInTop_5_1[7] , \wRegInTop_5_1[6] , \wRegInTop_5_1[5] , 
        \wRegInTop_5_1[4] , \wRegInTop_5_1[3] , \wRegInTop_5_1[2] , 
        \wRegInTop_5_1[1] , \wRegInTop_5_1[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_28 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink60[31] , \ScanLink60[30] , \ScanLink60[29] , 
        \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , \ScanLink60[25] , 
        \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , \ScanLink60[21] , 
        \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , \ScanLink60[17] , 
        \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , \ScanLink60[13] , 
        \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , \ScanLink60[9] , 
        \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , \ScanLink60[5] , 
        \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , \ScanLink60[1] , 
        \ScanLink60[0] }), .ScanOut({\ScanLink59[31] , \ScanLink59[30] , 
        \ScanLink59[29] , \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , 
        \ScanLink59[25] , \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , 
        \ScanLink59[21] , \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , 
        \ScanLink59[17] , \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , 
        \ScanLink59[13] , \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , 
        \ScanLink59[9] , \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , 
        \ScanLink59[5] , \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , 
        \ScanLink59[1] , \ScanLink59[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_28[31] , \wRegOut_5_28[30] , 
        \wRegOut_5_28[29] , \wRegOut_5_28[28] , \wRegOut_5_28[27] , 
        \wRegOut_5_28[26] , \wRegOut_5_28[25] , \wRegOut_5_28[24] , 
        \wRegOut_5_28[23] , \wRegOut_5_28[22] , \wRegOut_5_28[21] , 
        \wRegOut_5_28[20] , \wRegOut_5_28[19] , \wRegOut_5_28[18] , 
        \wRegOut_5_28[17] , \wRegOut_5_28[16] , \wRegOut_5_28[15] , 
        \wRegOut_5_28[14] , \wRegOut_5_28[13] , \wRegOut_5_28[12] , 
        \wRegOut_5_28[11] , \wRegOut_5_28[10] , \wRegOut_5_28[9] , 
        \wRegOut_5_28[8] , \wRegOut_5_28[7] , \wRegOut_5_28[6] , 
        \wRegOut_5_28[5] , \wRegOut_5_28[4] , \wRegOut_5_28[3] , 
        \wRegOut_5_28[2] , \wRegOut_5_28[1] , \wRegOut_5_28[0] }), .Enable1(
        \wRegEnTop_5_28[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_28[31] , 
        \wRegInTop_5_28[30] , \wRegInTop_5_28[29] , \wRegInTop_5_28[28] , 
        \wRegInTop_5_28[27] , \wRegInTop_5_28[26] , \wRegInTop_5_28[25] , 
        \wRegInTop_5_28[24] , \wRegInTop_5_28[23] , \wRegInTop_5_28[22] , 
        \wRegInTop_5_28[21] , \wRegInTop_5_28[20] , \wRegInTop_5_28[19] , 
        \wRegInTop_5_28[18] , \wRegInTop_5_28[17] , \wRegInTop_5_28[16] , 
        \wRegInTop_5_28[15] , \wRegInTop_5_28[14] , \wRegInTop_5_28[13] , 
        \wRegInTop_5_28[12] , \wRegInTop_5_28[11] , \wRegInTop_5_28[10] , 
        \wRegInTop_5_28[9] , \wRegInTop_5_28[8] , \wRegInTop_5_28[7] , 
        \wRegInTop_5_28[6] , \wRegInTop_5_28[5] , \wRegInTop_5_28[4] , 
        \wRegInTop_5_28[3] , \wRegInTop_5_28[2] , \wRegInTop_5_28[1] , 
        \wRegInTop_5_28[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_3[0] ), .P_In({\wRegOut_4_3[31] , 
        \wRegOut_4_3[30] , \wRegOut_4_3[29] , \wRegOut_4_3[28] , 
        \wRegOut_4_3[27] , \wRegOut_4_3[26] , \wRegOut_4_3[25] , 
        \wRegOut_4_3[24] , \wRegOut_4_3[23] , \wRegOut_4_3[22] , 
        \wRegOut_4_3[21] , \wRegOut_4_3[20] , \wRegOut_4_3[19] , 
        \wRegOut_4_3[18] , \wRegOut_4_3[17] , \wRegOut_4_3[16] , 
        \wRegOut_4_3[15] , \wRegOut_4_3[14] , \wRegOut_4_3[13] , 
        \wRegOut_4_3[12] , \wRegOut_4_3[11] , \wRegOut_4_3[10] , 
        \wRegOut_4_3[9] , \wRegOut_4_3[8] , \wRegOut_4_3[7] , \wRegOut_4_3[6] , 
        \wRegOut_4_3[5] , \wRegOut_4_3[4] , \wRegOut_4_3[3] , \wRegOut_4_3[2] , 
        \wRegOut_4_3[1] , \wRegOut_4_3[0] }), .P_Out({\wRegInBot_4_3[31] , 
        \wRegInBot_4_3[30] , \wRegInBot_4_3[29] , \wRegInBot_4_3[28] , 
        \wRegInBot_4_3[27] , \wRegInBot_4_3[26] , \wRegInBot_4_3[25] , 
        \wRegInBot_4_3[24] , \wRegInBot_4_3[23] , \wRegInBot_4_3[22] , 
        \wRegInBot_4_3[21] , \wRegInBot_4_3[20] , \wRegInBot_4_3[19] , 
        \wRegInBot_4_3[18] , \wRegInBot_4_3[17] , \wRegInBot_4_3[16] , 
        \wRegInBot_4_3[15] , \wRegInBot_4_3[14] , \wRegInBot_4_3[13] , 
        \wRegInBot_4_3[12] , \wRegInBot_4_3[11] , \wRegInBot_4_3[10] , 
        \wRegInBot_4_3[9] , \wRegInBot_4_3[8] , \wRegInBot_4_3[7] , 
        \wRegInBot_4_3[6] , \wRegInBot_4_3[5] , \wRegInBot_4_3[4] , 
        \wRegInBot_4_3[3] , \wRegInBot_4_3[2] , \wRegInBot_4_3[1] , 
        \wRegInBot_4_3[0] }), .L_WR(\wRegEnTop_5_6[0] ), .L_In({
        \wRegOut_5_6[31] , \wRegOut_5_6[30] , \wRegOut_5_6[29] , 
        \wRegOut_5_6[28] , \wRegOut_5_6[27] , \wRegOut_5_6[26] , 
        \wRegOut_5_6[25] , \wRegOut_5_6[24] , \wRegOut_5_6[23] , 
        \wRegOut_5_6[22] , \wRegOut_5_6[21] , \wRegOut_5_6[20] , 
        \wRegOut_5_6[19] , \wRegOut_5_6[18] , \wRegOut_5_6[17] , 
        \wRegOut_5_6[16] , \wRegOut_5_6[15] , \wRegOut_5_6[14] , 
        \wRegOut_5_6[13] , \wRegOut_5_6[12] , \wRegOut_5_6[11] , 
        \wRegOut_5_6[10] , \wRegOut_5_6[9] , \wRegOut_5_6[8] , 
        \wRegOut_5_6[7] , \wRegOut_5_6[6] , \wRegOut_5_6[5] , \wRegOut_5_6[4] , 
        \wRegOut_5_6[3] , \wRegOut_5_6[2] , \wRegOut_5_6[1] , \wRegOut_5_6[0] 
        }), .L_Out({\wRegInTop_5_6[31] , \wRegInTop_5_6[30] , 
        \wRegInTop_5_6[29] , \wRegInTop_5_6[28] , \wRegInTop_5_6[27] , 
        \wRegInTop_5_6[26] , \wRegInTop_5_6[25] , \wRegInTop_5_6[24] , 
        \wRegInTop_5_6[23] , \wRegInTop_5_6[22] , \wRegInTop_5_6[21] , 
        \wRegInTop_5_6[20] , \wRegInTop_5_6[19] , \wRegInTop_5_6[18] , 
        \wRegInTop_5_6[17] , \wRegInTop_5_6[16] , \wRegInTop_5_6[15] , 
        \wRegInTop_5_6[14] , \wRegInTop_5_6[13] , \wRegInTop_5_6[12] , 
        \wRegInTop_5_6[11] , \wRegInTop_5_6[10] , \wRegInTop_5_6[9] , 
        \wRegInTop_5_6[8] , \wRegInTop_5_6[7] , \wRegInTop_5_6[6] , 
        \wRegInTop_5_6[5] , \wRegInTop_5_6[4] , \wRegInTop_5_6[3] , 
        \wRegInTop_5_6[2] , \wRegInTop_5_6[1] , \wRegInTop_5_6[0] }), .R_WR(
        \wRegEnTop_5_7[0] ), .R_In({\wRegOut_5_7[31] , \wRegOut_5_7[30] , 
        \wRegOut_5_7[29] , \wRegOut_5_7[28] , \wRegOut_5_7[27] , 
        \wRegOut_5_7[26] , \wRegOut_5_7[25] , \wRegOut_5_7[24] , 
        \wRegOut_5_7[23] , \wRegOut_5_7[22] , \wRegOut_5_7[21] , 
        \wRegOut_5_7[20] , \wRegOut_5_7[19] , \wRegOut_5_7[18] , 
        \wRegOut_5_7[17] , \wRegOut_5_7[16] , \wRegOut_5_7[15] , 
        \wRegOut_5_7[14] , \wRegOut_5_7[13] , \wRegOut_5_7[12] , 
        \wRegOut_5_7[11] , \wRegOut_5_7[10] , \wRegOut_5_7[9] , 
        \wRegOut_5_7[8] , \wRegOut_5_7[7] , \wRegOut_5_7[6] , \wRegOut_5_7[5] , 
        \wRegOut_5_7[4] , \wRegOut_5_7[3] , \wRegOut_5_7[2] , \wRegOut_5_7[1] , 
        \wRegOut_5_7[0] }), .R_Out({\wRegInTop_5_7[31] , \wRegInTop_5_7[30] , 
        \wRegInTop_5_7[29] , \wRegInTop_5_7[28] , \wRegInTop_5_7[27] , 
        \wRegInTop_5_7[26] , \wRegInTop_5_7[25] , \wRegInTop_5_7[24] , 
        \wRegInTop_5_7[23] , \wRegInTop_5_7[22] , \wRegInTop_5_7[21] , 
        \wRegInTop_5_7[20] , \wRegInTop_5_7[19] , \wRegInTop_5_7[18] , 
        \wRegInTop_5_7[17] , \wRegInTop_5_7[16] , \wRegInTop_5_7[15] , 
        \wRegInTop_5_7[14] , \wRegInTop_5_7[13] , \wRegInTop_5_7[12] , 
        \wRegInTop_5_7[11] , \wRegInTop_5_7[10] , \wRegInTop_5_7[9] , 
        \wRegInTop_5_7[8] , \wRegInTop_5_7[7] , \wRegInTop_5_7[6] , 
        \wRegInTop_5_7[5] , \wRegInTop_5_7[4] , \wRegInTop_5_7[3] , 
        \wRegInTop_5_7[2] , \wRegInTop_5_7[1] , \wRegInTop_5_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink24[31] , \ScanLink24[30] , \ScanLink24[29] , 
        \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , \ScanLink24[25] , 
        \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , \ScanLink24[21] , 
        \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , \ScanLink24[17] , 
        \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , \ScanLink24[13] , 
        \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , \ScanLink24[9] , 
        \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , \ScanLink24[5] , 
        \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , \ScanLink24[1] , 
        \ScanLink24[0] }), .ScanOut({\ScanLink23[31] , \ScanLink23[30] , 
        \ScanLink23[29] , \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , 
        \ScanLink23[25] , \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , 
        \ScanLink23[21] , \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , 
        \ScanLink23[17] , \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , 
        \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , 
        \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , 
        \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , 
        \ScanLink23[1] , \ScanLink23[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_8[31] , \wRegOut_4_8[30] , \wRegOut_4_8[29] , 
        \wRegOut_4_8[28] , \wRegOut_4_8[27] , \wRegOut_4_8[26] , 
        \wRegOut_4_8[25] , \wRegOut_4_8[24] , \wRegOut_4_8[23] , 
        \wRegOut_4_8[22] , \wRegOut_4_8[21] , \wRegOut_4_8[20] , 
        \wRegOut_4_8[19] , \wRegOut_4_8[18] , \wRegOut_4_8[17] , 
        \wRegOut_4_8[16] , \wRegOut_4_8[15] , \wRegOut_4_8[14] , 
        \wRegOut_4_8[13] , \wRegOut_4_8[12] , \wRegOut_4_8[11] , 
        \wRegOut_4_8[10] , \wRegOut_4_8[9] , \wRegOut_4_8[8] , 
        \wRegOut_4_8[7] , \wRegOut_4_8[6] , \wRegOut_4_8[5] , \wRegOut_4_8[4] , 
        \wRegOut_4_8[3] , \wRegOut_4_8[2] , \wRegOut_4_8[1] , \wRegOut_4_8[0] 
        }), .Enable1(\wRegEnTop_4_8[0] ), .Enable2(\wRegEnBot_4_8[0] ), .In1({
        \wRegInTop_4_8[31] , \wRegInTop_4_8[30] , \wRegInTop_4_8[29] , 
        \wRegInTop_4_8[28] , \wRegInTop_4_8[27] , \wRegInTop_4_8[26] , 
        \wRegInTop_4_8[25] , \wRegInTop_4_8[24] , \wRegInTop_4_8[23] , 
        \wRegInTop_4_8[22] , \wRegInTop_4_8[21] , \wRegInTop_4_8[20] , 
        \wRegInTop_4_8[19] , \wRegInTop_4_8[18] , \wRegInTop_4_8[17] , 
        \wRegInTop_4_8[16] , \wRegInTop_4_8[15] , \wRegInTop_4_8[14] , 
        \wRegInTop_4_8[13] , \wRegInTop_4_8[12] , \wRegInTop_4_8[11] , 
        \wRegInTop_4_8[10] , \wRegInTop_4_8[9] , \wRegInTop_4_8[8] , 
        \wRegInTop_4_8[7] , \wRegInTop_4_8[6] , \wRegInTop_4_8[5] , 
        \wRegInTop_4_8[4] , \wRegInTop_4_8[3] , \wRegInTop_4_8[2] , 
        \wRegInTop_4_8[1] , \wRegInTop_4_8[0] }), .In2({\wRegInBot_4_8[31] , 
        \wRegInBot_4_8[30] , \wRegInBot_4_8[29] , \wRegInBot_4_8[28] , 
        \wRegInBot_4_8[27] , \wRegInBot_4_8[26] , \wRegInBot_4_8[25] , 
        \wRegInBot_4_8[24] , \wRegInBot_4_8[23] , \wRegInBot_4_8[22] , 
        \wRegInBot_4_8[21] , \wRegInBot_4_8[20] , \wRegInBot_4_8[19] , 
        \wRegInBot_4_8[18] , \wRegInBot_4_8[17] , \wRegInBot_4_8[16] , 
        \wRegInBot_4_8[15] , \wRegInBot_4_8[14] , \wRegInBot_4_8[13] , 
        \wRegInBot_4_8[12] , \wRegInBot_4_8[11] , \wRegInBot_4_8[10] , 
        \wRegInBot_4_8[9] , \wRegInBot_4_8[8] , \wRegInBot_4_8[7] , 
        \wRegInBot_4_8[6] , \wRegInBot_4_8[5] , \wRegInBot_4_8[4] , 
        \wRegInBot_4_8[3] , \wRegInBot_4_8[2] , \wRegInBot_4_8[1] , 
        \wRegInBot_4_8[0] }) );
    BHeap_Node_WIDTH32 BHN_2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_2[0] ), .P_WR(\wRegEnBot_2_0[0] ), .P_In({\wRegOut_2_0[31] , 
        \wRegOut_2_0[30] , \wRegOut_2_0[29] , \wRegOut_2_0[28] , 
        \wRegOut_2_0[27] , \wRegOut_2_0[26] , \wRegOut_2_0[25] , 
        \wRegOut_2_0[24] , \wRegOut_2_0[23] , \wRegOut_2_0[22] , 
        \wRegOut_2_0[21] , \wRegOut_2_0[20] , \wRegOut_2_0[19] , 
        \wRegOut_2_0[18] , \wRegOut_2_0[17] , \wRegOut_2_0[16] , 
        \wRegOut_2_0[15] , \wRegOut_2_0[14] , \wRegOut_2_0[13] , 
        \wRegOut_2_0[12] , \wRegOut_2_0[11] , \wRegOut_2_0[10] , 
        \wRegOut_2_0[9] , \wRegOut_2_0[8] , \wRegOut_2_0[7] , \wRegOut_2_0[6] , 
        \wRegOut_2_0[5] , \wRegOut_2_0[4] , \wRegOut_2_0[3] , \wRegOut_2_0[2] , 
        \wRegOut_2_0[1] , \wRegOut_2_0[0] }), .P_Out({\wRegInBot_2_0[31] , 
        \wRegInBot_2_0[30] , \wRegInBot_2_0[29] , \wRegInBot_2_0[28] , 
        \wRegInBot_2_0[27] , \wRegInBot_2_0[26] , \wRegInBot_2_0[25] , 
        \wRegInBot_2_0[24] , \wRegInBot_2_0[23] , \wRegInBot_2_0[22] , 
        \wRegInBot_2_0[21] , \wRegInBot_2_0[20] , \wRegInBot_2_0[19] , 
        \wRegInBot_2_0[18] , \wRegInBot_2_0[17] , \wRegInBot_2_0[16] , 
        \wRegInBot_2_0[15] , \wRegInBot_2_0[14] , \wRegInBot_2_0[13] , 
        \wRegInBot_2_0[12] , \wRegInBot_2_0[11] , \wRegInBot_2_0[10] , 
        \wRegInBot_2_0[9] , \wRegInBot_2_0[8] , \wRegInBot_2_0[7] , 
        \wRegInBot_2_0[6] , \wRegInBot_2_0[5] , \wRegInBot_2_0[4] , 
        \wRegInBot_2_0[3] , \wRegInBot_2_0[2] , \wRegInBot_2_0[1] , 
        \wRegInBot_2_0[0] }), .L_WR(\wRegEnTop_3_0[0] ), .L_In({
        \wRegOut_3_0[31] , \wRegOut_3_0[30] , \wRegOut_3_0[29] , 
        \wRegOut_3_0[28] , \wRegOut_3_0[27] , \wRegOut_3_0[26] , 
        \wRegOut_3_0[25] , \wRegOut_3_0[24] , \wRegOut_3_0[23] , 
        \wRegOut_3_0[22] , \wRegOut_3_0[21] , \wRegOut_3_0[20] , 
        \wRegOut_3_0[19] , \wRegOut_3_0[18] , \wRegOut_3_0[17] , 
        \wRegOut_3_0[16] , \wRegOut_3_0[15] , \wRegOut_3_0[14] , 
        \wRegOut_3_0[13] , \wRegOut_3_0[12] , \wRegOut_3_0[11] , 
        \wRegOut_3_0[10] , \wRegOut_3_0[9] , \wRegOut_3_0[8] , 
        \wRegOut_3_0[7] , \wRegOut_3_0[6] , \wRegOut_3_0[5] , \wRegOut_3_0[4] , 
        \wRegOut_3_0[3] , \wRegOut_3_0[2] , \wRegOut_3_0[1] , \wRegOut_3_0[0] 
        }), .L_Out({\wRegInTop_3_0[31] , \wRegInTop_3_0[30] , 
        \wRegInTop_3_0[29] , \wRegInTop_3_0[28] , \wRegInTop_3_0[27] , 
        \wRegInTop_3_0[26] , \wRegInTop_3_0[25] , \wRegInTop_3_0[24] , 
        \wRegInTop_3_0[23] , \wRegInTop_3_0[22] , \wRegInTop_3_0[21] , 
        \wRegInTop_3_0[20] , \wRegInTop_3_0[19] , \wRegInTop_3_0[18] , 
        \wRegInTop_3_0[17] , \wRegInTop_3_0[16] , \wRegInTop_3_0[15] , 
        \wRegInTop_3_0[14] , \wRegInTop_3_0[13] , \wRegInTop_3_0[12] , 
        \wRegInTop_3_0[11] , \wRegInTop_3_0[10] , \wRegInTop_3_0[9] , 
        \wRegInTop_3_0[8] , \wRegInTop_3_0[7] , \wRegInTop_3_0[6] , 
        \wRegInTop_3_0[5] , \wRegInTop_3_0[4] , \wRegInTop_3_0[3] , 
        \wRegInTop_3_0[2] , \wRegInTop_3_0[1] , \wRegInTop_3_0[0] }), .R_WR(
        \wRegEnTop_3_1[0] ), .R_In({\wRegOut_3_1[31] , \wRegOut_3_1[30] , 
        \wRegOut_3_1[29] , \wRegOut_3_1[28] , \wRegOut_3_1[27] , 
        \wRegOut_3_1[26] , \wRegOut_3_1[25] , \wRegOut_3_1[24] , 
        \wRegOut_3_1[23] , \wRegOut_3_1[22] , \wRegOut_3_1[21] , 
        \wRegOut_3_1[20] , \wRegOut_3_1[19] , \wRegOut_3_1[18] , 
        \wRegOut_3_1[17] , \wRegOut_3_1[16] , \wRegOut_3_1[15] , 
        \wRegOut_3_1[14] , \wRegOut_3_1[13] , \wRegOut_3_1[12] , 
        \wRegOut_3_1[11] , \wRegOut_3_1[10] , \wRegOut_3_1[9] , 
        \wRegOut_3_1[8] , \wRegOut_3_1[7] , \wRegOut_3_1[6] , \wRegOut_3_1[5] , 
        \wRegOut_3_1[4] , \wRegOut_3_1[3] , \wRegOut_3_1[2] , \wRegOut_3_1[1] , 
        \wRegOut_3_1[0] }), .R_Out({\wRegInTop_3_1[31] , \wRegInTop_3_1[30] , 
        \wRegInTop_3_1[29] , \wRegInTop_3_1[28] , \wRegInTop_3_1[27] , 
        \wRegInTop_3_1[26] , \wRegInTop_3_1[25] , \wRegInTop_3_1[24] , 
        \wRegInTop_3_1[23] , \wRegInTop_3_1[22] , \wRegInTop_3_1[21] , 
        \wRegInTop_3_1[20] , \wRegInTop_3_1[19] , \wRegInTop_3_1[18] , 
        \wRegInTop_3_1[17] , \wRegInTop_3_1[16] , \wRegInTop_3_1[15] , 
        \wRegInTop_3_1[14] , \wRegInTop_3_1[13] , \wRegInTop_3_1[12] , 
        \wRegInTop_3_1[11] , \wRegInTop_3_1[10] , \wRegInTop_3_1[9] , 
        \wRegInTop_3_1[8] , \wRegInTop_3_1[7] , \wRegInTop_3_1[6] , 
        \wRegInTop_3_1[5] , \wRegInTop_3_1[4] , \wRegInTop_3_1[3] , 
        \wRegInTop_3_1[2] , \wRegInTop_3_1[1] , \wRegInTop_3_1[0] }) );
    BHeap_CtrlReg_WIDTH32 BHCR_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_5[0] ), 
        .Out(\wCtrlOut_4[0] ), .Enable(\wEnable_4[0] ) );
    BHeap_Node_WIDTH32 BHN_3_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_0[0] ), .P_In({\wRegOut_3_0[31] , 
        \wRegOut_3_0[30] , \wRegOut_3_0[29] , \wRegOut_3_0[28] , 
        \wRegOut_3_0[27] , \wRegOut_3_0[26] , \wRegOut_3_0[25] , 
        \wRegOut_3_0[24] , \wRegOut_3_0[23] , \wRegOut_3_0[22] , 
        \wRegOut_3_0[21] , \wRegOut_3_0[20] , \wRegOut_3_0[19] , 
        \wRegOut_3_0[18] , \wRegOut_3_0[17] , \wRegOut_3_0[16] , 
        \wRegOut_3_0[15] , \wRegOut_3_0[14] , \wRegOut_3_0[13] , 
        \wRegOut_3_0[12] , \wRegOut_3_0[11] , \wRegOut_3_0[10] , 
        \wRegOut_3_0[9] , \wRegOut_3_0[8] , \wRegOut_3_0[7] , \wRegOut_3_0[6] , 
        \wRegOut_3_0[5] , \wRegOut_3_0[4] , \wRegOut_3_0[3] , \wRegOut_3_0[2] , 
        \wRegOut_3_0[1] , \wRegOut_3_0[0] }), .P_Out({\wRegInBot_3_0[31] , 
        \wRegInBot_3_0[30] , \wRegInBot_3_0[29] , \wRegInBot_3_0[28] , 
        \wRegInBot_3_0[27] , \wRegInBot_3_0[26] , \wRegInBot_3_0[25] , 
        \wRegInBot_3_0[24] , \wRegInBot_3_0[23] , \wRegInBot_3_0[22] , 
        \wRegInBot_3_0[21] , \wRegInBot_3_0[20] , \wRegInBot_3_0[19] , 
        \wRegInBot_3_0[18] , \wRegInBot_3_0[17] , \wRegInBot_3_0[16] , 
        \wRegInBot_3_0[15] , \wRegInBot_3_0[14] , \wRegInBot_3_0[13] , 
        \wRegInBot_3_0[12] , \wRegInBot_3_0[11] , \wRegInBot_3_0[10] , 
        \wRegInBot_3_0[9] , \wRegInBot_3_0[8] , \wRegInBot_3_0[7] , 
        \wRegInBot_3_0[6] , \wRegInBot_3_0[5] , \wRegInBot_3_0[4] , 
        \wRegInBot_3_0[3] , \wRegInBot_3_0[2] , \wRegInBot_3_0[1] , 
        \wRegInBot_3_0[0] }), .L_WR(\wRegEnTop_4_0[0] ), .L_In({
        \wRegOut_4_0[31] , \wRegOut_4_0[30] , \wRegOut_4_0[29] , 
        \wRegOut_4_0[28] , \wRegOut_4_0[27] , \wRegOut_4_0[26] , 
        \wRegOut_4_0[25] , \wRegOut_4_0[24] , \wRegOut_4_0[23] , 
        \wRegOut_4_0[22] , \wRegOut_4_0[21] , \wRegOut_4_0[20] , 
        \wRegOut_4_0[19] , \wRegOut_4_0[18] , \wRegOut_4_0[17] , 
        \wRegOut_4_0[16] , \wRegOut_4_0[15] , \wRegOut_4_0[14] , 
        \wRegOut_4_0[13] , \wRegOut_4_0[12] , \wRegOut_4_0[11] , 
        \wRegOut_4_0[10] , \wRegOut_4_0[9] , \wRegOut_4_0[8] , 
        \wRegOut_4_0[7] , \wRegOut_4_0[6] , \wRegOut_4_0[5] , \wRegOut_4_0[4] , 
        \wRegOut_4_0[3] , \wRegOut_4_0[2] , \wRegOut_4_0[1] , \wRegOut_4_0[0] 
        }), .L_Out({\wRegInTop_4_0[31] , \wRegInTop_4_0[30] , 
        \wRegInTop_4_0[29] , \wRegInTop_4_0[28] , \wRegInTop_4_0[27] , 
        \wRegInTop_4_0[26] , \wRegInTop_4_0[25] , \wRegInTop_4_0[24] , 
        \wRegInTop_4_0[23] , \wRegInTop_4_0[22] , \wRegInTop_4_0[21] , 
        \wRegInTop_4_0[20] , \wRegInTop_4_0[19] , \wRegInTop_4_0[18] , 
        \wRegInTop_4_0[17] , \wRegInTop_4_0[16] , \wRegInTop_4_0[15] , 
        \wRegInTop_4_0[14] , \wRegInTop_4_0[13] , \wRegInTop_4_0[12] , 
        \wRegInTop_4_0[11] , \wRegInTop_4_0[10] , \wRegInTop_4_0[9] , 
        \wRegInTop_4_0[8] , \wRegInTop_4_0[7] , \wRegInTop_4_0[6] , 
        \wRegInTop_4_0[5] , \wRegInTop_4_0[4] , \wRegInTop_4_0[3] , 
        \wRegInTop_4_0[2] , \wRegInTop_4_0[1] , \wRegInTop_4_0[0] }), .R_WR(
        \wRegEnTop_4_1[0] ), .R_In({\wRegOut_4_1[31] , \wRegOut_4_1[30] , 
        \wRegOut_4_1[29] , \wRegOut_4_1[28] , \wRegOut_4_1[27] , 
        \wRegOut_4_1[26] , \wRegOut_4_1[25] , \wRegOut_4_1[24] , 
        \wRegOut_4_1[23] , \wRegOut_4_1[22] , \wRegOut_4_1[21] , 
        \wRegOut_4_1[20] , \wRegOut_4_1[19] , \wRegOut_4_1[18] , 
        \wRegOut_4_1[17] , \wRegOut_4_1[16] , \wRegOut_4_1[15] , 
        \wRegOut_4_1[14] , \wRegOut_4_1[13] , \wRegOut_4_1[12] , 
        \wRegOut_4_1[11] , \wRegOut_4_1[10] , \wRegOut_4_1[9] , 
        \wRegOut_4_1[8] , \wRegOut_4_1[7] , \wRegOut_4_1[6] , \wRegOut_4_1[5] , 
        \wRegOut_4_1[4] , \wRegOut_4_1[3] , \wRegOut_4_1[2] , \wRegOut_4_1[1] , 
        \wRegOut_4_1[0] }), .R_Out({\wRegInTop_4_1[31] , \wRegInTop_4_1[30] , 
        \wRegInTop_4_1[29] , \wRegInTop_4_1[28] , \wRegInTop_4_1[27] , 
        \wRegInTop_4_1[26] , \wRegInTop_4_1[25] , \wRegInTop_4_1[24] , 
        \wRegInTop_4_1[23] , \wRegInTop_4_1[22] , \wRegInTop_4_1[21] , 
        \wRegInTop_4_1[20] , \wRegInTop_4_1[19] , \wRegInTop_4_1[18] , 
        \wRegInTop_4_1[17] , \wRegInTop_4_1[16] , \wRegInTop_4_1[15] , 
        \wRegInTop_4_1[14] , \wRegInTop_4_1[13] , \wRegInTop_4_1[12] , 
        \wRegInTop_4_1[11] , \wRegInTop_4_1[10] , \wRegInTop_4_1[9] , 
        \wRegInTop_4_1[8] , \wRegInTop_4_1[7] , \wRegInTop_4_1[6] , 
        \wRegInTop_4_1[5] , \wRegInTop_4_1[4] , \wRegInTop_4_1[3] , 
        \wRegInTop_4_1[2] , \wRegInTop_4_1[1] , \wRegInTop_4_1[0] }) );
    BHeap_Node_WIDTH32 BHN_4_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_13[0] ), .P_In({\wRegOut_4_13[31] , 
        \wRegOut_4_13[30] , \wRegOut_4_13[29] , \wRegOut_4_13[28] , 
        \wRegOut_4_13[27] , \wRegOut_4_13[26] , \wRegOut_4_13[25] , 
        \wRegOut_4_13[24] , \wRegOut_4_13[23] , \wRegOut_4_13[22] , 
        \wRegOut_4_13[21] , \wRegOut_4_13[20] , \wRegOut_4_13[19] , 
        \wRegOut_4_13[18] , \wRegOut_4_13[17] , \wRegOut_4_13[16] , 
        \wRegOut_4_13[15] , \wRegOut_4_13[14] , \wRegOut_4_13[13] , 
        \wRegOut_4_13[12] , \wRegOut_4_13[11] , \wRegOut_4_13[10] , 
        \wRegOut_4_13[9] , \wRegOut_4_13[8] , \wRegOut_4_13[7] , 
        \wRegOut_4_13[6] , \wRegOut_4_13[5] , \wRegOut_4_13[4] , 
        \wRegOut_4_13[3] , \wRegOut_4_13[2] , \wRegOut_4_13[1] , 
        \wRegOut_4_13[0] }), .P_Out({\wRegInBot_4_13[31] , 
        \wRegInBot_4_13[30] , \wRegInBot_4_13[29] , \wRegInBot_4_13[28] , 
        \wRegInBot_4_13[27] , \wRegInBot_4_13[26] , \wRegInBot_4_13[25] , 
        \wRegInBot_4_13[24] , \wRegInBot_4_13[23] , \wRegInBot_4_13[22] , 
        \wRegInBot_4_13[21] , \wRegInBot_4_13[20] , \wRegInBot_4_13[19] , 
        \wRegInBot_4_13[18] , \wRegInBot_4_13[17] , \wRegInBot_4_13[16] , 
        \wRegInBot_4_13[15] , \wRegInBot_4_13[14] , \wRegInBot_4_13[13] , 
        \wRegInBot_4_13[12] , \wRegInBot_4_13[11] , \wRegInBot_4_13[10] , 
        \wRegInBot_4_13[9] , \wRegInBot_4_13[8] , \wRegInBot_4_13[7] , 
        \wRegInBot_4_13[6] , \wRegInBot_4_13[5] , \wRegInBot_4_13[4] , 
        \wRegInBot_4_13[3] , \wRegInBot_4_13[2] , \wRegInBot_4_13[1] , 
        \wRegInBot_4_13[0] }), .L_WR(\wRegEnTop_5_26[0] ), .L_In({
        \wRegOut_5_26[31] , \wRegOut_5_26[30] , \wRegOut_5_26[29] , 
        \wRegOut_5_26[28] , \wRegOut_5_26[27] , \wRegOut_5_26[26] , 
        \wRegOut_5_26[25] , \wRegOut_5_26[24] , \wRegOut_5_26[23] , 
        \wRegOut_5_26[22] , \wRegOut_5_26[21] , \wRegOut_5_26[20] , 
        \wRegOut_5_26[19] , \wRegOut_5_26[18] , \wRegOut_5_26[17] , 
        \wRegOut_5_26[16] , \wRegOut_5_26[15] , \wRegOut_5_26[14] , 
        \wRegOut_5_26[13] , \wRegOut_5_26[12] , \wRegOut_5_26[11] , 
        \wRegOut_5_26[10] , \wRegOut_5_26[9] , \wRegOut_5_26[8] , 
        \wRegOut_5_26[7] , \wRegOut_5_26[6] , \wRegOut_5_26[5] , 
        \wRegOut_5_26[4] , \wRegOut_5_26[3] , \wRegOut_5_26[2] , 
        \wRegOut_5_26[1] , \wRegOut_5_26[0] }), .L_Out({\wRegInTop_5_26[31] , 
        \wRegInTop_5_26[30] , \wRegInTop_5_26[29] , \wRegInTop_5_26[28] , 
        \wRegInTop_5_26[27] , \wRegInTop_5_26[26] , \wRegInTop_5_26[25] , 
        \wRegInTop_5_26[24] , \wRegInTop_5_26[23] , \wRegInTop_5_26[22] , 
        \wRegInTop_5_26[21] , \wRegInTop_5_26[20] , \wRegInTop_5_26[19] , 
        \wRegInTop_5_26[18] , \wRegInTop_5_26[17] , \wRegInTop_5_26[16] , 
        \wRegInTop_5_26[15] , \wRegInTop_5_26[14] , \wRegInTop_5_26[13] , 
        \wRegInTop_5_26[12] , \wRegInTop_5_26[11] , \wRegInTop_5_26[10] , 
        \wRegInTop_5_26[9] , \wRegInTop_5_26[8] , \wRegInTop_5_26[7] , 
        \wRegInTop_5_26[6] , \wRegInTop_5_26[5] , \wRegInTop_5_26[4] , 
        \wRegInTop_5_26[3] , \wRegInTop_5_26[2] , \wRegInTop_5_26[1] , 
        \wRegInTop_5_26[0] }), .R_WR(\wRegEnTop_5_27[0] ), .R_In({
        \wRegOut_5_27[31] , \wRegOut_5_27[30] , \wRegOut_5_27[29] , 
        \wRegOut_5_27[28] , \wRegOut_5_27[27] , \wRegOut_5_27[26] , 
        \wRegOut_5_27[25] , \wRegOut_5_27[24] , \wRegOut_5_27[23] , 
        \wRegOut_5_27[22] , \wRegOut_5_27[21] , \wRegOut_5_27[20] , 
        \wRegOut_5_27[19] , \wRegOut_5_27[18] , \wRegOut_5_27[17] , 
        \wRegOut_5_27[16] , \wRegOut_5_27[15] , \wRegOut_5_27[14] , 
        \wRegOut_5_27[13] , \wRegOut_5_27[12] , \wRegOut_5_27[11] , 
        \wRegOut_5_27[10] , \wRegOut_5_27[9] , \wRegOut_5_27[8] , 
        \wRegOut_5_27[7] , \wRegOut_5_27[6] , \wRegOut_5_27[5] , 
        \wRegOut_5_27[4] , \wRegOut_5_27[3] , \wRegOut_5_27[2] , 
        \wRegOut_5_27[1] , \wRegOut_5_27[0] }), .R_Out({\wRegInTop_5_27[31] , 
        \wRegInTop_5_27[30] , \wRegInTop_5_27[29] , \wRegInTop_5_27[28] , 
        \wRegInTop_5_27[27] , \wRegInTop_5_27[26] , \wRegInTop_5_27[25] , 
        \wRegInTop_5_27[24] , \wRegInTop_5_27[23] , \wRegInTop_5_27[22] , 
        \wRegInTop_5_27[21] , \wRegInTop_5_27[20] , \wRegInTop_5_27[19] , 
        \wRegInTop_5_27[18] , \wRegInTop_5_27[17] , \wRegInTop_5_27[16] , 
        \wRegInTop_5_27[15] , \wRegInTop_5_27[14] , \wRegInTop_5_27[13] , 
        \wRegInTop_5_27[12] , \wRegInTop_5_27[11] , \wRegInTop_5_27[10] , 
        \wRegInTop_5_27[9] , \wRegInTop_5_27[8] , \wRegInTop_5_27[7] , 
        \wRegInTop_5_27[6] , \wRegInTop_5_27[5] , \wRegInTop_5_27[4] , 
        \wRegInTop_5_27[3] , \wRegInTop_5_27[2] , \wRegInTop_5_27[1] , 
        \wRegInTop_5_27[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_2_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink7[31] , \ScanLink7[30] , \ScanLink7[29] , 
        \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , \ScanLink7[25] , 
        \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , \ScanLink7[21] , 
        \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , \ScanLink7[17] , 
        \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , \ScanLink7[13] , 
        \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , \ScanLink7[9] , 
        \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , \ScanLink7[5] , 
        \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , \ScanLink7[1] , 
        \ScanLink7[0] }), .ScanOut({\ScanLink6[31] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , 
        \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , 
        \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , 
        \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , 
        \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , 
        \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_2_3[31] , \wRegOut_2_3[30] , \wRegOut_2_3[29] , 
        \wRegOut_2_3[28] , \wRegOut_2_3[27] , \wRegOut_2_3[26] , 
        \wRegOut_2_3[25] , \wRegOut_2_3[24] , \wRegOut_2_3[23] , 
        \wRegOut_2_3[22] , \wRegOut_2_3[21] , \wRegOut_2_3[20] , 
        \wRegOut_2_3[19] , \wRegOut_2_3[18] , \wRegOut_2_3[17] , 
        \wRegOut_2_3[16] , \wRegOut_2_3[15] , \wRegOut_2_3[14] , 
        \wRegOut_2_3[13] , \wRegOut_2_3[12] , \wRegOut_2_3[11] , 
        \wRegOut_2_3[10] , \wRegOut_2_3[9] , \wRegOut_2_3[8] , 
        \wRegOut_2_3[7] , \wRegOut_2_3[6] , \wRegOut_2_3[5] , \wRegOut_2_3[4] , 
        \wRegOut_2_3[3] , \wRegOut_2_3[2] , \wRegOut_2_3[1] , \wRegOut_2_3[0] 
        }), .Enable1(\wRegEnTop_2_3[0] ), .Enable2(\wRegEnBot_2_3[0] ), .In1({
        \wRegInTop_2_3[31] , \wRegInTop_2_3[30] , \wRegInTop_2_3[29] , 
        \wRegInTop_2_3[28] , \wRegInTop_2_3[27] , \wRegInTop_2_3[26] , 
        \wRegInTop_2_3[25] , \wRegInTop_2_3[24] , \wRegInTop_2_3[23] , 
        \wRegInTop_2_3[22] , \wRegInTop_2_3[21] , \wRegInTop_2_3[20] , 
        \wRegInTop_2_3[19] , \wRegInTop_2_3[18] , \wRegInTop_2_3[17] , 
        \wRegInTop_2_3[16] , \wRegInTop_2_3[15] , \wRegInTop_2_3[14] , 
        \wRegInTop_2_3[13] , \wRegInTop_2_3[12] , \wRegInTop_2_3[11] , 
        \wRegInTop_2_3[10] , \wRegInTop_2_3[9] , \wRegInTop_2_3[8] , 
        \wRegInTop_2_3[7] , \wRegInTop_2_3[6] , \wRegInTop_2_3[5] , 
        \wRegInTop_2_3[4] , \wRegInTop_2_3[3] , \wRegInTop_2_3[2] , 
        \wRegInTop_2_3[1] , \wRegInTop_2_3[0] }), .In2({\wRegInBot_2_3[31] , 
        \wRegInBot_2_3[30] , \wRegInBot_2_3[29] , \wRegInBot_2_3[28] , 
        \wRegInBot_2_3[27] , \wRegInBot_2_3[26] , \wRegInBot_2_3[25] , 
        \wRegInBot_2_3[24] , \wRegInBot_2_3[23] , \wRegInBot_2_3[22] , 
        \wRegInBot_2_3[21] , \wRegInBot_2_3[20] , \wRegInBot_2_3[19] , 
        \wRegInBot_2_3[18] , \wRegInBot_2_3[17] , \wRegInBot_2_3[16] , 
        \wRegInBot_2_3[15] , \wRegInBot_2_3[14] , \wRegInBot_2_3[13] , 
        \wRegInBot_2_3[12] , \wRegInBot_2_3[11] , \wRegInBot_2_3[10] , 
        \wRegInBot_2_3[9] , \wRegInBot_2_3[8] , \wRegInBot_2_3[7] , 
        \wRegInBot_2_3[6] , \wRegInBot_2_3[5] , \wRegInBot_2_3[4] , 
        \wRegInBot_2_3[3] , \wRegInBot_2_3[2] , \wRegInBot_2_3[1] , 
        \wRegInBot_2_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink16[31] , \ScanLink16[30] , \ScanLink16[29] , 
        \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , \ScanLink16[25] , 
        \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , \ScanLink16[21] , 
        \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , \ScanLink16[17] , 
        \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , \ScanLink16[13] , 
        \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , \ScanLink16[9] , 
        \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , \ScanLink16[5] , 
        \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , \ScanLink16[1] , 
        \ScanLink16[0] }), .ScanOut({\ScanLink15[31] , \ScanLink15[30] , 
        \ScanLink15[29] , \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , 
        \ScanLink15[25] , \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , 
        \ScanLink15[21] , \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , 
        \ScanLink15[17] , \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , 
        \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , 
        \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , 
        \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , 
        \ScanLink15[1] , \ScanLink15[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_0[31] , \wRegOut_4_0[30] , \wRegOut_4_0[29] , 
        \wRegOut_4_0[28] , \wRegOut_4_0[27] , \wRegOut_4_0[26] , 
        \wRegOut_4_0[25] , \wRegOut_4_0[24] , \wRegOut_4_0[23] , 
        \wRegOut_4_0[22] , \wRegOut_4_0[21] , \wRegOut_4_0[20] , 
        \wRegOut_4_0[19] , \wRegOut_4_0[18] , \wRegOut_4_0[17] , 
        \wRegOut_4_0[16] , \wRegOut_4_0[15] , \wRegOut_4_0[14] , 
        \wRegOut_4_0[13] , \wRegOut_4_0[12] , \wRegOut_4_0[11] , 
        \wRegOut_4_0[10] , \wRegOut_4_0[9] , \wRegOut_4_0[8] , 
        \wRegOut_4_0[7] , \wRegOut_4_0[6] , \wRegOut_4_0[5] , \wRegOut_4_0[4] , 
        \wRegOut_4_0[3] , \wRegOut_4_0[2] , \wRegOut_4_0[1] , \wRegOut_4_0[0] 
        }), .Enable1(\wRegEnTop_4_0[0] ), .Enable2(\wRegEnBot_4_0[0] ), .In1({
        \wRegInTop_4_0[31] , \wRegInTop_4_0[30] , \wRegInTop_4_0[29] , 
        \wRegInTop_4_0[28] , \wRegInTop_4_0[27] , \wRegInTop_4_0[26] , 
        \wRegInTop_4_0[25] , \wRegInTop_4_0[24] , \wRegInTop_4_0[23] , 
        \wRegInTop_4_0[22] , \wRegInTop_4_0[21] , \wRegInTop_4_0[20] , 
        \wRegInTop_4_0[19] , \wRegInTop_4_0[18] , \wRegInTop_4_0[17] , 
        \wRegInTop_4_0[16] , \wRegInTop_4_0[15] , \wRegInTop_4_0[14] , 
        \wRegInTop_4_0[13] , \wRegInTop_4_0[12] , \wRegInTop_4_0[11] , 
        \wRegInTop_4_0[10] , \wRegInTop_4_0[9] , \wRegInTop_4_0[8] , 
        \wRegInTop_4_0[7] , \wRegInTop_4_0[6] , \wRegInTop_4_0[5] , 
        \wRegInTop_4_0[4] , \wRegInTop_4_0[3] , \wRegInTop_4_0[2] , 
        \wRegInTop_4_0[1] , \wRegInTop_4_0[0] }), .In2({\wRegInBot_4_0[31] , 
        \wRegInBot_4_0[30] , \wRegInBot_4_0[29] , \wRegInBot_4_0[28] , 
        \wRegInBot_4_0[27] , \wRegInBot_4_0[26] , \wRegInBot_4_0[25] , 
        \wRegInBot_4_0[24] , \wRegInBot_4_0[23] , \wRegInBot_4_0[22] , 
        \wRegInBot_4_0[21] , \wRegInBot_4_0[20] , \wRegInBot_4_0[19] , 
        \wRegInBot_4_0[18] , \wRegInBot_4_0[17] , \wRegInBot_4_0[16] , 
        \wRegInBot_4_0[15] , \wRegInBot_4_0[14] , \wRegInBot_4_0[13] , 
        \wRegInBot_4_0[12] , \wRegInBot_4_0[11] , \wRegInBot_4_0[10] , 
        \wRegInBot_4_0[9] , \wRegInBot_4_0[8] , \wRegInBot_4_0[7] , 
        \wRegInBot_4_0[6] , \wRegInBot_4_0[5] , \wRegInBot_4_0[4] , 
        \wRegInBot_4_0[3] , \wRegInBot_4_0[2] , \wRegInBot_4_0[1] , 
        \wRegInBot_4_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink30[31] , \ScanLink30[30] , \ScanLink30[29] , 
        \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , \ScanLink30[25] , 
        \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , \ScanLink30[21] , 
        \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , \ScanLink30[17] , 
        \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , \ScanLink30[13] , 
        \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , \ScanLink30[9] , 
        \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , \ScanLink30[5] , 
        \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , \ScanLink30[1] , 
        \ScanLink30[0] }), .ScanOut({\ScanLink29[31] , \ScanLink29[30] , 
        \ScanLink29[29] , \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , 
        \ScanLink29[25] , \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , 
        \ScanLink29[21] , \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , 
        \ScanLink29[17] , \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , 
        \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , 
        \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , 
        \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , 
        \ScanLink29[1] , \ScanLink29[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_14[31] , \wRegOut_4_14[30] , 
        \wRegOut_4_14[29] , \wRegOut_4_14[28] , \wRegOut_4_14[27] , 
        \wRegOut_4_14[26] , \wRegOut_4_14[25] , \wRegOut_4_14[24] , 
        \wRegOut_4_14[23] , \wRegOut_4_14[22] , \wRegOut_4_14[21] , 
        \wRegOut_4_14[20] , \wRegOut_4_14[19] , \wRegOut_4_14[18] , 
        \wRegOut_4_14[17] , \wRegOut_4_14[16] , \wRegOut_4_14[15] , 
        \wRegOut_4_14[14] , \wRegOut_4_14[13] , \wRegOut_4_14[12] , 
        \wRegOut_4_14[11] , \wRegOut_4_14[10] , \wRegOut_4_14[9] , 
        \wRegOut_4_14[8] , \wRegOut_4_14[7] , \wRegOut_4_14[6] , 
        \wRegOut_4_14[5] , \wRegOut_4_14[4] , \wRegOut_4_14[3] , 
        \wRegOut_4_14[2] , \wRegOut_4_14[1] , \wRegOut_4_14[0] }), .Enable1(
        \wRegEnTop_4_14[0] ), .Enable2(\wRegEnBot_4_14[0] ), .In1({
        \wRegInTop_4_14[31] , \wRegInTop_4_14[30] , \wRegInTop_4_14[29] , 
        \wRegInTop_4_14[28] , \wRegInTop_4_14[27] , \wRegInTop_4_14[26] , 
        \wRegInTop_4_14[25] , \wRegInTop_4_14[24] , \wRegInTop_4_14[23] , 
        \wRegInTop_4_14[22] , \wRegInTop_4_14[21] , \wRegInTop_4_14[20] , 
        \wRegInTop_4_14[19] , \wRegInTop_4_14[18] , \wRegInTop_4_14[17] , 
        \wRegInTop_4_14[16] , \wRegInTop_4_14[15] , \wRegInTop_4_14[14] , 
        \wRegInTop_4_14[13] , \wRegInTop_4_14[12] , \wRegInTop_4_14[11] , 
        \wRegInTop_4_14[10] , \wRegInTop_4_14[9] , \wRegInTop_4_14[8] , 
        \wRegInTop_4_14[7] , \wRegInTop_4_14[6] , \wRegInTop_4_14[5] , 
        \wRegInTop_4_14[4] , \wRegInTop_4_14[3] , \wRegInTop_4_14[2] , 
        \wRegInTop_4_14[1] , \wRegInTop_4_14[0] }), .In2({\wRegInBot_4_14[31] , 
        \wRegInBot_4_14[30] , \wRegInBot_4_14[29] , \wRegInBot_4_14[28] , 
        \wRegInBot_4_14[27] , \wRegInBot_4_14[26] , \wRegInBot_4_14[25] , 
        \wRegInBot_4_14[24] , \wRegInBot_4_14[23] , \wRegInBot_4_14[22] , 
        \wRegInBot_4_14[21] , \wRegInBot_4_14[20] , \wRegInBot_4_14[19] , 
        \wRegInBot_4_14[18] , \wRegInBot_4_14[17] , \wRegInBot_4_14[16] , 
        \wRegInBot_4_14[15] , \wRegInBot_4_14[14] , \wRegInBot_4_14[13] , 
        \wRegInBot_4_14[12] , \wRegInBot_4_14[11] , \wRegInBot_4_14[10] , 
        \wRegInBot_4_14[9] , \wRegInBot_4_14[8] , \wRegInBot_4_14[7] , 
        \wRegInBot_4_14[6] , \wRegInBot_4_14[5] , \wRegInBot_4_14[4] , 
        \wRegInBot_4_14[3] , \wRegInBot_4_14[2] , \wRegInBot_4_14[1] , 
        \wRegInBot_4_14[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink32[31] , \ScanLink32[30] , \ScanLink32[29] , 
        \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , \ScanLink32[25] , 
        \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , \ScanLink32[21] , 
        \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , \ScanLink32[17] , 
        \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , \ScanLink32[13] , 
        \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , \ScanLink32[9] , 
        \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , \ScanLink32[5] , 
        \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , \ScanLink32[1] , 
        \ScanLink32[0] }), .ScanOut({\ScanLink31[31] , \ScanLink31[30] , 
        \ScanLink31[29] , \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , 
        \ScanLink31[25] , \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , 
        \ScanLink31[21] , \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , 
        \ScanLink31[17] , \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , 
        \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , 
        \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , 
        \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , 
        \ScanLink31[1] , \ScanLink31[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_0[31] , \wRegOut_5_0[30] , \wRegOut_5_0[29] , 
        \wRegOut_5_0[28] , \wRegOut_5_0[27] , \wRegOut_5_0[26] , 
        \wRegOut_5_0[25] , \wRegOut_5_0[24] , \wRegOut_5_0[23] , 
        \wRegOut_5_0[22] , \wRegOut_5_0[21] , \wRegOut_5_0[20] , 
        \wRegOut_5_0[19] , \wRegOut_5_0[18] , \wRegOut_5_0[17] , 
        \wRegOut_5_0[16] , \wRegOut_5_0[15] , \wRegOut_5_0[14] , 
        \wRegOut_5_0[13] , \wRegOut_5_0[12] , \wRegOut_5_0[11] , 
        \wRegOut_5_0[10] , \wRegOut_5_0[9] , \wRegOut_5_0[8] , 
        \wRegOut_5_0[7] , \wRegOut_5_0[6] , \wRegOut_5_0[5] , \wRegOut_5_0[4] , 
        \wRegOut_5_0[3] , \wRegOut_5_0[2] , \wRegOut_5_0[1] , \wRegOut_5_0[0] 
        }), .Enable1(\wRegEnTop_5_0[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_0[31] , \wRegInTop_5_0[30] , \wRegInTop_5_0[29] , 
        \wRegInTop_5_0[28] , \wRegInTop_5_0[27] , \wRegInTop_5_0[26] , 
        \wRegInTop_5_0[25] , \wRegInTop_5_0[24] , \wRegInTop_5_0[23] , 
        \wRegInTop_5_0[22] , \wRegInTop_5_0[21] , \wRegInTop_5_0[20] , 
        \wRegInTop_5_0[19] , \wRegInTop_5_0[18] , \wRegInTop_5_0[17] , 
        \wRegInTop_5_0[16] , \wRegInTop_5_0[15] , \wRegInTop_5_0[14] , 
        \wRegInTop_5_0[13] , \wRegInTop_5_0[12] , \wRegInTop_5_0[11] , 
        \wRegInTop_5_0[10] , \wRegInTop_5_0[9] , \wRegInTop_5_0[8] , 
        \wRegInTop_5_0[7] , \wRegInTop_5_0[6] , \wRegInTop_5_0[5] , 
        \wRegInTop_5_0[4] , \wRegInTop_5_0[3] , \wRegInTop_5_0[2] , 
        \wRegInTop_5_0[1] , \wRegInTop_5_0[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink40[31] , \ScanLink40[30] , \ScanLink40[29] , 
        \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , \ScanLink40[25] , 
        \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , \ScanLink40[21] , 
        \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , \ScanLink40[17] , 
        \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , \ScanLink40[13] , 
        \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , \ScanLink40[9] , 
        \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , \ScanLink40[5] , 
        \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , \ScanLink40[1] , 
        \ScanLink40[0] }), .ScanOut({\ScanLink39[31] , \ScanLink39[30] , 
        \ScanLink39[29] , \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , 
        \ScanLink39[25] , \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , 
        \ScanLink39[21] , \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , 
        \ScanLink39[17] , \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , 
        \ScanLink39[13] , \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , 
        \ScanLink39[9] , \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , 
        \ScanLink39[5] , \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , 
        \ScanLink39[1] , \ScanLink39[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_8[31] , \wRegOut_5_8[30] , \wRegOut_5_8[29] , 
        \wRegOut_5_8[28] , \wRegOut_5_8[27] , \wRegOut_5_8[26] , 
        \wRegOut_5_8[25] , \wRegOut_5_8[24] , \wRegOut_5_8[23] , 
        \wRegOut_5_8[22] , \wRegOut_5_8[21] , \wRegOut_5_8[20] , 
        \wRegOut_5_8[19] , \wRegOut_5_8[18] , \wRegOut_5_8[17] , 
        \wRegOut_5_8[16] , \wRegOut_5_8[15] , \wRegOut_5_8[14] , 
        \wRegOut_5_8[13] , \wRegOut_5_8[12] , \wRegOut_5_8[11] , 
        \wRegOut_5_8[10] , \wRegOut_5_8[9] , \wRegOut_5_8[8] , 
        \wRegOut_5_8[7] , \wRegOut_5_8[6] , \wRegOut_5_8[5] , \wRegOut_5_8[4] , 
        \wRegOut_5_8[3] , \wRegOut_5_8[2] , \wRegOut_5_8[1] , \wRegOut_5_8[0] 
        }), .Enable1(\wRegEnTop_5_8[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_8[31] , \wRegInTop_5_8[30] , \wRegInTop_5_8[29] , 
        \wRegInTop_5_8[28] , \wRegInTop_5_8[27] , \wRegInTop_5_8[26] , 
        \wRegInTop_5_8[25] , \wRegInTop_5_8[24] , \wRegInTop_5_8[23] , 
        \wRegInTop_5_8[22] , \wRegInTop_5_8[21] , \wRegInTop_5_8[20] , 
        \wRegInTop_5_8[19] , \wRegInTop_5_8[18] , \wRegInTop_5_8[17] , 
        \wRegInTop_5_8[16] , \wRegInTop_5_8[15] , \wRegInTop_5_8[14] , 
        \wRegInTop_5_8[13] , \wRegInTop_5_8[12] , \wRegInTop_5_8[11] , 
        \wRegInTop_5_8[10] , \wRegInTop_5_8[9] , \wRegInTop_5_8[8] , 
        \wRegInTop_5_8[7] , \wRegInTop_5_8[6] , \wRegInTop_5_8[5] , 
        \wRegInTop_5_8[4] , \wRegInTop_5_8[3] , \wRegInTop_5_8[2] , 
        \wRegInTop_5_8[1] , \wRegInTop_5_8[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_21 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink53[31] , \ScanLink53[30] , \ScanLink53[29] , 
        \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , \ScanLink53[25] , 
        \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , \ScanLink53[21] , 
        \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , \ScanLink53[17] , 
        \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , \ScanLink53[13] , 
        \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , \ScanLink53[9] , 
        \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , \ScanLink53[5] , 
        \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , \ScanLink53[1] , 
        \ScanLink53[0] }), .ScanOut({\ScanLink52[31] , \ScanLink52[30] , 
        \ScanLink52[29] , \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , 
        \ScanLink52[25] , \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , 
        \ScanLink52[21] , \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , 
        \ScanLink52[17] , \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , 
        \ScanLink52[13] , \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , 
        \ScanLink52[9] , \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , 
        \ScanLink52[5] , \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , 
        \ScanLink52[1] , \ScanLink52[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_21[31] , \wRegOut_5_21[30] , 
        \wRegOut_5_21[29] , \wRegOut_5_21[28] , \wRegOut_5_21[27] , 
        \wRegOut_5_21[26] , \wRegOut_5_21[25] , \wRegOut_5_21[24] , 
        \wRegOut_5_21[23] , \wRegOut_5_21[22] , \wRegOut_5_21[21] , 
        \wRegOut_5_21[20] , \wRegOut_5_21[19] , \wRegOut_5_21[18] , 
        \wRegOut_5_21[17] , \wRegOut_5_21[16] , \wRegOut_5_21[15] , 
        \wRegOut_5_21[14] , \wRegOut_5_21[13] , \wRegOut_5_21[12] , 
        \wRegOut_5_21[11] , \wRegOut_5_21[10] , \wRegOut_5_21[9] , 
        \wRegOut_5_21[8] , \wRegOut_5_21[7] , \wRegOut_5_21[6] , 
        \wRegOut_5_21[5] , \wRegOut_5_21[4] , \wRegOut_5_21[3] , 
        \wRegOut_5_21[2] , \wRegOut_5_21[1] , \wRegOut_5_21[0] }), .Enable1(
        \wRegEnTop_5_21[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_21[31] , 
        \wRegInTop_5_21[30] , \wRegInTop_5_21[29] , \wRegInTop_5_21[28] , 
        \wRegInTop_5_21[27] , \wRegInTop_5_21[26] , \wRegInTop_5_21[25] , 
        \wRegInTop_5_21[24] , \wRegInTop_5_21[23] , \wRegInTop_5_21[22] , 
        \wRegInTop_5_21[21] , \wRegInTop_5_21[20] , \wRegInTop_5_21[19] , 
        \wRegInTop_5_21[18] , \wRegInTop_5_21[17] , \wRegInTop_5_21[16] , 
        \wRegInTop_5_21[15] , \wRegInTop_5_21[14] , \wRegInTop_5_21[13] , 
        \wRegInTop_5_21[12] , \wRegInTop_5_21[11] , \wRegInTop_5_21[10] , 
        \wRegInTop_5_21[9] , \wRegInTop_5_21[8] , \wRegInTop_5_21[7] , 
        \wRegInTop_5_21[6] , \wRegInTop_5_21[5] , \wRegInTop_5_21[4] , 
        \wRegInTop_5_21[3] , \wRegInTop_5_21[2] , \wRegInTop_5_21[1] , 
        \wRegInTop_5_21[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_29 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink61[31] , \ScanLink61[30] , \ScanLink61[29] , 
        \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , \ScanLink61[25] , 
        \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , \ScanLink61[21] , 
        \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , \ScanLink61[17] , 
        \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , \ScanLink61[13] , 
        \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , \ScanLink61[9] , 
        \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , \ScanLink61[5] , 
        \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , \ScanLink61[1] , 
        \ScanLink61[0] }), .ScanOut({\ScanLink60[31] , \ScanLink60[30] , 
        \ScanLink60[29] , \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , 
        \ScanLink60[25] , \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , 
        \ScanLink60[21] , \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , 
        \ScanLink60[17] , \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , 
        \ScanLink60[13] , \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , 
        \ScanLink60[9] , \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , 
        \ScanLink60[5] , \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , 
        \ScanLink60[1] , \ScanLink60[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_29[31] , \wRegOut_5_29[30] , 
        \wRegOut_5_29[29] , \wRegOut_5_29[28] , \wRegOut_5_29[27] , 
        \wRegOut_5_29[26] , \wRegOut_5_29[25] , \wRegOut_5_29[24] , 
        \wRegOut_5_29[23] , \wRegOut_5_29[22] , \wRegOut_5_29[21] , 
        \wRegOut_5_29[20] , \wRegOut_5_29[19] , \wRegOut_5_29[18] , 
        \wRegOut_5_29[17] , \wRegOut_5_29[16] , \wRegOut_5_29[15] , 
        \wRegOut_5_29[14] , \wRegOut_5_29[13] , \wRegOut_5_29[12] , 
        \wRegOut_5_29[11] , \wRegOut_5_29[10] , \wRegOut_5_29[9] , 
        \wRegOut_5_29[8] , \wRegOut_5_29[7] , \wRegOut_5_29[6] , 
        \wRegOut_5_29[5] , \wRegOut_5_29[4] , \wRegOut_5_29[3] , 
        \wRegOut_5_29[2] , \wRegOut_5_29[1] , \wRegOut_5_29[0] }), .Enable1(
        \wRegEnTop_5_29[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_29[31] , 
        \wRegInTop_5_29[30] , \wRegInTop_5_29[29] , \wRegInTop_5_29[28] , 
        \wRegInTop_5_29[27] , \wRegInTop_5_29[26] , \wRegInTop_5_29[25] , 
        \wRegInTop_5_29[24] , \wRegInTop_5_29[23] , \wRegInTop_5_29[22] , 
        \wRegInTop_5_29[21] , \wRegInTop_5_29[20] , \wRegInTop_5_29[19] , 
        \wRegInTop_5_29[18] , \wRegInTop_5_29[17] , \wRegInTop_5_29[16] , 
        \wRegInTop_5_29[15] , \wRegInTop_5_29[14] , \wRegInTop_5_29[13] , 
        \wRegInTop_5_29[12] , \wRegInTop_5_29[11] , \wRegInTop_5_29[10] , 
        \wRegInTop_5_29[9] , \wRegInTop_5_29[8] , \wRegInTop_5_29[7] , 
        \wRegInTop_5_29[6] , \wRegInTop_5_29[5] , \wRegInTop_5_29[4] , 
        \wRegInTop_5_29[3] , \wRegInTop_5_29[2] , \wRegInTop_5_29[1] , 
        \wRegInTop_5_29[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink47[31] , \ScanLink47[30] , \ScanLink47[29] , 
        \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , \ScanLink47[25] , 
        \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , \ScanLink47[21] , 
        \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , \ScanLink47[17] , 
        \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , \ScanLink47[13] , 
        \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , \ScanLink47[9] , 
        \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , \ScanLink47[5] , 
        \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , \ScanLink47[1] , 
        \ScanLink47[0] }), .ScanOut({\ScanLink46[31] , \ScanLink46[30] , 
        \ScanLink46[29] , \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , 
        \ScanLink46[25] , \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , 
        \ScanLink46[21] , \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , 
        \ScanLink46[17] , \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , 
        \ScanLink46[13] , \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , 
        \ScanLink46[9] , \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , 
        \ScanLink46[5] , \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , 
        \ScanLink46[1] , \ScanLink46[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_15[31] , \wRegOut_5_15[30] , 
        \wRegOut_5_15[29] , \wRegOut_5_15[28] , \wRegOut_5_15[27] , 
        \wRegOut_5_15[26] , \wRegOut_5_15[25] , \wRegOut_5_15[24] , 
        \wRegOut_5_15[23] , \wRegOut_5_15[22] , \wRegOut_5_15[21] , 
        \wRegOut_5_15[20] , \wRegOut_5_15[19] , \wRegOut_5_15[18] , 
        \wRegOut_5_15[17] , \wRegOut_5_15[16] , \wRegOut_5_15[15] , 
        \wRegOut_5_15[14] , \wRegOut_5_15[13] , \wRegOut_5_15[12] , 
        \wRegOut_5_15[11] , \wRegOut_5_15[10] , \wRegOut_5_15[9] , 
        \wRegOut_5_15[8] , \wRegOut_5_15[7] , \wRegOut_5_15[6] , 
        \wRegOut_5_15[5] , \wRegOut_5_15[4] , \wRegOut_5_15[3] , 
        \wRegOut_5_15[2] , \wRegOut_5_15[1] , \wRegOut_5_15[0] }), .Enable1(
        \wRegEnTop_5_15[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_15[31] , 
        \wRegInTop_5_15[30] , \wRegInTop_5_15[29] , \wRegInTop_5_15[28] , 
        \wRegInTop_5_15[27] , \wRegInTop_5_15[26] , \wRegInTop_5_15[25] , 
        \wRegInTop_5_15[24] , \wRegInTop_5_15[23] , \wRegInTop_5_15[22] , 
        \wRegInTop_5_15[21] , \wRegInTop_5_15[20] , \wRegInTop_5_15[19] , 
        \wRegInTop_5_15[18] , \wRegInTop_5_15[17] , \wRegInTop_5_15[16] , 
        \wRegInTop_5_15[15] , \wRegInTop_5_15[14] , \wRegInTop_5_15[13] , 
        \wRegInTop_5_15[12] , \wRegInTop_5_15[11] , \wRegInTop_5_15[10] , 
        \wRegInTop_5_15[9] , \wRegInTop_5_15[8] , \wRegInTop_5_15[7] , 
        \wRegInTop_5_15[6] , \wRegInTop_5_15[5] , \wRegInTop_5_15[4] , 
        \wRegInTop_5_15[3] , \wRegInTop_5_15[2] , \wRegInTop_5_15[1] , 
        \wRegInTop_5_15[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_2[0] ), .P_In({\wRegOut_4_2[31] , 
        \wRegOut_4_2[30] , \wRegOut_4_2[29] , \wRegOut_4_2[28] , 
        \wRegOut_4_2[27] , \wRegOut_4_2[26] , \wRegOut_4_2[25] , 
        \wRegOut_4_2[24] , \wRegOut_4_2[23] , \wRegOut_4_2[22] , 
        \wRegOut_4_2[21] , \wRegOut_4_2[20] , \wRegOut_4_2[19] , 
        \wRegOut_4_2[18] , \wRegOut_4_2[17] , \wRegOut_4_2[16] , 
        \wRegOut_4_2[15] , \wRegOut_4_2[14] , \wRegOut_4_2[13] , 
        \wRegOut_4_2[12] , \wRegOut_4_2[11] , \wRegOut_4_2[10] , 
        \wRegOut_4_2[9] , \wRegOut_4_2[8] , \wRegOut_4_2[7] , \wRegOut_4_2[6] , 
        \wRegOut_4_2[5] , \wRegOut_4_2[4] , \wRegOut_4_2[3] , \wRegOut_4_2[2] , 
        \wRegOut_4_2[1] , \wRegOut_4_2[0] }), .P_Out({\wRegInBot_4_2[31] , 
        \wRegInBot_4_2[30] , \wRegInBot_4_2[29] , \wRegInBot_4_2[28] , 
        \wRegInBot_4_2[27] , \wRegInBot_4_2[26] , \wRegInBot_4_2[25] , 
        \wRegInBot_4_2[24] , \wRegInBot_4_2[23] , \wRegInBot_4_2[22] , 
        \wRegInBot_4_2[21] , \wRegInBot_4_2[20] , \wRegInBot_4_2[19] , 
        \wRegInBot_4_2[18] , \wRegInBot_4_2[17] , \wRegInBot_4_2[16] , 
        \wRegInBot_4_2[15] , \wRegInBot_4_2[14] , \wRegInBot_4_2[13] , 
        \wRegInBot_4_2[12] , \wRegInBot_4_2[11] , \wRegInBot_4_2[10] , 
        \wRegInBot_4_2[9] , \wRegInBot_4_2[8] , \wRegInBot_4_2[7] , 
        \wRegInBot_4_2[6] , \wRegInBot_4_2[5] , \wRegInBot_4_2[4] , 
        \wRegInBot_4_2[3] , \wRegInBot_4_2[2] , \wRegInBot_4_2[1] , 
        \wRegInBot_4_2[0] }), .L_WR(\wRegEnTop_5_4[0] ), .L_In({
        \wRegOut_5_4[31] , \wRegOut_5_4[30] , \wRegOut_5_4[29] , 
        \wRegOut_5_4[28] , \wRegOut_5_4[27] , \wRegOut_5_4[26] , 
        \wRegOut_5_4[25] , \wRegOut_5_4[24] , \wRegOut_5_4[23] , 
        \wRegOut_5_4[22] , \wRegOut_5_4[21] , \wRegOut_5_4[20] , 
        \wRegOut_5_4[19] , \wRegOut_5_4[18] , \wRegOut_5_4[17] , 
        \wRegOut_5_4[16] , \wRegOut_5_4[15] , \wRegOut_5_4[14] , 
        \wRegOut_5_4[13] , \wRegOut_5_4[12] , \wRegOut_5_4[11] , 
        \wRegOut_5_4[10] , \wRegOut_5_4[9] , \wRegOut_5_4[8] , 
        \wRegOut_5_4[7] , \wRegOut_5_4[6] , \wRegOut_5_4[5] , \wRegOut_5_4[4] , 
        \wRegOut_5_4[3] , \wRegOut_5_4[2] , \wRegOut_5_4[1] , \wRegOut_5_4[0] 
        }), .L_Out({\wRegInTop_5_4[31] , \wRegInTop_5_4[30] , 
        \wRegInTop_5_4[29] , \wRegInTop_5_4[28] , \wRegInTop_5_4[27] , 
        \wRegInTop_5_4[26] , \wRegInTop_5_4[25] , \wRegInTop_5_4[24] , 
        \wRegInTop_5_4[23] , \wRegInTop_5_4[22] , \wRegInTop_5_4[21] , 
        \wRegInTop_5_4[20] , \wRegInTop_5_4[19] , \wRegInTop_5_4[18] , 
        \wRegInTop_5_4[17] , \wRegInTop_5_4[16] , \wRegInTop_5_4[15] , 
        \wRegInTop_5_4[14] , \wRegInTop_5_4[13] , \wRegInTop_5_4[12] , 
        \wRegInTop_5_4[11] , \wRegInTop_5_4[10] , \wRegInTop_5_4[9] , 
        \wRegInTop_5_4[8] , \wRegInTop_5_4[7] , \wRegInTop_5_4[6] , 
        \wRegInTop_5_4[5] , \wRegInTop_5_4[4] , \wRegInTop_5_4[3] , 
        \wRegInTop_5_4[2] , \wRegInTop_5_4[1] , \wRegInTop_5_4[0] }), .R_WR(
        \wRegEnTop_5_5[0] ), .R_In({\wRegOut_5_5[31] , \wRegOut_5_5[30] , 
        \wRegOut_5_5[29] , \wRegOut_5_5[28] , \wRegOut_5_5[27] , 
        \wRegOut_5_5[26] , \wRegOut_5_5[25] , \wRegOut_5_5[24] , 
        \wRegOut_5_5[23] , \wRegOut_5_5[22] , \wRegOut_5_5[21] , 
        \wRegOut_5_5[20] , \wRegOut_5_5[19] , \wRegOut_5_5[18] , 
        \wRegOut_5_5[17] , \wRegOut_5_5[16] , \wRegOut_5_5[15] , 
        \wRegOut_5_5[14] , \wRegOut_5_5[13] , \wRegOut_5_5[12] , 
        \wRegOut_5_5[11] , \wRegOut_5_5[10] , \wRegOut_5_5[9] , 
        \wRegOut_5_5[8] , \wRegOut_5_5[7] , \wRegOut_5_5[6] , \wRegOut_5_5[5] , 
        \wRegOut_5_5[4] , \wRegOut_5_5[3] , \wRegOut_5_5[2] , \wRegOut_5_5[1] , 
        \wRegOut_5_5[0] }), .R_Out({\wRegInTop_5_5[31] , \wRegInTop_5_5[30] , 
        \wRegInTop_5_5[29] , \wRegInTop_5_5[28] , \wRegInTop_5_5[27] , 
        \wRegInTop_5_5[26] , \wRegInTop_5_5[25] , \wRegInTop_5_5[24] , 
        \wRegInTop_5_5[23] , \wRegInTop_5_5[22] , \wRegInTop_5_5[21] , 
        \wRegInTop_5_5[20] , \wRegInTop_5_5[19] , \wRegInTop_5_5[18] , 
        \wRegInTop_5_5[17] , \wRegInTop_5_5[16] , \wRegInTop_5_5[15] , 
        \wRegInTop_5_5[14] , \wRegInTop_5_5[13] , \wRegInTop_5_5[12] , 
        \wRegInTop_5_5[11] , \wRegInTop_5_5[10] , \wRegInTop_5_5[9] , 
        \wRegInTop_5_5[8] , \wRegInTop_5_5[7] , \wRegInTop_5_5[6] , 
        \wRegInTop_5_5[5] , \wRegInTop_5_5[4] , \wRegInTop_5_5[3] , 
        \wRegInTop_5_5[2] , \wRegInTop_5_5[1] , \wRegInTop_5_5[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink11[31] , \ScanLink11[30] , \ScanLink11[29] , 
        \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , \ScanLink11[25] , 
        \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , \ScanLink11[21] , 
        \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , \ScanLink11[17] , 
        \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , \ScanLink11[13] , 
        \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , \ScanLink11[9] , 
        \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , \ScanLink11[5] , 
        \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , \ScanLink11[1] , 
        \ScanLink11[0] }), .ScanOut({\ScanLink10[31] , \ScanLink10[30] , 
        \ScanLink10[29] , \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , 
        \ScanLink10[25] , \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , 
        \ScanLink10[21] , \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , 
        \ScanLink10[17] , \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , 
        \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , 
        \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , 
        \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , 
        \ScanLink10[1] , \ScanLink10[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_3[31] , \wRegOut_3_3[30] , \wRegOut_3_3[29] , 
        \wRegOut_3_3[28] , \wRegOut_3_3[27] , \wRegOut_3_3[26] , 
        \wRegOut_3_3[25] , \wRegOut_3_3[24] , \wRegOut_3_3[23] , 
        \wRegOut_3_3[22] , \wRegOut_3_3[21] , \wRegOut_3_3[20] , 
        \wRegOut_3_3[19] , \wRegOut_3_3[18] , \wRegOut_3_3[17] , 
        \wRegOut_3_3[16] , \wRegOut_3_3[15] , \wRegOut_3_3[14] , 
        \wRegOut_3_3[13] , \wRegOut_3_3[12] , \wRegOut_3_3[11] , 
        \wRegOut_3_3[10] , \wRegOut_3_3[9] , \wRegOut_3_3[8] , 
        \wRegOut_3_3[7] , \wRegOut_3_3[6] , \wRegOut_3_3[5] , \wRegOut_3_3[4] , 
        \wRegOut_3_3[3] , \wRegOut_3_3[2] , \wRegOut_3_3[1] , \wRegOut_3_3[0] 
        }), .Enable1(\wRegEnTop_3_3[0] ), .Enable2(\wRegEnBot_3_3[0] ), .In1({
        \wRegInTop_3_3[31] , \wRegInTop_3_3[30] , \wRegInTop_3_3[29] , 
        \wRegInTop_3_3[28] , \wRegInTop_3_3[27] , \wRegInTop_3_3[26] , 
        \wRegInTop_3_3[25] , \wRegInTop_3_3[24] , \wRegInTop_3_3[23] , 
        \wRegInTop_3_3[22] , \wRegInTop_3_3[21] , \wRegInTop_3_3[20] , 
        \wRegInTop_3_3[19] , \wRegInTop_3_3[18] , \wRegInTop_3_3[17] , 
        \wRegInTop_3_3[16] , \wRegInTop_3_3[15] , \wRegInTop_3_3[14] , 
        \wRegInTop_3_3[13] , \wRegInTop_3_3[12] , \wRegInTop_3_3[11] , 
        \wRegInTop_3_3[10] , \wRegInTop_3_3[9] , \wRegInTop_3_3[8] , 
        \wRegInTop_3_3[7] , \wRegInTop_3_3[6] , \wRegInTop_3_3[5] , 
        \wRegInTop_3_3[4] , \wRegInTop_3_3[3] , \wRegInTop_3_3[2] , 
        \wRegInTop_3_3[1] , \wRegInTop_3_3[0] }), .In2({\wRegInBot_3_3[31] , 
        \wRegInBot_3_3[30] , \wRegInBot_3_3[29] , \wRegInBot_3_3[28] , 
        \wRegInBot_3_3[27] , \wRegInBot_3_3[26] , \wRegInBot_3_3[25] , 
        \wRegInBot_3_3[24] , \wRegInBot_3_3[23] , \wRegInBot_3_3[22] , 
        \wRegInBot_3_3[21] , \wRegInBot_3_3[20] , \wRegInBot_3_3[19] , 
        \wRegInBot_3_3[18] , \wRegInBot_3_3[17] , \wRegInBot_3_3[16] , 
        \wRegInBot_3_3[15] , \wRegInBot_3_3[14] , \wRegInBot_3_3[13] , 
        \wRegInBot_3_3[12] , \wRegInBot_3_3[11] , \wRegInBot_3_3[10] , 
        \wRegInBot_3_3[9] , \wRegInBot_3_3[8] , \wRegInBot_3_3[7] , 
        \wRegInBot_3_3[6] , \wRegInBot_3_3[5] , \wRegInBot_3_3[4] , 
        \wRegInBot_3_3[3] , \wRegInBot_3_3[2] , \wRegInBot_3_3[1] , 
        \wRegInBot_3_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink41[31] , \ScanLink41[30] , \ScanLink41[29] , 
        \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , \ScanLink41[25] , 
        \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , \ScanLink41[21] , 
        \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , \ScanLink41[17] , 
        \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , \ScanLink41[13] , 
        \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , \ScanLink41[9] , 
        \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , \ScanLink41[5] , 
        \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , \ScanLink41[1] , 
        \ScanLink41[0] }), .ScanOut({\ScanLink40[31] , \ScanLink40[30] , 
        \ScanLink40[29] , \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , 
        \ScanLink40[25] , \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , 
        \ScanLink40[21] , \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , 
        \ScanLink40[17] , \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , 
        \ScanLink40[13] , \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , 
        \ScanLink40[9] , \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , 
        \ScanLink40[5] , \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , 
        \ScanLink40[1] , \ScanLink40[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_9[31] , \wRegOut_5_9[30] , \wRegOut_5_9[29] , 
        \wRegOut_5_9[28] , \wRegOut_5_9[27] , \wRegOut_5_9[26] , 
        \wRegOut_5_9[25] , \wRegOut_5_9[24] , \wRegOut_5_9[23] , 
        \wRegOut_5_9[22] , \wRegOut_5_9[21] , \wRegOut_5_9[20] , 
        \wRegOut_5_9[19] , \wRegOut_5_9[18] , \wRegOut_5_9[17] , 
        \wRegOut_5_9[16] , \wRegOut_5_9[15] , \wRegOut_5_9[14] , 
        \wRegOut_5_9[13] , \wRegOut_5_9[12] , \wRegOut_5_9[11] , 
        \wRegOut_5_9[10] , \wRegOut_5_9[9] , \wRegOut_5_9[8] , 
        \wRegOut_5_9[7] , \wRegOut_5_9[6] , \wRegOut_5_9[5] , \wRegOut_5_9[4] , 
        \wRegOut_5_9[3] , \wRegOut_5_9[2] , \wRegOut_5_9[1] , \wRegOut_5_9[0] 
        }), .Enable1(\wRegEnTop_5_9[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_9[31] , \wRegInTop_5_9[30] , \wRegInTop_5_9[29] , 
        \wRegInTop_5_9[28] , \wRegInTop_5_9[27] , \wRegInTop_5_9[26] , 
        \wRegInTop_5_9[25] , \wRegInTop_5_9[24] , \wRegInTop_5_9[23] , 
        \wRegInTop_5_9[22] , \wRegInTop_5_9[21] , \wRegInTop_5_9[20] , 
        \wRegInTop_5_9[19] , \wRegInTop_5_9[18] , \wRegInTop_5_9[17] , 
        \wRegInTop_5_9[16] , \wRegInTop_5_9[15] , \wRegInTop_5_9[14] , 
        \wRegInTop_5_9[13] , \wRegInTop_5_9[12] , \wRegInTop_5_9[11] , 
        \wRegInTop_5_9[10] , \wRegInTop_5_9[9] , \wRegInTop_5_9[8] , 
        \wRegInTop_5_9[7] , \wRegInTop_5_9[6] , \wRegInTop_5_9[5] , 
        \wRegInTop_5_9[4] , \wRegInTop_5_9[3] , \wRegInTop_5_9[2] , 
        \wRegInTop_5_9[1] , \wRegInTop_5_9[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_20 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink52[31] , \ScanLink52[30] , \ScanLink52[29] , 
        \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , \ScanLink52[25] , 
        \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , \ScanLink52[21] , 
        \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , \ScanLink52[17] , 
        \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , \ScanLink52[13] , 
        \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , \ScanLink52[9] , 
        \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , \ScanLink52[5] , 
        \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , \ScanLink52[1] , 
        \ScanLink52[0] }), .ScanOut({\ScanLink51[31] , \ScanLink51[30] , 
        \ScanLink51[29] , \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , 
        \ScanLink51[25] , \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , 
        \ScanLink51[21] , \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , 
        \ScanLink51[17] , \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , 
        \ScanLink51[13] , \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , 
        \ScanLink51[9] , \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , 
        \ScanLink51[5] , \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , 
        \ScanLink51[1] , \ScanLink51[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_20[31] , \wRegOut_5_20[30] , 
        \wRegOut_5_20[29] , \wRegOut_5_20[28] , \wRegOut_5_20[27] , 
        \wRegOut_5_20[26] , \wRegOut_5_20[25] , \wRegOut_5_20[24] , 
        \wRegOut_5_20[23] , \wRegOut_5_20[22] , \wRegOut_5_20[21] , 
        \wRegOut_5_20[20] , \wRegOut_5_20[19] , \wRegOut_5_20[18] , 
        \wRegOut_5_20[17] , \wRegOut_5_20[16] , \wRegOut_5_20[15] , 
        \wRegOut_5_20[14] , \wRegOut_5_20[13] , \wRegOut_5_20[12] , 
        \wRegOut_5_20[11] , \wRegOut_5_20[10] , \wRegOut_5_20[9] , 
        \wRegOut_5_20[8] , \wRegOut_5_20[7] , \wRegOut_5_20[6] , 
        \wRegOut_5_20[5] , \wRegOut_5_20[4] , \wRegOut_5_20[3] , 
        \wRegOut_5_20[2] , \wRegOut_5_20[1] , \wRegOut_5_20[0] }), .Enable1(
        \wRegEnTop_5_20[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_20[31] , 
        \wRegInTop_5_20[30] , \wRegInTop_5_20[29] , \wRegInTop_5_20[28] , 
        \wRegInTop_5_20[27] , \wRegInTop_5_20[26] , \wRegInTop_5_20[25] , 
        \wRegInTop_5_20[24] , \wRegInTop_5_20[23] , \wRegInTop_5_20[22] , 
        \wRegInTop_5_20[21] , \wRegInTop_5_20[20] , \wRegInTop_5_20[19] , 
        \wRegInTop_5_20[18] , \wRegInTop_5_20[17] , \wRegInTop_5_20[16] , 
        \wRegInTop_5_20[15] , \wRegInTop_5_20[14] , \wRegInTop_5_20[13] , 
        \wRegInTop_5_20[12] , \wRegInTop_5_20[11] , \wRegInTop_5_20[10] , 
        \wRegInTop_5_20[9] , \wRegInTop_5_20[8] , \wRegInTop_5_20[7] , 
        \wRegInTop_5_20[6] , \wRegInTop_5_20[5] , \wRegInTop_5_20[4] , 
        \wRegInTop_5_20[3] , \wRegInTop_5_20[2] , \wRegInTop_5_20[1] , 
        \wRegInTop_5_20[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_2_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_2[0] ), .P_WR(\wRegEnBot_2_1[0] ), .P_In({\wRegOut_2_1[31] , 
        \wRegOut_2_1[30] , \wRegOut_2_1[29] , \wRegOut_2_1[28] , 
        \wRegOut_2_1[27] , \wRegOut_2_1[26] , \wRegOut_2_1[25] , 
        \wRegOut_2_1[24] , \wRegOut_2_1[23] , \wRegOut_2_1[22] , 
        \wRegOut_2_1[21] , \wRegOut_2_1[20] , \wRegOut_2_1[19] , 
        \wRegOut_2_1[18] , \wRegOut_2_1[17] , \wRegOut_2_1[16] , 
        \wRegOut_2_1[15] , \wRegOut_2_1[14] , \wRegOut_2_1[13] , 
        \wRegOut_2_1[12] , \wRegOut_2_1[11] , \wRegOut_2_1[10] , 
        \wRegOut_2_1[9] , \wRegOut_2_1[8] , \wRegOut_2_1[7] , \wRegOut_2_1[6] , 
        \wRegOut_2_1[5] , \wRegOut_2_1[4] , \wRegOut_2_1[3] , \wRegOut_2_1[2] , 
        \wRegOut_2_1[1] , \wRegOut_2_1[0] }), .P_Out({\wRegInBot_2_1[31] , 
        \wRegInBot_2_1[30] , \wRegInBot_2_1[29] , \wRegInBot_2_1[28] , 
        \wRegInBot_2_1[27] , \wRegInBot_2_1[26] , \wRegInBot_2_1[25] , 
        \wRegInBot_2_1[24] , \wRegInBot_2_1[23] , \wRegInBot_2_1[22] , 
        \wRegInBot_2_1[21] , \wRegInBot_2_1[20] , \wRegInBot_2_1[19] , 
        \wRegInBot_2_1[18] , \wRegInBot_2_1[17] , \wRegInBot_2_1[16] , 
        \wRegInBot_2_1[15] , \wRegInBot_2_1[14] , \wRegInBot_2_1[13] , 
        \wRegInBot_2_1[12] , \wRegInBot_2_1[11] , \wRegInBot_2_1[10] , 
        \wRegInBot_2_1[9] , \wRegInBot_2_1[8] , \wRegInBot_2_1[7] , 
        \wRegInBot_2_1[6] , \wRegInBot_2_1[5] , \wRegInBot_2_1[4] , 
        \wRegInBot_2_1[3] , \wRegInBot_2_1[2] , \wRegInBot_2_1[1] , 
        \wRegInBot_2_1[0] }), .L_WR(\wRegEnTop_3_2[0] ), .L_In({
        \wRegOut_3_2[31] , \wRegOut_3_2[30] , \wRegOut_3_2[29] , 
        \wRegOut_3_2[28] , \wRegOut_3_2[27] , \wRegOut_3_2[26] , 
        \wRegOut_3_2[25] , \wRegOut_3_2[24] , \wRegOut_3_2[23] , 
        \wRegOut_3_2[22] , \wRegOut_3_2[21] , \wRegOut_3_2[20] , 
        \wRegOut_3_2[19] , \wRegOut_3_2[18] , \wRegOut_3_2[17] , 
        \wRegOut_3_2[16] , \wRegOut_3_2[15] , \wRegOut_3_2[14] , 
        \wRegOut_3_2[13] , \wRegOut_3_2[12] , \wRegOut_3_2[11] , 
        \wRegOut_3_2[10] , \wRegOut_3_2[9] , \wRegOut_3_2[8] , 
        \wRegOut_3_2[7] , \wRegOut_3_2[6] , \wRegOut_3_2[5] , \wRegOut_3_2[4] , 
        \wRegOut_3_2[3] , \wRegOut_3_2[2] , \wRegOut_3_2[1] , \wRegOut_3_2[0] 
        }), .L_Out({\wRegInTop_3_2[31] , \wRegInTop_3_2[30] , 
        \wRegInTop_3_2[29] , \wRegInTop_3_2[28] , \wRegInTop_3_2[27] , 
        \wRegInTop_3_2[26] , \wRegInTop_3_2[25] , \wRegInTop_3_2[24] , 
        \wRegInTop_3_2[23] , \wRegInTop_3_2[22] , \wRegInTop_3_2[21] , 
        \wRegInTop_3_2[20] , \wRegInTop_3_2[19] , \wRegInTop_3_2[18] , 
        \wRegInTop_3_2[17] , \wRegInTop_3_2[16] , \wRegInTop_3_2[15] , 
        \wRegInTop_3_2[14] , \wRegInTop_3_2[13] , \wRegInTop_3_2[12] , 
        \wRegInTop_3_2[11] , \wRegInTop_3_2[10] , \wRegInTop_3_2[9] , 
        \wRegInTop_3_2[8] , \wRegInTop_3_2[7] , \wRegInTop_3_2[6] , 
        \wRegInTop_3_2[5] , \wRegInTop_3_2[4] , \wRegInTop_3_2[3] , 
        \wRegInTop_3_2[2] , \wRegInTop_3_2[1] , \wRegInTop_3_2[0] }), .R_WR(
        \wRegEnTop_3_3[0] ), .R_In({\wRegOut_3_3[31] , \wRegOut_3_3[30] , 
        \wRegOut_3_3[29] , \wRegOut_3_3[28] , \wRegOut_3_3[27] , 
        \wRegOut_3_3[26] , \wRegOut_3_3[25] , \wRegOut_3_3[24] , 
        \wRegOut_3_3[23] , \wRegOut_3_3[22] , \wRegOut_3_3[21] , 
        \wRegOut_3_3[20] , \wRegOut_3_3[19] , \wRegOut_3_3[18] , 
        \wRegOut_3_3[17] , \wRegOut_3_3[16] , \wRegOut_3_3[15] , 
        \wRegOut_3_3[14] , \wRegOut_3_3[13] , \wRegOut_3_3[12] , 
        \wRegOut_3_3[11] , \wRegOut_3_3[10] , \wRegOut_3_3[9] , 
        \wRegOut_3_3[8] , \wRegOut_3_3[7] , \wRegOut_3_3[6] , \wRegOut_3_3[5] , 
        \wRegOut_3_3[4] , \wRegOut_3_3[3] , \wRegOut_3_3[2] , \wRegOut_3_3[1] , 
        \wRegOut_3_3[0] }), .R_Out({\wRegInTop_3_3[31] , \wRegInTop_3_3[30] , 
        \wRegInTop_3_3[29] , \wRegInTop_3_3[28] , \wRegInTop_3_3[27] , 
        \wRegInTop_3_3[26] , \wRegInTop_3_3[25] , \wRegInTop_3_3[24] , 
        \wRegInTop_3_3[23] , \wRegInTop_3_3[22] , \wRegInTop_3_3[21] , 
        \wRegInTop_3_3[20] , \wRegInTop_3_3[19] , \wRegInTop_3_3[18] , 
        \wRegInTop_3_3[17] , \wRegInTop_3_3[16] , \wRegInTop_3_3[15] , 
        \wRegInTop_3_3[14] , \wRegInTop_3_3[13] , \wRegInTop_3_3[12] , 
        \wRegInTop_3_3[11] , \wRegInTop_3_3[10] , \wRegInTop_3_3[9] , 
        \wRegInTop_3_3[8] , \wRegInTop_3_3[7] , \wRegInTop_3_3[6] , 
        \wRegInTop_3_3[5] , \wRegInTop_3_3[4] , \wRegInTop_3_3[3] , 
        \wRegInTop_3_3[2] , \wRegInTop_3_3[1] , \wRegInTop_3_3[0] }) );
    BHeap_Node_WIDTH32 BHN_3_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_1[0] ), .P_In({\wRegOut_3_1[31] , 
        \wRegOut_3_1[30] , \wRegOut_3_1[29] , \wRegOut_3_1[28] , 
        \wRegOut_3_1[27] , \wRegOut_3_1[26] , \wRegOut_3_1[25] , 
        \wRegOut_3_1[24] , \wRegOut_3_1[23] , \wRegOut_3_1[22] , 
        \wRegOut_3_1[21] , \wRegOut_3_1[20] , \wRegOut_3_1[19] , 
        \wRegOut_3_1[18] , \wRegOut_3_1[17] , \wRegOut_3_1[16] , 
        \wRegOut_3_1[15] , \wRegOut_3_1[14] , \wRegOut_3_1[13] , 
        \wRegOut_3_1[12] , \wRegOut_3_1[11] , \wRegOut_3_1[10] , 
        \wRegOut_3_1[9] , \wRegOut_3_1[8] , \wRegOut_3_1[7] , \wRegOut_3_1[6] , 
        \wRegOut_3_1[5] , \wRegOut_3_1[4] , \wRegOut_3_1[3] , \wRegOut_3_1[2] , 
        \wRegOut_3_1[1] , \wRegOut_3_1[0] }), .P_Out({\wRegInBot_3_1[31] , 
        \wRegInBot_3_1[30] , \wRegInBot_3_1[29] , \wRegInBot_3_1[28] , 
        \wRegInBot_3_1[27] , \wRegInBot_3_1[26] , \wRegInBot_3_1[25] , 
        \wRegInBot_3_1[24] , \wRegInBot_3_1[23] , \wRegInBot_3_1[22] , 
        \wRegInBot_3_1[21] , \wRegInBot_3_1[20] , \wRegInBot_3_1[19] , 
        \wRegInBot_3_1[18] , \wRegInBot_3_1[17] , \wRegInBot_3_1[16] , 
        \wRegInBot_3_1[15] , \wRegInBot_3_1[14] , \wRegInBot_3_1[13] , 
        \wRegInBot_3_1[12] , \wRegInBot_3_1[11] , \wRegInBot_3_1[10] , 
        \wRegInBot_3_1[9] , \wRegInBot_3_1[8] , \wRegInBot_3_1[7] , 
        \wRegInBot_3_1[6] , \wRegInBot_3_1[5] , \wRegInBot_3_1[4] , 
        \wRegInBot_3_1[3] , \wRegInBot_3_1[2] , \wRegInBot_3_1[1] , 
        \wRegInBot_3_1[0] }), .L_WR(\wRegEnTop_4_2[0] ), .L_In({
        \wRegOut_4_2[31] , \wRegOut_4_2[30] , \wRegOut_4_2[29] , 
        \wRegOut_4_2[28] , \wRegOut_4_2[27] , \wRegOut_4_2[26] , 
        \wRegOut_4_2[25] , \wRegOut_4_2[24] , \wRegOut_4_2[23] , 
        \wRegOut_4_2[22] , \wRegOut_4_2[21] , \wRegOut_4_2[20] , 
        \wRegOut_4_2[19] , \wRegOut_4_2[18] , \wRegOut_4_2[17] , 
        \wRegOut_4_2[16] , \wRegOut_4_2[15] , \wRegOut_4_2[14] , 
        \wRegOut_4_2[13] , \wRegOut_4_2[12] , \wRegOut_4_2[11] , 
        \wRegOut_4_2[10] , \wRegOut_4_2[9] , \wRegOut_4_2[8] , 
        \wRegOut_4_2[7] , \wRegOut_4_2[6] , \wRegOut_4_2[5] , \wRegOut_4_2[4] , 
        \wRegOut_4_2[3] , \wRegOut_4_2[2] , \wRegOut_4_2[1] , \wRegOut_4_2[0] 
        }), .L_Out({\wRegInTop_4_2[31] , \wRegInTop_4_2[30] , 
        \wRegInTop_4_2[29] , \wRegInTop_4_2[28] , \wRegInTop_4_2[27] , 
        \wRegInTop_4_2[26] , \wRegInTop_4_2[25] , \wRegInTop_4_2[24] , 
        \wRegInTop_4_2[23] , \wRegInTop_4_2[22] , \wRegInTop_4_2[21] , 
        \wRegInTop_4_2[20] , \wRegInTop_4_2[19] , \wRegInTop_4_2[18] , 
        \wRegInTop_4_2[17] , \wRegInTop_4_2[16] , \wRegInTop_4_2[15] , 
        \wRegInTop_4_2[14] , \wRegInTop_4_2[13] , \wRegInTop_4_2[12] , 
        \wRegInTop_4_2[11] , \wRegInTop_4_2[10] , \wRegInTop_4_2[9] , 
        \wRegInTop_4_2[8] , \wRegInTop_4_2[7] , \wRegInTop_4_2[6] , 
        \wRegInTop_4_2[5] , \wRegInTop_4_2[4] , \wRegInTop_4_2[3] , 
        \wRegInTop_4_2[2] , \wRegInTop_4_2[1] , \wRegInTop_4_2[0] }), .R_WR(
        \wRegEnTop_4_3[0] ), .R_In({\wRegOut_4_3[31] , \wRegOut_4_3[30] , 
        \wRegOut_4_3[29] , \wRegOut_4_3[28] , \wRegOut_4_3[27] , 
        \wRegOut_4_3[26] , \wRegOut_4_3[25] , \wRegOut_4_3[24] , 
        \wRegOut_4_3[23] , \wRegOut_4_3[22] , \wRegOut_4_3[21] , 
        \wRegOut_4_3[20] , \wRegOut_4_3[19] , \wRegOut_4_3[18] , 
        \wRegOut_4_3[17] , \wRegOut_4_3[16] , \wRegOut_4_3[15] , 
        \wRegOut_4_3[14] , \wRegOut_4_3[13] , \wRegOut_4_3[12] , 
        \wRegOut_4_3[11] , \wRegOut_4_3[10] , \wRegOut_4_3[9] , 
        \wRegOut_4_3[8] , \wRegOut_4_3[7] , \wRegOut_4_3[6] , \wRegOut_4_3[5] , 
        \wRegOut_4_3[4] , \wRegOut_4_3[3] , \wRegOut_4_3[2] , \wRegOut_4_3[1] , 
        \wRegOut_4_3[0] }), .R_Out({\wRegInTop_4_3[31] , \wRegInTop_4_3[30] , 
        \wRegInTop_4_3[29] , \wRegInTop_4_3[28] , \wRegInTop_4_3[27] , 
        \wRegInTop_4_3[26] , \wRegInTop_4_3[25] , \wRegInTop_4_3[24] , 
        \wRegInTop_4_3[23] , \wRegInTop_4_3[22] , \wRegInTop_4_3[21] , 
        \wRegInTop_4_3[20] , \wRegInTop_4_3[19] , \wRegInTop_4_3[18] , 
        \wRegInTop_4_3[17] , \wRegInTop_4_3[16] , \wRegInTop_4_3[15] , 
        \wRegInTop_4_3[14] , \wRegInTop_4_3[13] , \wRegInTop_4_3[12] , 
        \wRegInTop_4_3[11] , \wRegInTop_4_3[10] , \wRegInTop_4_3[9] , 
        \wRegInTop_4_3[8] , \wRegInTop_4_3[7] , \wRegInTop_4_3[6] , 
        \wRegInTop_4_3[5] , \wRegInTop_4_3[4] , \wRegInTop_4_3[3] , 
        \wRegInTop_4_3[2] , \wRegInTop_4_3[1] , \wRegInTop_4_3[0] }) );
    BHeap_Node_WIDTH32 BHN_4_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_12[0] ), .P_In({\wRegOut_4_12[31] , 
        \wRegOut_4_12[30] , \wRegOut_4_12[29] , \wRegOut_4_12[28] , 
        \wRegOut_4_12[27] , \wRegOut_4_12[26] , \wRegOut_4_12[25] , 
        \wRegOut_4_12[24] , \wRegOut_4_12[23] , \wRegOut_4_12[22] , 
        \wRegOut_4_12[21] , \wRegOut_4_12[20] , \wRegOut_4_12[19] , 
        \wRegOut_4_12[18] , \wRegOut_4_12[17] , \wRegOut_4_12[16] , 
        \wRegOut_4_12[15] , \wRegOut_4_12[14] , \wRegOut_4_12[13] , 
        \wRegOut_4_12[12] , \wRegOut_4_12[11] , \wRegOut_4_12[10] , 
        \wRegOut_4_12[9] , \wRegOut_4_12[8] , \wRegOut_4_12[7] , 
        \wRegOut_4_12[6] , \wRegOut_4_12[5] , \wRegOut_4_12[4] , 
        \wRegOut_4_12[3] , \wRegOut_4_12[2] , \wRegOut_4_12[1] , 
        \wRegOut_4_12[0] }), .P_Out({\wRegInBot_4_12[31] , 
        \wRegInBot_4_12[30] , \wRegInBot_4_12[29] , \wRegInBot_4_12[28] , 
        \wRegInBot_4_12[27] , \wRegInBot_4_12[26] , \wRegInBot_4_12[25] , 
        \wRegInBot_4_12[24] , \wRegInBot_4_12[23] , \wRegInBot_4_12[22] , 
        \wRegInBot_4_12[21] , \wRegInBot_4_12[20] , \wRegInBot_4_12[19] , 
        \wRegInBot_4_12[18] , \wRegInBot_4_12[17] , \wRegInBot_4_12[16] , 
        \wRegInBot_4_12[15] , \wRegInBot_4_12[14] , \wRegInBot_4_12[13] , 
        \wRegInBot_4_12[12] , \wRegInBot_4_12[11] , \wRegInBot_4_12[10] , 
        \wRegInBot_4_12[9] , \wRegInBot_4_12[8] , \wRegInBot_4_12[7] , 
        \wRegInBot_4_12[6] , \wRegInBot_4_12[5] , \wRegInBot_4_12[4] , 
        \wRegInBot_4_12[3] , \wRegInBot_4_12[2] , \wRegInBot_4_12[1] , 
        \wRegInBot_4_12[0] }), .L_WR(\wRegEnTop_5_24[0] ), .L_In({
        \wRegOut_5_24[31] , \wRegOut_5_24[30] , \wRegOut_5_24[29] , 
        \wRegOut_5_24[28] , \wRegOut_5_24[27] , \wRegOut_5_24[26] , 
        \wRegOut_5_24[25] , \wRegOut_5_24[24] , \wRegOut_5_24[23] , 
        \wRegOut_5_24[22] , \wRegOut_5_24[21] , \wRegOut_5_24[20] , 
        \wRegOut_5_24[19] , \wRegOut_5_24[18] , \wRegOut_5_24[17] , 
        \wRegOut_5_24[16] , \wRegOut_5_24[15] , \wRegOut_5_24[14] , 
        \wRegOut_5_24[13] , \wRegOut_5_24[12] , \wRegOut_5_24[11] , 
        \wRegOut_5_24[10] , \wRegOut_5_24[9] , \wRegOut_5_24[8] , 
        \wRegOut_5_24[7] , \wRegOut_5_24[6] , \wRegOut_5_24[5] , 
        \wRegOut_5_24[4] , \wRegOut_5_24[3] , \wRegOut_5_24[2] , 
        \wRegOut_5_24[1] , \wRegOut_5_24[0] }), .L_Out({\wRegInTop_5_24[31] , 
        \wRegInTop_5_24[30] , \wRegInTop_5_24[29] , \wRegInTop_5_24[28] , 
        \wRegInTop_5_24[27] , \wRegInTop_5_24[26] , \wRegInTop_5_24[25] , 
        \wRegInTop_5_24[24] , \wRegInTop_5_24[23] , \wRegInTop_5_24[22] , 
        \wRegInTop_5_24[21] , \wRegInTop_5_24[20] , \wRegInTop_5_24[19] , 
        \wRegInTop_5_24[18] , \wRegInTop_5_24[17] , \wRegInTop_5_24[16] , 
        \wRegInTop_5_24[15] , \wRegInTop_5_24[14] , \wRegInTop_5_24[13] , 
        \wRegInTop_5_24[12] , \wRegInTop_5_24[11] , \wRegInTop_5_24[10] , 
        \wRegInTop_5_24[9] , \wRegInTop_5_24[8] , \wRegInTop_5_24[7] , 
        \wRegInTop_5_24[6] , \wRegInTop_5_24[5] , \wRegInTop_5_24[4] , 
        \wRegInTop_5_24[3] , \wRegInTop_5_24[2] , \wRegInTop_5_24[1] , 
        \wRegInTop_5_24[0] }), .R_WR(\wRegEnTop_5_25[0] ), .R_In({
        \wRegOut_5_25[31] , \wRegOut_5_25[30] , \wRegOut_5_25[29] , 
        \wRegOut_5_25[28] , \wRegOut_5_25[27] , \wRegOut_5_25[26] , 
        \wRegOut_5_25[25] , \wRegOut_5_25[24] , \wRegOut_5_25[23] , 
        \wRegOut_5_25[22] , \wRegOut_5_25[21] , \wRegOut_5_25[20] , 
        \wRegOut_5_25[19] , \wRegOut_5_25[18] , \wRegOut_5_25[17] , 
        \wRegOut_5_25[16] , \wRegOut_5_25[15] , \wRegOut_5_25[14] , 
        \wRegOut_5_25[13] , \wRegOut_5_25[12] , \wRegOut_5_25[11] , 
        \wRegOut_5_25[10] , \wRegOut_5_25[9] , \wRegOut_5_25[8] , 
        \wRegOut_5_25[7] , \wRegOut_5_25[6] , \wRegOut_5_25[5] , 
        \wRegOut_5_25[4] , \wRegOut_5_25[3] , \wRegOut_5_25[2] , 
        \wRegOut_5_25[1] , \wRegOut_5_25[0] }), .R_Out({\wRegInTop_5_25[31] , 
        \wRegInTop_5_25[30] , \wRegInTop_5_25[29] , \wRegInTop_5_25[28] , 
        \wRegInTop_5_25[27] , \wRegInTop_5_25[26] , \wRegInTop_5_25[25] , 
        \wRegInTop_5_25[24] , \wRegInTop_5_25[23] , \wRegInTop_5_25[22] , 
        \wRegInTop_5_25[21] , \wRegInTop_5_25[20] , \wRegInTop_5_25[19] , 
        \wRegInTop_5_25[18] , \wRegInTop_5_25[17] , \wRegInTop_5_25[16] , 
        \wRegInTop_5_25[15] , \wRegInTop_5_25[14] , \wRegInTop_5_25[13] , 
        \wRegInTop_5_25[12] , \wRegInTop_5_25[11] , \wRegInTop_5_25[10] , 
        \wRegInTop_5_25[9] , \wRegInTop_5_25[8] , \wRegInTop_5_25[7] , 
        \wRegInTop_5_25[6] , \wRegInTop_5_25[5] , \wRegInTop_5_25[4] , 
        \wRegInTop_5_25[3] , \wRegInTop_5_25[2] , \wRegInTop_5_25[1] , 
        \wRegInTop_5_25[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink12[31] , \ScanLink12[30] , \ScanLink12[29] , 
        \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , \ScanLink12[25] , 
        \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , \ScanLink12[21] , 
        \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , \ScanLink12[17] , 
        \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , \ScanLink12[13] , 
        \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , \ScanLink12[9] , 
        \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , \ScanLink12[5] , 
        \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , \ScanLink12[1] , 
        \ScanLink12[0] }), .ScanOut({\ScanLink11[31] , \ScanLink11[30] , 
        \ScanLink11[29] , \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , 
        \ScanLink11[25] , \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , 
        \ScanLink11[21] , \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , 
        \ScanLink11[17] , \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , 
        \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , 
        \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , 
        \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , 
        \ScanLink11[1] , \ScanLink11[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_4[31] , \wRegOut_3_4[30] , \wRegOut_3_4[29] , 
        \wRegOut_3_4[28] , \wRegOut_3_4[27] , \wRegOut_3_4[26] , 
        \wRegOut_3_4[25] , \wRegOut_3_4[24] , \wRegOut_3_4[23] , 
        \wRegOut_3_4[22] , \wRegOut_3_4[21] , \wRegOut_3_4[20] , 
        \wRegOut_3_4[19] , \wRegOut_3_4[18] , \wRegOut_3_4[17] , 
        \wRegOut_3_4[16] , \wRegOut_3_4[15] , \wRegOut_3_4[14] , 
        \wRegOut_3_4[13] , \wRegOut_3_4[12] , \wRegOut_3_4[11] , 
        \wRegOut_3_4[10] , \wRegOut_3_4[9] , \wRegOut_3_4[8] , 
        \wRegOut_3_4[7] , \wRegOut_3_4[6] , \wRegOut_3_4[5] , \wRegOut_3_4[4] , 
        \wRegOut_3_4[3] , \wRegOut_3_4[2] , \wRegOut_3_4[1] , \wRegOut_3_4[0] 
        }), .Enable1(\wRegEnTop_3_4[0] ), .Enable2(\wRegEnBot_3_4[0] ), .In1({
        \wRegInTop_3_4[31] , \wRegInTop_3_4[30] , \wRegInTop_3_4[29] , 
        \wRegInTop_3_4[28] , \wRegInTop_3_4[27] , \wRegInTop_3_4[26] , 
        \wRegInTop_3_4[25] , \wRegInTop_3_4[24] , \wRegInTop_3_4[23] , 
        \wRegInTop_3_4[22] , \wRegInTop_3_4[21] , \wRegInTop_3_4[20] , 
        \wRegInTop_3_4[19] , \wRegInTop_3_4[18] , \wRegInTop_3_4[17] , 
        \wRegInTop_3_4[16] , \wRegInTop_3_4[15] , \wRegInTop_3_4[14] , 
        \wRegInTop_3_4[13] , \wRegInTop_3_4[12] , \wRegInTop_3_4[11] , 
        \wRegInTop_3_4[10] , \wRegInTop_3_4[9] , \wRegInTop_3_4[8] , 
        \wRegInTop_3_4[7] , \wRegInTop_3_4[6] , \wRegInTop_3_4[5] , 
        \wRegInTop_3_4[4] , \wRegInTop_3_4[3] , \wRegInTop_3_4[2] , 
        \wRegInTop_3_4[1] , \wRegInTop_3_4[0] }), .In2({\wRegInBot_3_4[31] , 
        \wRegInBot_3_4[30] , \wRegInBot_3_4[29] , \wRegInBot_3_4[28] , 
        \wRegInBot_3_4[27] , \wRegInBot_3_4[26] , \wRegInBot_3_4[25] , 
        \wRegInBot_3_4[24] , \wRegInBot_3_4[23] , \wRegInBot_3_4[22] , 
        \wRegInBot_3_4[21] , \wRegInBot_3_4[20] , \wRegInBot_3_4[19] , 
        \wRegInBot_3_4[18] , \wRegInBot_3_4[17] , \wRegInBot_3_4[16] , 
        \wRegInBot_3_4[15] , \wRegInBot_3_4[14] , \wRegInBot_3_4[13] , 
        \wRegInBot_3_4[12] , \wRegInBot_3_4[11] , \wRegInBot_3_4[10] , 
        \wRegInBot_3_4[9] , \wRegInBot_3_4[8] , \wRegInBot_3_4[7] , 
        \wRegInBot_3_4[6] , \wRegInBot_3_4[5] , \wRegInBot_3_4[4] , 
        \wRegInBot_3_4[3] , \wRegInBot_3_4[2] , \wRegInBot_3_4[1] , 
        \wRegInBot_3_4[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink25[31] , \ScanLink25[30] , \ScanLink25[29] , 
        \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , \ScanLink25[25] , 
        \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , \ScanLink25[21] , 
        \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , \ScanLink25[17] , 
        \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , \ScanLink25[13] , 
        \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , \ScanLink25[9] , 
        \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , \ScanLink25[5] , 
        \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , \ScanLink25[1] , 
        \ScanLink25[0] }), .ScanOut({\ScanLink24[31] , \ScanLink24[30] , 
        \ScanLink24[29] , \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , 
        \ScanLink24[25] , \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , 
        \ScanLink24[21] , \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , 
        \ScanLink24[17] , \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , 
        \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , 
        \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , 
        \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , 
        \ScanLink24[1] , \ScanLink24[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_9[31] , \wRegOut_4_9[30] , \wRegOut_4_9[29] , 
        \wRegOut_4_9[28] , \wRegOut_4_9[27] , \wRegOut_4_9[26] , 
        \wRegOut_4_9[25] , \wRegOut_4_9[24] , \wRegOut_4_9[23] , 
        \wRegOut_4_9[22] , \wRegOut_4_9[21] , \wRegOut_4_9[20] , 
        \wRegOut_4_9[19] , \wRegOut_4_9[18] , \wRegOut_4_9[17] , 
        \wRegOut_4_9[16] , \wRegOut_4_9[15] , \wRegOut_4_9[14] , 
        \wRegOut_4_9[13] , \wRegOut_4_9[12] , \wRegOut_4_9[11] , 
        \wRegOut_4_9[10] , \wRegOut_4_9[9] , \wRegOut_4_9[8] , 
        \wRegOut_4_9[7] , \wRegOut_4_9[6] , \wRegOut_4_9[5] , \wRegOut_4_9[4] , 
        \wRegOut_4_9[3] , \wRegOut_4_9[2] , \wRegOut_4_9[1] , \wRegOut_4_9[0] 
        }), .Enable1(\wRegEnTop_4_9[0] ), .Enable2(\wRegEnBot_4_9[0] ), .In1({
        \wRegInTop_4_9[31] , \wRegInTop_4_9[30] , \wRegInTop_4_9[29] , 
        \wRegInTop_4_9[28] , \wRegInTop_4_9[27] , \wRegInTop_4_9[26] , 
        \wRegInTop_4_9[25] , \wRegInTop_4_9[24] , \wRegInTop_4_9[23] , 
        \wRegInTop_4_9[22] , \wRegInTop_4_9[21] , \wRegInTop_4_9[20] , 
        \wRegInTop_4_9[19] , \wRegInTop_4_9[18] , \wRegInTop_4_9[17] , 
        \wRegInTop_4_9[16] , \wRegInTop_4_9[15] , \wRegInTop_4_9[14] , 
        \wRegInTop_4_9[13] , \wRegInTop_4_9[12] , \wRegInTop_4_9[11] , 
        \wRegInTop_4_9[10] , \wRegInTop_4_9[9] , \wRegInTop_4_9[8] , 
        \wRegInTop_4_9[7] , \wRegInTop_4_9[6] , \wRegInTop_4_9[5] , 
        \wRegInTop_4_9[4] , \wRegInTop_4_9[3] , \wRegInTop_4_9[2] , 
        \wRegInTop_4_9[1] , \wRegInTop_4_9[0] }), .In2({\wRegInBot_4_9[31] , 
        \wRegInBot_4_9[30] , \wRegInBot_4_9[29] , \wRegInBot_4_9[28] , 
        \wRegInBot_4_9[27] , \wRegInBot_4_9[26] , \wRegInBot_4_9[25] , 
        \wRegInBot_4_9[24] , \wRegInBot_4_9[23] , \wRegInBot_4_9[22] , 
        \wRegInBot_4_9[21] , \wRegInBot_4_9[20] , \wRegInBot_4_9[19] , 
        \wRegInBot_4_9[18] , \wRegInBot_4_9[17] , \wRegInBot_4_9[16] , 
        \wRegInBot_4_9[15] , \wRegInBot_4_9[14] , \wRegInBot_4_9[13] , 
        \wRegInBot_4_9[12] , \wRegInBot_4_9[11] , \wRegInBot_4_9[10] , 
        \wRegInBot_4_9[9] , \wRegInBot_4_9[8] , \wRegInBot_4_9[7] , 
        \wRegInBot_4_9[6] , \wRegInBot_4_9[5] , \wRegInBot_4_9[4] , 
        \wRegInBot_4_9[3] , \wRegInBot_4_9[2] , \wRegInBot_4_9[1] , 
        \wRegInBot_4_9[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink23[31] , \ScanLink23[30] , \ScanLink23[29] , 
        \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , \ScanLink23[25] , 
        \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , \ScanLink23[21] , 
        \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , \ScanLink23[17] , 
        \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , \ScanLink23[13] , 
        \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , \ScanLink23[9] , 
        \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , \ScanLink23[5] , 
        \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , \ScanLink23[1] , 
        \ScanLink23[0] }), .ScanOut({\ScanLink22[31] , \ScanLink22[30] , 
        \ScanLink22[29] , \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , 
        \ScanLink22[25] , \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , 
        \ScanLink22[21] , \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , 
        \ScanLink22[17] , \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , 
        \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , 
        \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , 
        \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , 
        \ScanLink22[1] , \ScanLink22[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_7[31] , \wRegOut_4_7[30] , \wRegOut_4_7[29] , 
        \wRegOut_4_7[28] , \wRegOut_4_7[27] , \wRegOut_4_7[26] , 
        \wRegOut_4_7[25] , \wRegOut_4_7[24] , \wRegOut_4_7[23] , 
        \wRegOut_4_7[22] , \wRegOut_4_7[21] , \wRegOut_4_7[20] , 
        \wRegOut_4_7[19] , \wRegOut_4_7[18] , \wRegOut_4_7[17] , 
        \wRegOut_4_7[16] , \wRegOut_4_7[15] , \wRegOut_4_7[14] , 
        \wRegOut_4_7[13] , \wRegOut_4_7[12] , \wRegOut_4_7[11] , 
        \wRegOut_4_7[10] , \wRegOut_4_7[9] , \wRegOut_4_7[8] , 
        \wRegOut_4_7[7] , \wRegOut_4_7[6] , \wRegOut_4_7[5] , \wRegOut_4_7[4] , 
        \wRegOut_4_7[3] , \wRegOut_4_7[2] , \wRegOut_4_7[1] , \wRegOut_4_7[0] 
        }), .Enable1(\wRegEnTop_4_7[0] ), .Enable2(\wRegEnBot_4_7[0] ), .In1({
        \wRegInTop_4_7[31] , \wRegInTop_4_7[30] , \wRegInTop_4_7[29] , 
        \wRegInTop_4_7[28] , \wRegInTop_4_7[27] , \wRegInTop_4_7[26] , 
        \wRegInTop_4_7[25] , \wRegInTop_4_7[24] , \wRegInTop_4_7[23] , 
        \wRegInTop_4_7[22] , \wRegInTop_4_7[21] , \wRegInTop_4_7[20] , 
        \wRegInTop_4_7[19] , \wRegInTop_4_7[18] , \wRegInTop_4_7[17] , 
        \wRegInTop_4_7[16] , \wRegInTop_4_7[15] , \wRegInTop_4_7[14] , 
        \wRegInTop_4_7[13] , \wRegInTop_4_7[12] , \wRegInTop_4_7[11] , 
        \wRegInTop_4_7[10] , \wRegInTop_4_7[9] , \wRegInTop_4_7[8] , 
        \wRegInTop_4_7[7] , \wRegInTop_4_7[6] , \wRegInTop_4_7[5] , 
        \wRegInTop_4_7[4] , \wRegInTop_4_7[3] , \wRegInTop_4_7[2] , 
        \wRegInTop_4_7[1] , \wRegInTop_4_7[0] }), .In2({\wRegInBot_4_7[31] , 
        \wRegInBot_4_7[30] , \wRegInBot_4_7[29] , \wRegInBot_4_7[28] , 
        \wRegInBot_4_7[27] , \wRegInBot_4_7[26] , \wRegInBot_4_7[25] , 
        \wRegInBot_4_7[24] , \wRegInBot_4_7[23] , \wRegInBot_4_7[22] , 
        \wRegInBot_4_7[21] , \wRegInBot_4_7[20] , \wRegInBot_4_7[19] , 
        \wRegInBot_4_7[18] , \wRegInBot_4_7[17] , \wRegInBot_4_7[16] , 
        \wRegInBot_4_7[15] , \wRegInBot_4_7[14] , \wRegInBot_4_7[13] , 
        \wRegInBot_4_7[12] , \wRegInBot_4_7[11] , \wRegInBot_4_7[10] , 
        \wRegInBot_4_7[9] , \wRegInBot_4_7[8] , \wRegInBot_4_7[7] , 
        \wRegInBot_4_7[6] , \wRegInBot_4_7[5] , \wRegInBot_4_7[4] , 
        \wRegInBot_4_7[3] , \wRegInBot_4_7[2] , \wRegInBot_4_7[1] , 
        \wRegInBot_4_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_27 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink59[31] , \ScanLink59[30] , \ScanLink59[29] , 
        \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , \ScanLink59[25] , 
        \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , \ScanLink59[21] , 
        \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , \ScanLink59[17] , 
        \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , \ScanLink59[13] , 
        \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , \ScanLink59[9] , 
        \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , \ScanLink59[5] , 
        \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , \ScanLink59[1] , 
        \ScanLink59[0] }), .ScanOut({\ScanLink58[31] , \ScanLink58[30] , 
        \ScanLink58[29] , \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , 
        \ScanLink58[25] , \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , 
        \ScanLink58[21] , \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , 
        \ScanLink58[17] , \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , 
        \ScanLink58[13] , \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , 
        \ScanLink58[9] , \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , 
        \ScanLink58[5] , \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , 
        \ScanLink58[1] , \ScanLink58[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_27[31] , \wRegOut_5_27[30] , 
        \wRegOut_5_27[29] , \wRegOut_5_27[28] , \wRegOut_5_27[27] , 
        \wRegOut_5_27[26] , \wRegOut_5_27[25] , \wRegOut_5_27[24] , 
        \wRegOut_5_27[23] , \wRegOut_5_27[22] , \wRegOut_5_27[21] , 
        \wRegOut_5_27[20] , \wRegOut_5_27[19] , \wRegOut_5_27[18] , 
        \wRegOut_5_27[17] , \wRegOut_5_27[16] , \wRegOut_5_27[15] , 
        \wRegOut_5_27[14] , \wRegOut_5_27[13] , \wRegOut_5_27[12] , 
        \wRegOut_5_27[11] , \wRegOut_5_27[10] , \wRegOut_5_27[9] , 
        \wRegOut_5_27[8] , \wRegOut_5_27[7] , \wRegOut_5_27[6] , 
        \wRegOut_5_27[5] , \wRegOut_5_27[4] , \wRegOut_5_27[3] , 
        \wRegOut_5_27[2] , \wRegOut_5_27[1] , \wRegOut_5_27[0] }), .Enable1(
        \wRegEnTop_5_27[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_27[31] , 
        \wRegInTop_5_27[30] , \wRegInTop_5_27[29] , \wRegInTop_5_27[28] , 
        \wRegInTop_5_27[27] , \wRegInTop_5_27[26] , \wRegInTop_5_27[25] , 
        \wRegInTop_5_27[24] , \wRegInTop_5_27[23] , \wRegInTop_5_27[22] , 
        \wRegInTop_5_27[21] , \wRegInTop_5_27[20] , \wRegInTop_5_27[19] , 
        \wRegInTop_5_27[18] , \wRegInTop_5_27[17] , \wRegInTop_5_27[16] , 
        \wRegInTop_5_27[15] , \wRegInTop_5_27[14] , \wRegInTop_5_27[13] , 
        \wRegInTop_5_27[12] , \wRegInTop_5_27[11] , \wRegInTop_5_27[10] , 
        \wRegInTop_5_27[9] , \wRegInTop_5_27[8] , \wRegInTop_5_27[7] , 
        \wRegInTop_5_27[6] , \wRegInTop_5_27[5] , \wRegInTop_5_27[4] , 
        \wRegInTop_5_27[3] , \wRegInTop_5_27[2] , \wRegInTop_5_27[1] , 
        \wRegInTop_5_27[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_6[0] ), .P_In({\wRegOut_3_6[31] , 
        \wRegOut_3_6[30] , \wRegOut_3_6[29] , \wRegOut_3_6[28] , 
        \wRegOut_3_6[27] , \wRegOut_3_6[26] , \wRegOut_3_6[25] , 
        \wRegOut_3_6[24] , \wRegOut_3_6[23] , \wRegOut_3_6[22] , 
        \wRegOut_3_6[21] , \wRegOut_3_6[20] , \wRegOut_3_6[19] , 
        \wRegOut_3_6[18] , \wRegOut_3_6[17] , \wRegOut_3_6[16] , 
        \wRegOut_3_6[15] , \wRegOut_3_6[14] , \wRegOut_3_6[13] , 
        \wRegOut_3_6[12] , \wRegOut_3_6[11] , \wRegOut_3_6[10] , 
        \wRegOut_3_6[9] , \wRegOut_3_6[8] , \wRegOut_3_6[7] , \wRegOut_3_6[6] , 
        \wRegOut_3_6[5] , \wRegOut_3_6[4] , \wRegOut_3_6[3] , \wRegOut_3_6[2] , 
        \wRegOut_3_6[1] , \wRegOut_3_6[0] }), .P_Out({\wRegInBot_3_6[31] , 
        \wRegInBot_3_6[30] , \wRegInBot_3_6[29] , \wRegInBot_3_6[28] , 
        \wRegInBot_3_6[27] , \wRegInBot_3_6[26] , \wRegInBot_3_6[25] , 
        \wRegInBot_3_6[24] , \wRegInBot_3_6[23] , \wRegInBot_3_6[22] , 
        \wRegInBot_3_6[21] , \wRegInBot_3_6[20] , \wRegInBot_3_6[19] , 
        \wRegInBot_3_6[18] , \wRegInBot_3_6[17] , \wRegInBot_3_6[16] , 
        \wRegInBot_3_6[15] , \wRegInBot_3_6[14] , \wRegInBot_3_6[13] , 
        \wRegInBot_3_6[12] , \wRegInBot_3_6[11] , \wRegInBot_3_6[10] , 
        \wRegInBot_3_6[9] , \wRegInBot_3_6[8] , \wRegInBot_3_6[7] , 
        \wRegInBot_3_6[6] , \wRegInBot_3_6[5] , \wRegInBot_3_6[4] , 
        \wRegInBot_3_6[3] , \wRegInBot_3_6[2] , \wRegInBot_3_6[1] , 
        \wRegInBot_3_6[0] }), .L_WR(\wRegEnTop_4_12[0] ), .L_In({
        \wRegOut_4_12[31] , \wRegOut_4_12[30] , \wRegOut_4_12[29] , 
        \wRegOut_4_12[28] , \wRegOut_4_12[27] , \wRegOut_4_12[26] , 
        \wRegOut_4_12[25] , \wRegOut_4_12[24] , \wRegOut_4_12[23] , 
        \wRegOut_4_12[22] , \wRegOut_4_12[21] , \wRegOut_4_12[20] , 
        \wRegOut_4_12[19] , \wRegOut_4_12[18] , \wRegOut_4_12[17] , 
        \wRegOut_4_12[16] , \wRegOut_4_12[15] , \wRegOut_4_12[14] , 
        \wRegOut_4_12[13] , \wRegOut_4_12[12] , \wRegOut_4_12[11] , 
        \wRegOut_4_12[10] , \wRegOut_4_12[9] , \wRegOut_4_12[8] , 
        \wRegOut_4_12[7] , \wRegOut_4_12[6] , \wRegOut_4_12[5] , 
        \wRegOut_4_12[4] , \wRegOut_4_12[3] , \wRegOut_4_12[2] , 
        \wRegOut_4_12[1] , \wRegOut_4_12[0] }), .L_Out({\wRegInTop_4_12[31] , 
        \wRegInTop_4_12[30] , \wRegInTop_4_12[29] , \wRegInTop_4_12[28] , 
        \wRegInTop_4_12[27] , \wRegInTop_4_12[26] , \wRegInTop_4_12[25] , 
        \wRegInTop_4_12[24] , \wRegInTop_4_12[23] , \wRegInTop_4_12[22] , 
        \wRegInTop_4_12[21] , \wRegInTop_4_12[20] , \wRegInTop_4_12[19] , 
        \wRegInTop_4_12[18] , \wRegInTop_4_12[17] , \wRegInTop_4_12[16] , 
        \wRegInTop_4_12[15] , \wRegInTop_4_12[14] , \wRegInTop_4_12[13] , 
        \wRegInTop_4_12[12] , \wRegInTop_4_12[11] , \wRegInTop_4_12[10] , 
        \wRegInTop_4_12[9] , \wRegInTop_4_12[8] , \wRegInTop_4_12[7] , 
        \wRegInTop_4_12[6] , \wRegInTop_4_12[5] , \wRegInTop_4_12[4] , 
        \wRegInTop_4_12[3] , \wRegInTop_4_12[2] , \wRegInTop_4_12[1] , 
        \wRegInTop_4_12[0] }), .R_WR(\wRegEnTop_4_13[0] ), .R_In({
        \wRegOut_4_13[31] , \wRegOut_4_13[30] , \wRegOut_4_13[29] , 
        \wRegOut_4_13[28] , \wRegOut_4_13[27] , \wRegOut_4_13[26] , 
        \wRegOut_4_13[25] , \wRegOut_4_13[24] , \wRegOut_4_13[23] , 
        \wRegOut_4_13[22] , \wRegOut_4_13[21] , \wRegOut_4_13[20] , 
        \wRegOut_4_13[19] , \wRegOut_4_13[18] , \wRegOut_4_13[17] , 
        \wRegOut_4_13[16] , \wRegOut_4_13[15] , \wRegOut_4_13[14] , 
        \wRegOut_4_13[13] , \wRegOut_4_13[12] , \wRegOut_4_13[11] , 
        \wRegOut_4_13[10] , \wRegOut_4_13[9] , \wRegOut_4_13[8] , 
        \wRegOut_4_13[7] , \wRegOut_4_13[6] , \wRegOut_4_13[5] , 
        \wRegOut_4_13[4] , \wRegOut_4_13[3] , \wRegOut_4_13[2] , 
        \wRegOut_4_13[1] , \wRegOut_4_13[0] }), .R_Out({\wRegInTop_4_13[31] , 
        \wRegInTop_4_13[30] , \wRegInTop_4_13[29] , \wRegInTop_4_13[28] , 
        \wRegInTop_4_13[27] , \wRegInTop_4_13[26] , \wRegInTop_4_13[25] , 
        \wRegInTop_4_13[24] , \wRegInTop_4_13[23] , \wRegInTop_4_13[22] , 
        \wRegInTop_4_13[21] , \wRegInTop_4_13[20] , \wRegInTop_4_13[19] , 
        \wRegInTop_4_13[18] , \wRegInTop_4_13[17] , \wRegInTop_4_13[16] , 
        \wRegInTop_4_13[15] , \wRegInTop_4_13[14] , \wRegInTop_4_13[13] , 
        \wRegInTop_4_13[12] , \wRegInTop_4_13[11] , \wRegInTop_4_13[10] , 
        \wRegInTop_4_13[9] , \wRegInTop_4_13[8] , \wRegInTop_4_13[7] , 
        \wRegInTop_4_13[6] , \wRegInTop_4_13[5] , \wRegInTop_4_13[4] , 
        \wRegInTop_4_13[3] , \wRegInTop_4_13[2] , \wRegInTop_4_13[1] , 
        \wRegInTop_4_13[0] }) );
    BHeap_CtrlReg_WIDTH32 BHCR_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_3[0] ), 
        .Out(\wCtrlOut_2[0] ), .Enable(\wEnable_2[0] ) );
    BHeap_Node_WIDTH32 BHN_4_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_15[0] ), .P_In({\wRegOut_4_15[31] , 
        \wRegOut_4_15[30] , \wRegOut_4_15[29] , \wRegOut_4_15[28] , 
        \wRegOut_4_15[27] , \wRegOut_4_15[26] , \wRegOut_4_15[25] , 
        \wRegOut_4_15[24] , \wRegOut_4_15[23] , \wRegOut_4_15[22] , 
        \wRegOut_4_15[21] , \wRegOut_4_15[20] , \wRegOut_4_15[19] , 
        \wRegOut_4_15[18] , \wRegOut_4_15[17] , \wRegOut_4_15[16] , 
        \wRegOut_4_15[15] , \wRegOut_4_15[14] , \wRegOut_4_15[13] , 
        \wRegOut_4_15[12] , \wRegOut_4_15[11] , \wRegOut_4_15[10] , 
        \wRegOut_4_15[9] , \wRegOut_4_15[8] , \wRegOut_4_15[7] , 
        \wRegOut_4_15[6] , \wRegOut_4_15[5] , \wRegOut_4_15[4] , 
        \wRegOut_4_15[3] , \wRegOut_4_15[2] , \wRegOut_4_15[1] , 
        \wRegOut_4_15[0] }), .P_Out({\wRegInBot_4_15[31] , 
        \wRegInBot_4_15[30] , \wRegInBot_4_15[29] , \wRegInBot_4_15[28] , 
        \wRegInBot_4_15[27] , \wRegInBot_4_15[26] , \wRegInBot_4_15[25] , 
        \wRegInBot_4_15[24] , \wRegInBot_4_15[23] , \wRegInBot_4_15[22] , 
        \wRegInBot_4_15[21] , \wRegInBot_4_15[20] , \wRegInBot_4_15[19] , 
        \wRegInBot_4_15[18] , \wRegInBot_4_15[17] , \wRegInBot_4_15[16] , 
        \wRegInBot_4_15[15] , \wRegInBot_4_15[14] , \wRegInBot_4_15[13] , 
        \wRegInBot_4_15[12] , \wRegInBot_4_15[11] , \wRegInBot_4_15[10] , 
        \wRegInBot_4_15[9] , \wRegInBot_4_15[8] , \wRegInBot_4_15[7] , 
        \wRegInBot_4_15[6] , \wRegInBot_4_15[5] , \wRegInBot_4_15[4] , 
        \wRegInBot_4_15[3] , \wRegInBot_4_15[2] , \wRegInBot_4_15[1] , 
        \wRegInBot_4_15[0] }), .L_WR(\wRegEnTop_5_30[0] ), .L_In({
        \wRegOut_5_30[31] , \wRegOut_5_30[30] , \wRegOut_5_30[29] , 
        \wRegOut_5_30[28] , \wRegOut_5_30[27] , \wRegOut_5_30[26] , 
        \wRegOut_5_30[25] , \wRegOut_5_30[24] , \wRegOut_5_30[23] , 
        \wRegOut_5_30[22] , \wRegOut_5_30[21] , \wRegOut_5_30[20] , 
        \wRegOut_5_30[19] , \wRegOut_5_30[18] , \wRegOut_5_30[17] , 
        \wRegOut_5_30[16] , \wRegOut_5_30[15] , \wRegOut_5_30[14] , 
        \wRegOut_5_30[13] , \wRegOut_5_30[12] , \wRegOut_5_30[11] , 
        \wRegOut_5_30[10] , \wRegOut_5_30[9] , \wRegOut_5_30[8] , 
        \wRegOut_5_30[7] , \wRegOut_5_30[6] , \wRegOut_5_30[5] , 
        \wRegOut_5_30[4] , \wRegOut_5_30[3] , \wRegOut_5_30[2] , 
        \wRegOut_5_30[1] , \wRegOut_5_30[0] }), .L_Out({\wRegInTop_5_30[31] , 
        \wRegInTop_5_30[30] , \wRegInTop_5_30[29] , \wRegInTop_5_30[28] , 
        \wRegInTop_5_30[27] , \wRegInTop_5_30[26] , \wRegInTop_5_30[25] , 
        \wRegInTop_5_30[24] , \wRegInTop_5_30[23] , \wRegInTop_5_30[22] , 
        \wRegInTop_5_30[21] , \wRegInTop_5_30[20] , \wRegInTop_5_30[19] , 
        \wRegInTop_5_30[18] , \wRegInTop_5_30[17] , \wRegInTop_5_30[16] , 
        \wRegInTop_5_30[15] , \wRegInTop_5_30[14] , \wRegInTop_5_30[13] , 
        \wRegInTop_5_30[12] , \wRegInTop_5_30[11] , \wRegInTop_5_30[10] , 
        \wRegInTop_5_30[9] , \wRegInTop_5_30[8] , \wRegInTop_5_30[7] , 
        \wRegInTop_5_30[6] , \wRegInTop_5_30[5] , \wRegInTop_5_30[4] , 
        \wRegInTop_5_30[3] , \wRegInTop_5_30[2] , \wRegInTop_5_30[1] , 
        \wRegInTop_5_30[0] }), .R_WR(\wRegEnTop_5_31[0] ), .R_In({
        \wRegOut_5_31[31] , \wRegOut_5_31[30] , \wRegOut_5_31[29] , 
        \wRegOut_5_31[28] , \wRegOut_5_31[27] , \wRegOut_5_31[26] , 
        \wRegOut_5_31[25] , \wRegOut_5_31[24] , \wRegOut_5_31[23] , 
        \wRegOut_5_31[22] , \wRegOut_5_31[21] , \wRegOut_5_31[20] , 
        \wRegOut_5_31[19] , \wRegOut_5_31[18] , \wRegOut_5_31[17] , 
        \wRegOut_5_31[16] , \wRegOut_5_31[15] , \wRegOut_5_31[14] , 
        \wRegOut_5_31[13] , \wRegOut_5_31[12] , \wRegOut_5_31[11] , 
        \wRegOut_5_31[10] , \wRegOut_5_31[9] , \wRegOut_5_31[8] , 
        \wRegOut_5_31[7] , \wRegOut_5_31[6] , \wRegOut_5_31[5] , 
        \wRegOut_5_31[4] , \wRegOut_5_31[3] , \wRegOut_5_31[2] , 
        \wRegOut_5_31[1] , \wRegOut_5_31[0] }), .R_Out({\wRegInTop_5_31[31] , 
        \wRegInTop_5_31[30] , \wRegInTop_5_31[29] , \wRegInTop_5_31[28] , 
        \wRegInTop_5_31[27] , \wRegInTop_5_31[26] , \wRegInTop_5_31[25] , 
        \wRegInTop_5_31[24] , \wRegInTop_5_31[23] , \wRegInTop_5_31[22] , 
        \wRegInTop_5_31[21] , \wRegInTop_5_31[20] , \wRegInTop_5_31[19] , 
        \wRegInTop_5_31[18] , \wRegInTop_5_31[17] , \wRegInTop_5_31[16] , 
        \wRegInTop_5_31[15] , \wRegInTop_5_31[14] , \wRegInTop_5_31[13] , 
        \wRegInTop_5_31[12] , \wRegInTop_5_31[11] , \wRegInTop_5_31[10] , 
        \wRegInTop_5_31[9] , \wRegInTop_5_31[8] , \wRegInTop_5_31[7] , 
        \wRegInTop_5_31[6] , \wRegInTop_5_31[5] , \wRegInTop_5_31[4] , 
        \wRegInTop_5_31[3] , \wRegInTop_5_31[2] , \wRegInTop_5_31[1] , 
        \wRegInTop_5_31[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink44[31] , \ScanLink44[30] , \ScanLink44[29] , 
        \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , \ScanLink44[25] , 
        \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , \ScanLink44[21] , 
        \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , \ScanLink44[17] , 
        \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , \ScanLink44[13] , 
        \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , \ScanLink44[9] , 
        \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , \ScanLink44[5] , 
        \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , \ScanLink44[1] , 
        \ScanLink44[0] }), .ScanOut({\ScanLink43[31] , \ScanLink43[30] , 
        \ScanLink43[29] , \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , 
        \ScanLink43[25] , \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , 
        \ScanLink43[21] , \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , 
        \ScanLink43[17] , \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , 
        \ScanLink43[13] , \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , 
        \ScanLink43[9] , \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , 
        \ScanLink43[5] , \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , 
        \ScanLink43[1] , \ScanLink43[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_12[31] , \wRegOut_5_12[30] , 
        \wRegOut_5_12[29] , \wRegOut_5_12[28] , \wRegOut_5_12[27] , 
        \wRegOut_5_12[26] , \wRegOut_5_12[25] , \wRegOut_5_12[24] , 
        \wRegOut_5_12[23] , \wRegOut_5_12[22] , \wRegOut_5_12[21] , 
        \wRegOut_5_12[20] , \wRegOut_5_12[19] , \wRegOut_5_12[18] , 
        \wRegOut_5_12[17] , \wRegOut_5_12[16] , \wRegOut_5_12[15] , 
        \wRegOut_5_12[14] , \wRegOut_5_12[13] , \wRegOut_5_12[12] , 
        \wRegOut_5_12[11] , \wRegOut_5_12[10] , \wRegOut_5_12[9] , 
        \wRegOut_5_12[8] , \wRegOut_5_12[7] , \wRegOut_5_12[6] , 
        \wRegOut_5_12[5] , \wRegOut_5_12[4] , \wRegOut_5_12[3] , 
        \wRegOut_5_12[2] , \wRegOut_5_12[1] , \wRegOut_5_12[0] }), .Enable1(
        \wRegEnTop_5_12[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_12[31] , 
        \wRegInTop_5_12[30] , \wRegInTop_5_12[29] , \wRegInTop_5_12[28] , 
        \wRegInTop_5_12[27] , \wRegInTop_5_12[26] , \wRegInTop_5_12[25] , 
        \wRegInTop_5_12[24] , \wRegInTop_5_12[23] , \wRegInTop_5_12[22] , 
        \wRegInTop_5_12[21] , \wRegInTop_5_12[20] , \wRegInTop_5_12[19] , 
        \wRegInTop_5_12[18] , \wRegInTop_5_12[17] , \wRegInTop_5_12[16] , 
        \wRegInTop_5_12[15] , \wRegInTop_5_12[14] , \wRegInTop_5_12[13] , 
        \wRegInTop_5_12[12] , \wRegInTop_5_12[11] , \wRegInTop_5_12[10] , 
        \wRegInTop_5_12[9] , \wRegInTop_5_12[8] , \wRegInTop_5_12[7] , 
        \wRegInTop_5_12[6] , \wRegInTop_5_12[5] , \wRegInTop_5_12[4] , 
        \wRegInTop_5_12[3] , \wRegInTop_5_12[2] , \wRegInTop_5_12[1] , 
        \wRegInTop_5_12[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_2_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink4[31] , \ScanLink4[30] , \ScanLink4[29] , 
        \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , \ScanLink4[25] , 
        \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , \ScanLink4[21] , 
        \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , \ScanLink4[17] , 
        \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , \ScanLink4[13] , 
        \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , \ScanLink4[9] , 
        \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , \ScanLink4[5] , 
        \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , \ScanLink4[1] , 
        \ScanLink4[0] }), .ScanOut({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_2_0[31] , \wRegOut_2_0[30] , \wRegOut_2_0[29] , 
        \wRegOut_2_0[28] , \wRegOut_2_0[27] , \wRegOut_2_0[26] , 
        \wRegOut_2_0[25] , \wRegOut_2_0[24] , \wRegOut_2_0[23] , 
        \wRegOut_2_0[22] , \wRegOut_2_0[21] , \wRegOut_2_0[20] , 
        \wRegOut_2_0[19] , \wRegOut_2_0[18] , \wRegOut_2_0[17] , 
        \wRegOut_2_0[16] , \wRegOut_2_0[15] , \wRegOut_2_0[14] , 
        \wRegOut_2_0[13] , \wRegOut_2_0[12] , \wRegOut_2_0[11] , 
        \wRegOut_2_0[10] , \wRegOut_2_0[9] , \wRegOut_2_0[8] , 
        \wRegOut_2_0[7] , \wRegOut_2_0[6] , \wRegOut_2_0[5] , \wRegOut_2_0[4] , 
        \wRegOut_2_0[3] , \wRegOut_2_0[2] , \wRegOut_2_0[1] , \wRegOut_2_0[0] 
        }), .Enable1(\wRegEnTop_2_0[0] ), .Enable2(\wRegEnBot_2_0[0] ), .In1({
        \wRegInTop_2_0[31] , \wRegInTop_2_0[30] , \wRegInTop_2_0[29] , 
        \wRegInTop_2_0[28] , \wRegInTop_2_0[27] , \wRegInTop_2_0[26] , 
        \wRegInTop_2_0[25] , \wRegInTop_2_0[24] , \wRegInTop_2_0[23] , 
        \wRegInTop_2_0[22] , \wRegInTop_2_0[21] , \wRegInTop_2_0[20] , 
        \wRegInTop_2_0[19] , \wRegInTop_2_0[18] , \wRegInTop_2_0[17] , 
        \wRegInTop_2_0[16] , \wRegInTop_2_0[15] , \wRegInTop_2_0[14] , 
        \wRegInTop_2_0[13] , \wRegInTop_2_0[12] , \wRegInTop_2_0[11] , 
        \wRegInTop_2_0[10] , \wRegInTop_2_0[9] , \wRegInTop_2_0[8] , 
        \wRegInTop_2_0[7] , \wRegInTop_2_0[6] , \wRegInTop_2_0[5] , 
        \wRegInTop_2_0[4] , \wRegInTop_2_0[3] , \wRegInTop_2_0[2] , 
        \wRegInTop_2_0[1] , \wRegInTop_2_0[0] }), .In2({\wRegInBot_2_0[31] , 
        \wRegInBot_2_0[30] , \wRegInBot_2_0[29] , \wRegInBot_2_0[28] , 
        \wRegInBot_2_0[27] , \wRegInBot_2_0[26] , \wRegInBot_2_0[25] , 
        \wRegInBot_2_0[24] , \wRegInBot_2_0[23] , \wRegInBot_2_0[22] , 
        \wRegInBot_2_0[21] , \wRegInBot_2_0[20] , \wRegInBot_2_0[19] , 
        \wRegInBot_2_0[18] , \wRegInBot_2_0[17] , \wRegInBot_2_0[16] , 
        \wRegInBot_2_0[15] , \wRegInBot_2_0[14] , \wRegInBot_2_0[13] , 
        \wRegInBot_2_0[12] , \wRegInBot_2_0[11] , \wRegInBot_2_0[10] , 
        \wRegInBot_2_0[9] , \wRegInBot_2_0[8] , \wRegInBot_2_0[7] , 
        \wRegInBot_2_0[6] , \wRegInBot_2_0[5] , \wRegInBot_2_0[4] , 
        \wRegInBot_2_0[3] , \wRegInBot_2_0[2] , \wRegInBot_2_0[1] , 
        \wRegInBot_2_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_2_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink5[31] , \ScanLink5[30] , \ScanLink5[29] , 
        \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , \ScanLink5[25] , 
        \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , \ScanLink5[21] , 
        \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , \ScanLink5[17] , 
        \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , \ScanLink5[13] , 
        \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , \ScanLink5[9] , 
        \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , \ScanLink5[5] , 
        \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , \ScanLink5[1] , 
        \ScanLink5[0] }), .ScanOut({\ScanLink4[31] , \ScanLink4[30] , 
        \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , 
        \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , 
        \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , 
        \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , 
        \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , 
        \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_2_1[31] , \wRegOut_2_1[30] , \wRegOut_2_1[29] , 
        \wRegOut_2_1[28] , \wRegOut_2_1[27] , \wRegOut_2_1[26] , 
        \wRegOut_2_1[25] , \wRegOut_2_1[24] , \wRegOut_2_1[23] , 
        \wRegOut_2_1[22] , \wRegOut_2_1[21] , \wRegOut_2_1[20] , 
        \wRegOut_2_1[19] , \wRegOut_2_1[18] , \wRegOut_2_1[17] , 
        \wRegOut_2_1[16] , \wRegOut_2_1[15] , \wRegOut_2_1[14] , 
        \wRegOut_2_1[13] , \wRegOut_2_1[12] , \wRegOut_2_1[11] , 
        \wRegOut_2_1[10] , \wRegOut_2_1[9] , \wRegOut_2_1[8] , 
        \wRegOut_2_1[7] , \wRegOut_2_1[6] , \wRegOut_2_1[5] , \wRegOut_2_1[4] , 
        \wRegOut_2_1[3] , \wRegOut_2_1[2] , \wRegOut_2_1[1] , \wRegOut_2_1[0] 
        }), .Enable1(\wRegEnTop_2_1[0] ), .Enable2(\wRegEnBot_2_1[0] ), .In1({
        \wRegInTop_2_1[31] , \wRegInTop_2_1[30] , \wRegInTop_2_1[29] , 
        \wRegInTop_2_1[28] , \wRegInTop_2_1[27] , \wRegInTop_2_1[26] , 
        \wRegInTop_2_1[25] , \wRegInTop_2_1[24] , \wRegInTop_2_1[23] , 
        \wRegInTop_2_1[22] , \wRegInTop_2_1[21] , \wRegInTop_2_1[20] , 
        \wRegInTop_2_1[19] , \wRegInTop_2_1[18] , \wRegInTop_2_1[17] , 
        \wRegInTop_2_1[16] , \wRegInTop_2_1[15] , \wRegInTop_2_1[14] , 
        \wRegInTop_2_1[13] , \wRegInTop_2_1[12] , \wRegInTop_2_1[11] , 
        \wRegInTop_2_1[10] , \wRegInTop_2_1[9] , \wRegInTop_2_1[8] , 
        \wRegInTop_2_1[7] , \wRegInTop_2_1[6] , \wRegInTop_2_1[5] , 
        \wRegInTop_2_1[4] , \wRegInTop_2_1[3] , \wRegInTop_2_1[2] , 
        \wRegInTop_2_1[1] , \wRegInTop_2_1[0] }), .In2({\wRegInBot_2_1[31] , 
        \wRegInBot_2_1[30] , \wRegInBot_2_1[29] , \wRegInBot_2_1[28] , 
        \wRegInBot_2_1[27] , \wRegInBot_2_1[26] , \wRegInBot_2_1[25] , 
        \wRegInBot_2_1[24] , \wRegInBot_2_1[23] , \wRegInBot_2_1[22] , 
        \wRegInBot_2_1[21] , \wRegInBot_2_1[20] , \wRegInBot_2_1[19] , 
        \wRegInBot_2_1[18] , \wRegInBot_2_1[17] , \wRegInBot_2_1[16] , 
        \wRegInBot_2_1[15] , \wRegInBot_2_1[14] , \wRegInBot_2_1[13] , 
        \wRegInBot_2_1[12] , \wRegInBot_2_1[11] , \wRegInBot_2_1[10] , 
        \wRegInBot_2_1[9] , \wRegInBot_2_1[8] , \wRegInBot_2_1[7] , 
        \wRegInBot_2_1[6] , \wRegInBot_2_1[5] , \wRegInBot_2_1[4] , 
        \wRegInBot_2_1[3] , \wRegInBot_2_1[2] , \wRegInBot_2_1[1] , 
        \wRegInBot_2_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink9[31] , \ScanLink9[30] , \ScanLink9[29] , 
        \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , \ScanLink9[25] , 
        \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , \ScanLink9[21] , 
        \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , \ScanLink9[17] , 
        \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , \ScanLink9[13] , 
        \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , \ScanLink9[9] , 
        \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , \ScanLink9[5] , 
        \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , \ScanLink9[1] , 
        \ScanLink9[0] }), .ScanOut({\ScanLink8[31] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , 
        \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , 
        \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , 
        \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , 
        \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , 
        \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_1[31] , \wRegOut_3_1[30] , \wRegOut_3_1[29] , 
        \wRegOut_3_1[28] , \wRegOut_3_1[27] , \wRegOut_3_1[26] , 
        \wRegOut_3_1[25] , \wRegOut_3_1[24] , \wRegOut_3_1[23] , 
        \wRegOut_3_1[22] , \wRegOut_3_1[21] , \wRegOut_3_1[20] , 
        \wRegOut_3_1[19] , \wRegOut_3_1[18] , \wRegOut_3_1[17] , 
        \wRegOut_3_1[16] , \wRegOut_3_1[15] , \wRegOut_3_1[14] , 
        \wRegOut_3_1[13] , \wRegOut_3_1[12] , \wRegOut_3_1[11] , 
        \wRegOut_3_1[10] , \wRegOut_3_1[9] , \wRegOut_3_1[8] , 
        \wRegOut_3_1[7] , \wRegOut_3_1[6] , \wRegOut_3_1[5] , \wRegOut_3_1[4] , 
        \wRegOut_3_1[3] , \wRegOut_3_1[2] , \wRegOut_3_1[1] , \wRegOut_3_1[0] 
        }), .Enable1(\wRegEnTop_3_1[0] ), .Enable2(\wRegEnBot_3_1[0] ), .In1({
        \wRegInTop_3_1[31] , \wRegInTop_3_1[30] , \wRegInTop_3_1[29] , 
        \wRegInTop_3_1[28] , \wRegInTop_3_1[27] , \wRegInTop_3_1[26] , 
        \wRegInTop_3_1[25] , \wRegInTop_3_1[24] , \wRegInTop_3_1[23] , 
        \wRegInTop_3_1[22] , \wRegInTop_3_1[21] , \wRegInTop_3_1[20] , 
        \wRegInTop_3_1[19] , \wRegInTop_3_1[18] , \wRegInTop_3_1[17] , 
        \wRegInTop_3_1[16] , \wRegInTop_3_1[15] , \wRegInTop_3_1[14] , 
        \wRegInTop_3_1[13] , \wRegInTop_3_1[12] , \wRegInTop_3_1[11] , 
        \wRegInTop_3_1[10] , \wRegInTop_3_1[9] , \wRegInTop_3_1[8] , 
        \wRegInTop_3_1[7] , \wRegInTop_3_1[6] , \wRegInTop_3_1[5] , 
        \wRegInTop_3_1[4] , \wRegInTop_3_1[3] , \wRegInTop_3_1[2] , 
        \wRegInTop_3_1[1] , \wRegInTop_3_1[0] }), .In2({\wRegInBot_3_1[31] , 
        \wRegInBot_3_1[30] , \wRegInBot_3_1[29] , \wRegInBot_3_1[28] , 
        \wRegInBot_3_1[27] , \wRegInBot_3_1[26] , \wRegInBot_3_1[25] , 
        \wRegInBot_3_1[24] , \wRegInBot_3_1[23] , \wRegInBot_3_1[22] , 
        \wRegInBot_3_1[21] , \wRegInBot_3_1[20] , \wRegInBot_3_1[19] , 
        \wRegInBot_3_1[18] , \wRegInBot_3_1[17] , \wRegInBot_3_1[16] , 
        \wRegInBot_3_1[15] , \wRegInBot_3_1[14] , \wRegInBot_3_1[13] , 
        \wRegInBot_3_1[12] , \wRegInBot_3_1[11] , \wRegInBot_3_1[10] , 
        \wRegInBot_3_1[9] , \wRegInBot_3_1[8] , \wRegInBot_3_1[7] , 
        \wRegInBot_3_1[6] , \wRegInBot_3_1[5] , \wRegInBot_3_1[4] , 
        \wRegInBot_3_1[3] , \wRegInBot_3_1[2] , \wRegInBot_3_1[1] , 
        \wRegInBot_3_1[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink14[31] , \ScanLink14[30] , \ScanLink14[29] , 
        \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , \ScanLink14[25] , 
        \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , \ScanLink14[21] , 
        \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , \ScanLink14[17] , 
        \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , \ScanLink14[13] , 
        \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , \ScanLink14[9] , 
        \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , \ScanLink14[5] , 
        \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , \ScanLink14[1] , 
        \ScanLink14[0] }), .ScanOut({\ScanLink13[31] , \ScanLink13[30] , 
        \ScanLink13[29] , \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , 
        \ScanLink13[25] , \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , 
        \ScanLink13[21] , \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , 
        \ScanLink13[17] , \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , 
        \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , 
        \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , 
        \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , 
        \ScanLink13[1] , \ScanLink13[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_6[31] , \wRegOut_3_6[30] , \wRegOut_3_6[29] , 
        \wRegOut_3_6[28] , \wRegOut_3_6[27] , \wRegOut_3_6[26] , 
        \wRegOut_3_6[25] , \wRegOut_3_6[24] , \wRegOut_3_6[23] , 
        \wRegOut_3_6[22] , \wRegOut_3_6[21] , \wRegOut_3_6[20] , 
        \wRegOut_3_6[19] , \wRegOut_3_6[18] , \wRegOut_3_6[17] , 
        \wRegOut_3_6[16] , \wRegOut_3_6[15] , \wRegOut_3_6[14] , 
        \wRegOut_3_6[13] , \wRegOut_3_6[12] , \wRegOut_3_6[11] , 
        \wRegOut_3_6[10] , \wRegOut_3_6[9] , \wRegOut_3_6[8] , 
        \wRegOut_3_6[7] , \wRegOut_3_6[6] , \wRegOut_3_6[5] , \wRegOut_3_6[4] , 
        \wRegOut_3_6[3] , \wRegOut_3_6[2] , \wRegOut_3_6[1] , \wRegOut_3_6[0] 
        }), .Enable1(\wRegEnTop_3_6[0] ), .Enable2(\wRegEnBot_3_6[0] ), .In1({
        \wRegInTop_3_6[31] , \wRegInTop_3_6[30] , \wRegInTop_3_6[29] , 
        \wRegInTop_3_6[28] , \wRegInTop_3_6[27] , \wRegInTop_3_6[26] , 
        \wRegInTop_3_6[25] , \wRegInTop_3_6[24] , \wRegInTop_3_6[23] , 
        \wRegInTop_3_6[22] , \wRegInTop_3_6[21] , \wRegInTop_3_6[20] , 
        \wRegInTop_3_6[19] , \wRegInTop_3_6[18] , \wRegInTop_3_6[17] , 
        \wRegInTop_3_6[16] , \wRegInTop_3_6[15] , \wRegInTop_3_6[14] , 
        \wRegInTop_3_6[13] , \wRegInTop_3_6[12] , \wRegInTop_3_6[11] , 
        \wRegInTop_3_6[10] , \wRegInTop_3_6[9] , \wRegInTop_3_6[8] , 
        \wRegInTop_3_6[7] , \wRegInTop_3_6[6] , \wRegInTop_3_6[5] , 
        \wRegInTop_3_6[4] , \wRegInTop_3_6[3] , \wRegInTop_3_6[2] , 
        \wRegInTop_3_6[1] , \wRegInTop_3_6[0] }), .In2({\wRegInBot_3_6[31] , 
        \wRegInBot_3_6[30] , \wRegInBot_3_6[29] , \wRegInBot_3_6[28] , 
        \wRegInBot_3_6[27] , \wRegInBot_3_6[26] , \wRegInBot_3_6[25] , 
        \wRegInBot_3_6[24] , \wRegInBot_3_6[23] , \wRegInBot_3_6[22] , 
        \wRegInBot_3_6[21] , \wRegInBot_3_6[20] , \wRegInBot_3_6[19] , 
        \wRegInBot_3_6[18] , \wRegInBot_3_6[17] , \wRegInBot_3_6[16] , 
        \wRegInBot_3_6[15] , \wRegInBot_3_6[14] , \wRegInBot_3_6[13] , 
        \wRegInBot_3_6[12] , \wRegInBot_3_6[11] , \wRegInBot_3_6[10] , 
        \wRegInBot_3_6[9] , \wRegInBot_3_6[8] , \wRegInBot_3_6[7] , 
        \wRegInBot_3_6[6] , \wRegInBot_3_6[5] , \wRegInBot_3_6[4] , 
        \wRegInBot_3_6[3] , \wRegInBot_3_6[2] , \wRegInBot_3_6[1] , 
        \wRegInBot_3_6[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink29[31] , \ScanLink29[30] , \ScanLink29[29] , 
        \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , \ScanLink29[25] , 
        \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , \ScanLink29[21] , 
        \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , \ScanLink29[17] , 
        \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , \ScanLink29[13] , 
        \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , \ScanLink29[9] , 
        \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , \ScanLink29[5] , 
        \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , \ScanLink29[1] , 
        \ScanLink29[0] }), .ScanOut({\ScanLink28[31] , \ScanLink28[30] , 
        \ScanLink28[29] , \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , 
        \ScanLink28[25] , \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , 
        \ScanLink28[21] , \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , 
        \ScanLink28[17] , \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , 
        \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , 
        \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , 
        \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , 
        \ScanLink28[1] , \ScanLink28[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_13[31] , \wRegOut_4_13[30] , 
        \wRegOut_4_13[29] , \wRegOut_4_13[28] , \wRegOut_4_13[27] , 
        \wRegOut_4_13[26] , \wRegOut_4_13[25] , \wRegOut_4_13[24] , 
        \wRegOut_4_13[23] , \wRegOut_4_13[22] , \wRegOut_4_13[21] , 
        \wRegOut_4_13[20] , \wRegOut_4_13[19] , \wRegOut_4_13[18] , 
        \wRegOut_4_13[17] , \wRegOut_4_13[16] , \wRegOut_4_13[15] , 
        \wRegOut_4_13[14] , \wRegOut_4_13[13] , \wRegOut_4_13[12] , 
        \wRegOut_4_13[11] , \wRegOut_4_13[10] , \wRegOut_4_13[9] , 
        \wRegOut_4_13[8] , \wRegOut_4_13[7] , \wRegOut_4_13[6] , 
        \wRegOut_4_13[5] , \wRegOut_4_13[4] , \wRegOut_4_13[3] , 
        \wRegOut_4_13[2] , \wRegOut_4_13[1] , \wRegOut_4_13[0] }), .Enable1(
        \wRegEnTop_4_13[0] ), .Enable2(\wRegEnBot_4_13[0] ), .In1({
        \wRegInTop_4_13[31] , \wRegInTop_4_13[30] , \wRegInTop_4_13[29] , 
        \wRegInTop_4_13[28] , \wRegInTop_4_13[27] , \wRegInTop_4_13[26] , 
        \wRegInTop_4_13[25] , \wRegInTop_4_13[24] , \wRegInTop_4_13[23] , 
        \wRegInTop_4_13[22] , \wRegInTop_4_13[21] , \wRegInTop_4_13[20] , 
        \wRegInTop_4_13[19] , \wRegInTop_4_13[18] , \wRegInTop_4_13[17] , 
        \wRegInTop_4_13[16] , \wRegInTop_4_13[15] , \wRegInTop_4_13[14] , 
        \wRegInTop_4_13[13] , \wRegInTop_4_13[12] , \wRegInTop_4_13[11] , 
        \wRegInTop_4_13[10] , \wRegInTop_4_13[9] , \wRegInTop_4_13[8] , 
        \wRegInTop_4_13[7] , \wRegInTop_4_13[6] , \wRegInTop_4_13[5] , 
        \wRegInTop_4_13[4] , \wRegInTop_4_13[3] , \wRegInTop_4_13[2] , 
        \wRegInTop_4_13[1] , \wRegInTop_4_13[0] }), .In2({\wRegInBot_4_13[31] , 
        \wRegInBot_4_13[30] , \wRegInBot_4_13[29] , \wRegInBot_4_13[28] , 
        \wRegInBot_4_13[27] , \wRegInBot_4_13[26] , \wRegInBot_4_13[25] , 
        \wRegInBot_4_13[24] , \wRegInBot_4_13[23] , \wRegInBot_4_13[22] , 
        \wRegInBot_4_13[21] , \wRegInBot_4_13[20] , \wRegInBot_4_13[19] , 
        \wRegInBot_4_13[18] , \wRegInBot_4_13[17] , \wRegInBot_4_13[16] , 
        \wRegInBot_4_13[15] , \wRegInBot_4_13[14] , \wRegInBot_4_13[13] , 
        \wRegInBot_4_13[12] , \wRegInBot_4_13[11] , \wRegInBot_4_13[10] , 
        \wRegInBot_4_13[9] , \wRegInBot_4_13[8] , \wRegInBot_4_13[7] , 
        \wRegInBot_4_13[6] , \wRegInBot_4_13[5] , \wRegInBot_4_13[4] , 
        \wRegInBot_4_13[3] , \wRegInBot_4_13[2] , \wRegInBot_4_13[1] , 
        \wRegInBot_4_13[0] }) );
    BHeap_Node_WIDTH32 BHN_4_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_5[0] ), .P_In({\wRegOut_4_5[31] , 
        \wRegOut_4_5[30] , \wRegOut_4_5[29] , \wRegOut_4_5[28] , 
        \wRegOut_4_5[27] , \wRegOut_4_5[26] , \wRegOut_4_5[25] , 
        \wRegOut_4_5[24] , \wRegOut_4_5[23] , \wRegOut_4_5[22] , 
        \wRegOut_4_5[21] , \wRegOut_4_5[20] , \wRegOut_4_5[19] , 
        \wRegOut_4_5[18] , \wRegOut_4_5[17] , \wRegOut_4_5[16] , 
        \wRegOut_4_5[15] , \wRegOut_4_5[14] , \wRegOut_4_5[13] , 
        \wRegOut_4_5[12] , \wRegOut_4_5[11] , \wRegOut_4_5[10] , 
        \wRegOut_4_5[9] , \wRegOut_4_5[8] , \wRegOut_4_5[7] , \wRegOut_4_5[6] , 
        \wRegOut_4_5[5] , \wRegOut_4_5[4] , \wRegOut_4_5[3] , \wRegOut_4_5[2] , 
        \wRegOut_4_5[1] , \wRegOut_4_5[0] }), .P_Out({\wRegInBot_4_5[31] , 
        \wRegInBot_4_5[30] , \wRegInBot_4_5[29] , \wRegInBot_4_5[28] , 
        \wRegInBot_4_5[27] , \wRegInBot_4_5[26] , \wRegInBot_4_5[25] , 
        \wRegInBot_4_5[24] , \wRegInBot_4_5[23] , \wRegInBot_4_5[22] , 
        \wRegInBot_4_5[21] , \wRegInBot_4_5[20] , \wRegInBot_4_5[19] , 
        \wRegInBot_4_5[18] , \wRegInBot_4_5[17] , \wRegInBot_4_5[16] , 
        \wRegInBot_4_5[15] , \wRegInBot_4_5[14] , \wRegInBot_4_5[13] , 
        \wRegInBot_4_5[12] , \wRegInBot_4_5[11] , \wRegInBot_4_5[10] , 
        \wRegInBot_4_5[9] , \wRegInBot_4_5[8] , \wRegInBot_4_5[7] , 
        \wRegInBot_4_5[6] , \wRegInBot_4_5[5] , \wRegInBot_4_5[4] , 
        \wRegInBot_4_5[3] , \wRegInBot_4_5[2] , \wRegInBot_4_5[1] , 
        \wRegInBot_4_5[0] }), .L_WR(\wRegEnTop_5_10[0] ), .L_In({
        \wRegOut_5_10[31] , \wRegOut_5_10[30] , \wRegOut_5_10[29] , 
        \wRegOut_5_10[28] , \wRegOut_5_10[27] , \wRegOut_5_10[26] , 
        \wRegOut_5_10[25] , \wRegOut_5_10[24] , \wRegOut_5_10[23] , 
        \wRegOut_5_10[22] , \wRegOut_5_10[21] , \wRegOut_5_10[20] , 
        \wRegOut_5_10[19] , \wRegOut_5_10[18] , \wRegOut_5_10[17] , 
        \wRegOut_5_10[16] , \wRegOut_5_10[15] , \wRegOut_5_10[14] , 
        \wRegOut_5_10[13] , \wRegOut_5_10[12] , \wRegOut_5_10[11] , 
        \wRegOut_5_10[10] , \wRegOut_5_10[9] , \wRegOut_5_10[8] , 
        \wRegOut_5_10[7] , \wRegOut_5_10[6] , \wRegOut_5_10[5] , 
        \wRegOut_5_10[4] , \wRegOut_5_10[3] , \wRegOut_5_10[2] , 
        \wRegOut_5_10[1] , \wRegOut_5_10[0] }), .L_Out({\wRegInTop_5_10[31] , 
        \wRegInTop_5_10[30] , \wRegInTop_5_10[29] , \wRegInTop_5_10[28] , 
        \wRegInTop_5_10[27] , \wRegInTop_5_10[26] , \wRegInTop_5_10[25] , 
        \wRegInTop_5_10[24] , \wRegInTop_5_10[23] , \wRegInTop_5_10[22] , 
        \wRegInTop_5_10[21] , \wRegInTop_5_10[20] , \wRegInTop_5_10[19] , 
        \wRegInTop_5_10[18] , \wRegInTop_5_10[17] , \wRegInTop_5_10[16] , 
        \wRegInTop_5_10[15] , \wRegInTop_5_10[14] , \wRegInTop_5_10[13] , 
        \wRegInTop_5_10[12] , \wRegInTop_5_10[11] , \wRegInTop_5_10[10] , 
        \wRegInTop_5_10[9] , \wRegInTop_5_10[8] , \wRegInTop_5_10[7] , 
        \wRegInTop_5_10[6] , \wRegInTop_5_10[5] , \wRegInTop_5_10[4] , 
        \wRegInTop_5_10[3] , \wRegInTop_5_10[2] , \wRegInTop_5_10[1] , 
        \wRegInTop_5_10[0] }), .R_WR(\wRegEnTop_5_11[0] ), .R_In({
        \wRegOut_5_11[31] , \wRegOut_5_11[30] , \wRegOut_5_11[29] , 
        \wRegOut_5_11[28] , \wRegOut_5_11[27] , \wRegOut_5_11[26] , 
        \wRegOut_5_11[25] , \wRegOut_5_11[24] , \wRegOut_5_11[23] , 
        \wRegOut_5_11[22] , \wRegOut_5_11[21] , \wRegOut_5_11[20] , 
        \wRegOut_5_11[19] , \wRegOut_5_11[18] , \wRegOut_5_11[17] , 
        \wRegOut_5_11[16] , \wRegOut_5_11[15] , \wRegOut_5_11[14] , 
        \wRegOut_5_11[13] , \wRegOut_5_11[12] , \wRegOut_5_11[11] , 
        \wRegOut_5_11[10] , \wRegOut_5_11[9] , \wRegOut_5_11[8] , 
        \wRegOut_5_11[7] , \wRegOut_5_11[6] , \wRegOut_5_11[5] , 
        \wRegOut_5_11[4] , \wRegOut_5_11[3] , \wRegOut_5_11[2] , 
        \wRegOut_5_11[1] , \wRegOut_5_11[0] }), .R_Out({\wRegInTop_5_11[31] , 
        \wRegInTop_5_11[30] , \wRegInTop_5_11[29] , \wRegInTop_5_11[28] , 
        \wRegInTop_5_11[27] , \wRegInTop_5_11[26] , \wRegInTop_5_11[25] , 
        \wRegInTop_5_11[24] , \wRegInTop_5_11[23] , \wRegInTop_5_11[22] , 
        \wRegInTop_5_11[21] , \wRegInTop_5_11[20] , \wRegInTop_5_11[19] , 
        \wRegInTop_5_11[18] , \wRegInTop_5_11[17] , \wRegInTop_5_11[16] , 
        \wRegInTop_5_11[15] , \wRegInTop_5_11[14] , \wRegInTop_5_11[13] , 
        \wRegInTop_5_11[12] , \wRegInTop_5_11[11] , \wRegInTop_5_11[10] , 
        \wRegInTop_5_11[9] , \wRegInTop_5_11[8] , \wRegInTop_5_11[7] , 
        \wRegInTop_5_11[6] , \wRegInTop_5_11[5] , \wRegInTop_5_11[4] , 
        \wRegInTop_5_11[3] , \wRegInTop_5_11[2] , \wRegInTop_5_11[1] , 
        \wRegInTop_5_11[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink39[31] , \ScanLink39[30] , \ScanLink39[29] , 
        \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , \ScanLink39[25] , 
        \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , \ScanLink39[21] , 
        \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , \ScanLink39[17] , 
        \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , \ScanLink39[13] , 
        \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , \ScanLink39[9] , 
        \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , \ScanLink39[5] , 
        \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , \ScanLink39[1] , 
        \ScanLink39[0] }), .ScanOut({\ScanLink38[31] , \ScanLink38[30] , 
        \ScanLink38[29] , \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , 
        \ScanLink38[25] , \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , 
        \ScanLink38[21] , \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , 
        \ScanLink38[17] , \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , 
        \ScanLink38[13] , \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , 
        \ScanLink38[9] , \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , 
        \ScanLink38[5] , \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , 
        \ScanLink38[1] , \ScanLink38[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_7[31] , \wRegOut_5_7[30] , \wRegOut_5_7[29] , 
        \wRegOut_5_7[28] , \wRegOut_5_7[27] , \wRegOut_5_7[26] , 
        \wRegOut_5_7[25] , \wRegOut_5_7[24] , \wRegOut_5_7[23] , 
        \wRegOut_5_7[22] , \wRegOut_5_7[21] , \wRegOut_5_7[20] , 
        \wRegOut_5_7[19] , \wRegOut_5_7[18] , \wRegOut_5_7[17] , 
        \wRegOut_5_7[16] , \wRegOut_5_7[15] , \wRegOut_5_7[14] , 
        \wRegOut_5_7[13] , \wRegOut_5_7[12] , \wRegOut_5_7[11] , 
        \wRegOut_5_7[10] , \wRegOut_5_7[9] , \wRegOut_5_7[8] , 
        \wRegOut_5_7[7] , \wRegOut_5_7[6] , \wRegOut_5_7[5] , \wRegOut_5_7[4] , 
        \wRegOut_5_7[3] , \wRegOut_5_7[2] , \wRegOut_5_7[1] , \wRegOut_5_7[0] 
        }), .Enable1(\wRegEnTop_5_7[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_7[31] , \wRegInTop_5_7[30] , \wRegInTop_5_7[29] , 
        \wRegInTop_5_7[28] , \wRegInTop_5_7[27] , \wRegInTop_5_7[26] , 
        \wRegInTop_5_7[25] , \wRegInTop_5_7[24] , \wRegInTop_5_7[23] , 
        \wRegInTop_5_7[22] , \wRegInTop_5_7[21] , \wRegInTop_5_7[20] , 
        \wRegInTop_5_7[19] , \wRegInTop_5_7[18] , \wRegInTop_5_7[17] , 
        \wRegInTop_5_7[16] , \wRegInTop_5_7[15] , \wRegInTop_5_7[14] , 
        \wRegInTop_5_7[13] , \wRegInTop_5_7[12] , \wRegInTop_5_7[11] , 
        \wRegInTop_5_7[10] , \wRegInTop_5_7[9] , \wRegInTop_5_7[8] , 
        \wRegInTop_5_7[7] , \wRegInTop_5_7[6] , \wRegInTop_5_7[5] , 
        \wRegInTop_5_7[4] , \wRegInTop_5_7[3] , \wRegInTop_5_7[2] , 
        \wRegInTop_5_7[1] , \wRegInTop_5_7[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_19 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink51[31] , \ScanLink51[30] , \ScanLink51[29] , 
        \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , \ScanLink51[25] , 
        \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , \ScanLink51[21] , 
        \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , \ScanLink51[17] , 
        \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , \ScanLink51[13] , 
        \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , \ScanLink51[9] , 
        \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , \ScanLink51[5] , 
        \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , \ScanLink51[1] , 
        \ScanLink51[0] }), .ScanOut({\ScanLink50[31] , \ScanLink50[30] , 
        \ScanLink50[29] , \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , 
        \ScanLink50[25] , \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , 
        \ScanLink50[21] , \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , 
        \ScanLink50[17] , \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , 
        \ScanLink50[13] , \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , 
        \ScanLink50[9] , \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , 
        \ScanLink50[5] , \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , 
        \ScanLink50[1] , \ScanLink50[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_19[31] , \wRegOut_5_19[30] , 
        \wRegOut_5_19[29] , \wRegOut_5_19[28] , \wRegOut_5_19[27] , 
        \wRegOut_5_19[26] , \wRegOut_5_19[25] , \wRegOut_5_19[24] , 
        \wRegOut_5_19[23] , \wRegOut_5_19[22] , \wRegOut_5_19[21] , 
        \wRegOut_5_19[20] , \wRegOut_5_19[19] , \wRegOut_5_19[18] , 
        \wRegOut_5_19[17] , \wRegOut_5_19[16] , \wRegOut_5_19[15] , 
        \wRegOut_5_19[14] , \wRegOut_5_19[13] , \wRegOut_5_19[12] , 
        \wRegOut_5_19[11] , \wRegOut_5_19[10] , \wRegOut_5_19[9] , 
        \wRegOut_5_19[8] , \wRegOut_5_19[7] , \wRegOut_5_19[6] , 
        \wRegOut_5_19[5] , \wRegOut_5_19[4] , \wRegOut_5_19[3] , 
        \wRegOut_5_19[2] , \wRegOut_5_19[1] , \wRegOut_5_19[0] }), .Enable1(
        \wRegEnTop_5_19[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_19[31] , 
        \wRegInTop_5_19[30] , \wRegInTop_5_19[29] , \wRegInTop_5_19[28] , 
        \wRegInTop_5_19[27] , \wRegInTop_5_19[26] , \wRegInTop_5_19[25] , 
        \wRegInTop_5_19[24] , \wRegInTop_5_19[23] , \wRegInTop_5_19[22] , 
        \wRegInTop_5_19[21] , \wRegInTop_5_19[20] , \wRegInTop_5_19[19] , 
        \wRegInTop_5_19[18] , \wRegInTop_5_19[17] , \wRegInTop_5_19[16] , 
        \wRegInTop_5_19[15] , \wRegInTop_5_19[14] , \wRegInTop_5_19[13] , 
        \wRegInTop_5_19[12] , \wRegInTop_5_19[11] , \wRegInTop_5_19[10] , 
        \wRegInTop_5_19[9] , \wRegInTop_5_19[8] , \wRegInTop_5_19[7] , 
        \wRegInTop_5_19[6] , \wRegInTop_5_19[5] , \wRegInTop_5_19[4] , 
        \wRegInTop_5_19[3] , \wRegInTop_5_19[2] , \wRegInTop_5_19[1] , 
        \wRegInTop_5_19[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_25 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink57[31] , \ScanLink57[30] , \ScanLink57[29] , 
        \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , \ScanLink57[25] , 
        \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , \ScanLink57[21] , 
        \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , \ScanLink57[17] , 
        \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , \ScanLink57[13] , 
        \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , \ScanLink57[9] , 
        \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , \ScanLink57[5] , 
        \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , \ScanLink57[1] , 
        \ScanLink57[0] }), .ScanOut({\ScanLink56[31] , \ScanLink56[30] , 
        \ScanLink56[29] , \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , 
        \ScanLink56[25] , \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , 
        \ScanLink56[21] , \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , 
        \ScanLink56[17] , \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , 
        \ScanLink56[13] , \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , 
        \ScanLink56[9] , \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , 
        \ScanLink56[5] , \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , 
        \ScanLink56[1] , \ScanLink56[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_25[31] , \wRegOut_5_25[30] , 
        \wRegOut_5_25[29] , \wRegOut_5_25[28] , \wRegOut_5_25[27] , 
        \wRegOut_5_25[26] , \wRegOut_5_25[25] , \wRegOut_5_25[24] , 
        \wRegOut_5_25[23] , \wRegOut_5_25[22] , \wRegOut_5_25[21] , 
        \wRegOut_5_25[20] , \wRegOut_5_25[19] , \wRegOut_5_25[18] , 
        \wRegOut_5_25[17] , \wRegOut_5_25[16] , \wRegOut_5_25[15] , 
        \wRegOut_5_25[14] , \wRegOut_5_25[13] , \wRegOut_5_25[12] , 
        \wRegOut_5_25[11] , \wRegOut_5_25[10] , \wRegOut_5_25[9] , 
        \wRegOut_5_25[8] , \wRegOut_5_25[7] , \wRegOut_5_25[6] , 
        \wRegOut_5_25[5] , \wRegOut_5_25[4] , \wRegOut_5_25[3] , 
        \wRegOut_5_25[2] , \wRegOut_5_25[1] , \wRegOut_5_25[0] }), .Enable1(
        \wRegEnTop_5_25[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_25[31] , 
        \wRegInTop_5_25[30] , \wRegInTop_5_25[29] , \wRegInTop_5_25[28] , 
        \wRegInTop_5_25[27] , \wRegInTop_5_25[26] , \wRegInTop_5_25[25] , 
        \wRegInTop_5_25[24] , \wRegInTop_5_25[23] , \wRegInTop_5_25[22] , 
        \wRegInTop_5_25[21] , \wRegInTop_5_25[20] , \wRegInTop_5_25[19] , 
        \wRegInTop_5_25[18] , \wRegInTop_5_25[17] , \wRegInTop_5_25[16] , 
        \wRegInTop_5_25[15] , \wRegInTop_5_25[14] , \wRegInTop_5_25[13] , 
        \wRegInTop_5_25[12] , \wRegInTop_5_25[11] , \wRegInTop_5_25[10] , 
        \wRegInTop_5_25[9] , \wRegInTop_5_25[8] , \wRegInTop_5_25[7] , 
        \wRegInTop_5_25[6] , \wRegInTop_5_25[5] , \wRegInTop_5_25[4] , 
        \wRegInTop_5_25[3] , \wRegInTop_5_25[2] , \wRegInTop_5_25[1] , 
        \wRegInTop_5_25[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_4[0] ), .P_In({\wRegOut_3_4[31] , 
        \wRegOut_3_4[30] , \wRegOut_3_4[29] , \wRegOut_3_4[28] , 
        \wRegOut_3_4[27] , \wRegOut_3_4[26] , \wRegOut_3_4[25] , 
        \wRegOut_3_4[24] , \wRegOut_3_4[23] , \wRegOut_3_4[22] , 
        \wRegOut_3_4[21] , \wRegOut_3_4[20] , \wRegOut_3_4[19] , 
        \wRegOut_3_4[18] , \wRegOut_3_4[17] , \wRegOut_3_4[16] , 
        \wRegOut_3_4[15] , \wRegOut_3_4[14] , \wRegOut_3_4[13] , 
        \wRegOut_3_4[12] , \wRegOut_3_4[11] , \wRegOut_3_4[10] , 
        \wRegOut_3_4[9] , \wRegOut_3_4[8] , \wRegOut_3_4[7] , \wRegOut_3_4[6] , 
        \wRegOut_3_4[5] , \wRegOut_3_4[4] , \wRegOut_3_4[3] , \wRegOut_3_4[2] , 
        \wRegOut_3_4[1] , \wRegOut_3_4[0] }), .P_Out({\wRegInBot_3_4[31] , 
        \wRegInBot_3_4[30] , \wRegInBot_3_4[29] , \wRegInBot_3_4[28] , 
        \wRegInBot_3_4[27] , \wRegInBot_3_4[26] , \wRegInBot_3_4[25] , 
        \wRegInBot_3_4[24] , \wRegInBot_3_4[23] , \wRegInBot_3_4[22] , 
        \wRegInBot_3_4[21] , \wRegInBot_3_4[20] , \wRegInBot_3_4[19] , 
        \wRegInBot_3_4[18] , \wRegInBot_3_4[17] , \wRegInBot_3_4[16] , 
        \wRegInBot_3_4[15] , \wRegInBot_3_4[14] , \wRegInBot_3_4[13] , 
        \wRegInBot_3_4[12] , \wRegInBot_3_4[11] , \wRegInBot_3_4[10] , 
        \wRegInBot_3_4[9] , \wRegInBot_3_4[8] , \wRegInBot_3_4[7] , 
        \wRegInBot_3_4[6] , \wRegInBot_3_4[5] , \wRegInBot_3_4[4] , 
        \wRegInBot_3_4[3] , \wRegInBot_3_4[2] , \wRegInBot_3_4[1] , 
        \wRegInBot_3_4[0] }), .L_WR(\wRegEnTop_4_8[0] ), .L_In({
        \wRegOut_4_8[31] , \wRegOut_4_8[30] , \wRegOut_4_8[29] , 
        \wRegOut_4_8[28] , \wRegOut_4_8[27] , \wRegOut_4_8[26] , 
        \wRegOut_4_8[25] , \wRegOut_4_8[24] , \wRegOut_4_8[23] , 
        \wRegOut_4_8[22] , \wRegOut_4_8[21] , \wRegOut_4_8[20] , 
        \wRegOut_4_8[19] , \wRegOut_4_8[18] , \wRegOut_4_8[17] , 
        \wRegOut_4_8[16] , \wRegOut_4_8[15] , \wRegOut_4_8[14] , 
        \wRegOut_4_8[13] , \wRegOut_4_8[12] , \wRegOut_4_8[11] , 
        \wRegOut_4_8[10] , \wRegOut_4_8[9] , \wRegOut_4_8[8] , 
        \wRegOut_4_8[7] , \wRegOut_4_8[6] , \wRegOut_4_8[5] , \wRegOut_4_8[4] , 
        \wRegOut_4_8[3] , \wRegOut_4_8[2] , \wRegOut_4_8[1] , \wRegOut_4_8[0] 
        }), .L_Out({\wRegInTop_4_8[31] , \wRegInTop_4_8[30] , 
        \wRegInTop_4_8[29] , \wRegInTop_4_8[28] , \wRegInTop_4_8[27] , 
        \wRegInTop_4_8[26] , \wRegInTop_4_8[25] , \wRegInTop_4_8[24] , 
        \wRegInTop_4_8[23] , \wRegInTop_4_8[22] , \wRegInTop_4_8[21] , 
        \wRegInTop_4_8[20] , \wRegInTop_4_8[19] , \wRegInTop_4_8[18] , 
        \wRegInTop_4_8[17] , \wRegInTop_4_8[16] , \wRegInTop_4_8[15] , 
        \wRegInTop_4_8[14] , \wRegInTop_4_8[13] , \wRegInTop_4_8[12] , 
        \wRegInTop_4_8[11] , \wRegInTop_4_8[10] , \wRegInTop_4_8[9] , 
        \wRegInTop_4_8[8] , \wRegInTop_4_8[7] , \wRegInTop_4_8[6] , 
        \wRegInTop_4_8[5] , \wRegInTop_4_8[4] , \wRegInTop_4_8[3] , 
        \wRegInTop_4_8[2] , \wRegInTop_4_8[1] , \wRegInTop_4_8[0] }), .R_WR(
        \wRegEnTop_4_9[0] ), .R_In({\wRegOut_4_9[31] , \wRegOut_4_9[30] , 
        \wRegOut_4_9[29] , \wRegOut_4_9[28] , \wRegOut_4_9[27] , 
        \wRegOut_4_9[26] , \wRegOut_4_9[25] , \wRegOut_4_9[24] , 
        \wRegOut_4_9[23] , \wRegOut_4_9[22] , \wRegOut_4_9[21] , 
        \wRegOut_4_9[20] , \wRegOut_4_9[19] , \wRegOut_4_9[18] , 
        \wRegOut_4_9[17] , \wRegOut_4_9[16] , \wRegOut_4_9[15] , 
        \wRegOut_4_9[14] , \wRegOut_4_9[13] , \wRegOut_4_9[12] , 
        \wRegOut_4_9[11] , \wRegOut_4_9[10] , \wRegOut_4_9[9] , 
        \wRegOut_4_9[8] , \wRegOut_4_9[7] , \wRegOut_4_9[6] , \wRegOut_4_9[5] , 
        \wRegOut_4_9[4] , \wRegOut_4_9[3] , \wRegOut_4_9[2] , \wRegOut_4_9[1] , 
        \wRegOut_4_9[0] }), .R_Out({\wRegInTop_4_9[31] , \wRegInTop_4_9[30] , 
        \wRegInTop_4_9[29] , \wRegInTop_4_9[28] , \wRegInTop_4_9[27] , 
        \wRegInTop_4_9[26] , \wRegInTop_4_9[25] , \wRegInTop_4_9[24] , 
        \wRegInTop_4_9[23] , \wRegInTop_4_9[22] , \wRegInTop_4_9[21] , 
        \wRegInTop_4_9[20] , \wRegInTop_4_9[19] , \wRegInTop_4_9[18] , 
        \wRegInTop_4_9[17] , \wRegInTop_4_9[16] , \wRegInTop_4_9[15] , 
        \wRegInTop_4_9[14] , \wRegInTop_4_9[13] , \wRegInTop_4_9[12] , 
        \wRegInTop_4_9[11] , \wRegInTop_4_9[10] , \wRegInTop_4_9[9] , 
        \wRegInTop_4_9[8] , \wRegInTop_4_9[7] , \wRegInTop_4_9[6] , 
        \wRegInTop_4_9[5] , \wRegInTop_4_9[4] , \wRegInTop_4_9[3] , 
        \wRegInTop_4_9[2] , \wRegInTop_4_9[1] , \wRegInTop_4_9[0] }) );
    BHeap_CtrlReg_WIDTH32 BHCR_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_1[0] ), 
        .Out(\wCtrlOut_0[0] ), .Enable(\wEnable_0[0] ) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink18[31] , \ScanLink18[30] , \ScanLink18[29] , 
        \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , \ScanLink18[25] , 
        \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , \ScanLink18[21] , 
        \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , \ScanLink18[17] , 
        \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , \ScanLink18[13] , 
        \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , \ScanLink18[9] , 
        \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , \ScanLink18[5] , 
        \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , \ScanLink18[1] , 
        \ScanLink18[0] }), .ScanOut({\ScanLink17[31] , \ScanLink17[30] , 
        \ScanLink17[29] , \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , 
        \ScanLink17[25] , \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , 
        \ScanLink17[21] , \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , 
        \ScanLink17[17] , \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , 
        \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , 
        \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , 
        \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , 
        \ScanLink17[1] , \ScanLink17[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_2[31] , \wRegOut_4_2[30] , \wRegOut_4_2[29] , 
        \wRegOut_4_2[28] , \wRegOut_4_2[27] , \wRegOut_4_2[26] , 
        \wRegOut_4_2[25] , \wRegOut_4_2[24] , \wRegOut_4_2[23] , 
        \wRegOut_4_2[22] , \wRegOut_4_2[21] , \wRegOut_4_2[20] , 
        \wRegOut_4_2[19] , \wRegOut_4_2[18] , \wRegOut_4_2[17] , 
        \wRegOut_4_2[16] , \wRegOut_4_2[15] , \wRegOut_4_2[14] , 
        \wRegOut_4_2[13] , \wRegOut_4_2[12] , \wRegOut_4_2[11] , 
        \wRegOut_4_2[10] , \wRegOut_4_2[9] , \wRegOut_4_2[8] , 
        \wRegOut_4_2[7] , \wRegOut_4_2[6] , \wRegOut_4_2[5] , \wRegOut_4_2[4] , 
        \wRegOut_4_2[3] , \wRegOut_4_2[2] , \wRegOut_4_2[1] , \wRegOut_4_2[0] 
        }), .Enable1(\wRegEnTop_4_2[0] ), .Enable2(\wRegEnBot_4_2[0] ), .In1({
        \wRegInTop_4_2[31] , \wRegInTop_4_2[30] , \wRegInTop_4_2[29] , 
        \wRegInTop_4_2[28] , \wRegInTop_4_2[27] , \wRegInTop_4_2[26] , 
        \wRegInTop_4_2[25] , \wRegInTop_4_2[24] , \wRegInTop_4_2[23] , 
        \wRegInTop_4_2[22] , \wRegInTop_4_2[21] , \wRegInTop_4_2[20] , 
        \wRegInTop_4_2[19] , \wRegInTop_4_2[18] , \wRegInTop_4_2[17] , 
        \wRegInTop_4_2[16] , \wRegInTop_4_2[15] , \wRegInTop_4_2[14] , 
        \wRegInTop_4_2[13] , \wRegInTop_4_2[12] , \wRegInTop_4_2[11] , 
        \wRegInTop_4_2[10] , \wRegInTop_4_2[9] , \wRegInTop_4_2[8] , 
        \wRegInTop_4_2[7] , \wRegInTop_4_2[6] , \wRegInTop_4_2[5] , 
        \wRegInTop_4_2[4] , \wRegInTop_4_2[3] , \wRegInTop_4_2[2] , 
        \wRegInTop_4_2[1] , \wRegInTop_4_2[0] }), .In2({\wRegInBot_4_2[31] , 
        \wRegInBot_4_2[30] , \wRegInBot_4_2[29] , \wRegInBot_4_2[28] , 
        \wRegInBot_4_2[27] , \wRegInBot_4_2[26] , \wRegInBot_4_2[25] , 
        \wRegInBot_4_2[24] , \wRegInBot_4_2[23] , \wRegInBot_4_2[22] , 
        \wRegInBot_4_2[21] , \wRegInBot_4_2[20] , \wRegInBot_4_2[19] , 
        \wRegInBot_4_2[18] , \wRegInBot_4_2[17] , \wRegInBot_4_2[16] , 
        \wRegInBot_4_2[15] , \wRegInBot_4_2[14] , \wRegInBot_4_2[13] , 
        \wRegInBot_4_2[12] , \wRegInBot_4_2[11] , \wRegInBot_4_2[10] , 
        \wRegInBot_4_2[9] , \wRegInBot_4_2[8] , \wRegInBot_4_2[7] , 
        \wRegInBot_4_2[6] , \wRegInBot_4_2[5] , \wRegInBot_4_2[4] , 
        \wRegInBot_4_2[3] , \wRegInBot_4_2[2] , \wRegInBot_4_2[1] , 
        \wRegInBot_4_2[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink21[31] , \ScanLink21[30] , \ScanLink21[29] , 
        \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , \ScanLink21[25] , 
        \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , \ScanLink21[21] , 
        \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , \ScanLink21[17] , 
        \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , \ScanLink21[13] , 
        \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , \ScanLink21[9] , 
        \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , \ScanLink21[5] , 
        \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , \ScanLink21[1] , 
        \ScanLink21[0] }), .ScanOut({\ScanLink20[31] , \ScanLink20[30] , 
        \ScanLink20[29] , \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , 
        \ScanLink20[25] , \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , 
        \ScanLink20[21] , \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , 
        \ScanLink20[17] , \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , 
        \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , 
        \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , 
        \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , 
        \ScanLink20[1] , \ScanLink20[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_5[31] , \wRegOut_4_5[30] , \wRegOut_4_5[29] , 
        \wRegOut_4_5[28] , \wRegOut_4_5[27] , \wRegOut_4_5[26] , 
        \wRegOut_4_5[25] , \wRegOut_4_5[24] , \wRegOut_4_5[23] , 
        \wRegOut_4_5[22] , \wRegOut_4_5[21] , \wRegOut_4_5[20] , 
        \wRegOut_4_5[19] , \wRegOut_4_5[18] , \wRegOut_4_5[17] , 
        \wRegOut_4_5[16] , \wRegOut_4_5[15] , \wRegOut_4_5[14] , 
        \wRegOut_4_5[13] , \wRegOut_4_5[12] , \wRegOut_4_5[11] , 
        \wRegOut_4_5[10] , \wRegOut_4_5[9] , \wRegOut_4_5[8] , 
        \wRegOut_4_5[7] , \wRegOut_4_5[6] , \wRegOut_4_5[5] , \wRegOut_4_5[4] , 
        \wRegOut_4_5[3] , \wRegOut_4_5[2] , \wRegOut_4_5[1] , \wRegOut_4_5[0] 
        }), .Enable1(\wRegEnTop_4_5[0] ), .Enable2(\wRegEnBot_4_5[0] ), .In1({
        \wRegInTop_4_5[31] , \wRegInTop_4_5[30] , \wRegInTop_4_5[29] , 
        \wRegInTop_4_5[28] , \wRegInTop_4_5[27] , \wRegInTop_4_5[26] , 
        \wRegInTop_4_5[25] , \wRegInTop_4_5[24] , \wRegInTop_4_5[23] , 
        \wRegInTop_4_5[22] , \wRegInTop_4_5[21] , \wRegInTop_4_5[20] , 
        \wRegInTop_4_5[19] , \wRegInTop_4_5[18] , \wRegInTop_4_5[17] , 
        \wRegInTop_4_5[16] , \wRegInTop_4_5[15] , \wRegInTop_4_5[14] , 
        \wRegInTop_4_5[13] , \wRegInTop_4_5[12] , \wRegInTop_4_5[11] , 
        \wRegInTop_4_5[10] , \wRegInTop_4_5[9] , \wRegInTop_4_5[8] , 
        \wRegInTop_4_5[7] , \wRegInTop_4_5[6] , \wRegInTop_4_5[5] , 
        \wRegInTop_4_5[4] , \wRegInTop_4_5[3] , \wRegInTop_4_5[2] , 
        \wRegInTop_4_5[1] , \wRegInTop_4_5[0] }), .In2({\wRegInBot_4_5[31] , 
        \wRegInBot_4_5[30] , \wRegInBot_4_5[29] , \wRegInBot_4_5[28] , 
        \wRegInBot_4_5[27] , \wRegInBot_4_5[26] , \wRegInBot_4_5[25] , 
        \wRegInBot_4_5[24] , \wRegInBot_4_5[23] , \wRegInBot_4_5[22] , 
        \wRegInBot_4_5[21] , \wRegInBot_4_5[20] , \wRegInBot_4_5[19] , 
        \wRegInBot_4_5[18] , \wRegInBot_4_5[17] , \wRegInBot_4_5[16] , 
        \wRegInBot_4_5[15] , \wRegInBot_4_5[14] , \wRegInBot_4_5[13] , 
        \wRegInBot_4_5[12] , \wRegInBot_4_5[11] , \wRegInBot_4_5[10] , 
        \wRegInBot_4_5[9] , \wRegInBot_4_5[8] , \wRegInBot_4_5[7] , 
        \wRegInBot_4_5[6] , \wRegInBot_4_5[5] , \wRegInBot_4_5[4] , 
        \wRegInBot_4_5[3] , \wRegInBot_4_5[2] , \wRegInBot_4_5[1] , 
        \wRegInBot_4_5[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink27[31] , \ScanLink27[30] , \ScanLink27[29] , 
        \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , \ScanLink27[25] , 
        \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , \ScanLink27[21] , 
        \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , \ScanLink27[17] , 
        \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , \ScanLink27[13] , 
        \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , \ScanLink27[9] , 
        \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , \ScanLink27[5] , 
        \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , \ScanLink27[1] , 
        \ScanLink27[0] }), .ScanOut({\ScanLink26[31] , \ScanLink26[30] , 
        \ScanLink26[29] , \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , 
        \ScanLink26[25] , \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , 
        \ScanLink26[21] , \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , 
        \ScanLink26[17] , \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , 
        \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , 
        \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , 
        \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , 
        \ScanLink26[1] , \ScanLink26[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_11[31] , \wRegOut_4_11[30] , 
        \wRegOut_4_11[29] , \wRegOut_4_11[28] , \wRegOut_4_11[27] , 
        \wRegOut_4_11[26] , \wRegOut_4_11[25] , \wRegOut_4_11[24] , 
        \wRegOut_4_11[23] , \wRegOut_4_11[22] , \wRegOut_4_11[21] , 
        \wRegOut_4_11[20] , \wRegOut_4_11[19] , \wRegOut_4_11[18] , 
        \wRegOut_4_11[17] , \wRegOut_4_11[16] , \wRegOut_4_11[15] , 
        \wRegOut_4_11[14] , \wRegOut_4_11[13] , \wRegOut_4_11[12] , 
        \wRegOut_4_11[11] , \wRegOut_4_11[10] , \wRegOut_4_11[9] , 
        \wRegOut_4_11[8] , \wRegOut_4_11[7] , \wRegOut_4_11[6] , 
        \wRegOut_4_11[5] , \wRegOut_4_11[4] , \wRegOut_4_11[3] , 
        \wRegOut_4_11[2] , \wRegOut_4_11[1] , \wRegOut_4_11[0] }), .Enable1(
        \wRegEnTop_4_11[0] ), .Enable2(\wRegEnBot_4_11[0] ), .In1({
        \wRegInTop_4_11[31] , \wRegInTop_4_11[30] , \wRegInTop_4_11[29] , 
        \wRegInTop_4_11[28] , \wRegInTop_4_11[27] , \wRegInTop_4_11[26] , 
        \wRegInTop_4_11[25] , \wRegInTop_4_11[24] , \wRegInTop_4_11[23] , 
        \wRegInTop_4_11[22] , \wRegInTop_4_11[21] , \wRegInTop_4_11[20] , 
        \wRegInTop_4_11[19] , \wRegInTop_4_11[18] , \wRegInTop_4_11[17] , 
        \wRegInTop_4_11[16] , \wRegInTop_4_11[15] , \wRegInTop_4_11[14] , 
        \wRegInTop_4_11[13] , \wRegInTop_4_11[12] , \wRegInTop_4_11[11] , 
        \wRegInTop_4_11[10] , \wRegInTop_4_11[9] , \wRegInTop_4_11[8] , 
        \wRegInTop_4_11[7] , \wRegInTop_4_11[6] , \wRegInTop_4_11[5] , 
        \wRegInTop_4_11[4] , \wRegInTop_4_11[3] , \wRegInTop_4_11[2] , 
        \wRegInTop_4_11[1] , \wRegInTop_4_11[0] }), .In2({\wRegInBot_4_11[31] , 
        \wRegInBot_4_11[30] , \wRegInBot_4_11[29] , \wRegInBot_4_11[28] , 
        \wRegInBot_4_11[27] , \wRegInBot_4_11[26] , \wRegInBot_4_11[25] , 
        \wRegInBot_4_11[24] , \wRegInBot_4_11[23] , \wRegInBot_4_11[22] , 
        \wRegInBot_4_11[21] , \wRegInBot_4_11[20] , \wRegInBot_4_11[19] , 
        \wRegInBot_4_11[18] , \wRegInBot_4_11[17] , \wRegInBot_4_11[16] , 
        \wRegInBot_4_11[15] , \wRegInBot_4_11[14] , \wRegInBot_4_11[13] , 
        \wRegInBot_4_11[12] , \wRegInBot_4_11[11] , \wRegInBot_4_11[10] , 
        \wRegInBot_4_11[9] , \wRegInBot_4_11[8] , \wRegInBot_4_11[7] , 
        \wRegInBot_4_11[6] , \wRegInBot_4_11[5] , \wRegInBot_4_11[4] , 
        \wRegInBot_4_11[3] , \wRegInBot_4_11[2] , \wRegInBot_4_11[1] , 
        \wRegInBot_4_11[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink37[31] , \ScanLink37[30] , \ScanLink37[29] , 
        \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , \ScanLink37[25] , 
        \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , \ScanLink37[21] , 
        \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , \ScanLink37[17] , 
        \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , \ScanLink37[13] , 
        \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , \ScanLink37[9] , 
        \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , \ScanLink37[5] , 
        \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , \ScanLink37[1] , 
        \ScanLink37[0] }), .ScanOut({\ScanLink36[31] , \ScanLink36[30] , 
        \ScanLink36[29] , \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , 
        \ScanLink36[25] , \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , 
        \ScanLink36[21] , \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , 
        \ScanLink36[17] , \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , 
        \ScanLink36[13] , \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , 
        \ScanLink36[9] , \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , 
        \ScanLink36[5] , \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , 
        \ScanLink36[1] , \ScanLink36[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_5[31] , \wRegOut_5_5[30] , \wRegOut_5_5[29] , 
        \wRegOut_5_5[28] , \wRegOut_5_5[27] , \wRegOut_5_5[26] , 
        \wRegOut_5_5[25] , \wRegOut_5_5[24] , \wRegOut_5_5[23] , 
        \wRegOut_5_5[22] , \wRegOut_5_5[21] , \wRegOut_5_5[20] , 
        \wRegOut_5_5[19] , \wRegOut_5_5[18] , \wRegOut_5_5[17] , 
        \wRegOut_5_5[16] , \wRegOut_5_5[15] , \wRegOut_5_5[14] , 
        \wRegOut_5_5[13] , \wRegOut_5_5[12] , \wRegOut_5_5[11] , 
        \wRegOut_5_5[10] , \wRegOut_5_5[9] , \wRegOut_5_5[8] , 
        \wRegOut_5_5[7] , \wRegOut_5_5[6] , \wRegOut_5_5[5] , \wRegOut_5_5[4] , 
        \wRegOut_5_5[3] , \wRegOut_5_5[2] , \wRegOut_5_5[1] , \wRegOut_5_5[0] 
        }), .Enable1(\wRegEnTop_5_5[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_5[31] , \wRegInTop_5_5[30] , \wRegInTop_5_5[29] , 
        \wRegInTop_5_5[28] , \wRegInTop_5_5[27] , \wRegInTop_5_5[26] , 
        \wRegInTop_5_5[25] , \wRegInTop_5_5[24] , \wRegInTop_5_5[23] , 
        \wRegInTop_5_5[22] , \wRegInTop_5_5[21] , \wRegInTop_5_5[20] , 
        \wRegInTop_5_5[19] , \wRegInTop_5_5[18] , \wRegInTop_5_5[17] , 
        \wRegInTop_5_5[16] , \wRegInTop_5_5[15] , \wRegInTop_5_5[14] , 
        \wRegInTop_5_5[13] , \wRegInTop_5_5[12] , \wRegInTop_5_5[11] , 
        \wRegInTop_5_5[10] , \wRegInTop_5_5[9] , \wRegInTop_5_5[8] , 
        \wRegInTop_5_5[7] , \wRegInTop_5_5[6] , \wRegInTop_5_5[5] , 
        \wRegInTop_5_5[4] , \wRegInTop_5_5[3] , \wRegInTop_5_5[2] , 
        \wRegInTop_5_5[1] , \wRegInTop_5_5[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_1[0] ), .P_WR(\wRegEnBot_1_1[0] ), .P_In({\wRegOut_1_1[31] , 
        \wRegOut_1_1[30] , \wRegOut_1_1[29] , \wRegOut_1_1[28] , 
        \wRegOut_1_1[27] , \wRegOut_1_1[26] , \wRegOut_1_1[25] , 
        \wRegOut_1_1[24] , \wRegOut_1_1[23] , \wRegOut_1_1[22] , 
        \wRegOut_1_1[21] , \wRegOut_1_1[20] , \wRegOut_1_1[19] , 
        \wRegOut_1_1[18] , \wRegOut_1_1[17] , \wRegOut_1_1[16] , 
        \wRegOut_1_1[15] , \wRegOut_1_1[14] , \wRegOut_1_1[13] , 
        \wRegOut_1_1[12] , \wRegOut_1_1[11] , \wRegOut_1_1[10] , 
        \wRegOut_1_1[9] , \wRegOut_1_1[8] , \wRegOut_1_1[7] , \wRegOut_1_1[6] , 
        \wRegOut_1_1[5] , \wRegOut_1_1[4] , \wRegOut_1_1[3] , \wRegOut_1_1[2] , 
        \wRegOut_1_1[1] , \wRegOut_1_1[0] }), .P_Out({\wRegInBot_1_1[31] , 
        \wRegInBot_1_1[30] , \wRegInBot_1_1[29] , \wRegInBot_1_1[28] , 
        \wRegInBot_1_1[27] , \wRegInBot_1_1[26] , \wRegInBot_1_1[25] , 
        \wRegInBot_1_1[24] , \wRegInBot_1_1[23] , \wRegInBot_1_1[22] , 
        \wRegInBot_1_1[21] , \wRegInBot_1_1[20] , \wRegInBot_1_1[19] , 
        \wRegInBot_1_1[18] , \wRegInBot_1_1[17] , \wRegInBot_1_1[16] , 
        \wRegInBot_1_1[15] , \wRegInBot_1_1[14] , \wRegInBot_1_1[13] , 
        \wRegInBot_1_1[12] , \wRegInBot_1_1[11] , \wRegInBot_1_1[10] , 
        \wRegInBot_1_1[9] , \wRegInBot_1_1[8] , \wRegInBot_1_1[7] , 
        \wRegInBot_1_1[6] , \wRegInBot_1_1[5] , \wRegInBot_1_1[4] , 
        \wRegInBot_1_1[3] , \wRegInBot_1_1[2] , \wRegInBot_1_1[1] , 
        \wRegInBot_1_1[0] }), .L_WR(\wRegEnTop_2_2[0] ), .L_In({
        \wRegOut_2_2[31] , \wRegOut_2_2[30] , \wRegOut_2_2[29] , 
        \wRegOut_2_2[28] , \wRegOut_2_2[27] , \wRegOut_2_2[26] , 
        \wRegOut_2_2[25] , \wRegOut_2_2[24] , \wRegOut_2_2[23] , 
        \wRegOut_2_2[22] , \wRegOut_2_2[21] , \wRegOut_2_2[20] , 
        \wRegOut_2_2[19] , \wRegOut_2_2[18] , \wRegOut_2_2[17] , 
        \wRegOut_2_2[16] , \wRegOut_2_2[15] , \wRegOut_2_2[14] , 
        \wRegOut_2_2[13] , \wRegOut_2_2[12] , \wRegOut_2_2[11] , 
        \wRegOut_2_2[10] , \wRegOut_2_2[9] , \wRegOut_2_2[8] , 
        \wRegOut_2_2[7] , \wRegOut_2_2[6] , \wRegOut_2_2[5] , \wRegOut_2_2[4] , 
        \wRegOut_2_2[3] , \wRegOut_2_2[2] , \wRegOut_2_2[1] , \wRegOut_2_2[0] 
        }), .L_Out({\wRegInTop_2_2[31] , \wRegInTop_2_2[30] , 
        \wRegInTop_2_2[29] , \wRegInTop_2_2[28] , \wRegInTop_2_2[27] , 
        \wRegInTop_2_2[26] , \wRegInTop_2_2[25] , \wRegInTop_2_2[24] , 
        \wRegInTop_2_2[23] , \wRegInTop_2_2[22] , \wRegInTop_2_2[21] , 
        \wRegInTop_2_2[20] , \wRegInTop_2_2[19] , \wRegInTop_2_2[18] , 
        \wRegInTop_2_2[17] , \wRegInTop_2_2[16] , \wRegInTop_2_2[15] , 
        \wRegInTop_2_2[14] , \wRegInTop_2_2[13] , \wRegInTop_2_2[12] , 
        \wRegInTop_2_2[11] , \wRegInTop_2_2[10] , \wRegInTop_2_2[9] , 
        \wRegInTop_2_2[8] , \wRegInTop_2_2[7] , \wRegInTop_2_2[6] , 
        \wRegInTop_2_2[5] , \wRegInTop_2_2[4] , \wRegInTop_2_2[3] , 
        \wRegInTop_2_2[2] , \wRegInTop_2_2[1] , \wRegInTop_2_2[0] }), .R_WR(
        \wRegEnTop_2_3[0] ), .R_In({\wRegOut_2_3[31] , \wRegOut_2_3[30] , 
        \wRegOut_2_3[29] , \wRegOut_2_3[28] , \wRegOut_2_3[27] , 
        \wRegOut_2_3[26] , \wRegOut_2_3[25] , \wRegOut_2_3[24] , 
        \wRegOut_2_3[23] , \wRegOut_2_3[22] , \wRegOut_2_3[21] , 
        \wRegOut_2_3[20] , \wRegOut_2_3[19] , \wRegOut_2_3[18] , 
        \wRegOut_2_3[17] , \wRegOut_2_3[16] , \wRegOut_2_3[15] , 
        \wRegOut_2_3[14] , \wRegOut_2_3[13] , \wRegOut_2_3[12] , 
        \wRegOut_2_3[11] , \wRegOut_2_3[10] , \wRegOut_2_3[9] , 
        \wRegOut_2_3[8] , \wRegOut_2_3[7] , \wRegOut_2_3[6] , \wRegOut_2_3[5] , 
        \wRegOut_2_3[4] , \wRegOut_2_3[3] , \wRegOut_2_3[2] , \wRegOut_2_3[1] , 
        \wRegOut_2_3[0] }), .R_Out({\wRegInTop_2_3[31] , \wRegInTop_2_3[30] , 
        \wRegInTop_2_3[29] , \wRegInTop_2_3[28] , \wRegInTop_2_3[27] , 
        \wRegInTop_2_3[26] , \wRegInTop_2_3[25] , \wRegInTop_2_3[24] , 
        \wRegInTop_2_3[23] , \wRegInTop_2_3[22] , \wRegInTop_2_3[21] , 
        \wRegInTop_2_3[20] , \wRegInTop_2_3[19] , \wRegInTop_2_3[18] , 
        \wRegInTop_2_3[17] , \wRegInTop_2_3[16] , \wRegInTop_2_3[15] , 
        \wRegInTop_2_3[14] , \wRegInTop_2_3[13] , \wRegInTop_2_3[12] , 
        \wRegInTop_2_3[11] , \wRegInTop_2_3[10] , \wRegInTop_2_3[9] , 
        \wRegInTop_2_3[8] , \wRegInTop_2_3[7] , \wRegInTop_2_3[6] , 
        \wRegInTop_2_3[5] , \wRegInTop_2_3[4] , \wRegInTop_2_3[3] , 
        \wRegInTop_2_3[2] , \wRegInTop_2_3[1] , \wRegInTop_2_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink42[31] , \ScanLink42[30] , \ScanLink42[29] , 
        \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , \ScanLink42[25] , 
        \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , \ScanLink42[21] , 
        \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , \ScanLink42[17] , 
        \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , \ScanLink42[13] , 
        \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , \ScanLink42[9] , 
        \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , \ScanLink42[5] , 
        \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , \ScanLink42[1] , 
        \ScanLink42[0] }), .ScanOut({\ScanLink41[31] , \ScanLink41[30] , 
        \ScanLink41[29] , \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , 
        \ScanLink41[25] , \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , 
        \ScanLink41[21] , \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , 
        \ScanLink41[17] , \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , 
        \ScanLink41[13] , \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , 
        \ScanLink41[9] , \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , 
        \ScanLink41[5] , \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , 
        \ScanLink41[1] , \ScanLink41[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_10[31] , \wRegOut_5_10[30] , 
        \wRegOut_5_10[29] , \wRegOut_5_10[28] , \wRegOut_5_10[27] , 
        \wRegOut_5_10[26] , \wRegOut_5_10[25] , \wRegOut_5_10[24] , 
        \wRegOut_5_10[23] , \wRegOut_5_10[22] , \wRegOut_5_10[21] , 
        \wRegOut_5_10[20] , \wRegOut_5_10[19] , \wRegOut_5_10[18] , 
        \wRegOut_5_10[17] , \wRegOut_5_10[16] , \wRegOut_5_10[15] , 
        \wRegOut_5_10[14] , \wRegOut_5_10[13] , \wRegOut_5_10[12] , 
        \wRegOut_5_10[11] , \wRegOut_5_10[10] , \wRegOut_5_10[9] , 
        \wRegOut_5_10[8] , \wRegOut_5_10[7] , \wRegOut_5_10[6] , 
        \wRegOut_5_10[5] , \wRegOut_5_10[4] , \wRegOut_5_10[3] , 
        \wRegOut_5_10[2] , \wRegOut_5_10[1] , \wRegOut_5_10[0] }), .Enable1(
        \wRegEnTop_5_10[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_10[31] , 
        \wRegInTop_5_10[30] , \wRegInTop_5_10[29] , \wRegInTop_5_10[28] , 
        \wRegInTop_5_10[27] , \wRegInTop_5_10[26] , \wRegInTop_5_10[25] , 
        \wRegInTop_5_10[24] , \wRegInTop_5_10[23] , \wRegInTop_5_10[22] , 
        \wRegInTop_5_10[21] , \wRegInTop_5_10[20] , \wRegInTop_5_10[19] , 
        \wRegInTop_5_10[18] , \wRegInTop_5_10[17] , \wRegInTop_5_10[16] , 
        \wRegInTop_5_10[15] , \wRegInTop_5_10[14] , \wRegInTop_5_10[13] , 
        \wRegInTop_5_10[12] , \wRegInTop_5_10[11] , \wRegInTop_5_10[10] , 
        \wRegInTop_5_10[9] , \wRegInTop_5_10[8] , \wRegInTop_5_10[7] , 
        \wRegInTop_5_10[6] , \wRegInTop_5_10[5] , \wRegInTop_5_10[4] , 
        \wRegInTop_5_10[3] , \wRegInTop_5_10[2] , \wRegInTop_5_10[1] , 
        \wRegInTop_5_10[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_7[0] ), .P_In({\wRegOut_4_7[31] , 
        \wRegOut_4_7[30] , \wRegOut_4_7[29] , \wRegOut_4_7[28] , 
        \wRegOut_4_7[27] , \wRegOut_4_7[26] , \wRegOut_4_7[25] , 
        \wRegOut_4_7[24] , \wRegOut_4_7[23] , \wRegOut_4_7[22] , 
        \wRegOut_4_7[21] , \wRegOut_4_7[20] , \wRegOut_4_7[19] , 
        \wRegOut_4_7[18] , \wRegOut_4_7[17] , \wRegOut_4_7[16] , 
        \wRegOut_4_7[15] , \wRegOut_4_7[14] , \wRegOut_4_7[13] , 
        \wRegOut_4_7[12] , \wRegOut_4_7[11] , \wRegOut_4_7[10] , 
        \wRegOut_4_7[9] , \wRegOut_4_7[8] , \wRegOut_4_7[7] , \wRegOut_4_7[6] , 
        \wRegOut_4_7[5] , \wRegOut_4_7[4] , \wRegOut_4_7[3] , \wRegOut_4_7[2] , 
        \wRegOut_4_7[1] , \wRegOut_4_7[0] }), .P_Out({\wRegInBot_4_7[31] , 
        \wRegInBot_4_7[30] , \wRegInBot_4_7[29] , \wRegInBot_4_7[28] , 
        \wRegInBot_4_7[27] , \wRegInBot_4_7[26] , \wRegInBot_4_7[25] , 
        \wRegInBot_4_7[24] , \wRegInBot_4_7[23] , \wRegInBot_4_7[22] , 
        \wRegInBot_4_7[21] , \wRegInBot_4_7[20] , \wRegInBot_4_7[19] , 
        \wRegInBot_4_7[18] , \wRegInBot_4_7[17] , \wRegInBot_4_7[16] , 
        \wRegInBot_4_7[15] , \wRegInBot_4_7[14] , \wRegInBot_4_7[13] , 
        \wRegInBot_4_7[12] , \wRegInBot_4_7[11] , \wRegInBot_4_7[10] , 
        \wRegInBot_4_7[9] , \wRegInBot_4_7[8] , \wRegInBot_4_7[7] , 
        \wRegInBot_4_7[6] , \wRegInBot_4_7[5] , \wRegInBot_4_7[4] , 
        \wRegInBot_4_7[3] , \wRegInBot_4_7[2] , \wRegInBot_4_7[1] , 
        \wRegInBot_4_7[0] }), .L_WR(\wRegEnTop_5_14[0] ), .L_In({
        \wRegOut_5_14[31] , \wRegOut_5_14[30] , \wRegOut_5_14[29] , 
        \wRegOut_5_14[28] , \wRegOut_5_14[27] , \wRegOut_5_14[26] , 
        \wRegOut_5_14[25] , \wRegOut_5_14[24] , \wRegOut_5_14[23] , 
        \wRegOut_5_14[22] , \wRegOut_5_14[21] , \wRegOut_5_14[20] , 
        \wRegOut_5_14[19] , \wRegOut_5_14[18] , \wRegOut_5_14[17] , 
        \wRegOut_5_14[16] , \wRegOut_5_14[15] , \wRegOut_5_14[14] , 
        \wRegOut_5_14[13] , \wRegOut_5_14[12] , \wRegOut_5_14[11] , 
        \wRegOut_5_14[10] , \wRegOut_5_14[9] , \wRegOut_5_14[8] , 
        \wRegOut_5_14[7] , \wRegOut_5_14[6] , \wRegOut_5_14[5] , 
        \wRegOut_5_14[4] , \wRegOut_5_14[3] , \wRegOut_5_14[2] , 
        \wRegOut_5_14[1] , \wRegOut_5_14[0] }), .L_Out({\wRegInTop_5_14[31] , 
        \wRegInTop_5_14[30] , \wRegInTop_5_14[29] , \wRegInTop_5_14[28] , 
        \wRegInTop_5_14[27] , \wRegInTop_5_14[26] , \wRegInTop_5_14[25] , 
        \wRegInTop_5_14[24] , \wRegInTop_5_14[23] , \wRegInTop_5_14[22] , 
        \wRegInTop_5_14[21] , \wRegInTop_5_14[20] , \wRegInTop_5_14[19] , 
        \wRegInTop_5_14[18] , \wRegInTop_5_14[17] , \wRegInTop_5_14[16] , 
        \wRegInTop_5_14[15] , \wRegInTop_5_14[14] , \wRegInTop_5_14[13] , 
        \wRegInTop_5_14[12] , \wRegInTop_5_14[11] , \wRegInTop_5_14[10] , 
        \wRegInTop_5_14[9] , \wRegInTop_5_14[8] , \wRegInTop_5_14[7] , 
        \wRegInTop_5_14[6] , \wRegInTop_5_14[5] , \wRegInTop_5_14[4] , 
        \wRegInTop_5_14[3] , \wRegInTop_5_14[2] , \wRegInTop_5_14[1] , 
        \wRegInTop_5_14[0] }), .R_WR(\wRegEnTop_5_15[0] ), .R_In({
        \wRegOut_5_15[31] , \wRegOut_5_15[30] , \wRegOut_5_15[29] , 
        \wRegOut_5_15[28] , \wRegOut_5_15[27] , \wRegOut_5_15[26] , 
        \wRegOut_5_15[25] , \wRegOut_5_15[24] , \wRegOut_5_15[23] , 
        \wRegOut_5_15[22] , \wRegOut_5_15[21] , \wRegOut_5_15[20] , 
        \wRegOut_5_15[19] , \wRegOut_5_15[18] , \wRegOut_5_15[17] , 
        \wRegOut_5_15[16] , \wRegOut_5_15[15] , \wRegOut_5_15[14] , 
        \wRegOut_5_15[13] , \wRegOut_5_15[12] , \wRegOut_5_15[11] , 
        \wRegOut_5_15[10] , \wRegOut_5_15[9] , \wRegOut_5_15[8] , 
        \wRegOut_5_15[7] , \wRegOut_5_15[6] , \wRegOut_5_15[5] , 
        \wRegOut_5_15[4] , \wRegOut_5_15[3] , \wRegOut_5_15[2] , 
        \wRegOut_5_15[1] , \wRegOut_5_15[0] }), .R_Out({\wRegInTop_5_15[31] , 
        \wRegInTop_5_15[30] , \wRegInTop_5_15[29] , \wRegInTop_5_15[28] , 
        \wRegInTop_5_15[27] , \wRegInTop_5_15[26] , \wRegInTop_5_15[25] , 
        \wRegInTop_5_15[24] , \wRegInTop_5_15[23] , \wRegInTop_5_15[22] , 
        \wRegInTop_5_15[21] , \wRegInTop_5_15[20] , \wRegInTop_5_15[19] , 
        \wRegInTop_5_15[18] , \wRegInTop_5_15[17] , \wRegInTop_5_15[16] , 
        \wRegInTop_5_15[15] , \wRegInTop_5_15[14] , \wRegInTop_5_15[13] , 
        \wRegInTop_5_15[12] , \wRegInTop_5_15[11] , \wRegInTop_5_15[10] , 
        \wRegInTop_5_15[9] , \wRegInTop_5_15[8] , \wRegInTop_5_15[7] , 
        \wRegInTop_5_15[6] , \wRegInTop_5_15[5] , \wRegInTop_5_15[4] , 
        \wRegInTop_5_15[3] , \wRegInTop_5_15[2] , \wRegInTop_5_15[1] , 
        \wRegInTop_5_15[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink34[31] , \ScanLink34[30] , \ScanLink34[29] , 
        \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , \ScanLink34[25] , 
        \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , \ScanLink34[21] , 
        \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , \ScanLink34[17] , 
        \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , \ScanLink34[13] , 
        \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , \ScanLink34[9] , 
        \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , \ScanLink34[5] , 
        \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , \ScanLink34[1] , 
        \ScanLink34[0] }), .ScanOut({\ScanLink33[31] , \ScanLink33[30] , 
        \ScanLink33[29] , \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , 
        \ScanLink33[25] , \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , 
        \ScanLink33[21] , \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , 
        \ScanLink33[17] , \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , 
        \ScanLink33[13] , \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , 
        \ScanLink33[9] , \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , 
        \ScanLink33[5] , \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , 
        \ScanLink33[1] , \ScanLink33[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_2[31] , \wRegOut_5_2[30] , \wRegOut_5_2[29] , 
        \wRegOut_5_2[28] , \wRegOut_5_2[27] , \wRegOut_5_2[26] , 
        \wRegOut_5_2[25] , \wRegOut_5_2[24] , \wRegOut_5_2[23] , 
        \wRegOut_5_2[22] , \wRegOut_5_2[21] , \wRegOut_5_2[20] , 
        \wRegOut_5_2[19] , \wRegOut_5_2[18] , \wRegOut_5_2[17] , 
        \wRegOut_5_2[16] , \wRegOut_5_2[15] , \wRegOut_5_2[14] , 
        \wRegOut_5_2[13] , \wRegOut_5_2[12] , \wRegOut_5_2[11] , 
        \wRegOut_5_2[10] , \wRegOut_5_2[9] , \wRegOut_5_2[8] , 
        \wRegOut_5_2[7] , \wRegOut_5_2[6] , \wRegOut_5_2[5] , \wRegOut_5_2[4] , 
        \wRegOut_5_2[3] , \wRegOut_5_2[2] , \wRegOut_5_2[1] , \wRegOut_5_2[0] 
        }), .Enable1(\wRegEnTop_5_2[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_2[31] , \wRegInTop_5_2[30] , \wRegInTop_5_2[29] , 
        \wRegInTop_5_2[28] , \wRegInTop_5_2[27] , \wRegInTop_5_2[26] , 
        \wRegInTop_5_2[25] , \wRegInTop_5_2[24] , \wRegInTop_5_2[23] , 
        \wRegInTop_5_2[22] , \wRegInTop_5_2[21] , \wRegInTop_5_2[20] , 
        \wRegInTop_5_2[19] , \wRegInTop_5_2[18] , \wRegInTop_5_2[17] , 
        \wRegInTop_5_2[16] , \wRegInTop_5_2[15] , \wRegInTop_5_2[14] , 
        \wRegInTop_5_2[13] , \wRegInTop_5_2[12] , \wRegInTop_5_2[11] , 
        \wRegInTop_5_2[10] , \wRegInTop_5_2[9] , \wRegInTop_5_2[8] , 
        \wRegInTop_5_2[7] , \wRegInTop_5_2[6] , \wRegInTop_5_2[5] , 
        \wRegInTop_5_2[4] , \wRegInTop_5_2[3] , \wRegInTop_5_2[2] , 
        \wRegInTop_5_2[1] , \wRegInTop_5_2[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_17 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink49[31] , \ScanLink49[30] , \ScanLink49[29] , 
        \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , \ScanLink49[25] , 
        \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , \ScanLink49[21] , 
        \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , \ScanLink49[17] , 
        \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , \ScanLink49[13] , 
        \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , \ScanLink49[9] , 
        \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , \ScanLink49[5] , 
        \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , \ScanLink49[1] , 
        \ScanLink49[0] }), .ScanOut({\ScanLink48[31] , \ScanLink48[30] , 
        \ScanLink48[29] , \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , 
        \ScanLink48[25] , \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , 
        \ScanLink48[21] , \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , 
        \ScanLink48[17] , \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , 
        \ScanLink48[13] , \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , 
        \ScanLink48[9] , \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , 
        \ScanLink48[5] , \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , 
        \ScanLink48[1] , \ScanLink48[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_17[31] , \wRegOut_5_17[30] , 
        \wRegOut_5_17[29] , \wRegOut_5_17[28] , \wRegOut_5_17[27] , 
        \wRegOut_5_17[26] , \wRegOut_5_17[25] , \wRegOut_5_17[24] , 
        \wRegOut_5_17[23] , \wRegOut_5_17[22] , \wRegOut_5_17[21] , 
        \wRegOut_5_17[20] , \wRegOut_5_17[19] , \wRegOut_5_17[18] , 
        \wRegOut_5_17[17] , \wRegOut_5_17[16] , \wRegOut_5_17[15] , 
        \wRegOut_5_17[14] , \wRegOut_5_17[13] , \wRegOut_5_17[12] , 
        \wRegOut_5_17[11] , \wRegOut_5_17[10] , \wRegOut_5_17[9] , 
        \wRegOut_5_17[8] , \wRegOut_5_17[7] , \wRegOut_5_17[6] , 
        \wRegOut_5_17[5] , \wRegOut_5_17[4] , \wRegOut_5_17[3] , 
        \wRegOut_5_17[2] , \wRegOut_5_17[1] , \wRegOut_5_17[0] }), .Enable1(
        \wRegEnTop_5_17[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_17[31] , 
        \wRegInTop_5_17[30] , \wRegInTop_5_17[29] , \wRegInTop_5_17[28] , 
        \wRegInTop_5_17[27] , \wRegInTop_5_17[26] , \wRegInTop_5_17[25] , 
        \wRegInTop_5_17[24] , \wRegInTop_5_17[23] , \wRegInTop_5_17[22] , 
        \wRegInTop_5_17[21] , \wRegInTop_5_17[20] , \wRegInTop_5_17[19] , 
        \wRegInTop_5_17[18] , \wRegInTop_5_17[17] , \wRegInTop_5_17[16] , 
        \wRegInTop_5_17[15] , \wRegInTop_5_17[14] , \wRegInTop_5_17[13] , 
        \wRegInTop_5_17[12] , \wRegInTop_5_17[11] , \wRegInTop_5_17[10] , 
        \wRegInTop_5_17[9] , \wRegInTop_5_17[8] , \wRegInTop_5_17[7] , 
        \wRegInTop_5_17[6] , \wRegInTop_5_17[5] , \wRegInTop_5_17[4] , 
        \wRegInTop_5_17[3] , \wRegInTop_5_17[2] , \wRegInTop_5_17[1] , 
        \wRegInTop_5_17[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_30 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink62[31] , \ScanLink62[30] , \ScanLink62[29] , 
        \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , \ScanLink62[25] , 
        \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , \ScanLink62[21] , 
        \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , \ScanLink62[17] , 
        \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , \ScanLink62[13] , 
        \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , \ScanLink62[9] , 
        \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , \ScanLink62[5] , 
        \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , \ScanLink62[1] , 
        \ScanLink62[0] }), .ScanOut({\ScanLink61[31] , \ScanLink61[30] , 
        \ScanLink61[29] , \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , 
        \ScanLink61[25] , \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , 
        \ScanLink61[21] , \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , 
        \ScanLink61[17] , \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , 
        \ScanLink61[13] , \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , 
        \ScanLink61[9] , \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , 
        \ScanLink61[5] , \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , 
        \ScanLink61[1] , \ScanLink61[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_30[31] , \wRegOut_5_30[30] , 
        \wRegOut_5_30[29] , \wRegOut_5_30[28] , \wRegOut_5_30[27] , 
        \wRegOut_5_30[26] , \wRegOut_5_30[25] , \wRegOut_5_30[24] , 
        \wRegOut_5_30[23] , \wRegOut_5_30[22] , \wRegOut_5_30[21] , 
        \wRegOut_5_30[20] , \wRegOut_5_30[19] , \wRegOut_5_30[18] , 
        \wRegOut_5_30[17] , \wRegOut_5_30[16] , \wRegOut_5_30[15] , 
        \wRegOut_5_30[14] , \wRegOut_5_30[13] , \wRegOut_5_30[12] , 
        \wRegOut_5_30[11] , \wRegOut_5_30[10] , \wRegOut_5_30[9] , 
        \wRegOut_5_30[8] , \wRegOut_5_30[7] , \wRegOut_5_30[6] , 
        \wRegOut_5_30[5] , \wRegOut_5_30[4] , \wRegOut_5_30[3] , 
        \wRegOut_5_30[2] , \wRegOut_5_30[1] , \wRegOut_5_30[0] }), .Enable1(
        \wRegEnTop_5_30[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_30[31] , 
        \wRegInTop_5_30[30] , \wRegInTop_5_30[29] , \wRegInTop_5_30[28] , 
        \wRegInTop_5_30[27] , \wRegInTop_5_30[26] , \wRegInTop_5_30[25] , 
        \wRegInTop_5_30[24] , \wRegInTop_5_30[23] , \wRegInTop_5_30[22] , 
        \wRegInTop_5_30[21] , \wRegInTop_5_30[20] , \wRegInTop_5_30[19] , 
        \wRegInTop_5_30[18] , \wRegInTop_5_30[17] , \wRegInTop_5_30[16] , 
        \wRegInTop_5_30[15] , \wRegInTop_5_30[14] , \wRegInTop_5_30[13] , 
        \wRegInTop_5_30[12] , \wRegInTop_5_30[11] , \wRegInTop_5_30[10] , 
        \wRegInTop_5_30[9] , \wRegInTop_5_30[8] , \wRegInTop_5_30[7] , 
        \wRegInTop_5_30[6] , \wRegInTop_5_30[5] , \wRegInTop_5_30[4] , 
        \wRegInTop_5_30[3] , \wRegInTop_5_30[2] , \wRegInTop_5_30[1] , 
        \wRegInTop_5_30[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_0[0] ), .P_In({\wRegOut_4_0[31] , 
        \wRegOut_4_0[30] , \wRegOut_4_0[29] , \wRegOut_4_0[28] , 
        \wRegOut_4_0[27] , \wRegOut_4_0[26] , \wRegOut_4_0[25] , 
        \wRegOut_4_0[24] , \wRegOut_4_0[23] , \wRegOut_4_0[22] , 
        \wRegOut_4_0[21] , \wRegOut_4_0[20] , \wRegOut_4_0[19] , 
        \wRegOut_4_0[18] , \wRegOut_4_0[17] , \wRegOut_4_0[16] , 
        \wRegOut_4_0[15] , \wRegOut_4_0[14] , \wRegOut_4_0[13] , 
        \wRegOut_4_0[12] , \wRegOut_4_0[11] , \wRegOut_4_0[10] , 
        \wRegOut_4_0[9] , \wRegOut_4_0[8] , \wRegOut_4_0[7] , \wRegOut_4_0[6] , 
        \wRegOut_4_0[5] , \wRegOut_4_0[4] , \wRegOut_4_0[3] , \wRegOut_4_0[2] , 
        \wRegOut_4_0[1] , \wRegOut_4_0[0] }), .P_Out({\wRegInBot_4_0[31] , 
        \wRegInBot_4_0[30] , \wRegInBot_4_0[29] , \wRegInBot_4_0[28] , 
        \wRegInBot_4_0[27] , \wRegInBot_4_0[26] , \wRegInBot_4_0[25] , 
        \wRegInBot_4_0[24] , \wRegInBot_4_0[23] , \wRegInBot_4_0[22] , 
        \wRegInBot_4_0[21] , \wRegInBot_4_0[20] , \wRegInBot_4_0[19] , 
        \wRegInBot_4_0[18] , \wRegInBot_4_0[17] , \wRegInBot_4_0[16] , 
        \wRegInBot_4_0[15] , \wRegInBot_4_0[14] , \wRegInBot_4_0[13] , 
        \wRegInBot_4_0[12] , \wRegInBot_4_0[11] , \wRegInBot_4_0[10] , 
        \wRegInBot_4_0[9] , \wRegInBot_4_0[8] , \wRegInBot_4_0[7] , 
        \wRegInBot_4_0[6] , \wRegInBot_4_0[5] , \wRegInBot_4_0[4] , 
        \wRegInBot_4_0[3] , \wRegInBot_4_0[2] , \wRegInBot_4_0[1] , 
        \wRegInBot_4_0[0] }), .L_WR(\wRegEnTop_5_0[0] ), .L_In({
        \wRegOut_5_0[31] , \wRegOut_5_0[30] , \wRegOut_5_0[29] , 
        \wRegOut_5_0[28] , \wRegOut_5_0[27] , \wRegOut_5_0[26] , 
        \wRegOut_5_0[25] , \wRegOut_5_0[24] , \wRegOut_5_0[23] , 
        \wRegOut_5_0[22] , \wRegOut_5_0[21] , \wRegOut_5_0[20] , 
        \wRegOut_5_0[19] , \wRegOut_5_0[18] , \wRegOut_5_0[17] , 
        \wRegOut_5_0[16] , \wRegOut_5_0[15] , \wRegOut_5_0[14] , 
        \wRegOut_5_0[13] , \wRegOut_5_0[12] , \wRegOut_5_0[11] , 
        \wRegOut_5_0[10] , \wRegOut_5_0[9] , \wRegOut_5_0[8] , 
        \wRegOut_5_0[7] , \wRegOut_5_0[6] , \wRegOut_5_0[5] , \wRegOut_5_0[4] , 
        \wRegOut_5_0[3] , \wRegOut_5_0[2] , \wRegOut_5_0[1] , \wRegOut_5_0[0] 
        }), .L_Out({\wRegInTop_5_0[31] , \wRegInTop_5_0[30] , 
        \wRegInTop_5_0[29] , \wRegInTop_5_0[28] , \wRegInTop_5_0[27] , 
        \wRegInTop_5_0[26] , \wRegInTop_5_0[25] , \wRegInTop_5_0[24] , 
        \wRegInTop_5_0[23] , \wRegInTop_5_0[22] , \wRegInTop_5_0[21] , 
        \wRegInTop_5_0[20] , \wRegInTop_5_0[19] , \wRegInTop_5_0[18] , 
        \wRegInTop_5_0[17] , \wRegInTop_5_0[16] , \wRegInTop_5_0[15] , 
        \wRegInTop_5_0[14] , \wRegInTop_5_0[13] , \wRegInTop_5_0[12] , 
        \wRegInTop_5_0[11] , \wRegInTop_5_0[10] , \wRegInTop_5_0[9] , 
        \wRegInTop_5_0[8] , \wRegInTop_5_0[7] , \wRegInTop_5_0[6] , 
        \wRegInTop_5_0[5] , \wRegInTop_5_0[4] , \wRegInTop_5_0[3] , 
        \wRegInTop_5_0[2] , \wRegInTop_5_0[1] , \wRegInTop_5_0[0] }), .R_WR(
        \wRegEnTop_5_1[0] ), .R_In({\wRegOut_5_1[31] , \wRegOut_5_1[30] , 
        \wRegOut_5_1[29] , \wRegOut_5_1[28] , \wRegOut_5_1[27] , 
        \wRegOut_5_1[26] , \wRegOut_5_1[25] , \wRegOut_5_1[24] , 
        \wRegOut_5_1[23] , \wRegOut_5_1[22] , \wRegOut_5_1[21] , 
        \wRegOut_5_1[20] , \wRegOut_5_1[19] , \wRegOut_5_1[18] , 
        \wRegOut_5_1[17] , \wRegOut_5_1[16] , \wRegOut_5_1[15] , 
        \wRegOut_5_1[14] , \wRegOut_5_1[13] , \wRegOut_5_1[12] , 
        \wRegOut_5_1[11] , \wRegOut_5_1[10] , \wRegOut_5_1[9] , 
        \wRegOut_5_1[8] , \wRegOut_5_1[7] , \wRegOut_5_1[6] , \wRegOut_5_1[5] , 
        \wRegOut_5_1[4] , \wRegOut_5_1[3] , \wRegOut_5_1[2] , \wRegOut_5_1[1] , 
        \wRegOut_5_1[0] }), .R_Out({\wRegInTop_5_1[31] , \wRegInTop_5_1[30] , 
        \wRegInTop_5_1[29] , \wRegInTop_5_1[28] , \wRegInTop_5_1[27] , 
        \wRegInTop_5_1[26] , \wRegInTop_5_1[25] , \wRegInTop_5_1[24] , 
        \wRegInTop_5_1[23] , \wRegInTop_5_1[22] , \wRegInTop_5_1[21] , 
        \wRegInTop_5_1[20] , \wRegInTop_5_1[19] , \wRegInTop_5_1[18] , 
        \wRegInTop_5_1[17] , \wRegInTop_5_1[16] , \wRegInTop_5_1[15] , 
        \wRegInTop_5_1[14] , \wRegInTop_5_1[13] , \wRegInTop_5_1[12] , 
        \wRegInTop_5_1[11] , \wRegInTop_5_1[10] , \wRegInTop_5_1[9] , 
        \wRegInTop_5_1[8] , \wRegInTop_5_1[7] , \wRegInTop_5_1[6] , 
        \wRegInTop_5_1[5] , \wRegInTop_5_1[4] , \wRegInTop_5_1[3] , 
        \wRegInTop_5_1[2] , \wRegInTop_5_1[1] , \wRegInTop_5_1[0] }) );
    BHeap_Node_WIDTH32 BHN_2_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_2[0] ), .P_WR(\wRegEnBot_2_3[0] ), .P_In({\wRegOut_2_3[31] , 
        \wRegOut_2_3[30] , \wRegOut_2_3[29] , \wRegOut_2_3[28] , 
        \wRegOut_2_3[27] , \wRegOut_2_3[26] , \wRegOut_2_3[25] , 
        \wRegOut_2_3[24] , \wRegOut_2_3[23] , \wRegOut_2_3[22] , 
        \wRegOut_2_3[21] , \wRegOut_2_3[20] , \wRegOut_2_3[19] , 
        \wRegOut_2_3[18] , \wRegOut_2_3[17] , \wRegOut_2_3[16] , 
        \wRegOut_2_3[15] , \wRegOut_2_3[14] , \wRegOut_2_3[13] , 
        \wRegOut_2_3[12] , \wRegOut_2_3[11] , \wRegOut_2_3[10] , 
        \wRegOut_2_3[9] , \wRegOut_2_3[8] , \wRegOut_2_3[7] , \wRegOut_2_3[6] , 
        \wRegOut_2_3[5] , \wRegOut_2_3[4] , \wRegOut_2_3[3] , \wRegOut_2_3[2] , 
        \wRegOut_2_3[1] , \wRegOut_2_3[0] }), .P_Out({\wRegInBot_2_3[31] , 
        \wRegInBot_2_3[30] , \wRegInBot_2_3[29] , \wRegInBot_2_3[28] , 
        \wRegInBot_2_3[27] , \wRegInBot_2_3[26] , \wRegInBot_2_3[25] , 
        \wRegInBot_2_3[24] , \wRegInBot_2_3[23] , \wRegInBot_2_3[22] , 
        \wRegInBot_2_3[21] , \wRegInBot_2_3[20] , \wRegInBot_2_3[19] , 
        \wRegInBot_2_3[18] , \wRegInBot_2_3[17] , \wRegInBot_2_3[16] , 
        \wRegInBot_2_3[15] , \wRegInBot_2_3[14] , \wRegInBot_2_3[13] , 
        \wRegInBot_2_3[12] , \wRegInBot_2_3[11] , \wRegInBot_2_3[10] , 
        \wRegInBot_2_3[9] , \wRegInBot_2_3[8] , \wRegInBot_2_3[7] , 
        \wRegInBot_2_3[6] , \wRegInBot_2_3[5] , \wRegInBot_2_3[4] , 
        \wRegInBot_2_3[3] , \wRegInBot_2_3[2] , \wRegInBot_2_3[1] , 
        \wRegInBot_2_3[0] }), .L_WR(\wRegEnTop_3_6[0] ), .L_In({
        \wRegOut_3_6[31] , \wRegOut_3_6[30] , \wRegOut_3_6[29] , 
        \wRegOut_3_6[28] , \wRegOut_3_6[27] , \wRegOut_3_6[26] , 
        \wRegOut_3_6[25] , \wRegOut_3_6[24] , \wRegOut_3_6[23] , 
        \wRegOut_3_6[22] , \wRegOut_3_6[21] , \wRegOut_3_6[20] , 
        \wRegOut_3_6[19] , \wRegOut_3_6[18] , \wRegOut_3_6[17] , 
        \wRegOut_3_6[16] , \wRegOut_3_6[15] , \wRegOut_3_6[14] , 
        \wRegOut_3_6[13] , \wRegOut_3_6[12] , \wRegOut_3_6[11] , 
        \wRegOut_3_6[10] , \wRegOut_3_6[9] , \wRegOut_3_6[8] , 
        \wRegOut_3_6[7] , \wRegOut_3_6[6] , \wRegOut_3_6[5] , \wRegOut_3_6[4] , 
        \wRegOut_3_6[3] , \wRegOut_3_6[2] , \wRegOut_3_6[1] , \wRegOut_3_6[0] 
        }), .L_Out({\wRegInTop_3_6[31] , \wRegInTop_3_6[30] , 
        \wRegInTop_3_6[29] , \wRegInTop_3_6[28] , \wRegInTop_3_6[27] , 
        \wRegInTop_3_6[26] , \wRegInTop_3_6[25] , \wRegInTop_3_6[24] , 
        \wRegInTop_3_6[23] , \wRegInTop_3_6[22] , \wRegInTop_3_6[21] , 
        \wRegInTop_3_6[20] , \wRegInTop_3_6[19] , \wRegInTop_3_6[18] , 
        \wRegInTop_3_6[17] , \wRegInTop_3_6[16] , \wRegInTop_3_6[15] , 
        \wRegInTop_3_6[14] , \wRegInTop_3_6[13] , \wRegInTop_3_6[12] , 
        \wRegInTop_3_6[11] , \wRegInTop_3_6[10] , \wRegInTop_3_6[9] , 
        \wRegInTop_3_6[8] , \wRegInTop_3_6[7] , \wRegInTop_3_6[6] , 
        \wRegInTop_3_6[5] , \wRegInTop_3_6[4] , \wRegInTop_3_6[3] , 
        \wRegInTop_3_6[2] , \wRegInTop_3_6[1] , \wRegInTop_3_6[0] }), .R_WR(
        \wRegEnTop_3_7[0] ), .R_In({\wRegOut_3_7[31] , \wRegOut_3_7[30] , 
        \wRegOut_3_7[29] , \wRegOut_3_7[28] , \wRegOut_3_7[27] , 
        \wRegOut_3_7[26] , \wRegOut_3_7[25] , \wRegOut_3_7[24] , 
        \wRegOut_3_7[23] , \wRegOut_3_7[22] , \wRegOut_3_7[21] , 
        \wRegOut_3_7[20] , \wRegOut_3_7[19] , \wRegOut_3_7[18] , 
        \wRegOut_3_7[17] , \wRegOut_3_7[16] , \wRegOut_3_7[15] , 
        \wRegOut_3_7[14] , \wRegOut_3_7[13] , \wRegOut_3_7[12] , 
        \wRegOut_3_7[11] , \wRegOut_3_7[10] , \wRegOut_3_7[9] , 
        \wRegOut_3_7[8] , \wRegOut_3_7[7] , \wRegOut_3_7[6] , \wRegOut_3_7[5] , 
        \wRegOut_3_7[4] , \wRegOut_3_7[3] , \wRegOut_3_7[2] , \wRegOut_3_7[1] , 
        \wRegOut_3_7[0] }), .R_Out({\wRegInTop_3_7[31] , \wRegInTop_3_7[30] , 
        \wRegInTop_3_7[29] , \wRegInTop_3_7[28] , \wRegInTop_3_7[27] , 
        \wRegInTop_3_7[26] , \wRegInTop_3_7[25] , \wRegInTop_3_7[24] , 
        \wRegInTop_3_7[23] , \wRegInTop_3_7[22] , \wRegInTop_3_7[21] , 
        \wRegInTop_3_7[20] , \wRegInTop_3_7[19] , \wRegInTop_3_7[18] , 
        \wRegInTop_3_7[17] , \wRegInTop_3_7[16] , \wRegInTop_3_7[15] , 
        \wRegInTop_3_7[14] , \wRegInTop_3_7[13] , \wRegInTop_3_7[12] , 
        \wRegInTop_3_7[11] , \wRegInTop_3_7[10] , \wRegInTop_3_7[9] , 
        \wRegInTop_3_7[8] , \wRegInTop_3_7[7] , \wRegInTop_3_7[6] , 
        \wRegInTop_3_7[5] , \wRegInTop_3_7[4] , \wRegInTop_3_7[3] , 
        \wRegInTop_3_7[2] , \wRegInTop_3_7[1] , \wRegInTop_3_7[0] }) );
    BHeap_Node_WIDTH32 BHN_3_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_3[0] ), .P_In({\wRegOut_3_3[31] , 
        \wRegOut_3_3[30] , \wRegOut_3_3[29] , \wRegOut_3_3[28] , 
        \wRegOut_3_3[27] , \wRegOut_3_3[26] , \wRegOut_3_3[25] , 
        \wRegOut_3_3[24] , \wRegOut_3_3[23] , \wRegOut_3_3[22] , 
        \wRegOut_3_3[21] , \wRegOut_3_3[20] , \wRegOut_3_3[19] , 
        \wRegOut_3_3[18] , \wRegOut_3_3[17] , \wRegOut_3_3[16] , 
        \wRegOut_3_3[15] , \wRegOut_3_3[14] , \wRegOut_3_3[13] , 
        \wRegOut_3_3[12] , \wRegOut_3_3[11] , \wRegOut_3_3[10] , 
        \wRegOut_3_3[9] , \wRegOut_3_3[8] , \wRegOut_3_3[7] , \wRegOut_3_3[6] , 
        \wRegOut_3_3[5] , \wRegOut_3_3[4] , \wRegOut_3_3[3] , \wRegOut_3_3[2] , 
        \wRegOut_3_3[1] , \wRegOut_3_3[0] }), .P_Out({\wRegInBot_3_3[31] , 
        \wRegInBot_3_3[30] , \wRegInBot_3_3[29] , \wRegInBot_3_3[28] , 
        \wRegInBot_3_3[27] , \wRegInBot_3_3[26] , \wRegInBot_3_3[25] , 
        \wRegInBot_3_3[24] , \wRegInBot_3_3[23] , \wRegInBot_3_3[22] , 
        \wRegInBot_3_3[21] , \wRegInBot_3_3[20] , \wRegInBot_3_3[19] , 
        \wRegInBot_3_3[18] , \wRegInBot_3_3[17] , \wRegInBot_3_3[16] , 
        \wRegInBot_3_3[15] , \wRegInBot_3_3[14] , \wRegInBot_3_3[13] , 
        \wRegInBot_3_3[12] , \wRegInBot_3_3[11] , \wRegInBot_3_3[10] , 
        \wRegInBot_3_3[9] , \wRegInBot_3_3[8] , \wRegInBot_3_3[7] , 
        \wRegInBot_3_3[6] , \wRegInBot_3_3[5] , \wRegInBot_3_3[4] , 
        \wRegInBot_3_3[3] , \wRegInBot_3_3[2] , \wRegInBot_3_3[1] , 
        \wRegInBot_3_3[0] }), .L_WR(\wRegEnTop_4_6[0] ), .L_In({
        \wRegOut_4_6[31] , \wRegOut_4_6[30] , \wRegOut_4_6[29] , 
        \wRegOut_4_6[28] , \wRegOut_4_6[27] , \wRegOut_4_6[26] , 
        \wRegOut_4_6[25] , \wRegOut_4_6[24] , \wRegOut_4_6[23] , 
        \wRegOut_4_6[22] , \wRegOut_4_6[21] , \wRegOut_4_6[20] , 
        \wRegOut_4_6[19] , \wRegOut_4_6[18] , \wRegOut_4_6[17] , 
        \wRegOut_4_6[16] , \wRegOut_4_6[15] , \wRegOut_4_6[14] , 
        \wRegOut_4_6[13] , \wRegOut_4_6[12] , \wRegOut_4_6[11] , 
        \wRegOut_4_6[10] , \wRegOut_4_6[9] , \wRegOut_4_6[8] , 
        \wRegOut_4_6[7] , \wRegOut_4_6[6] , \wRegOut_4_6[5] , \wRegOut_4_6[4] , 
        \wRegOut_4_6[3] , \wRegOut_4_6[2] , \wRegOut_4_6[1] , \wRegOut_4_6[0] 
        }), .L_Out({\wRegInTop_4_6[31] , \wRegInTop_4_6[30] , 
        \wRegInTop_4_6[29] , \wRegInTop_4_6[28] , \wRegInTop_4_6[27] , 
        \wRegInTop_4_6[26] , \wRegInTop_4_6[25] , \wRegInTop_4_6[24] , 
        \wRegInTop_4_6[23] , \wRegInTop_4_6[22] , \wRegInTop_4_6[21] , 
        \wRegInTop_4_6[20] , \wRegInTop_4_6[19] , \wRegInTop_4_6[18] , 
        \wRegInTop_4_6[17] , \wRegInTop_4_6[16] , \wRegInTop_4_6[15] , 
        \wRegInTop_4_6[14] , \wRegInTop_4_6[13] , \wRegInTop_4_6[12] , 
        \wRegInTop_4_6[11] , \wRegInTop_4_6[10] , \wRegInTop_4_6[9] , 
        \wRegInTop_4_6[8] , \wRegInTop_4_6[7] , \wRegInTop_4_6[6] , 
        \wRegInTop_4_6[5] , \wRegInTop_4_6[4] , \wRegInTop_4_6[3] , 
        \wRegInTop_4_6[2] , \wRegInTop_4_6[1] , \wRegInTop_4_6[0] }), .R_WR(
        \wRegEnTop_4_7[0] ), .R_In({\wRegOut_4_7[31] , \wRegOut_4_7[30] , 
        \wRegOut_4_7[29] , \wRegOut_4_7[28] , \wRegOut_4_7[27] , 
        \wRegOut_4_7[26] , \wRegOut_4_7[25] , \wRegOut_4_7[24] , 
        \wRegOut_4_7[23] , \wRegOut_4_7[22] , \wRegOut_4_7[21] , 
        \wRegOut_4_7[20] , \wRegOut_4_7[19] , \wRegOut_4_7[18] , 
        \wRegOut_4_7[17] , \wRegOut_4_7[16] , \wRegOut_4_7[15] , 
        \wRegOut_4_7[14] , \wRegOut_4_7[13] , \wRegOut_4_7[12] , 
        \wRegOut_4_7[11] , \wRegOut_4_7[10] , \wRegOut_4_7[9] , 
        \wRegOut_4_7[8] , \wRegOut_4_7[7] , \wRegOut_4_7[6] , \wRegOut_4_7[5] , 
        \wRegOut_4_7[4] , \wRegOut_4_7[3] , \wRegOut_4_7[2] , \wRegOut_4_7[1] , 
        \wRegOut_4_7[0] }), .R_Out({\wRegInTop_4_7[31] , \wRegInTop_4_7[30] , 
        \wRegInTop_4_7[29] , \wRegInTop_4_7[28] , \wRegInTop_4_7[27] , 
        \wRegInTop_4_7[26] , \wRegInTop_4_7[25] , \wRegInTop_4_7[24] , 
        \wRegInTop_4_7[23] , \wRegInTop_4_7[22] , \wRegInTop_4_7[21] , 
        \wRegInTop_4_7[20] , \wRegInTop_4_7[19] , \wRegInTop_4_7[18] , 
        \wRegInTop_4_7[17] , \wRegInTop_4_7[16] , \wRegInTop_4_7[15] , 
        \wRegInTop_4_7[14] , \wRegInTop_4_7[13] , \wRegInTop_4_7[12] , 
        \wRegInTop_4_7[11] , \wRegInTop_4_7[10] , \wRegInTop_4_7[9] , 
        \wRegInTop_4_7[8] , \wRegInTop_4_7[7] , \wRegInTop_4_7[6] , 
        \wRegInTop_4_7[5] , \wRegInTop_4_7[4] , \wRegInTop_4_7[3] , 
        \wRegInTop_4_7[2] , \wRegInTop_4_7[1] , \wRegInTop_4_7[0] }) );
    BHeap_Node_WIDTH32 BHN_4_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_9[0] ), .P_In({\wRegOut_4_9[31] , 
        \wRegOut_4_9[30] , \wRegOut_4_9[29] , \wRegOut_4_9[28] , 
        \wRegOut_4_9[27] , \wRegOut_4_9[26] , \wRegOut_4_9[25] , 
        \wRegOut_4_9[24] , \wRegOut_4_9[23] , \wRegOut_4_9[22] , 
        \wRegOut_4_9[21] , \wRegOut_4_9[20] , \wRegOut_4_9[19] , 
        \wRegOut_4_9[18] , \wRegOut_4_9[17] , \wRegOut_4_9[16] , 
        \wRegOut_4_9[15] , \wRegOut_4_9[14] , \wRegOut_4_9[13] , 
        \wRegOut_4_9[12] , \wRegOut_4_9[11] , \wRegOut_4_9[10] , 
        \wRegOut_4_9[9] , \wRegOut_4_9[8] , \wRegOut_4_9[7] , \wRegOut_4_9[6] , 
        \wRegOut_4_9[5] , \wRegOut_4_9[4] , \wRegOut_4_9[3] , \wRegOut_4_9[2] , 
        \wRegOut_4_9[1] , \wRegOut_4_9[0] }), .P_Out({\wRegInBot_4_9[31] , 
        \wRegInBot_4_9[30] , \wRegInBot_4_9[29] , \wRegInBot_4_9[28] , 
        \wRegInBot_4_9[27] , \wRegInBot_4_9[26] , \wRegInBot_4_9[25] , 
        \wRegInBot_4_9[24] , \wRegInBot_4_9[23] , \wRegInBot_4_9[22] , 
        \wRegInBot_4_9[21] , \wRegInBot_4_9[20] , \wRegInBot_4_9[19] , 
        \wRegInBot_4_9[18] , \wRegInBot_4_9[17] , \wRegInBot_4_9[16] , 
        \wRegInBot_4_9[15] , \wRegInBot_4_9[14] , \wRegInBot_4_9[13] , 
        \wRegInBot_4_9[12] , \wRegInBot_4_9[11] , \wRegInBot_4_9[10] , 
        \wRegInBot_4_9[9] , \wRegInBot_4_9[8] , \wRegInBot_4_9[7] , 
        \wRegInBot_4_9[6] , \wRegInBot_4_9[5] , \wRegInBot_4_9[4] , 
        \wRegInBot_4_9[3] , \wRegInBot_4_9[2] , \wRegInBot_4_9[1] , 
        \wRegInBot_4_9[0] }), .L_WR(\wRegEnTop_5_18[0] ), .L_In({
        \wRegOut_5_18[31] , \wRegOut_5_18[30] , \wRegOut_5_18[29] , 
        \wRegOut_5_18[28] , \wRegOut_5_18[27] , \wRegOut_5_18[26] , 
        \wRegOut_5_18[25] , \wRegOut_5_18[24] , \wRegOut_5_18[23] , 
        \wRegOut_5_18[22] , \wRegOut_5_18[21] , \wRegOut_5_18[20] , 
        \wRegOut_5_18[19] , \wRegOut_5_18[18] , \wRegOut_5_18[17] , 
        \wRegOut_5_18[16] , \wRegOut_5_18[15] , \wRegOut_5_18[14] , 
        \wRegOut_5_18[13] , \wRegOut_5_18[12] , \wRegOut_5_18[11] , 
        \wRegOut_5_18[10] , \wRegOut_5_18[9] , \wRegOut_5_18[8] , 
        \wRegOut_5_18[7] , \wRegOut_5_18[6] , \wRegOut_5_18[5] , 
        \wRegOut_5_18[4] , \wRegOut_5_18[3] , \wRegOut_5_18[2] , 
        \wRegOut_5_18[1] , \wRegOut_5_18[0] }), .L_Out({\wRegInTop_5_18[31] , 
        \wRegInTop_5_18[30] , \wRegInTop_5_18[29] , \wRegInTop_5_18[28] , 
        \wRegInTop_5_18[27] , \wRegInTop_5_18[26] , \wRegInTop_5_18[25] , 
        \wRegInTop_5_18[24] , \wRegInTop_5_18[23] , \wRegInTop_5_18[22] , 
        \wRegInTop_5_18[21] , \wRegInTop_5_18[20] , \wRegInTop_5_18[19] , 
        \wRegInTop_5_18[18] , \wRegInTop_5_18[17] , \wRegInTop_5_18[16] , 
        \wRegInTop_5_18[15] , \wRegInTop_5_18[14] , \wRegInTop_5_18[13] , 
        \wRegInTop_5_18[12] , \wRegInTop_5_18[11] , \wRegInTop_5_18[10] , 
        \wRegInTop_5_18[9] , \wRegInTop_5_18[8] , \wRegInTop_5_18[7] , 
        \wRegInTop_5_18[6] , \wRegInTop_5_18[5] , \wRegInTop_5_18[4] , 
        \wRegInTop_5_18[3] , \wRegInTop_5_18[2] , \wRegInTop_5_18[1] , 
        \wRegInTop_5_18[0] }), .R_WR(\wRegEnTop_5_19[0] ), .R_In({
        \wRegOut_5_19[31] , \wRegOut_5_19[30] , \wRegOut_5_19[29] , 
        \wRegOut_5_19[28] , \wRegOut_5_19[27] , \wRegOut_5_19[26] , 
        \wRegOut_5_19[25] , \wRegOut_5_19[24] , \wRegOut_5_19[23] , 
        \wRegOut_5_19[22] , \wRegOut_5_19[21] , \wRegOut_5_19[20] , 
        \wRegOut_5_19[19] , \wRegOut_5_19[18] , \wRegOut_5_19[17] , 
        \wRegOut_5_19[16] , \wRegOut_5_19[15] , \wRegOut_5_19[14] , 
        \wRegOut_5_19[13] , \wRegOut_5_19[12] , \wRegOut_5_19[11] , 
        \wRegOut_5_19[10] , \wRegOut_5_19[9] , \wRegOut_5_19[8] , 
        \wRegOut_5_19[7] , \wRegOut_5_19[6] , \wRegOut_5_19[5] , 
        \wRegOut_5_19[4] , \wRegOut_5_19[3] , \wRegOut_5_19[2] , 
        \wRegOut_5_19[1] , \wRegOut_5_19[0] }), .R_Out({\wRegInTop_5_19[31] , 
        \wRegInTop_5_19[30] , \wRegInTop_5_19[29] , \wRegInTop_5_19[28] , 
        \wRegInTop_5_19[27] , \wRegInTop_5_19[26] , \wRegInTop_5_19[25] , 
        \wRegInTop_5_19[24] , \wRegInTop_5_19[23] , \wRegInTop_5_19[22] , 
        \wRegInTop_5_19[21] , \wRegInTop_5_19[20] , \wRegInTop_5_19[19] , 
        \wRegInTop_5_19[18] , \wRegInTop_5_19[17] , \wRegInTop_5_19[16] , 
        \wRegInTop_5_19[15] , \wRegInTop_5_19[14] , \wRegInTop_5_19[13] , 
        \wRegInTop_5_19[12] , \wRegInTop_5_19[11] , \wRegInTop_5_19[10] , 
        \wRegInTop_5_19[9] , \wRegInTop_5_19[8] , \wRegInTop_5_19[7] , 
        \wRegInTop_5_19[6] , \wRegInTop_5_19[5] , \wRegInTop_5_19[4] , 
        \wRegInTop_5_19[3] , \wRegInTop_5_19[2] , \wRegInTop_5_19[1] , 
        \wRegInTop_5_19[0] }) );
    BHeap_Node_WIDTH32 BHN_4_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_10[0] ), .P_In({\wRegOut_4_10[31] , 
        \wRegOut_4_10[30] , \wRegOut_4_10[29] , \wRegOut_4_10[28] , 
        \wRegOut_4_10[27] , \wRegOut_4_10[26] , \wRegOut_4_10[25] , 
        \wRegOut_4_10[24] , \wRegOut_4_10[23] , \wRegOut_4_10[22] , 
        \wRegOut_4_10[21] , \wRegOut_4_10[20] , \wRegOut_4_10[19] , 
        \wRegOut_4_10[18] , \wRegOut_4_10[17] , \wRegOut_4_10[16] , 
        \wRegOut_4_10[15] , \wRegOut_4_10[14] , \wRegOut_4_10[13] , 
        \wRegOut_4_10[12] , \wRegOut_4_10[11] , \wRegOut_4_10[10] , 
        \wRegOut_4_10[9] , \wRegOut_4_10[8] , \wRegOut_4_10[7] , 
        \wRegOut_4_10[6] , \wRegOut_4_10[5] , \wRegOut_4_10[4] , 
        \wRegOut_4_10[3] , \wRegOut_4_10[2] , \wRegOut_4_10[1] , 
        \wRegOut_4_10[0] }), .P_Out({\wRegInBot_4_10[31] , 
        \wRegInBot_4_10[30] , \wRegInBot_4_10[29] , \wRegInBot_4_10[28] , 
        \wRegInBot_4_10[27] , \wRegInBot_4_10[26] , \wRegInBot_4_10[25] , 
        \wRegInBot_4_10[24] , \wRegInBot_4_10[23] , \wRegInBot_4_10[22] , 
        \wRegInBot_4_10[21] , \wRegInBot_4_10[20] , \wRegInBot_4_10[19] , 
        \wRegInBot_4_10[18] , \wRegInBot_4_10[17] , \wRegInBot_4_10[16] , 
        \wRegInBot_4_10[15] , \wRegInBot_4_10[14] , \wRegInBot_4_10[13] , 
        \wRegInBot_4_10[12] , \wRegInBot_4_10[11] , \wRegInBot_4_10[10] , 
        \wRegInBot_4_10[9] , \wRegInBot_4_10[8] , \wRegInBot_4_10[7] , 
        \wRegInBot_4_10[6] , \wRegInBot_4_10[5] , \wRegInBot_4_10[4] , 
        \wRegInBot_4_10[3] , \wRegInBot_4_10[2] , \wRegInBot_4_10[1] , 
        \wRegInBot_4_10[0] }), .L_WR(\wRegEnTop_5_20[0] ), .L_In({
        \wRegOut_5_20[31] , \wRegOut_5_20[30] , \wRegOut_5_20[29] , 
        \wRegOut_5_20[28] , \wRegOut_5_20[27] , \wRegOut_5_20[26] , 
        \wRegOut_5_20[25] , \wRegOut_5_20[24] , \wRegOut_5_20[23] , 
        \wRegOut_5_20[22] , \wRegOut_5_20[21] , \wRegOut_5_20[20] , 
        \wRegOut_5_20[19] , \wRegOut_5_20[18] , \wRegOut_5_20[17] , 
        \wRegOut_5_20[16] , \wRegOut_5_20[15] , \wRegOut_5_20[14] , 
        \wRegOut_5_20[13] , \wRegOut_5_20[12] , \wRegOut_5_20[11] , 
        \wRegOut_5_20[10] , \wRegOut_5_20[9] , \wRegOut_5_20[8] , 
        \wRegOut_5_20[7] , \wRegOut_5_20[6] , \wRegOut_5_20[5] , 
        \wRegOut_5_20[4] , \wRegOut_5_20[3] , \wRegOut_5_20[2] , 
        \wRegOut_5_20[1] , \wRegOut_5_20[0] }), .L_Out({\wRegInTop_5_20[31] , 
        \wRegInTop_5_20[30] , \wRegInTop_5_20[29] , \wRegInTop_5_20[28] , 
        \wRegInTop_5_20[27] , \wRegInTop_5_20[26] , \wRegInTop_5_20[25] , 
        \wRegInTop_5_20[24] , \wRegInTop_5_20[23] , \wRegInTop_5_20[22] , 
        \wRegInTop_5_20[21] , \wRegInTop_5_20[20] , \wRegInTop_5_20[19] , 
        \wRegInTop_5_20[18] , \wRegInTop_5_20[17] , \wRegInTop_5_20[16] , 
        \wRegInTop_5_20[15] , \wRegInTop_5_20[14] , \wRegInTop_5_20[13] , 
        \wRegInTop_5_20[12] , \wRegInTop_5_20[11] , \wRegInTop_5_20[10] , 
        \wRegInTop_5_20[9] , \wRegInTop_5_20[8] , \wRegInTop_5_20[7] , 
        \wRegInTop_5_20[6] , \wRegInTop_5_20[5] , \wRegInTop_5_20[4] , 
        \wRegInTop_5_20[3] , \wRegInTop_5_20[2] , \wRegInTop_5_20[1] , 
        \wRegInTop_5_20[0] }), .R_WR(\wRegEnTop_5_21[0] ), .R_In({
        \wRegOut_5_21[31] , \wRegOut_5_21[30] , \wRegOut_5_21[29] , 
        \wRegOut_5_21[28] , \wRegOut_5_21[27] , \wRegOut_5_21[26] , 
        \wRegOut_5_21[25] , \wRegOut_5_21[24] , \wRegOut_5_21[23] , 
        \wRegOut_5_21[22] , \wRegOut_5_21[21] , \wRegOut_5_21[20] , 
        \wRegOut_5_21[19] , \wRegOut_5_21[18] , \wRegOut_5_21[17] , 
        \wRegOut_5_21[16] , \wRegOut_5_21[15] , \wRegOut_5_21[14] , 
        \wRegOut_5_21[13] , \wRegOut_5_21[12] , \wRegOut_5_21[11] , 
        \wRegOut_5_21[10] , \wRegOut_5_21[9] , \wRegOut_5_21[8] , 
        \wRegOut_5_21[7] , \wRegOut_5_21[6] , \wRegOut_5_21[5] , 
        \wRegOut_5_21[4] , \wRegOut_5_21[3] , \wRegOut_5_21[2] , 
        \wRegOut_5_21[1] , \wRegOut_5_21[0] }), .R_Out({\wRegInTop_5_21[31] , 
        \wRegInTop_5_21[30] , \wRegInTop_5_21[29] , \wRegInTop_5_21[28] , 
        \wRegInTop_5_21[27] , \wRegInTop_5_21[26] , \wRegInTop_5_21[25] , 
        \wRegInTop_5_21[24] , \wRegInTop_5_21[23] , \wRegInTop_5_21[22] , 
        \wRegInTop_5_21[21] , \wRegInTop_5_21[20] , \wRegInTop_5_21[19] , 
        \wRegInTop_5_21[18] , \wRegInTop_5_21[17] , \wRegInTop_5_21[16] , 
        \wRegInTop_5_21[15] , \wRegInTop_5_21[14] , \wRegInTop_5_21[13] , 
        \wRegInTop_5_21[12] , \wRegInTop_5_21[11] , \wRegInTop_5_21[10] , 
        \wRegInTop_5_21[9] , \wRegInTop_5_21[8] , \wRegInTop_5_21[7] , 
        \wRegInTop_5_21[6] , \wRegInTop_5_21[5] , \wRegInTop_5_21[4] , 
        \wRegInTop_5_21[3] , \wRegInTop_5_21[2] , \wRegInTop_5_21[1] , 
        \wRegInTop_5_21[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink19[31] , \ScanLink19[30] , \ScanLink19[29] , 
        \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , \ScanLink19[25] , 
        \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , \ScanLink19[21] , 
        \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , \ScanLink19[17] , 
        \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , \ScanLink19[13] , 
        \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , \ScanLink19[9] , 
        \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , \ScanLink19[5] , 
        \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , \ScanLink19[1] , 
        \ScanLink19[0] }), .ScanOut({\ScanLink18[31] , \ScanLink18[30] , 
        \ScanLink18[29] , \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , 
        \ScanLink18[25] , \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , 
        \ScanLink18[21] , \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , 
        \ScanLink18[17] , \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , 
        \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , 
        \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , 
        \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , 
        \ScanLink18[1] , \ScanLink18[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_3[31] , \wRegOut_4_3[30] , \wRegOut_4_3[29] , 
        \wRegOut_4_3[28] , \wRegOut_4_3[27] , \wRegOut_4_3[26] , 
        \wRegOut_4_3[25] , \wRegOut_4_3[24] , \wRegOut_4_3[23] , 
        \wRegOut_4_3[22] , \wRegOut_4_3[21] , \wRegOut_4_3[20] , 
        \wRegOut_4_3[19] , \wRegOut_4_3[18] , \wRegOut_4_3[17] , 
        \wRegOut_4_3[16] , \wRegOut_4_3[15] , \wRegOut_4_3[14] , 
        \wRegOut_4_3[13] , \wRegOut_4_3[12] , \wRegOut_4_3[11] , 
        \wRegOut_4_3[10] , \wRegOut_4_3[9] , \wRegOut_4_3[8] , 
        \wRegOut_4_3[7] , \wRegOut_4_3[6] , \wRegOut_4_3[5] , \wRegOut_4_3[4] , 
        \wRegOut_4_3[3] , \wRegOut_4_3[2] , \wRegOut_4_3[1] , \wRegOut_4_3[0] 
        }), .Enable1(\wRegEnTop_4_3[0] ), .Enable2(\wRegEnBot_4_3[0] ), .In1({
        \wRegInTop_4_3[31] , \wRegInTop_4_3[30] , \wRegInTop_4_3[29] , 
        \wRegInTop_4_3[28] , \wRegInTop_4_3[27] , \wRegInTop_4_3[26] , 
        \wRegInTop_4_3[25] , \wRegInTop_4_3[24] , \wRegInTop_4_3[23] , 
        \wRegInTop_4_3[22] , \wRegInTop_4_3[21] , \wRegInTop_4_3[20] , 
        \wRegInTop_4_3[19] , \wRegInTop_4_3[18] , \wRegInTop_4_3[17] , 
        \wRegInTop_4_3[16] , \wRegInTop_4_3[15] , \wRegInTop_4_3[14] , 
        \wRegInTop_4_3[13] , \wRegInTop_4_3[12] , \wRegInTop_4_3[11] , 
        \wRegInTop_4_3[10] , \wRegInTop_4_3[9] , \wRegInTop_4_3[8] , 
        \wRegInTop_4_3[7] , \wRegInTop_4_3[6] , \wRegInTop_4_3[5] , 
        \wRegInTop_4_3[4] , \wRegInTop_4_3[3] , \wRegInTop_4_3[2] , 
        \wRegInTop_4_3[1] , \wRegInTop_4_3[0] }), .In2({\wRegInBot_4_3[31] , 
        \wRegInBot_4_3[30] , \wRegInBot_4_3[29] , \wRegInBot_4_3[28] , 
        \wRegInBot_4_3[27] , \wRegInBot_4_3[26] , \wRegInBot_4_3[25] , 
        \wRegInBot_4_3[24] , \wRegInBot_4_3[23] , \wRegInBot_4_3[22] , 
        \wRegInBot_4_3[21] , \wRegInBot_4_3[20] , \wRegInBot_4_3[19] , 
        \wRegInBot_4_3[18] , \wRegInBot_4_3[17] , \wRegInBot_4_3[16] , 
        \wRegInBot_4_3[15] , \wRegInBot_4_3[14] , \wRegInBot_4_3[13] , 
        \wRegInBot_4_3[12] , \wRegInBot_4_3[11] , \wRegInBot_4_3[10] , 
        \wRegInBot_4_3[9] , \wRegInBot_4_3[8] , \wRegInBot_4_3[7] , 
        \wRegInBot_4_3[6] , \wRegInBot_4_3[5] , \wRegInBot_4_3[4] , 
        \wRegInBot_4_3[3] , \wRegInBot_4_3[2] , \wRegInBot_4_3[1] , 
        \wRegInBot_4_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink35[31] , \ScanLink35[30] , \ScanLink35[29] , 
        \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , \ScanLink35[25] , 
        \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , \ScanLink35[21] , 
        \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , \ScanLink35[17] , 
        \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , \ScanLink35[13] , 
        \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , \ScanLink35[9] , 
        \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , \ScanLink35[5] , 
        \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , \ScanLink35[1] , 
        \ScanLink35[0] }), .ScanOut({\ScanLink34[31] , \ScanLink34[30] , 
        \ScanLink34[29] , \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , 
        \ScanLink34[25] , \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , 
        \ScanLink34[21] , \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , 
        \ScanLink34[17] , \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , 
        \ScanLink34[13] , \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , 
        \ScanLink34[9] , \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , 
        \ScanLink34[5] , \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , 
        \ScanLink34[1] , \ScanLink34[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_3[31] , \wRegOut_5_3[30] , \wRegOut_5_3[29] , 
        \wRegOut_5_3[28] , \wRegOut_5_3[27] , \wRegOut_5_3[26] , 
        \wRegOut_5_3[25] , \wRegOut_5_3[24] , \wRegOut_5_3[23] , 
        \wRegOut_5_3[22] , \wRegOut_5_3[21] , \wRegOut_5_3[20] , 
        \wRegOut_5_3[19] , \wRegOut_5_3[18] , \wRegOut_5_3[17] , 
        \wRegOut_5_3[16] , \wRegOut_5_3[15] , \wRegOut_5_3[14] , 
        \wRegOut_5_3[13] , \wRegOut_5_3[12] , \wRegOut_5_3[11] , 
        \wRegOut_5_3[10] , \wRegOut_5_3[9] , \wRegOut_5_3[8] , 
        \wRegOut_5_3[7] , \wRegOut_5_3[6] , \wRegOut_5_3[5] , \wRegOut_5_3[4] , 
        \wRegOut_5_3[3] , \wRegOut_5_3[2] , \wRegOut_5_3[1] , \wRegOut_5_3[0] 
        }), .Enable1(\wRegEnTop_5_3[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_3[31] , \wRegInTop_5_3[30] , \wRegInTop_5_3[29] , 
        \wRegInTop_5_3[28] , \wRegInTop_5_3[27] , \wRegInTop_5_3[26] , 
        \wRegInTop_5_3[25] , \wRegInTop_5_3[24] , \wRegInTop_5_3[23] , 
        \wRegInTop_5_3[22] , \wRegInTop_5_3[21] , \wRegInTop_5_3[20] , 
        \wRegInTop_5_3[19] , \wRegInTop_5_3[18] , \wRegInTop_5_3[17] , 
        \wRegInTop_5_3[16] , \wRegInTop_5_3[15] , \wRegInTop_5_3[14] , 
        \wRegInTop_5_3[13] , \wRegInTop_5_3[12] , \wRegInTop_5_3[11] , 
        \wRegInTop_5_3[10] , \wRegInTop_5_3[9] , \wRegInTop_5_3[8] , 
        \wRegInTop_5_3[7] , \wRegInTop_5_3[6] , \wRegInTop_5_3[5] , 
        \wRegInTop_5_3[4] , \wRegInTop_5_3[3] , \wRegInTop_5_3[2] , 
        \wRegInTop_5_3[1] , \wRegInTop_5_3[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_22 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink54[31] , \ScanLink54[30] , \ScanLink54[29] , 
        \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , \ScanLink54[25] , 
        \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , \ScanLink54[21] , 
        \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , \ScanLink54[17] , 
        \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , \ScanLink54[13] , 
        \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , \ScanLink54[9] , 
        \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , \ScanLink54[5] , 
        \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , \ScanLink54[1] , 
        \ScanLink54[0] }), .ScanOut({\ScanLink53[31] , \ScanLink53[30] , 
        \ScanLink53[29] , \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , 
        \ScanLink53[25] , \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , 
        \ScanLink53[21] , \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , 
        \ScanLink53[17] , \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , 
        \ScanLink53[13] , \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , 
        \ScanLink53[9] , \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , 
        \ScanLink53[5] , \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , 
        \ScanLink53[1] , \ScanLink53[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_22[31] , \wRegOut_5_22[30] , 
        \wRegOut_5_22[29] , \wRegOut_5_22[28] , \wRegOut_5_22[27] , 
        \wRegOut_5_22[26] , \wRegOut_5_22[25] , \wRegOut_5_22[24] , 
        \wRegOut_5_22[23] , \wRegOut_5_22[22] , \wRegOut_5_22[21] , 
        \wRegOut_5_22[20] , \wRegOut_5_22[19] , \wRegOut_5_22[18] , 
        \wRegOut_5_22[17] , \wRegOut_5_22[16] , \wRegOut_5_22[15] , 
        \wRegOut_5_22[14] , \wRegOut_5_22[13] , \wRegOut_5_22[12] , 
        \wRegOut_5_22[11] , \wRegOut_5_22[10] , \wRegOut_5_22[9] , 
        \wRegOut_5_22[8] , \wRegOut_5_22[7] , \wRegOut_5_22[6] , 
        \wRegOut_5_22[5] , \wRegOut_5_22[4] , \wRegOut_5_22[3] , 
        \wRegOut_5_22[2] , \wRegOut_5_22[1] , \wRegOut_5_22[0] }), .Enable1(
        \wRegEnTop_5_22[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_22[31] , 
        \wRegInTop_5_22[30] , \wRegInTop_5_22[29] , \wRegInTop_5_22[28] , 
        \wRegInTop_5_22[27] , \wRegInTop_5_22[26] , \wRegInTop_5_22[25] , 
        \wRegInTop_5_22[24] , \wRegInTop_5_22[23] , \wRegInTop_5_22[22] , 
        \wRegInTop_5_22[21] , \wRegInTop_5_22[20] , \wRegInTop_5_22[19] , 
        \wRegInTop_5_22[18] , \wRegInTop_5_22[17] , \wRegInTop_5_22[16] , 
        \wRegInTop_5_22[15] , \wRegInTop_5_22[14] , \wRegInTop_5_22[13] , 
        \wRegInTop_5_22[12] , \wRegInTop_5_22[11] , \wRegInTop_5_22[10] , 
        \wRegInTop_5_22[9] , \wRegInTop_5_22[8] , \wRegInTop_5_22[7] , 
        \wRegInTop_5_22[6] , \wRegInTop_5_22[5] , \wRegInTop_5_22[4] , 
        \wRegInTop_5_22[3] , \wRegInTop_5_22[2] , \wRegInTop_5_22[1] , 
        \wRegInTop_5_22[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_4_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_1[0] ), .P_In({\wRegOut_4_1[31] , 
        \wRegOut_4_1[30] , \wRegOut_4_1[29] , \wRegOut_4_1[28] , 
        \wRegOut_4_1[27] , \wRegOut_4_1[26] , \wRegOut_4_1[25] , 
        \wRegOut_4_1[24] , \wRegOut_4_1[23] , \wRegOut_4_1[22] , 
        \wRegOut_4_1[21] , \wRegOut_4_1[20] , \wRegOut_4_1[19] , 
        \wRegOut_4_1[18] , \wRegOut_4_1[17] , \wRegOut_4_1[16] , 
        \wRegOut_4_1[15] , \wRegOut_4_1[14] , \wRegOut_4_1[13] , 
        \wRegOut_4_1[12] , \wRegOut_4_1[11] , \wRegOut_4_1[10] , 
        \wRegOut_4_1[9] , \wRegOut_4_1[8] , \wRegOut_4_1[7] , \wRegOut_4_1[6] , 
        \wRegOut_4_1[5] , \wRegOut_4_1[4] , \wRegOut_4_1[3] , \wRegOut_4_1[2] , 
        \wRegOut_4_1[1] , \wRegOut_4_1[0] }), .P_Out({\wRegInBot_4_1[31] , 
        \wRegInBot_4_1[30] , \wRegInBot_4_1[29] , \wRegInBot_4_1[28] , 
        \wRegInBot_4_1[27] , \wRegInBot_4_1[26] , \wRegInBot_4_1[25] , 
        \wRegInBot_4_1[24] , \wRegInBot_4_1[23] , \wRegInBot_4_1[22] , 
        \wRegInBot_4_1[21] , \wRegInBot_4_1[20] , \wRegInBot_4_1[19] , 
        \wRegInBot_4_1[18] , \wRegInBot_4_1[17] , \wRegInBot_4_1[16] , 
        \wRegInBot_4_1[15] , \wRegInBot_4_1[14] , \wRegInBot_4_1[13] , 
        \wRegInBot_4_1[12] , \wRegInBot_4_1[11] , \wRegInBot_4_1[10] , 
        \wRegInBot_4_1[9] , \wRegInBot_4_1[8] , \wRegInBot_4_1[7] , 
        \wRegInBot_4_1[6] , \wRegInBot_4_1[5] , \wRegInBot_4_1[4] , 
        \wRegInBot_4_1[3] , \wRegInBot_4_1[2] , \wRegInBot_4_1[1] , 
        \wRegInBot_4_1[0] }), .L_WR(\wRegEnTop_5_2[0] ), .L_In({
        \wRegOut_5_2[31] , \wRegOut_5_2[30] , \wRegOut_5_2[29] , 
        \wRegOut_5_2[28] , \wRegOut_5_2[27] , \wRegOut_5_2[26] , 
        \wRegOut_5_2[25] , \wRegOut_5_2[24] , \wRegOut_5_2[23] , 
        \wRegOut_5_2[22] , \wRegOut_5_2[21] , \wRegOut_5_2[20] , 
        \wRegOut_5_2[19] , \wRegOut_5_2[18] , \wRegOut_5_2[17] , 
        \wRegOut_5_2[16] , \wRegOut_5_2[15] , \wRegOut_5_2[14] , 
        \wRegOut_5_2[13] , \wRegOut_5_2[12] , \wRegOut_5_2[11] , 
        \wRegOut_5_2[10] , \wRegOut_5_2[9] , \wRegOut_5_2[8] , 
        \wRegOut_5_2[7] , \wRegOut_5_2[6] , \wRegOut_5_2[5] , \wRegOut_5_2[4] , 
        \wRegOut_5_2[3] , \wRegOut_5_2[2] , \wRegOut_5_2[1] , \wRegOut_5_2[0] 
        }), .L_Out({\wRegInTop_5_2[31] , \wRegInTop_5_2[30] , 
        \wRegInTop_5_2[29] , \wRegInTop_5_2[28] , \wRegInTop_5_2[27] , 
        \wRegInTop_5_2[26] , \wRegInTop_5_2[25] , \wRegInTop_5_2[24] , 
        \wRegInTop_5_2[23] , \wRegInTop_5_2[22] , \wRegInTop_5_2[21] , 
        \wRegInTop_5_2[20] , \wRegInTop_5_2[19] , \wRegInTop_5_2[18] , 
        \wRegInTop_5_2[17] , \wRegInTop_5_2[16] , \wRegInTop_5_2[15] , 
        \wRegInTop_5_2[14] , \wRegInTop_5_2[13] , \wRegInTop_5_2[12] , 
        \wRegInTop_5_2[11] , \wRegInTop_5_2[10] , \wRegInTop_5_2[9] , 
        \wRegInTop_5_2[8] , \wRegInTop_5_2[7] , \wRegInTop_5_2[6] , 
        \wRegInTop_5_2[5] , \wRegInTop_5_2[4] , \wRegInTop_5_2[3] , 
        \wRegInTop_5_2[2] , \wRegInTop_5_2[1] , \wRegInTop_5_2[0] }), .R_WR(
        \wRegEnTop_5_3[0] ), .R_In({\wRegOut_5_3[31] , \wRegOut_5_3[30] , 
        \wRegOut_5_3[29] , \wRegOut_5_3[28] , \wRegOut_5_3[27] , 
        \wRegOut_5_3[26] , \wRegOut_5_3[25] , \wRegOut_5_3[24] , 
        \wRegOut_5_3[23] , \wRegOut_5_3[22] , \wRegOut_5_3[21] , 
        \wRegOut_5_3[20] , \wRegOut_5_3[19] , \wRegOut_5_3[18] , 
        \wRegOut_5_3[17] , \wRegOut_5_3[16] , \wRegOut_5_3[15] , 
        \wRegOut_5_3[14] , \wRegOut_5_3[13] , \wRegOut_5_3[12] , 
        \wRegOut_5_3[11] , \wRegOut_5_3[10] , \wRegOut_5_3[9] , 
        \wRegOut_5_3[8] , \wRegOut_5_3[7] , \wRegOut_5_3[6] , \wRegOut_5_3[5] , 
        \wRegOut_5_3[4] , \wRegOut_5_3[3] , \wRegOut_5_3[2] , \wRegOut_5_3[1] , 
        \wRegOut_5_3[0] }), .R_Out({\wRegInTop_5_3[31] , \wRegInTop_5_3[30] , 
        \wRegInTop_5_3[29] , \wRegInTop_5_3[28] , \wRegInTop_5_3[27] , 
        \wRegInTop_5_3[26] , \wRegInTop_5_3[25] , \wRegInTop_5_3[24] , 
        \wRegInTop_5_3[23] , \wRegInTop_5_3[22] , \wRegInTop_5_3[21] , 
        \wRegInTop_5_3[20] , \wRegInTop_5_3[19] , \wRegInTop_5_3[18] , 
        \wRegInTop_5_3[17] , \wRegInTop_5_3[16] , \wRegInTop_5_3[15] , 
        \wRegInTop_5_3[14] , \wRegInTop_5_3[13] , \wRegInTop_5_3[12] , 
        \wRegInTop_5_3[11] , \wRegInTop_5_3[10] , \wRegInTop_5_3[9] , 
        \wRegInTop_5_3[8] , \wRegInTop_5_3[7] , \wRegInTop_5_3[6] , 
        \wRegInTop_5_3[5] , \wRegInTop_5_3[4] , \wRegInTop_5_3[3] , 
        \wRegInTop_5_3[2] , \wRegInTop_5_3[1] , \wRegInTop_5_3[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_16 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink48[31] , \ScanLink48[30] , \ScanLink48[29] , 
        \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , \ScanLink48[25] , 
        \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , \ScanLink48[21] , 
        \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , \ScanLink48[17] , 
        \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , \ScanLink48[13] , 
        \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , \ScanLink48[9] , 
        \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , \ScanLink48[5] , 
        \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , \ScanLink48[1] , 
        \ScanLink48[0] }), .ScanOut({\ScanLink47[31] , \ScanLink47[30] , 
        \ScanLink47[29] , \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , 
        \ScanLink47[25] , \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , 
        \ScanLink47[21] , \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , 
        \ScanLink47[17] , \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , 
        \ScanLink47[13] , \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , 
        \ScanLink47[9] , \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , 
        \ScanLink47[5] , \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , 
        \ScanLink47[1] , \ScanLink47[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_16[31] , \wRegOut_5_16[30] , 
        \wRegOut_5_16[29] , \wRegOut_5_16[28] , \wRegOut_5_16[27] , 
        \wRegOut_5_16[26] , \wRegOut_5_16[25] , \wRegOut_5_16[24] , 
        \wRegOut_5_16[23] , \wRegOut_5_16[22] , \wRegOut_5_16[21] , 
        \wRegOut_5_16[20] , \wRegOut_5_16[19] , \wRegOut_5_16[18] , 
        \wRegOut_5_16[17] , \wRegOut_5_16[16] , \wRegOut_5_16[15] , 
        \wRegOut_5_16[14] , \wRegOut_5_16[13] , \wRegOut_5_16[12] , 
        \wRegOut_5_16[11] , \wRegOut_5_16[10] , \wRegOut_5_16[9] , 
        \wRegOut_5_16[8] , \wRegOut_5_16[7] , \wRegOut_5_16[6] , 
        \wRegOut_5_16[5] , \wRegOut_5_16[4] , \wRegOut_5_16[3] , 
        \wRegOut_5_16[2] , \wRegOut_5_16[1] , \wRegOut_5_16[0] }), .Enable1(
        \wRegEnTop_5_16[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_16[31] , 
        \wRegInTop_5_16[30] , \wRegInTop_5_16[29] , \wRegInTop_5_16[28] , 
        \wRegInTop_5_16[27] , \wRegInTop_5_16[26] , \wRegInTop_5_16[25] , 
        \wRegInTop_5_16[24] , \wRegInTop_5_16[23] , \wRegInTop_5_16[22] , 
        \wRegInTop_5_16[21] , \wRegInTop_5_16[20] , \wRegInTop_5_16[19] , 
        \wRegInTop_5_16[18] , \wRegInTop_5_16[17] , \wRegInTop_5_16[16] , 
        \wRegInTop_5_16[15] , \wRegInTop_5_16[14] , \wRegInTop_5_16[13] , 
        \wRegInTop_5_16[12] , \wRegInTop_5_16[11] , \wRegInTop_5_16[10] , 
        \wRegInTop_5_16[9] , \wRegInTop_5_16[8] , \wRegInTop_5_16[7] , 
        \wRegInTop_5_16[6] , \wRegInTop_5_16[5] , \wRegInTop_5_16[4] , 
        \wRegInTop_5_16[3] , \wRegInTop_5_16[2] , \wRegInTop_5_16[1] , 
        \wRegInTop_5_16[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_31 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink63[31] , \ScanLink63[30] , \ScanLink63[29] , 
        \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , \ScanLink63[25] , 
        \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , \ScanLink63[21] , 
        \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , \ScanLink63[17] , 
        \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , \ScanLink63[13] , 
        \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , \ScanLink63[9] , 
        \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , \ScanLink63[5] , 
        \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , \ScanLink63[1] , 
        \ScanLink63[0] }), .ScanOut({\ScanLink62[31] , \ScanLink62[30] , 
        \ScanLink62[29] , \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , 
        \ScanLink62[25] , \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , 
        \ScanLink62[21] , \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , 
        \ScanLink62[17] , \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , 
        \ScanLink62[13] , \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , 
        \ScanLink62[9] , \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , 
        \ScanLink62[5] , \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , 
        \ScanLink62[1] , \ScanLink62[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_31[31] , \wRegOut_5_31[30] , 
        \wRegOut_5_31[29] , \wRegOut_5_31[28] , \wRegOut_5_31[27] , 
        \wRegOut_5_31[26] , \wRegOut_5_31[25] , \wRegOut_5_31[24] , 
        \wRegOut_5_31[23] , \wRegOut_5_31[22] , \wRegOut_5_31[21] , 
        \wRegOut_5_31[20] , \wRegOut_5_31[19] , \wRegOut_5_31[18] , 
        \wRegOut_5_31[17] , \wRegOut_5_31[16] , \wRegOut_5_31[15] , 
        \wRegOut_5_31[14] , \wRegOut_5_31[13] , \wRegOut_5_31[12] , 
        \wRegOut_5_31[11] , \wRegOut_5_31[10] , \wRegOut_5_31[9] , 
        \wRegOut_5_31[8] , \wRegOut_5_31[7] , \wRegOut_5_31[6] , 
        \wRegOut_5_31[5] , \wRegOut_5_31[4] , \wRegOut_5_31[3] , 
        \wRegOut_5_31[2] , \wRegOut_5_31[1] , \wRegOut_5_31[0] }), .Enable1(
        \wRegEnTop_5_31[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_31[31] , 
        \wRegInTop_5_31[30] , \wRegInTop_5_31[29] , \wRegInTop_5_31[28] , 
        \wRegInTop_5_31[27] , \wRegInTop_5_31[26] , \wRegInTop_5_31[25] , 
        \wRegInTop_5_31[24] , \wRegInTop_5_31[23] , \wRegInTop_5_31[22] , 
        \wRegInTop_5_31[21] , \wRegInTop_5_31[20] , \wRegInTop_5_31[19] , 
        \wRegInTop_5_31[18] , \wRegInTop_5_31[17] , \wRegInTop_5_31[16] , 
        \wRegInTop_5_31[15] , \wRegInTop_5_31[14] , \wRegInTop_5_31[13] , 
        \wRegInTop_5_31[12] , \wRegInTop_5_31[11] , \wRegInTop_5_31[10] , 
        \wRegInTop_5_31[9] , \wRegInTop_5_31[8] , \wRegInTop_5_31[7] , 
        \wRegInTop_5_31[6] , \wRegInTop_5_31[5] , \wRegInTop_5_31[4] , 
        \wRegInTop_5_31[3] , \wRegInTop_5_31[2] , \wRegInTop_5_31[1] , 
        \wRegInTop_5_31[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink8[31] , \ScanLink8[30] , \ScanLink8[29] , 
        \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , \ScanLink8[25] , 
        \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , \ScanLink8[21] , 
        \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , \ScanLink8[17] , 
        \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , \ScanLink8[13] , 
        \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , \ScanLink8[9] , 
        \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , \ScanLink8[5] , 
        \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , \ScanLink8[1] , 
        \ScanLink8[0] }), .ScanOut({\ScanLink7[31] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , 
        \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , 
        \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , 
        \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , 
        \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , 
        \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_0[31] , \wRegOut_3_0[30] , \wRegOut_3_0[29] , 
        \wRegOut_3_0[28] , \wRegOut_3_0[27] , \wRegOut_3_0[26] , 
        \wRegOut_3_0[25] , \wRegOut_3_0[24] , \wRegOut_3_0[23] , 
        \wRegOut_3_0[22] , \wRegOut_3_0[21] , \wRegOut_3_0[20] , 
        \wRegOut_3_0[19] , \wRegOut_3_0[18] , \wRegOut_3_0[17] , 
        \wRegOut_3_0[16] , \wRegOut_3_0[15] , \wRegOut_3_0[14] , 
        \wRegOut_3_0[13] , \wRegOut_3_0[12] , \wRegOut_3_0[11] , 
        \wRegOut_3_0[10] , \wRegOut_3_0[9] , \wRegOut_3_0[8] , 
        \wRegOut_3_0[7] , \wRegOut_3_0[6] , \wRegOut_3_0[5] , \wRegOut_3_0[4] , 
        \wRegOut_3_0[3] , \wRegOut_3_0[2] , \wRegOut_3_0[1] , \wRegOut_3_0[0] 
        }), .Enable1(\wRegEnTop_3_0[0] ), .Enable2(\wRegEnBot_3_0[0] ), .In1({
        \wRegInTop_3_0[31] , \wRegInTop_3_0[30] , \wRegInTop_3_0[29] , 
        \wRegInTop_3_0[28] , \wRegInTop_3_0[27] , \wRegInTop_3_0[26] , 
        \wRegInTop_3_0[25] , \wRegInTop_3_0[24] , \wRegInTop_3_0[23] , 
        \wRegInTop_3_0[22] , \wRegInTop_3_0[21] , \wRegInTop_3_0[20] , 
        \wRegInTop_3_0[19] , \wRegInTop_3_0[18] , \wRegInTop_3_0[17] , 
        \wRegInTop_3_0[16] , \wRegInTop_3_0[15] , \wRegInTop_3_0[14] , 
        \wRegInTop_3_0[13] , \wRegInTop_3_0[12] , \wRegInTop_3_0[11] , 
        \wRegInTop_3_0[10] , \wRegInTop_3_0[9] , \wRegInTop_3_0[8] , 
        \wRegInTop_3_0[7] , \wRegInTop_3_0[6] , \wRegInTop_3_0[5] , 
        \wRegInTop_3_0[4] , \wRegInTop_3_0[3] , \wRegInTop_3_0[2] , 
        \wRegInTop_3_0[1] , \wRegInTop_3_0[0] }), .In2({\wRegInBot_3_0[31] , 
        \wRegInBot_3_0[30] , \wRegInBot_3_0[29] , \wRegInBot_3_0[28] , 
        \wRegInBot_3_0[27] , \wRegInBot_3_0[26] , \wRegInBot_3_0[25] , 
        \wRegInBot_3_0[24] , \wRegInBot_3_0[23] , \wRegInBot_3_0[22] , 
        \wRegInBot_3_0[21] , \wRegInBot_3_0[20] , \wRegInBot_3_0[19] , 
        \wRegInBot_3_0[18] , \wRegInBot_3_0[17] , \wRegInBot_3_0[16] , 
        \wRegInBot_3_0[15] , \wRegInBot_3_0[14] , \wRegInBot_3_0[13] , 
        \wRegInBot_3_0[12] , \wRegInBot_3_0[11] , \wRegInBot_3_0[10] , 
        \wRegInBot_3_0[9] , \wRegInBot_3_0[8] , \wRegInBot_3_0[7] , 
        \wRegInBot_3_0[6] , \wRegInBot_3_0[5] , \wRegInBot_3_0[4] , 
        \wRegInBot_3_0[3] , \wRegInBot_3_0[2] , \wRegInBot_3_0[1] , 
        \wRegInBot_3_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_23 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink55[31] , \ScanLink55[30] , \ScanLink55[29] , 
        \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , \ScanLink55[25] , 
        \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , \ScanLink55[21] , 
        \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , \ScanLink55[17] , 
        \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , \ScanLink55[13] , 
        \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , \ScanLink55[9] , 
        \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , \ScanLink55[5] , 
        \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , \ScanLink55[1] , 
        \ScanLink55[0] }), .ScanOut({\ScanLink54[31] , \ScanLink54[30] , 
        \ScanLink54[29] , \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , 
        \ScanLink54[25] , \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , 
        \ScanLink54[21] , \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , 
        \ScanLink54[17] , \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , 
        \ScanLink54[13] , \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , 
        \ScanLink54[9] , \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , 
        \ScanLink54[5] , \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , 
        \ScanLink54[1] , \ScanLink54[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_23[31] , \wRegOut_5_23[30] , 
        \wRegOut_5_23[29] , \wRegOut_5_23[28] , \wRegOut_5_23[27] , 
        \wRegOut_5_23[26] , \wRegOut_5_23[25] , \wRegOut_5_23[24] , 
        \wRegOut_5_23[23] , \wRegOut_5_23[22] , \wRegOut_5_23[21] , 
        \wRegOut_5_23[20] , \wRegOut_5_23[19] , \wRegOut_5_23[18] , 
        \wRegOut_5_23[17] , \wRegOut_5_23[16] , \wRegOut_5_23[15] , 
        \wRegOut_5_23[14] , \wRegOut_5_23[13] , \wRegOut_5_23[12] , 
        \wRegOut_5_23[11] , \wRegOut_5_23[10] , \wRegOut_5_23[9] , 
        \wRegOut_5_23[8] , \wRegOut_5_23[7] , \wRegOut_5_23[6] , 
        \wRegOut_5_23[5] , \wRegOut_5_23[4] , \wRegOut_5_23[3] , 
        \wRegOut_5_23[2] , \wRegOut_5_23[1] , \wRegOut_5_23[0] }), .Enable1(
        \wRegEnTop_5_23[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_23[31] , 
        \wRegInTop_5_23[30] , \wRegInTop_5_23[29] , \wRegInTop_5_23[28] , 
        \wRegInTop_5_23[27] , \wRegInTop_5_23[26] , \wRegInTop_5_23[25] , 
        \wRegInTop_5_23[24] , \wRegInTop_5_23[23] , \wRegInTop_5_23[22] , 
        \wRegInTop_5_23[21] , \wRegInTop_5_23[20] , \wRegInTop_5_23[19] , 
        \wRegInTop_5_23[18] , \wRegInTop_5_23[17] , \wRegInTop_5_23[16] , 
        \wRegInTop_5_23[15] , \wRegInTop_5_23[14] , \wRegInTop_5_23[13] , 
        \wRegInTop_5_23[12] , \wRegInTop_5_23[11] , \wRegInTop_5_23[10] , 
        \wRegInTop_5_23[9] , \wRegInTop_5_23[8] , \wRegInTop_5_23[7] , 
        \wRegInTop_5_23[6] , \wRegInTop_5_23[5] , \wRegInTop_5_23[4] , 
        \wRegInTop_5_23[3] , \wRegInTop_5_23[2] , \wRegInTop_5_23[1] , 
        \wRegInTop_5_23[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_2[0] ), .P_WR(\wRegEnBot_2_2[0] ), .P_In({\wRegOut_2_2[31] , 
        \wRegOut_2_2[30] , \wRegOut_2_2[29] , \wRegOut_2_2[28] , 
        \wRegOut_2_2[27] , \wRegOut_2_2[26] , \wRegOut_2_2[25] , 
        \wRegOut_2_2[24] , \wRegOut_2_2[23] , \wRegOut_2_2[22] , 
        \wRegOut_2_2[21] , \wRegOut_2_2[20] , \wRegOut_2_2[19] , 
        \wRegOut_2_2[18] , \wRegOut_2_2[17] , \wRegOut_2_2[16] , 
        \wRegOut_2_2[15] , \wRegOut_2_2[14] , \wRegOut_2_2[13] , 
        \wRegOut_2_2[12] , \wRegOut_2_2[11] , \wRegOut_2_2[10] , 
        \wRegOut_2_2[9] , \wRegOut_2_2[8] , \wRegOut_2_2[7] , \wRegOut_2_2[6] , 
        \wRegOut_2_2[5] , \wRegOut_2_2[4] , \wRegOut_2_2[3] , \wRegOut_2_2[2] , 
        \wRegOut_2_2[1] , \wRegOut_2_2[0] }), .P_Out({\wRegInBot_2_2[31] , 
        \wRegInBot_2_2[30] , \wRegInBot_2_2[29] , \wRegInBot_2_2[28] , 
        \wRegInBot_2_2[27] , \wRegInBot_2_2[26] , \wRegInBot_2_2[25] , 
        \wRegInBot_2_2[24] , \wRegInBot_2_2[23] , \wRegInBot_2_2[22] , 
        \wRegInBot_2_2[21] , \wRegInBot_2_2[20] , \wRegInBot_2_2[19] , 
        \wRegInBot_2_2[18] , \wRegInBot_2_2[17] , \wRegInBot_2_2[16] , 
        \wRegInBot_2_2[15] , \wRegInBot_2_2[14] , \wRegInBot_2_2[13] , 
        \wRegInBot_2_2[12] , \wRegInBot_2_2[11] , \wRegInBot_2_2[10] , 
        \wRegInBot_2_2[9] , \wRegInBot_2_2[8] , \wRegInBot_2_2[7] , 
        \wRegInBot_2_2[6] , \wRegInBot_2_2[5] , \wRegInBot_2_2[4] , 
        \wRegInBot_2_2[3] , \wRegInBot_2_2[2] , \wRegInBot_2_2[1] , 
        \wRegInBot_2_2[0] }), .L_WR(\wRegEnTop_3_4[0] ), .L_In({
        \wRegOut_3_4[31] , \wRegOut_3_4[30] , \wRegOut_3_4[29] , 
        \wRegOut_3_4[28] , \wRegOut_3_4[27] , \wRegOut_3_4[26] , 
        \wRegOut_3_4[25] , \wRegOut_3_4[24] , \wRegOut_3_4[23] , 
        \wRegOut_3_4[22] , \wRegOut_3_4[21] , \wRegOut_3_4[20] , 
        \wRegOut_3_4[19] , \wRegOut_3_4[18] , \wRegOut_3_4[17] , 
        \wRegOut_3_4[16] , \wRegOut_3_4[15] , \wRegOut_3_4[14] , 
        \wRegOut_3_4[13] , \wRegOut_3_4[12] , \wRegOut_3_4[11] , 
        \wRegOut_3_4[10] , \wRegOut_3_4[9] , \wRegOut_3_4[8] , 
        \wRegOut_3_4[7] , \wRegOut_3_4[6] , \wRegOut_3_4[5] , \wRegOut_3_4[4] , 
        \wRegOut_3_4[3] , \wRegOut_3_4[2] , \wRegOut_3_4[1] , \wRegOut_3_4[0] 
        }), .L_Out({\wRegInTop_3_4[31] , \wRegInTop_3_4[30] , 
        \wRegInTop_3_4[29] , \wRegInTop_3_4[28] , \wRegInTop_3_4[27] , 
        \wRegInTop_3_4[26] , \wRegInTop_3_4[25] , \wRegInTop_3_4[24] , 
        \wRegInTop_3_4[23] , \wRegInTop_3_4[22] , \wRegInTop_3_4[21] , 
        \wRegInTop_3_4[20] , \wRegInTop_3_4[19] , \wRegInTop_3_4[18] , 
        \wRegInTop_3_4[17] , \wRegInTop_3_4[16] , \wRegInTop_3_4[15] , 
        \wRegInTop_3_4[14] , \wRegInTop_3_4[13] , \wRegInTop_3_4[12] , 
        \wRegInTop_3_4[11] , \wRegInTop_3_4[10] , \wRegInTop_3_4[9] , 
        \wRegInTop_3_4[8] , \wRegInTop_3_4[7] , \wRegInTop_3_4[6] , 
        \wRegInTop_3_4[5] , \wRegInTop_3_4[4] , \wRegInTop_3_4[3] , 
        \wRegInTop_3_4[2] , \wRegInTop_3_4[1] , \wRegInTop_3_4[0] }), .R_WR(
        \wRegEnTop_3_5[0] ), .R_In({\wRegOut_3_5[31] , \wRegOut_3_5[30] , 
        \wRegOut_3_5[29] , \wRegOut_3_5[28] , \wRegOut_3_5[27] , 
        \wRegOut_3_5[26] , \wRegOut_3_5[25] , \wRegOut_3_5[24] , 
        \wRegOut_3_5[23] , \wRegOut_3_5[22] , \wRegOut_3_5[21] , 
        \wRegOut_3_5[20] , \wRegOut_3_5[19] , \wRegOut_3_5[18] , 
        \wRegOut_3_5[17] , \wRegOut_3_5[16] , \wRegOut_3_5[15] , 
        \wRegOut_3_5[14] , \wRegOut_3_5[13] , \wRegOut_3_5[12] , 
        \wRegOut_3_5[11] , \wRegOut_3_5[10] , \wRegOut_3_5[9] , 
        \wRegOut_3_5[8] , \wRegOut_3_5[7] , \wRegOut_3_5[6] , \wRegOut_3_5[5] , 
        \wRegOut_3_5[4] , \wRegOut_3_5[3] , \wRegOut_3_5[2] , \wRegOut_3_5[1] , 
        \wRegOut_3_5[0] }), .R_Out({\wRegInTop_3_5[31] , \wRegInTop_3_5[30] , 
        \wRegInTop_3_5[29] , \wRegInTop_3_5[28] , \wRegInTop_3_5[27] , 
        \wRegInTop_3_5[26] , \wRegInTop_3_5[25] , \wRegInTop_3_5[24] , 
        \wRegInTop_3_5[23] , \wRegInTop_3_5[22] , \wRegInTop_3_5[21] , 
        \wRegInTop_3_5[20] , \wRegInTop_3_5[19] , \wRegInTop_3_5[18] , 
        \wRegInTop_3_5[17] , \wRegInTop_3_5[16] , \wRegInTop_3_5[15] , 
        \wRegInTop_3_5[14] , \wRegInTop_3_5[13] , \wRegInTop_3_5[12] , 
        \wRegInTop_3_5[11] , \wRegInTop_3_5[10] , \wRegInTop_3_5[9] , 
        \wRegInTop_3_5[8] , \wRegInTop_3_5[7] , \wRegInTop_3_5[6] , 
        \wRegInTop_3_5[5] , \wRegInTop_3_5[4] , \wRegInTop_3_5[3] , 
        \wRegInTop_3_5[2] , \wRegInTop_3_5[1] , \wRegInTop_3_5[0] }) );
    BHeap_Node_WIDTH32 BHN_3_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_2[0] ), .P_In({\wRegOut_3_2[31] , 
        \wRegOut_3_2[30] , \wRegOut_3_2[29] , \wRegOut_3_2[28] , 
        \wRegOut_3_2[27] , \wRegOut_3_2[26] , \wRegOut_3_2[25] , 
        \wRegOut_3_2[24] , \wRegOut_3_2[23] , \wRegOut_3_2[22] , 
        \wRegOut_3_2[21] , \wRegOut_3_2[20] , \wRegOut_3_2[19] , 
        \wRegOut_3_2[18] , \wRegOut_3_2[17] , \wRegOut_3_2[16] , 
        \wRegOut_3_2[15] , \wRegOut_3_2[14] , \wRegOut_3_2[13] , 
        \wRegOut_3_2[12] , \wRegOut_3_2[11] , \wRegOut_3_2[10] , 
        \wRegOut_3_2[9] , \wRegOut_3_2[8] , \wRegOut_3_2[7] , \wRegOut_3_2[6] , 
        \wRegOut_3_2[5] , \wRegOut_3_2[4] , \wRegOut_3_2[3] , \wRegOut_3_2[2] , 
        \wRegOut_3_2[1] , \wRegOut_3_2[0] }), .P_Out({\wRegInBot_3_2[31] , 
        \wRegInBot_3_2[30] , \wRegInBot_3_2[29] , \wRegInBot_3_2[28] , 
        \wRegInBot_3_2[27] , \wRegInBot_3_2[26] , \wRegInBot_3_2[25] , 
        \wRegInBot_3_2[24] , \wRegInBot_3_2[23] , \wRegInBot_3_2[22] , 
        \wRegInBot_3_2[21] , \wRegInBot_3_2[20] , \wRegInBot_3_2[19] , 
        \wRegInBot_3_2[18] , \wRegInBot_3_2[17] , \wRegInBot_3_2[16] , 
        \wRegInBot_3_2[15] , \wRegInBot_3_2[14] , \wRegInBot_3_2[13] , 
        \wRegInBot_3_2[12] , \wRegInBot_3_2[11] , \wRegInBot_3_2[10] , 
        \wRegInBot_3_2[9] , \wRegInBot_3_2[8] , \wRegInBot_3_2[7] , 
        \wRegInBot_3_2[6] , \wRegInBot_3_2[5] , \wRegInBot_3_2[4] , 
        \wRegInBot_3_2[3] , \wRegInBot_3_2[2] , \wRegInBot_3_2[1] , 
        \wRegInBot_3_2[0] }), .L_WR(\wRegEnTop_4_4[0] ), .L_In({
        \wRegOut_4_4[31] , \wRegOut_4_4[30] , \wRegOut_4_4[29] , 
        \wRegOut_4_4[28] , \wRegOut_4_4[27] , \wRegOut_4_4[26] , 
        \wRegOut_4_4[25] , \wRegOut_4_4[24] , \wRegOut_4_4[23] , 
        \wRegOut_4_4[22] , \wRegOut_4_4[21] , \wRegOut_4_4[20] , 
        \wRegOut_4_4[19] , \wRegOut_4_4[18] , \wRegOut_4_4[17] , 
        \wRegOut_4_4[16] , \wRegOut_4_4[15] , \wRegOut_4_4[14] , 
        \wRegOut_4_4[13] , \wRegOut_4_4[12] , \wRegOut_4_4[11] , 
        \wRegOut_4_4[10] , \wRegOut_4_4[9] , \wRegOut_4_4[8] , 
        \wRegOut_4_4[7] , \wRegOut_4_4[6] , \wRegOut_4_4[5] , \wRegOut_4_4[4] , 
        \wRegOut_4_4[3] , \wRegOut_4_4[2] , \wRegOut_4_4[1] , \wRegOut_4_4[0] 
        }), .L_Out({\wRegInTop_4_4[31] , \wRegInTop_4_4[30] , 
        \wRegInTop_4_4[29] , \wRegInTop_4_4[28] , \wRegInTop_4_4[27] , 
        \wRegInTop_4_4[26] , \wRegInTop_4_4[25] , \wRegInTop_4_4[24] , 
        \wRegInTop_4_4[23] , \wRegInTop_4_4[22] , \wRegInTop_4_4[21] , 
        \wRegInTop_4_4[20] , \wRegInTop_4_4[19] , \wRegInTop_4_4[18] , 
        \wRegInTop_4_4[17] , \wRegInTop_4_4[16] , \wRegInTop_4_4[15] , 
        \wRegInTop_4_4[14] , \wRegInTop_4_4[13] , \wRegInTop_4_4[12] , 
        \wRegInTop_4_4[11] , \wRegInTop_4_4[10] , \wRegInTop_4_4[9] , 
        \wRegInTop_4_4[8] , \wRegInTop_4_4[7] , \wRegInTop_4_4[6] , 
        \wRegInTop_4_4[5] , \wRegInTop_4_4[4] , \wRegInTop_4_4[3] , 
        \wRegInTop_4_4[2] , \wRegInTop_4_4[1] , \wRegInTop_4_4[0] }), .R_WR(
        \wRegEnTop_4_5[0] ), .R_In({\wRegOut_4_5[31] , \wRegOut_4_5[30] , 
        \wRegOut_4_5[29] , \wRegOut_4_5[28] , \wRegOut_4_5[27] , 
        \wRegOut_4_5[26] , \wRegOut_4_5[25] , \wRegOut_4_5[24] , 
        \wRegOut_4_5[23] , \wRegOut_4_5[22] , \wRegOut_4_5[21] , 
        \wRegOut_4_5[20] , \wRegOut_4_5[19] , \wRegOut_4_5[18] , 
        \wRegOut_4_5[17] , \wRegOut_4_5[16] , \wRegOut_4_5[15] , 
        \wRegOut_4_5[14] , \wRegOut_4_5[13] , \wRegOut_4_5[12] , 
        \wRegOut_4_5[11] , \wRegOut_4_5[10] , \wRegOut_4_5[9] , 
        \wRegOut_4_5[8] , \wRegOut_4_5[7] , \wRegOut_4_5[6] , \wRegOut_4_5[5] , 
        \wRegOut_4_5[4] , \wRegOut_4_5[3] , \wRegOut_4_5[2] , \wRegOut_4_5[1] , 
        \wRegOut_4_5[0] }), .R_Out({\wRegInTop_4_5[31] , \wRegInTop_4_5[30] , 
        \wRegInTop_4_5[29] , \wRegInTop_4_5[28] , \wRegInTop_4_5[27] , 
        \wRegInTop_4_5[26] , \wRegInTop_4_5[25] , \wRegInTop_4_5[24] , 
        \wRegInTop_4_5[23] , \wRegInTop_4_5[22] , \wRegInTop_4_5[21] , 
        \wRegInTop_4_5[20] , \wRegInTop_4_5[19] , \wRegInTop_4_5[18] , 
        \wRegInTop_4_5[17] , \wRegInTop_4_5[16] , \wRegInTop_4_5[15] , 
        \wRegInTop_4_5[14] , \wRegInTop_4_5[13] , \wRegInTop_4_5[12] , 
        \wRegInTop_4_5[11] , \wRegInTop_4_5[10] , \wRegInTop_4_5[9] , 
        \wRegInTop_4_5[8] , \wRegInTop_4_5[7] , \wRegInTop_4_5[6] , 
        \wRegInTop_4_5[5] , \wRegInTop_4_5[4] , \wRegInTop_4_5[3] , 
        \wRegInTop_4_5[2] , \wRegInTop_4_5[1] , \wRegInTop_4_5[0] }) );
    BHeap_Node_WIDTH32 BHN_4_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_8[0] ), .P_In({\wRegOut_4_8[31] , 
        \wRegOut_4_8[30] , \wRegOut_4_8[29] , \wRegOut_4_8[28] , 
        \wRegOut_4_8[27] , \wRegOut_4_8[26] , \wRegOut_4_8[25] , 
        \wRegOut_4_8[24] , \wRegOut_4_8[23] , \wRegOut_4_8[22] , 
        \wRegOut_4_8[21] , \wRegOut_4_8[20] , \wRegOut_4_8[19] , 
        \wRegOut_4_8[18] , \wRegOut_4_8[17] , \wRegOut_4_8[16] , 
        \wRegOut_4_8[15] , \wRegOut_4_8[14] , \wRegOut_4_8[13] , 
        \wRegOut_4_8[12] , \wRegOut_4_8[11] , \wRegOut_4_8[10] , 
        \wRegOut_4_8[9] , \wRegOut_4_8[8] , \wRegOut_4_8[7] , \wRegOut_4_8[6] , 
        \wRegOut_4_8[5] , \wRegOut_4_8[4] , \wRegOut_4_8[3] , \wRegOut_4_8[2] , 
        \wRegOut_4_8[1] , \wRegOut_4_8[0] }), .P_Out({\wRegInBot_4_8[31] , 
        \wRegInBot_4_8[30] , \wRegInBot_4_8[29] , \wRegInBot_4_8[28] , 
        \wRegInBot_4_8[27] , \wRegInBot_4_8[26] , \wRegInBot_4_8[25] , 
        \wRegInBot_4_8[24] , \wRegInBot_4_8[23] , \wRegInBot_4_8[22] , 
        \wRegInBot_4_8[21] , \wRegInBot_4_8[20] , \wRegInBot_4_8[19] , 
        \wRegInBot_4_8[18] , \wRegInBot_4_8[17] , \wRegInBot_4_8[16] , 
        \wRegInBot_4_8[15] , \wRegInBot_4_8[14] , \wRegInBot_4_8[13] , 
        \wRegInBot_4_8[12] , \wRegInBot_4_8[11] , \wRegInBot_4_8[10] , 
        \wRegInBot_4_8[9] , \wRegInBot_4_8[8] , \wRegInBot_4_8[7] , 
        \wRegInBot_4_8[6] , \wRegInBot_4_8[5] , \wRegInBot_4_8[4] , 
        \wRegInBot_4_8[3] , \wRegInBot_4_8[2] , \wRegInBot_4_8[1] , 
        \wRegInBot_4_8[0] }), .L_WR(\wRegEnTop_5_16[0] ), .L_In({
        \wRegOut_5_16[31] , \wRegOut_5_16[30] , \wRegOut_5_16[29] , 
        \wRegOut_5_16[28] , \wRegOut_5_16[27] , \wRegOut_5_16[26] , 
        \wRegOut_5_16[25] , \wRegOut_5_16[24] , \wRegOut_5_16[23] , 
        \wRegOut_5_16[22] , \wRegOut_5_16[21] , \wRegOut_5_16[20] , 
        \wRegOut_5_16[19] , \wRegOut_5_16[18] , \wRegOut_5_16[17] , 
        \wRegOut_5_16[16] , \wRegOut_5_16[15] , \wRegOut_5_16[14] , 
        \wRegOut_5_16[13] , \wRegOut_5_16[12] , \wRegOut_5_16[11] , 
        \wRegOut_5_16[10] , \wRegOut_5_16[9] , \wRegOut_5_16[8] , 
        \wRegOut_5_16[7] , \wRegOut_5_16[6] , \wRegOut_5_16[5] , 
        \wRegOut_5_16[4] , \wRegOut_5_16[3] , \wRegOut_5_16[2] , 
        \wRegOut_5_16[1] , \wRegOut_5_16[0] }), .L_Out({\wRegInTop_5_16[31] , 
        \wRegInTop_5_16[30] , \wRegInTop_5_16[29] , \wRegInTop_5_16[28] , 
        \wRegInTop_5_16[27] , \wRegInTop_5_16[26] , \wRegInTop_5_16[25] , 
        \wRegInTop_5_16[24] , \wRegInTop_5_16[23] , \wRegInTop_5_16[22] , 
        \wRegInTop_5_16[21] , \wRegInTop_5_16[20] , \wRegInTop_5_16[19] , 
        \wRegInTop_5_16[18] , \wRegInTop_5_16[17] , \wRegInTop_5_16[16] , 
        \wRegInTop_5_16[15] , \wRegInTop_5_16[14] , \wRegInTop_5_16[13] , 
        \wRegInTop_5_16[12] , \wRegInTop_5_16[11] , \wRegInTop_5_16[10] , 
        \wRegInTop_5_16[9] , \wRegInTop_5_16[8] , \wRegInTop_5_16[7] , 
        \wRegInTop_5_16[6] , \wRegInTop_5_16[5] , \wRegInTop_5_16[4] , 
        \wRegInTop_5_16[3] , \wRegInTop_5_16[2] , \wRegInTop_5_16[1] , 
        \wRegInTop_5_16[0] }), .R_WR(\wRegEnTop_5_17[0] ), .R_In({
        \wRegOut_5_17[31] , \wRegOut_5_17[30] , \wRegOut_5_17[29] , 
        \wRegOut_5_17[28] , \wRegOut_5_17[27] , \wRegOut_5_17[26] , 
        \wRegOut_5_17[25] , \wRegOut_5_17[24] , \wRegOut_5_17[23] , 
        \wRegOut_5_17[22] , \wRegOut_5_17[21] , \wRegOut_5_17[20] , 
        \wRegOut_5_17[19] , \wRegOut_5_17[18] , \wRegOut_5_17[17] , 
        \wRegOut_5_17[16] , \wRegOut_5_17[15] , \wRegOut_5_17[14] , 
        \wRegOut_5_17[13] , \wRegOut_5_17[12] , \wRegOut_5_17[11] , 
        \wRegOut_5_17[10] , \wRegOut_5_17[9] , \wRegOut_5_17[8] , 
        \wRegOut_5_17[7] , \wRegOut_5_17[6] , \wRegOut_5_17[5] , 
        \wRegOut_5_17[4] , \wRegOut_5_17[3] , \wRegOut_5_17[2] , 
        \wRegOut_5_17[1] , \wRegOut_5_17[0] }), .R_Out({\wRegInTop_5_17[31] , 
        \wRegInTop_5_17[30] , \wRegInTop_5_17[29] , \wRegInTop_5_17[28] , 
        \wRegInTop_5_17[27] , \wRegInTop_5_17[26] , \wRegInTop_5_17[25] , 
        \wRegInTop_5_17[24] , \wRegInTop_5_17[23] , \wRegInTop_5_17[22] , 
        \wRegInTop_5_17[21] , \wRegInTop_5_17[20] , \wRegInTop_5_17[19] , 
        \wRegInTop_5_17[18] , \wRegInTop_5_17[17] , \wRegInTop_5_17[16] , 
        \wRegInTop_5_17[15] , \wRegInTop_5_17[14] , \wRegInTop_5_17[13] , 
        \wRegInTop_5_17[12] , \wRegInTop_5_17[11] , \wRegInTop_5_17[10] , 
        \wRegInTop_5_17[9] , \wRegInTop_5_17[8] , \wRegInTop_5_17[7] , 
        \wRegInTop_5_17[6] , \wRegInTop_5_17[5] , \wRegInTop_5_17[4] , 
        \wRegInTop_5_17[3] , \wRegInTop_5_17[2] , \wRegInTop_5_17[1] , 
        \wRegInTop_5_17[0] }) );
    BHeap_Node_WIDTH32 BHN_4_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_11[0] ), .P_In({\wRegOut_4_11[31] , 
        \wRegOut_4_11[30] , \wRegOut_4_11[29] , \wRegOut_4_11[28] , 
        \wRegOut_4_11[27] , \wRegOut_4_11[26] , \wRegOut_4_11[25] , 
        \wRegOut_4_11[24] , \wRegOut_4_11[23] , \wRegOut_4_11[22] , 
        \wRegOut_4_11[21] , \wRegOut_4_11[20] , \wRegOut_4_11[19] , 
        \wRegOut_4_11[18] , \wRegOut_4_11[17] , \wRegOut_4_11[16] , 
        \wRegOut_4_11[15] , \wRegOut_4_11[14] , \wRegOut_4_11[13] , 
        \wRegOut_4_11[12] , \wRegOut_4_11[11] , \wRegOut_4_11[10] , 
        \wRegOut_4_11[9] , \wRegOut_4_11[8] , \wRegOut_4_11[7] , 
        \wRegOut_4_11[6] , \wRegOut_4_11[5] , \wRegOut_4_11[4] , 
        \wRegOut_4_11[3] , \wRegOut_4_11[2] , \wRegOut_4_11[1] , 
        \wRegOut_4_11[0] }), .P_Out({\wRegInBot_4_11[31] , 
        \wRegInBot_4_11[30] , \wRegInBot_4_11[29] , \wRegInBot_4_11[28] , 
        \wRegInBot_4_11[27] , \wRegInBot_4_11[26] , \wRegInBot_4_11[25] , 
        \wRegInBot_4_11[24] , \wRegInBot_4_11[23] , \wRegInBot_4_11[22] , 
        \wRegInBot_4_11[21] , \wRegInBot_4_11[20] , \wRegInBot_4_11[19] , 
        \wRegInBot_4_11[18] , \wRegInBot_4_11[17] , \wRegInBot_4_11[16] , 
        \wRegInBot_4_11[15] , \wRegInBot_4_11[14] , \wRegInBot_4_11[13] , 
        \wRegInBot_4_11[12] , \wRegInBot_4_11[11] , \wRegInBot_4_11[10] , 
        \wRegInBot_4_11[9] , \wRegInBot_4_11[8] , \wRegInBot_4_11[7] , 
        \wRegInBot_4_11[6] , \wRegInBot_4_11[5] , \wRegInBot_4_11[4] , 
        \wRegInBot_4_11[3] , \wRegInBot_4_11[2] , \wRegInBot_4_11[1] , 
        \wRegInBot_4_11[0] }), .L_WR(\wRegEnTop_5_22[0] ), .L_In({
        \wRegOut_5_22[31] , \wRegOut_5_22[30] , \wRegOut_5_22[29] , 
        \wRegOut_5_22[28] , \wRegOut_5_22[27] , \wRegOut_5_22[26] , 
        \wRegOut_5_22[25] , \wRegOut_5_22[24] , \wRegOut_5_22[23] , 
        \wRegOut_5_22[22] , \wRegOut_5_22[21] , \wRegOut_5_22[20] , 
        \wRegOut_5_22[19] , \wRegOut_5_22[18] , \wRegOut_5_22[17] , 
        \wRegOut_5_22[16] , \wRegOut_5_22[15] , \wRegOut_5_22[14] , 
        \wRegOut_5_22[13] , \wRegOut_5_22[12] , \wRegOut_5_22[11] , 
        \wRegOut_5_22[10] , \wRegOut_5_22[9] , \wRegOut_5_22[8] , 
        \wRegOut_5_22[7] , \wRegOut_5_22[6] , \wRegOut_5_22[5] , 
        \wRegOut_5_22[4] , \wRegOut_5_22[3] , \wRegOut_5_22[2] , 
        \wRegOut_5_22[1] , \wRegOut_5_22[0] }), .L_Out({\wRegInTop_5_22[31] , 
        \wRegInTop_5_22[30] , \wRegInTop_5_22[29] , \wRegInTop_5_22[28] , 
        \wRegInTop_5_22[27] , \wRegInTop_5_22[26] , \wRegInTop_5_22[25] , 
        \wRegInTop_5_22[24] , \wRegInTop_5_22[23] , \wRegInTop_5_22[22] , 
        \wRegInTop_5_22[21] , \wRegInTop_5_22[20] , \wRegInTop_5_22[19] , 
        \wRegInTop_5_22[18] , \wRegInTop_5_22[17] , \wRegInTop_5_22[16] , 
        \wRegInTop_5_22[15] , \wRegInTop_5_22[14] , \wRegInTop_5_22[13] , 
        \wRegInTop_5_22[12] , \wRegInTop_5_22[11] , \wRegInTop_5_22[10] , 
        \wRegInTop_5_22[9] , \wRegInTop_5_22[8] , \wRegInTop_5_22[7] , 
        \wRegInTop_5_22[6] , \wRegInTop_5_22[5] , \wRegInTop_5_22[4] , 
        \wRegInTop_5_22[3] , \wRegInTop_5_22[2] , \wRegInTop_5_22[1] , 
        \wRegInTop_5_22[0] }), .R_WR(\wRegEnTop_5_23[0] ), .R_In({
        \wRegOut_5_23[31] , \wRegOut_5_23[30] , \wRegOut_5_23[29] , 
        \wRegOut_5_23[28] , \wRegOut_5_23[27] , \wRegOut_5_23[26] , 
        \wRegOut_5_23[25] , \wRegOut_5_23[24] , \wRegOut_5_23[23] , 
        \wRegOut_5_23[22] , \wRegOut_5_23[21] , \wRegOut_5_23[20] , 
        \wRegOut_5_23[19] , \wRegOut_5_23[18] , \wRegOut_5_23[17] , 
        \wRegOut_5_23[16] , \wRegOut_5_23[15] , \wRegOut_5_23[14] , 
        \wRegOut_5_23[13] , \wRegOut_5_23[12] , \wRegOut_5_23[11] , 
        \wRegOut_5_23[10] , \wRegOut_5_23[9] , \wRegOut_5_23[8] , 
        \wRegOut_5_23[7] , \wRegOut_5_23[6] , \wRegOut_5_23[5] , 
        \wRegOut_5_23[4] , \wRegOut_5_23[3] , \wRegOut_5_23[2] , 
        \wRegOut_5_23[1] , \wRegOut_5_23[0] }), .R_Out({\wRegInTop_5_23[31] , 
        \wRegInTop_5_23[30] , \wRegInTop_5_23[29] , \wRegInTop_5_23[28] , 
        \wRegInTop_5_23[27] , \wRegInTop_5_23[26] , \wRegInTop_5_23[25] , 
        \wRegInTop_5_23[24] , \wRegInTop_5_23[23] , \wRegInTop_5_23[22] , 
        \wRegInTop_5_23[21] , \wRegInTop_5_23[20] , \wRegInTop_5_23[19] , 
        \wRegInTop_5_23[18] , \wRegInTop_5_23[17] , \wRegInTop_5_23[16] , 
        \wRegInTop_5_23[15] , \wRegInTop_5_23[14] , \wRegInTop_5_23[13] , 
        \wRegInTop_5_23[12] , \wRegInTop_5_23[11] , \wRegInTop_5_23[10] , 
        \wRegInTop_5_23[9] , \wRegInTop_5_23[8] , \wRegInTop_5_23[7] , 
        \wRegInTop_5_23[6] , \wRegInTop_5_23[5] , \wRegInTop_5_23[4] , 
        \wRegInTop_5_23[3] , \wRegInTop_5_23[2] , \wRegInTop_5_23[1] , 
        \wRegInTop_5_23[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_3_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink15[31] , \ScanLink15[30] , \ScanLink15[29] , 
        \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , \ScanLink15[25] , 
        \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , \ScanLink15[21] , 
        \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , \ScanLink15[17] , 
        \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , \ScanLink15[13] , 
        \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , \ScanLink15[9] , 
        \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , \ScanLink15[5] , 
        \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , \ScanLink15[1] , 
        \ScanLink15[0] }), .ScanOut({\ScanLink14[31] , \ScanLink14[30] , 
        \ScanLink14[29] , \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , 
        \ScanLink14[25] , \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , 
        \ScanLink14[21] , \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , 
        \ScanLink14[17] , \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , 
        \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , 
        \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , 
        \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , 
        \ScanLink14[1] , \ScanLink14[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_3_7[31] , \wRegOut_3_7[30] , \wRegOut_3_7[29] , 
        \wRegOut_3_7[28] , \wRegOut_3_7[27] , \wRegOut_3_7[26] , 
        \wRegOut_3_7[25] , \wRegOut_3_7[24] , \wRegOut_3_7[23] , 
        \wRegOut_3_7[22] , \wRegOut_3_7[21] , \wRegOut_3_7[20] , 
        \wRegOut_3_7[19] , \wRegOut_3_7[18] , \wRegOut_3_7[17] , 
        \wRegOut_3_7[16] , \wRegOut_3_7[15] , \wRegOut_3_7[14] , 
        \wRegOut_3_7[13] , \wRegOut_3_7[12] , \wRegOut_3_7[11] , 
        \wRegOut_3_7[10] , \wRegOut_3_7[9] , \wRegOut_3_7[8] , 
        \wRegOut_3_7[7] , \wRegOut_3_7[6] , \wRegOut_3_7[5] , \wRegOut_3_7[4] , 
        \wRegOut_3_7[3] , \wRegOut_3_7[2] , \wRegOut_3_7[1] , \wRegOut_3_7[0] 
        }), .Enable1(\wRegEnTop_3_7[0] ), .Enable2(\wRegEnBot_3_7[0] ), .In1({
        \wRegInTop_3_7[31] , \wRegInTop_3_7[30] , \wRegInTop_3_7[29] , 
        \wRegInTop_3_7[28] , \wRegInTop_3_7[27] , \wRegInTop_3_7[26] , 
        \wRegInTop_3_7[25] , \wRegInTop_3_7[24] , \wRegInTop_3_7[23] , 
        \wRegInTop_3_7[22] , \wRegInTop_3_7[21] , \wRegInTop_3_7[20] , 
        \wRegInTop_3_7[19] , \wRegInTop_3_7[18] , \wRegInTop_3_7[17] , 
        \wRegInTop_3_7[16] , \wRegInTop_3_7[15] , \wRegInTop_3_7[14] , 
        \wRegInTop_3_7[13] , \wRegInTop_3_7[12] , \wRegInTop_3_7[11] , 
        \wRegInTop_3_7[10] , \wRegInTop_3_7[9] , \wRegInTop_3_7[8] , 
        \wRegInTop_3_7[7] , \wRegInTop_3_7[6] , \wRegInTop_3_7[5] , 
        \wRegInTop_3_7[4] , \wRegInTop_3_7[3] , \wRegInTop_3_7[2] , 
        \wRegInTop_3_7[1] , \wRegInTop_3_7[0] }), .In2({\wRegInBot_3_7[31] , 
        \wRegInBot_3_7[30] , \wRegInBot_3_7[29] , \wRegInBot_3_7[28] , 
        \wRegInBot_3_7[27] , \wRegInBot_3_7[26] , \wRegInBot_3_7[25] , 
        \wRegInBot_3_7[24] , \wRegInBot_3_7[23] , \wRegInBot_3_7[22] , 
        \wRegInBot_3_7[21] , \wRegInBot_3_7[20] , \wRegInBot_3_7[19] , 
        \wRegInBot_3_7[18] , \wRegInBot_3_7[17] , \wRegInBot_3_7[16] , 
        \wRegInBot_3_7[15] , \wRegInBot_3_7[14] , \wRegInBot_3_7[13] , 
        \wRegInBot_3_7[12] , \wRegInBot_3_7[11] , \wRegInBot_3_7[10] , 
        \wRegInBot_3_7[9] , \wRegInBot_3_7[8] , \wRegInBot_3_7[7] , 
        \wRegInBot_3_7[6] , \wRegInBot_3_7[5] , \wRegInBot_3_7[4] , 
        \wRegInBot_3_7[3] , \wRegInBot_3_7[2] , \wRegInBot_3_7[1] , 
        \wRegInBot_3_7[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_18 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink50[31] , \ScanLink50[30] , \ScanLink50[29] , 
        \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , \ScanLink50[25] , 
        \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , \ScanLink50[21] , 
        \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , \ScanLink50[17] , 
        \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , \ScanLink50[13] , 
        \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , \ScanLink50[9] , 
        \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , \ScanLink50[5] , 
        \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , \ScanLink50[1] , 
        \ScanLink50[0] }), .ScanOut({\ScanLink49[31] , \ScanLink49[30] , 
        \ScanLink49[29] , \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , 
        \ScanLink49[25] , \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , 
        \ScanLink49[21] , \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , 
        \ScanLink49[17] , \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , 
        \ScanLink49[13] , \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , 
        \ScanLink49[9] , \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , 
        \ScanLink49[5] , \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , 
        \ScanLink49[1] , \ScanLink49[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_18[31] , \wRegOut_5_18[30] , 
        \wRegOut_5_18[29] , \wRegOut_5_18[28] , \wRegOut_5_18[27] , 
        \wRegOut_5_18[26] , \wRegOut_5_18[25] , \wRegOut_5_18[24] , 
        \wRegOut_5_18[23] , \wRegOut_5_18[22] , \wRegOut_5_18[21] , 
        \wRegOut_5_18[20] , \wRegOut_5_18[19] , \wRegOut_5_18[18] , 
        \wRegOut_5_18[17] , \wRegOut_5_18[16] , \wRegOut_5_18[15] , 
        \wRegOut_5_18[14] , \wRegOut_5_18[13] , \wRegOut_5_18[12] , 
        \wRegOut_5_18[11] , \wRegOut_5_18[10] , \wRegOut_5_18[9] , 
        \wRegOut_5_18[8] , \wRegOut_5_18[7] , \wRegOut_5_18[6] , 
        \wRegOut_5_18[5] , \wRegOut_5_18[4] , \wRegOut_5_18[3] , 
        \wRegOut_5_18[2] , \wRegOut_5_18[1] , \wRegOut_5_18[0] }), .Enable1(
        \wRegEnTop_5_18[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_18[31] , 
        \wRegInTop_5_18[30] , \wRegInTop_5_18[29] , \wRegInTop_5_18[28] , 
        \wRegInTop_5_18[27] , \wRegInTop_5_18[26] , \wRegInTop_5_18[25] , 
        \wRegInTop_5_18[24] , \wRegInTop_5_18[23] , \wRegInTop_5_18[22] , 
        \wRegInTop_5_18[21] , \wRegInTop_5_18[20] , \wRegInTop_5_18[19] , 
        \wRegInTop_5_18[18] , \wRegInTop_5_18[17] , \wRegInTop_5_18[16] , 
        \wRegInTop_5_18[15] , \wRegInTop_5_18[14] , \wRegInTop_5_18[13] , 
        \wRegInTop_5_18[12] , \wRegInTop_5_18[11] , \wRegInTop_5_18[10] , 
        \wRegInTop_5_18[9] , \wRegInTop_5_18[8] , \wRegInTop_5_18[7] , 
        \wRegInTop_5_18[6] , \wRegInTop_5_18[5] , \wRegInTop_5_18[4] , 
        \wRegInTop_5_18[3] , \wRegInTop_5_18[2] , \wRegInTop_5_18[1] , 
        \wRegInTop_5_18[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink20[31] , \ScanLink20[30] , \ScanLink20[29] , 
        \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , \ScanLink20[25] , 
        \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , \ScanLink20[21] , 
        \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , \ScanLink20[17] , 
        \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , \ScanLink20[13] , 
        \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , \ScanLink20[9] , 
        \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , \ScanLink20[5] , 
        \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , \ScanLink20[1] , 
        \ScanLink20[0] }), .ScanOut({\ScanLink19[31] , \ScanLink19[30] , 
        \ScanLink19[29] , \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , 
        \ScanLink19[25] , \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , 
        \ScanLink19[21] , \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , 
        \ScanLink19[17] , \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , 
        \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , 
        \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , 
        \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , 
        \ScanLink19[1] , \ScanLink19[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_4[31] , \wRegOut_4_4[30] , \wRegOut_4_4[29] , 
        \wRegOut_4_4[28] , \wRegOut_4_4[27] , \wRegOut_4_4[26] , 
        \wRegOut_4_4[25] , \wRegOut_4_4[24] , \wRegOut_4_4[23] , 
        \wRegOut_4_4[22] , \wRegOut_4_4[21] , \wRegOut_4_4[20] , 
        \wRegOut_4_4[19] , \wRegOut_4_4[18] , \wRegOut_4_4[17] , 
        \wRegOut_4_4[16] , \wRegOut_4_4[15] , \wRegOut_4_4[14] , 
        \wRegOut_4_4[13] , \wRegOut_4_4[12] , \wRegOut_4_4[11] , 
        \wRegOut_4_4[10] , \wRegOut_4_4[9] , \wRegOut_4_4[8] , 
        \wRegOut_4_4[7] , \wRegOut_4_4[6] , \wRegOut_4_4[5] , \wRegOut_4_4[4] , 
        \wRegOut_4_4[3] , \wRegOut_4_4[2] , \wRegOut_4_4[1] , \wRegOut_4_4[0] 
        }), .Enable1(\wRegEnTop_4_4[0] ), .Enable2(\wRegEnBot_4_4[0] ), .In1({
        \wRegInTop_4_4[31] , \wRegInTop_4_4[30] , \wRegInTop_4_4[29] , 
        \wRegInTop_4_4[28] , \wRegInTop_4_4[27] , \wRegInTop_4_4[26] , 
        \wRegInTop_4_4[25] , \wRegInTop_4_4[24] , \wRegInTop_4_4[23] , 
        \wRegInTop_4_4[22] , \wRegInTop_4_4[21] , \wRegInTop_4_4[20] , 
        \wRegInTop_4_4[19] , \wRegInTop_4_4[18] , \wRegInTop_4_4[17] , 
        \wRegInTop_4_4[16] , \wRegInTop_4_4[15] , \wRegInTop_4_4[14] , 
        \wRegInTop_4_4[13] , \wRegInTop_4_4[12] , \wRegInTop_4_4[11] , 
        \wRegInTop_4_4[10] , \wRegInTop_4_4[9] , \wRegInTop_4_4[8] , 
        \wRegInTop_4_4[7] , \wRegInTop_4_4[6] , \wRegInTop_4_4[5] , 
        \wRegInTop_4_4[4] , \wRegInTop_4_4[3] , \wRegInTop_4_4[2] , 
        \wRegInTop_4_4[1] , \wRegInTop_4_4[0] }), .In2({\wRegInBot_4_4[31] , 
        \wRegInBot_4_4[30] , \wRegInBot_4_4[29] , \wRegInBot_4_4[28] , 
        \wRegInBot_4_4[27] , \wRegInBot_4_4[26] , \wRegInBot_4_4[25] , 
        \wRegInBot_4_4[24] , \wRegInBot_4_4[23] , \wRegInBot_4_4[22] , 
        \wRegInBot_4_4[21] , \wRegInBot_4_4[20] , \wRegInBot_4_4[19] , 
        \wRegInBot_4_4[18] , \wRegInBot_4_4[17] , \wRegInBot_4_4[16] , 
        \wRegInBot_4_4[15] , \wRegInBot_4_4[14] , \wRegInBot_4_4[13] , 
        \wRegInBot_4_4[12] , \wRegInBot_4_4[11] , \wRegInBot_4_4[10] , 
        \wRegInBot_4_4[9] , \wRegInBot_4_4[8] , \wRegInBot_4_4[7] , 
        \wRegInBot_4_4[6] , \wRegInBot_4_4[5] , \wRegInBot_4_4[4] , 
        \wRegInBot_4_4[3] , \wRegInBot_4_4[2] , \wRegInBot_4_4[1] , 
        \wRegInBot_4_4[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink43[31] , \ScanLink43[30] , \ScanLink43[29] , 
        \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , \ScanLink43[25] , 
        \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , \ScanLink43[21] , 
        \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , \ScanLink43[17] , 
        \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , \ScanLink43[13] , 
        \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , \ScanLink43[9] , 
        \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , \ScanLink43[5] , 
        \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , \ScanLink43[1] , 
        \ScanLink43[0] }), .ScanOut({\ScanLink42[31] , \ScanLink42[30] , 
        \ScanLink42[29] , \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , 
        \ScanLink42[25] , \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , 
        \ScanLink42[21] , \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , 
        \ScanLink42[17] , \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , 
        \ScanLink42[13] , \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , 
        \ScanLink42[9] , \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , 
        \ScanLink42[5] , \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , 
        \ScanLink42[1] , \ScanLink42[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_11[31] , \wRegOut_5_11[30] , 
        \wRegOut_5_11[29] , \wRegOut_5_11[28] , \wRegOut_5_11[27] , 
        \wRegOut_5_11[26] , \wRegOut_5_11[25] , \wRegOut_5_11[24] , 
        \wRegOut_5_11[23] , \wRegOut_5_11[22] , \wRegOut_5_11[21] , 
        \wRegOut_5_11[20] , \wRegOut_5_11[19] , \wRegOut_5_11[18] , 
        \wRegOut_5_11[17] , \wRegOut_5_11[16] , \wRegOut_5_11[15] , 
        \wRegOut_5_11[14] , \wRegOut_5_11[13] , \wRegOut_5_11[12] , 
        \wRegOut_5_11[11] , \wRegOut_5_11[10] , \wRegOut_5_11[9] , 
        \wRegOut_5_11[8] , \wRegOut_5_11[7] , \wRegOut_5_11[6] , 
        \wRegOut_5_11[5] , \wRegOut_5_11[4] , \wRegOut_5_11[3] , 
        \wRegOut_5_11[2] , \wRegOut_5_11[1] , \wRegOut_5_11[0] }), .Enable1(
        \wRegEnTop_5_11[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_11[31] , 
        \wRegInTop_5_11[30] , \wRegInTop_5_11[29] , \wRegInTop_5_11[28] , 
        \wRegInTop_5_11[27] , \wRegInTop_5_11[26] , \wRegInTop_5_11[25] , 
        \wRegInTop_5_11[24] , \wRegInTop_5_11[23] , \wRegInTop_5_11[22] , 
        \wRegInTop_5_11[21] , \wRegInTop_5_11[20] , \wRegInTop_5_11[19] , 
        \wRegInTop_5_11[18] , \wRegInTop_5_11[17] , \wRegInTop_5_11[16] , 
        \wRegInTop_5_11[15] , \wRegInTop_5_11[14] , \wRegInTop_5_11[13] , 
        \wRegInTop_5_11[12] , \wRegInTop_5_11[11] , \wRegInTop_5_11[10] , 
        \wRegInTop_5_11[9] , \wRegInTop_5_11[8] , \wRegInTop_5_11[7] , 
        \wRegInTop_5_11[6] , \wRegInTop_5_11[5] , \wRegInTop_5_11[4] , 
        \wRegInTop_5_11[3] , \wRegInTop_5_11[2] , \wRegInTop_5_11[1] , 
        \wRegInTop_5_11[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_24 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink56[31] , \ScanLink56[30] , \ScanLink56[29] , 
        \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , \ScanLink56[25] , 
        \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , \ScanLink56[21] , 
        \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , \ScanLink56[17] , 
        \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , \ScanLink56[13] , 
        \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , \ScanLink56[9] , 
        \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , \ScanLink56[5] , 
        \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , \ScanLink56[1] , 
        \ScanLink56[0] }), .ScanOut({\ScanLink55[31] , \ScanLink55[30] , 
        \ScanLink55[29] , \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , 
        \ScanLink55[25] , \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , 
        \ScanLink55[21] , \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , 
        \ScanLink55[17] , \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , 
        \ScanLink55[13] , \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , 
        \ScanLink55[9] , \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , 
        \ScanLink55[5] , \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , 
        \ScanLink55[1] , \ScanLink55[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_24[31] , \wRegOut_5_24[30] , 
        \wRegOut_5_24[29] , \wRegOut_5_24[28] , \wRegOut_5_24[27] , 
        \wRegOut_5_24[26] , \wRegOut_5_24[25] , \wRegOut_5_24[24] , 
        \wRegOut_5_24[23] , \wRegOut_5_24[22] , \wRegOut_5_24[21] , 
        \wRegOut_5_24[20] , \wRegOut_5_24[19] , \wRegOut_5_24[18] , 
        \wRegOut_5_24[17] , \wRegOut_5_24[16] , \wRegOut_5_24[15] , 
        \wRegOut_5_24[14] , \wRegOut_5_24[13] , \wRegOut_5_24[12] , 
        \wRegOut_5_24[11] , \wRegOut_5_24[10] , \wRegOut_5_24[9] , 
        \wRegOut_5_24[8] , \wRegOut_5_24[7] , \wRegOut_5_24[6] , 
        \wRegOut_5_24[5] , \wRegOut_5_24[4] , \wRegOut_5_24[3] , 
        \wRegOut_5_24[2] , \wRegOut_5_24[1] , \wRegOut_5_24[0] }), .Enable1(
        \wRegEnTop_5_24[0] ), .Enable2(1'b0), .In1({\wRegInTop_5_24[31] , 
        \wRegInTop_5_24[30] , \wRegInTop_5_24[29] , \wRegInTop_5_24[28] , 
        \wRegInTop_5_24[27] , \wRegInTop_5_24[26] , \wRegInTop_5_24[25] , 
        \wRegInTop_5_24[24] , \wRegInTop_5_24[23] , \wRegInTop_5_24[22] , 
        \wRegInTop_5_24[21] , \wRegInTop_5_24[20] , \wRegInTop_5_24[19] , 
        \wRegInTop_5_24[18] , \wRegInTop_5_24[17] , \wRegInTop_5_24[16] , 
        \wRegInTop_5_24[15] , \wRegInTop_5_24[14] , \wRegInTop_5_24[13] , 
        \wRegInTop_5_24[12] , \wRegInTop_5_24[11] , \wRegInTop_5_24[10] , 
        \wRegInTop_5_24[9] , \wRegInTop_5_24[8] , \wRegInTop_5_24[7] , 
        \wRegInTop_5_24[6] , \wRegInTop_5_24[5] , \wRegInTop_5_24[4] , 
        \wRegInTop_5_24[3] , \wRegInTop_5_24[2] , \wRegInTop_5_24[1] , 
        \wRegInTop_5_24[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
    BHeap_Node_WIDTH32 BHN_3_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_3[0] ), .P_WR(\wRegEnBot_3_5[0] ), .P_In({\wRegOut_3_5[31] , 
        \wRegOut_3_5[30] , \wRegOut_3_5[29] , \wRegOut_3_5[28] , 
        \wRegOut_3_5[27] , \wRegOut_3_5[26] , \wRegOut_3_5[25] , 
        \wRegOut_3_5[24] , \wRegOut_3_5[23] , \wRegOut_3_5[22] , 
        \wRegOut_3_5[21] , \wRegOut_3_5[20] , \wRegOut_3_5[19] , 
        \wRegOut_3_5[18] , \wRegOut_3_5[17] , \wRegOut_3_5[16] , 
        \wRegOut_3_5[15] , \wRegOut_3_5[14] , \wRegOut_3_5[13] , 
        \wRegOut_3_5[12] , \wRegOut_3_5[11] , \wRegOut_3_5[10] , 
        \wRegOut_3_5[9] , \wRegOut_3_5[8] , \wRegOut_3_5[7] , \wRegOut_3_5[6] , 
        \wRegOut_3_5[5] , \wRegOut_3_5[4] , \wRegOut_3_5[3] , \wRegOut_3_5[2] , 
        \wRegOut_3_5[1] , \wRegOut_3_5[0] }), .P_Out({\wRegInBot_3_5[31] , 
        \wRegInBot_3_5[30] , \wRegInBot_3_5[29] , \wRegInBot_3_5[28] , 
        \wRegInBot_3_5[27] , \wRegInBot_3_5[26] , \wRegInBot_3_5[25] , 
        \wRegInBot_3_5[24] , \wRegInBot_3_5[23] , \wRegInBot_3_5[22] , 
        \wRegInBot_3_5[21] , \wRegInBot_3_5[20] , \wRegInBot_3_5[19] , 
        \wRegInBot_3_5[18] , \wRegInBot_3_5[17] , \wRegInBot_3_5[16] , 
        \wRegInBot_3_5[15] , \wRegInBot_3_5[14] , \wRegInBot_3_5[13] , 
        \wRegInBot_3_5[12] , \wRegInBot_3_5[11] , \wRegInBot_3_5[10] , 
        \wRegInBot_3_5[9] , \wRegInBot_3_5[8] , \wRegInBot_3_5[7] , 
        \wRegInBot_3_5[6] , \wRegInBot_3_5[5] , \wRegInBot_3_5[4] , 
        \wRegInBot_3_5[3] , \wRegInBot_3_5[2] , \wRegInBot_3_5[1] , 
        \wRegInBot_3_5[0] }), .L_WR(\wRegEnTop_4_10[0] ), .L_In({
        \wRegOut_4_10[31] , \wRegOut_4_10[30] , \wRegOut_4_10[29] , 
        \wRegOut_4_10[28] , \wRegOut_4_10[27] , \wRegOut_4_10[26] , 
        \wRegOut_4_10[25] , \wRegOut_4_10[24] , \wRegOut_4_10[23] , 
        \wRegOut_4_10[22] , \wRegOut_4_10[21] , \wRegOut_4_10[20] , 
        \wRegOut_4_10[19] , \wRegOut_4_10[18] , \wRegOut_4_10[17] , 
        \wRegOut_4_10[16] , \wRegOut_4_10[15] , \wRegOut_4_10[14] , 
        \wRegOut_4_10[13] , \wRegOut_4_10[12] , \wRegOut_4_10[11] , 
        \wRegOut_4_10[10] , \wRegOut_4_10[9] , \wRegOut_4_10[8] , 
        \wRegOut_4_10[7] , \wRegOut_4_10[6] , \wRegOut_4_10[5] , 
        \wRegOut_4_10[4] , \wRegOut_4_10[3] , \wRegOut_4_10[2] , 
        \wRegOut_4_10[1] , \wRegOut_4_10[0] }), .L_Out({\wRegInTop_4_10[31] , 
        \wRegInTop_4_10[30] , \wRegInTop_4_10[29] , \wRegInTop_4_10[28] , 
        \wRegInTop_4_10[27] , \wRegInTop_4_10[26] , \wRegInTop_4_10[25] , 
        \wRegInTop_4_10[24] , \wRegInTop_4_10[23] , \wRegInTop_4_10[22] , 
        \wRegInTop_4_10[21] , \wRegInTop_4_10[20] , \wRegInTop_4_10[19] , 
        \wRegInTop_4_10[18] , \wRegInTop_4_10[17] , \wRegInTop_4_10[16] , 
        \wRegInTop_4_10[15] , \wRegInTop_4_10[14] , \wRegInTop_4_10[13] , 
        \wRegInTop_4_10[12] , \wRegInTop_4_10[11] , \wRegInTop_4_10[10] , 
        \wRegInTop_4_10[9] , \wRegInTop_4_10[8] , \wRegInTop_4_10[7] , 
        \wRegInTop_4_10[6] , \wRegInTop_4_10[5] , \wRegInTop_4_10[4] , 
        \wRegInTop_4_10[3] , \wRegInTop_4_10[2] , \wRegInTop_4_10[1] , 
        \wRegInTop_4_10[0] }), .R_WR(\wRegEnTop_4_11[0] ), .R_In({
        \wRegOut_4_11[31] , \wRegOut_4_11[30] , \wRegOut_4_11[29] , 
        \wRegOut_4_11[28] , \wRegOut_4_11[27] , \wRegOut_4_11[26] , 
        \wRegOut_4_11[25] , \wRegOut_4_11[24] , \wRegOut_4_11[23] , 
        \wRegOut_4_11[22] , \wRegOut_4_11[21] , \wRegOut_4_11[20] , 
        \wRegOut_4_11[19] , \wRegOut_4_11[18] , \wRegOut_4_11[17] , 
        \wRegOut_4_11[16] , \wRegOut_4_11[15] , \wRegOut_4_11[14] , 
        \wRegOut_4_11[13] , \wRegOut_4_11[12] , \wRegOut_4_11[11] , 
        \wRegOut_4_11[10] , \wRegOut_4_11[9] , \wRegOut_4_11[8] , 
        \wRegOut_4_11[7] , \wRegOut_4_11[6] , \wRegOut_4_11[5] , 
        \wRegOut_4_11[4] , \wRegOut_4_11[3] , \wRegOut_4_11[2] , 
        \wRegOut_4_11[1] , \wRegOut_4_11[0] }), .R_Out({\wRegInTop_4_11[31] , 
        \wRegInTop_4_11[30] , \wRegInTop_4_11[29] , \wRegInTop_4_11[28] , 
        \wRegInTop_4_11[27] , \wRegInTop_4_11[26] , \wRegInTop_4_11[25] , 
        \wRegInTop_4_11[24] , \wRegInTop_4_11[23] , \wRegInTop_4_11[22] , 
        \wRegInTop_4_11[21] , \wRegInTop_4_11[20] , \wRegInTop_4_11[19] , 
        \wRegInTop_4_11[18] , \wRegInTop_4_11[17] , \wRegInTop_4_11[16] , 
        \wRegInTop_4_11[15] , \wRegInTop_4_11[14] , \wRegInTop_4_11[13] , 
        \wRegInTop_4_11[12] , \wRegInTop_4_11[11] , \wRegInTop_4_11[10] , 
        \wRegInTop_4_11[9] , \wRegInTop_4_11[8] , \wRegInTop_4_11[7] , 
        \wRegInTop_4_11[6] , \wRegInTop_4_11[5] , \wRegInTop_4_11[4] , 
        \wRegInTop_4_11[3] , \wRegInTop_4_11[2] , \wRegInTop_4_11[1] , 
        \wRegInTop_4_11[0] }) );
    BHeap_CtrlReg_WIDTH32 BHCR_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_2[0] ), 
        .Out(\wCtrlOut_1[0] ), .Enable(\wEnable_1[0] ) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_4_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink26[31] , \ScanLink26[30] , \ScanLink26[29] , 
        \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , \ScanLink26[25] , 
        \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , \ScanLink26[21] , 
        \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , \ScanLink26[17] , 
        \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , \ScanLink26[13] , 
        \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , \ScanLink26[9] , 
        \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , \ScanLink26[5] , 
        \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , \ScanLink26[1] , 
        \ScanLink26[0] }), .ScanOut({\ScanLink25[31] , \ScanLink25[30] , 
        \ScanLink25[29] , \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , 
        \ScanLink25[25] , \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , 
        \ScanLink25[21] , \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , 
        \ScanLink25[17] , \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , 
        \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , 
        \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , 
        \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , 
        \ScanLink25[1] , \ScanLink25[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_4_10[31] , \wRegOut_4_10[30] , 
        \wRegOut_4_10[29] , \wRegOut_4_10[28] , \wRegOut_4_10[27] , 
        \wRegOut_4_10[26] , \wRegOut_4_10[25] , \wRegOut_4_10[24] , 
        \wRegOut_4_10[23] , \wRegOut_4_10[22] , \wRegOut_4_10[21] , 
        \wRegOut_4_10[20] , \wRegOut_4_10[19] , \wRegOut_4_10[18] , 
        \wRegOut_4_10[17] , \wRegOut_4_10[16] , \wRegOut_4_10[15] , 
        \wRegOut_4_10[14] , \wRegOut_4_10[13] , \wRegOut_4_10[12] , 
        \wRegOut_4_10[11] , \wRegOut_4_10[10] , \wRegOut_4_10[9] , 
        \wRegOut_4_10[8] , \wRegOut_4_10[7] , \wRegOut_4_10[6] , 
        \wRegOut_4_10[5] , \wRegOut_4_10[4] , \wRegOut_4_10[3] , 
        \wRegOut_4_10[2] , \wRegOut_4_10[1] , \wRegOut_4_10[0] }), .Enable1(
        \wRegEnTop_4_10[0] ), .Enable2(\wRegEnBot_4_10[0] ), .In1({
        \wRegInTop_4_10[31] , \wRegInTop_4_10[30] , \wRegInTop_4_10[29] , 
        \wRegInTop_4_10[28] , \wRegInTop_4_10[27] , \wRegInTop_4_10[26] , 
        \wRegInTop_4_10[25] , \wRegInTop_4_10[24] , \wRegInTop_4_10[23] , 
        \wRegInTop_4_10[22] , \wRegInTop_4_10[21] , \wRegInTop_4_10[20] , 
        \wRegInTop_4_10[19] , \wRegInTop_4_10[18] , \wRegInTop_4_10[17] , 
        \wRegInTop_4_10[16] , \wRegInTop_4_10[15] , \wRegInTop_4_10[14] , 
        \wRegInTop_4_10[13] , \wRegInTop_4_10[12] , \wRegInTop_4_10[11] , 
        \wRegInTop_4_10[10] , \wRegInTop_4_10[9] , \wRegInTop_4_10[8] , 
        \wRegInTop_4_10[7] , \wRegInTop_4_10[6] , \wRegInTop_4_10[5] , 
        \wRegInTop_4_10[4] , \wRegInTop_4_10[3] , \wRegInTop_4_10[2] , 
        \wRegInTop_4_10[1] , \wRegInTop_4_10[0] }), .In2({\wRegInBot_4_10[31] , 
        \wRegInBot_4_10[30] , \wRegInBot_4_10[29] , \wRegInBot_4_10[28] , 
        \wRegInBot_4_10[27] , \wRegInBot_4_10[26] , \wRegInBot_4_10[25] , 
        \wRegInBot_4_10[24] , \wRegInBot_4_10[23] , \wRegInBot_4_10[22] , 
        \wRegInBot_4_10[21] , \wRegInBot_4_10[20] , \wRegInBot_4_10[19] , 
        \wRegInBot_4_10[18] , \wRegInBot_4_10[17] , \wRegInBot_4_10[16] , 
        \wRegInBot_4_10[15] , \wRegInBot_4_10[14] , \wRegInBot_4_10[13] , 
        \wRegInBot_4_10[12] , \wRegInBot_4_10[11] , \wRegInBot_4_10[10] , 
        \wRegInBot_4_10[9] , \wRegInBot_4_10[8] , \wRegInBot_4_10[7] , 
        \wRegInBot_4_10[6] , \wRegInBot_4_10[5] , \wRegInBot_4_10[4] , 
        \wRegInBot_4_10[3] , \wRegInBot_4_10[2] , \wRegInBot_4_10[1] , 
        \wRegInBot_4_10[0] }) );
    BHeap_Node_WIDTH32 BHN_0_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_0[0] ), .P_WR(\wRegEnBot_0_0[0] ), .P_In({\wRegOut_0_0[31] , 
        \wRegOut_0_0[30] , \wRegOut_0_0[29] , \wRegOut_0_0[28] , 
        \wRegOut_0_0[27] , \wRegOut_0_0[26] , \wRegOut_0_0[25] , 
        \wRegOut_0_0[24] , \wRegOut_0_0[23] , \wRegOut_0_0[22] , 
        \wRegOut_0_0[21] , \wRegOut_0_0[20] , \wRegOut_0_0[19] , 
        \wRegOut_0_0[18] , \wRegOut_0_0[17] , \wRegOut_0_0[16] , 
        \wRegOut_0_0[15] , \wRegOut_0_0[14] , \wRegOut_0_0[13] , 
        \wRegOut_0_0[12] , \wRegOut_0_0[11] , \wRegOut_0_0[10] , 
        \wRegOut_0_0[9] , \wRegOut_0_0[8] , \wRegOut_0_0[7] , \wRegOut_0_0[6] , 
        \wRegOut_0_0[5] , \wRegOut_0_0[4] , \wRegOut_0_0[3] , \wRegOut_0_0[2] , 
        \wRegOut_0_0[1] , \wRegOut_0_0[0] }), .P_Out({\wRegInBot_0_0[31] , 
        \wRegInBot_0_0[30] , \wRegInBot_0_0[29] , \wRegInBot_0_0[28] , 
        \wRegInBot_0_0[27] , \wRegInBot_0_0[26] , \wRegInBot_0_0[25] , 
        \wRegInBot_0_0[24] , \wRegInBot_0_0[23] , \wRegInBot_0_0[22] , 
        \wRegInBot_0_0[21] , \wRegInBot_0_0[20] , \wRegInBot_0_0[19] , 
        \wRegInBot_0_0[18] , \wRegInBot_0_0[17] , \wRegInBot_0_0[16] , 
        \wRegInBot_0_0[15] , \wRegInBot_0_0[14] , \wRegInBot_0_0[13] , 
        \wRegInBot_0_0[12] , \wRegInBot_0_0[11] , \wRegInBot_0_0[10] , 
        \wRegInBot_0_0[9] , \wRegInBot_0_0[8] , \wRegInBot_0_0[7] , 
        \wRegInBot_0_0[6] , \wRegInBot_0_0[5] , \wRegInBot_0_0[4] , 
        \wRegInBot_0_0[3] , \wRegInBot_0_0[2] , \wRegInBot_0_0[1] , 
        \wRegInBot_0_0[0] }), .L_WR(\wRegEnTop_1_0[0] ), .L_In({
        \wRegOut_1_0[31] , \wRegOut_1_0[30] , \wRegOut_1_0[29] , 
        \wRegOut_1_0[28] , \wRegOut_1_0[27] , \wRegOut_1_0[26] , 
        \wRegOut_1_0[25] , \wRegOut_1_0[24] , \wRegOut_1_0[23] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[21] , \wRegOut_1_0[20] , 
        \wRegOut_1_0[19] , \wRegOut_1_0[18] , \wRegOut_1_0[17] , 
        \wRegOut_1_0[16] , \wRegOut_1_0[15] , \wRegOut_1_0[14] , 
        \wRegOut_1_0[13] , \wRegOut_1_0[12] , \wRegOut_1_0[11] , 
        \wRegOut_1_0[10] , \wRegOut_1_0[9] , \wRegOut_1_0[8] , 
        \wRegOut_1_0[7] , \wRegOut_1_0[6] , \wRegOut_1_0[5] , \wRegOut_1_0[4] , 
        \wRegOut_1_0[3] , \wRegOut_1_0[2] , \wRegOut_1_0[1] , \wRegOut_1_0[0] 
        }), .L_Out({\wRegInTop_1_0[31] , \wRegInTop_1_0[30] , 
        \wRegInTop_1_0[29] , \wRegInTop_1_0[28] , \wRegInTop_1_0[27] , 
        \wRegInTop_1_0[26] , \wRegInTop_1_0[25] , \wRegInTop_1_0[24] , 
        \wRegInTop_1_0[23] , \wRegInTop_1_0[22] , \wRegInTop_1_0[21] , 
        \wRegInTop_1_0[20] , \wRegInTop_1_0[19] , \wRegInTop_1_0[18] , 
        \wRegInTop_1_0[17] , \wRegInTop_1_0[16] , \wRegInTop_1_0[15] , 
        \wRegInTop_1_0[14] , \wRegInTop_1_0[13] , \wRegInTop_1_0[12] , 
        \wRegInTop_1_0[11] , \wRegInTop_1_0[10] , \wRegInTop_1_0[9] , 
        \wRegInTop_1_0[8] , \wRegInTop_1_0[7] , \wRegInTop_1_0[6] , 
        \wRegInTop_1_0[5] , \wRegInTop_1_0[4] , \wRegInTop_1_0[3] , 
        \wRegInTop_1_0[2] , \wRegInTop_1_0[1] , \wRegInTop_1_0[0] }), .R_WR(
        \wRegEnTop_1_1[0] ), .R_In({\wRegOut_1_1[31] , \wRegOut_1_1[30] , 
        \wRegOut_1_1[29] , \wRegOut_1_1[28] , \wRegOut_1_1[27] , 
        \wRegOut_1_1[26] , \wRegOut_1_1[25] , \wRegOut_1_1[24] , 
        \wRegOut_1_1[23] , \wRegOut_1_1[22] , \wRegOut_1_1[21] , 
        \wRegOut_1_1[20] , \wRegOut_1_1[19] , \wRegOut_1_1[18] , 
        \wRegOut_1_1[17] , \wRegOut_1_1[16] , \wRegOut_1_1[15] , 
        \wRegOut_1_1[14] , \wRegOut_1_1[13] , \wRegOut_1_1[12] , 
        \wRegOut_1_1[11] , \wRegOut_1_1[10] , \wRegOut_1_1[9] , 
        \wRegOut_1_1[8] , \wRegOut_1_1[7] , \wRegOut_1_1[6] , \wRegOut_1_1[5] , 
        \wRegOut_1_1[4] , \wRegOut_1_1[3] , \wRegOut_1_1[2] , \wRegOut_1_1[1] , 
        \wRegOut_1_1[0] }), .R_Out({\wRegInTop_1_1[31] , \wRegInTop_1_1[30] , 
        \wRegInTop_1_1[29] , \wRegInTop_1_1[28] , \wRegInTop_1_1[27] , 
        \wRegInTop_1_1[26] , \wRegInTop_1_1[25] , \wRegInTop_1_1[24] , 
        \wRegInTop_1_1[23] , \wRegInTop_1_1[22] , \wRegInTop_1_1[21] , 
        \wRegInTop_1_1[20] , \wRegInTop_1_1[19] , \wRegInTop_1_1[18] , 
        \wRegInTop_1_1[17] , \wRegInTop_1_1[16] , \wRegInTop_1_1[15] , 
        \wRegInTop_1_1[14] , \wRegInTop_1_1[13] , \wRegInTop_1_1[12] , 
        \wRegInTop_1_1[11] , \wRegInTop_1_1[10] , \wRegInTop_1_1[9] , 
        \wRegInTop_1_1[8] , \wRegInTop_1_1[7] , \wRegInTop_1_1[6] , 
        \wRegInTop_1_1[5] , \wRegInTop_1_1[4] , \wRegInTop_1_1[3] , 
        \wRegInTop_1_1[2] , \wRegInTop_1_1[1] , \wRegInTop_1_1[0] }) );
    BHeap_Control_CWIDTH3_IDWIDTH1_WIDTH32_SCAN1 BHC ( .Clk(Clk), .Reset(Reset
        ), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink0[31] , \ScanLink0[30] , \ScanLink0[29] , 
        \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , \ScanLink0[25] , 
        \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , \ScanLink0[21] , 
        \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , \ScanLink0[17] , 
        \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , \ScanLink0[13] , 
        \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , \ScanLink0[9] , 
        \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , \ScanLink0[5] , 
        \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , \ScanLink0[1] , 
        \ScanLink0[0] }), .ScanOut({\ScanLink63[31] , \ScanLink63[30] , 
        \ScanLink63[29] , \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , 
        \ScanLink63[25] , \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , 
        \ScanLink63[21] , \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , 
        \ScanLink63[17] , \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , 
        \ScanLink63[13] , \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , 
        \ScanLink63[9] , \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , 
        \ScanLink63[5] , \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , 
        \ScanLink63[1] , \ScanLink63[0] }), .ScanEnable(\ScanEnable[0] ), 
        .ScanId(1'b0), .Id(1'b1), .Go(\wCtrlOut_5[0] ), .Done(\wCtrlOut_0[0] )
         );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_5_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink36[31] , \ScanLink36[30] , \ScanLink36[29] , 
        \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , \ScanLink36[25] , 
        \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , \ScanLink36[21] , 
        \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , \ScanLink36[17] , 
        \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , \ScanLink36[13] , 
        \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , \ScanLink36[9] , 
        \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , \ScanLink36[5] , 
        \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , \ScanLink36[1] , 
        \ScanLink36[0] }), .ScanOut({\ScanLink35[31] , \ScanLink35[30] , 
        \ScanLink35[29] , \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , 
        \ScanLink35[25] , \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , 
        \ScanLink35[21] , \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , 
        \ScanLink35[17] , \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , 
        \ScanLink35[13] , \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , 
        \ScanLink35[9] , \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , 
        \ScanLink35[5] , \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , 
        \ScanLink35[1] , \ScanLink35[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_5_4[31] , \wRegOut_5_4[30] , \wRegOut_5_4[29] , 
        \wRegOut_5_4[28] , \wRegOut_5_4[27] , \wRegOut_5_4[26] , 
        \wRegOut_5_4[25] , \wRegOut_5_4[24] , \wRegOut_5_4[23] , 
        \wRegOut_5_4[22] , \wRegOut_5_4[21] , \wRegOut_5_4[20] , 
        \wRegOut_5_4[19] , \wRegOut_5_4[18] , \wRegOut_5_4[17] , 
        \wRegOut_5_4[16] , \wRegOut_5_4[15] , \wRegOut_5_4[14] , 
        \wRegOut_5_4[13] , \wRegOut_5_4[12] , \wRegOut_5_4[11] , 
        \wRegOut_5_4[10] , \wRegOut_5_4[9] , \wRegOut_5_4[8] , 
        \wRegOut_5_4[7] , \wRegOut_5_4[6] , \wRegOut_5_4[5] , \wRegOut_5_4[4] , 
        \wRegOut_5_4[3] , \wRegOut_5_4[2] , \wRegOut_5_4[1] , \wRegOut_5_4[0] 
        }), .Enable1(\wRegEnTop_5_4[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_5_4[31] , \wRegInTop_5_4[30] , \wRegInTop_5_4[29] , 
        \wRegInTop_5_4[28] , \wRegInTop_5_4[27] , \wRegInTop_5_4[26] , 
        \wRegInTop_5_4[25] , \wRegInTop_5_4[24] , \wRegInTop_5_4[23] , 
        \wRegInTop_5_4[22] , \wRegInTop_5_4[21] , \wRegInTop_5_4[20] , 
        \wRegInTop_5_4[19] , \wRegInTop_5_4[18] , \wRegInTop_5_4[17] , 
        \wRegInTop_5_4[16] , \wRegInTop_5_4[15] , \wRegInTop_5_4[14] , 
        \wRegInTop_5_4[13] , \wRegInTop_5_4[12] , \wRegInTop_5_4[11] , 
        \wRegInTop_5_4[10] , \wRegInTop_5_4[9] , \wRegInTop_5_4[8] , 
        \wRegInTop_5_4[7] , \wRegInTop_5_4[6] , \wRegInTop_5_4[5] , 
        \wRegInTop_5_4[4] , \wRegInTop_5_4[3] , \wRegInTop_5_4[2] , 
        \wRegInTop_5_4[1] , \wRegInTop_5_4[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_1[0] ), .P_WR(\wRegEnBot_1_0[0] ), .P_In({\wRegOut_1_0[31] , 
        \wRegOut_1_0[30] , \wRegOut_1_0[29] , \wRegOut_1_0[28] , 
        \wRegOut_1_0[27] , \wRegOut_1_0[26] , \wRegOut_1_0[25] , 
        \wRegOut_1_0[24] , \wRegOut_1_0[23] , \wRegOut_1_0[22] , 
        \wRegOut_1_0[21] , \wRegOut_1_0[20] , \wRegOut_1_0[19] , 
        \wRegOut_1_0[18] , \wRegOut_1_0[17] , \wRegOut_1_0[16] , 
        \wRegOut_1_0[15] , \wRegOut_1_0[14] , \wRegOut_1_0[13] , 
        \wRegOut_1_0[12] , \wRegOut_1_0[11] , \wRegOut_1_0[10] , 
        \wRegOut_1_0[9] , \wRegOut_1_0[8] , \wRegOut_1_0[7] , \wRegOut_1_0[6] , 
        \wRegOut_1_0[5] , \wRegOut_1_0[4] , \wRegOut_1_0[3] , \wRegOut_1_0[2] , 
        \wRegOut_1_0[1] , \wRegOut_1_0[0] }), .P_Out({\wRegInBot_1_0[31] , 
        \wRegInBot_1_0[30] , \wRegInBot_1_0[29] , \wRegInBot_1_0[28] , 
        \wRegInBot_1_0[27] , \wRegInBot_1_0[26] , \wRegInBot_1_0[25] , 
        \wRegInBot_1_0[24] , \wRegInBot_1_0[23] , \wRegInBot_1_0[22] , 
        \wRegInBot_1_0[21] , \wRegInBot_1_0[20] , \wRegInBot_1_0[19] , 
        \wRegInBot_1_0[18] , \wRegInBot_1_0[17] , \wRegInBot_1_0[16] , 
        \wRegInBot_1_0[15] , \wRegInBot_1_0[14] , \wRegInBot_1_0[13] , 
        \wRegInBot_1_0[12] , \wRegInBot_1_0[11] , \wRegInBot_1_0[10] , 
        \wRegInBot_1_0[9] , \wRegInBot_1_0[8] , \wRegInBot_1_0[7] , 
        \wRegInBot_1_0[6] , \wRegInBot_1_0[5] , \wRegInBot_1_0[4] , 
        \wRegInBot_1_0[3] , \wRegInBot_1_0[2] , \wRegInBot_1_0[1] , 
        \wRegInBot_1_0[0] }), .L_WR(\wRegEnTop_2_0[0] ), .L_In({
        \wRegOut_2_0[31] , \wRegOut_2_0[30] , \wRegOut_2_0[29] , 
        \wRegOut_2_0[28] , \wRegOut_2_0[27] , \wRegOut_2_0[26] , 
        \wRegOut_2_0[25] , \wRegOut_2_0[24] , \wRegOut_2_0[23] , 
        \wRegOut_2_0[22] , \wRegOut_2_0[21] , \wRegOut_2_0[20] , 
        \wRegOut_2_0[19] , \wRegOut_2_0[18] , \wRegOut_2_0[17] , 
        \wRegOut_2_0[16] , \wRegOut_2_0[15] , \wRegOut_2_0[14] , 
        \wRegOut_2_0[13] , \wRegOut_2_0[12] , \wRegOut_2_0[11] , 
        \wRegOut_2_0[10] , \wRegOut_2_0[9] , \wRegOut_2_0[8] , 
        \wRegOut_2_0[7] , \wRegOut_2_0[6] , \wRegOut_2_0[5] , \wRegOut_2_0[4] , 
        \wRegOut_2_0[3] , \wRegOut_2_0[2] , \wRegOut_2_0[1] , \wRegOut_2_0[0] 
        }), .L_Out({\wRegInTop_2_0[31] , \wRegInTop_2_0[30] , 
        \wRegInTop_2_0[29] , \wRegInTop_2_0[28] , \wRegInTop_2_0[27] , 
        \wRegInTop_2_0[26] , \wRegInTop_2_0[25] , \wRegInTop_2_0[24] , 
        \wRegInTop_2_0[23] , \wRegInTop_2_0[22] , \wRegInTop_2_0[21] , 
        \wRegInTop_2_0[20] , \wRegInTop_2_0[19] , \wRegInTop_2_0[18] , 
        \wRegInTop_2_0[17] , \wRegInTop_2_0[16] , \wRegInTop_2_0[15] , 
        \wRegInTop_2_0[14] , \wRegInTop_2_0[13] , \wRegInTop_2_0[12] , 
        \wRegInTop_2_0[11] , \wRegInTop_2_0[10] , \wRegInTop_2_0[9] , 
        \wRegInTop_2_0[8] , \wRegInTop_2_0[7] , \wRegInTop_2_0[6] , 
        \wRegInTop_2_0[5] , \wRegInTop_2_0[4] , \wRegInTop_2_0[3] , 
        \wRegInTop_2_0[2] , \wRegInTop_2_0[1] , \wRegInTop_2_0[0] }), .R_WR(
        \wRegEnTop_2_1[0] ), .R_In({\wRegOut_2_1[31] , \wRegOut_2_1[30] , 
        \wRegOut_2_1[29] , \wRegOut_2_1[28] , \wRegOut_2_1[27] , 
        \wRegOut_2_1[26] , \wRegOut_2_1[25] , \wRegOut_2_1[24] , 
        \wRegOut_2_1[23] , \wRegOut_2_1[22] , \wRegOut_2_1[21] , 
        \wRegOut_2_1[20] , \wRegOut_2_1[19] , \wRegOut_2_1[18] , 
        \wRegOut_2_1[17] , \wRegOut_2_1[16] , \wRegOut_2_1[15] , 
        \wRegOut_2_1[14] , \wRegOut_2_1[13] , \wRegOut_2_1[12] , 
        \wRegOut_2_1[11] , \wRegOut_2_1[10] , \wRegOut_2_1[9] , 
        \wRegOut_2_1[8] , \wRegOut_2_1[7] , \wRegOut_2_1[6] , \wRegOut_2_1[5] , 
        \wRegOut_2_1[4] , \wRegOut_2_1[3] , \wRegOut_2_1[2] , \wRegOut_2_1[1] , 
        \wRegOut_2_1[0] }), .R_Out({\wRegInTop_2_1[31] , \wRegInTop_2_1[30] , 
        \wRegInTop_2_1[29] , \wRegInTop_2_1[28] , \wRegInTop_2_1[27] , 
        \wRegInTop_2_1[26] , \wRegInTop_2_1[25] , \wRegInTop_2_1[24] , 
        \wRegInTop_2_1[23] , \wRegInTop_2_1[22] , \wRegInTop_2_1[21] , 
        \wRegInTop_2_1[20] , \wRegInTop_2_1[19] , \wRegInTop_2_1[18] , 
        \wRegInTop_2_1[17] , \wRegInTop_2_1[16] , \wRegInTop_2_1[15] , 
        \wRegInTop_2_1[14] , \wRegInTop_2_1[13] , \wRegInTop_2_1[12] , 
        \wRegInTop_2_1[11] , \wRegInTop_2_1[10] , \wRegInTop_2_1[9] , 
        \wRegInTop_2_1[8] , \wRegInTop_2_1[7] , \wRegInTop_2_1[6] , 
        \wRegInTop_2_1[5] , \wRegInTop_2_1[4] , \wRegInTop_2_1[3] , 
        \wRegInTop_2_1[2] , \wRegInTop_2_1[1] , \wRegInTop_2_1[0] }) );
    BHeap_Node_WIDTH32 BHN_4_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_4[0] ), .P_WR(\wRegEnBot_4_6[0] ), .P_In({\wRegOut_4_6[31] , 
        \wRegOut_4_6[30] , \wRegOut_4_6[29] , \wRegOut_4_6[28] , 
        \wRegOut_4_6[27] , \wRegOut_4_6[26] , \wRegOut_4_6[25] , 
        \wRegOut_4_6[24] , \wRegOut_4_6[23] , \wRegOut_4_6[22] , 
        \wRegOut_4_6[21] , \wRegOut_4_6[20] , \wRegOut_4_6[19] , 
        \wRegOut_4_6[18] , \wRegOut_4_6[17] , \wRegOut_4_6[16] , 
        \wRegOut_4_6[15] , \wRegOut_4_6[14] , \wRegOut_4_6[13] , 
        \wRegOut_4_6[12] , \wRegOut_4_6[11] , \wRegOut_4_6[10] , 
        \wRegOut_4_6[9] , \wRegOut_4_6[8] , \wRegOut_4_6[7] , \wRegOut_4_6[6] , 
        \wRegOut_4_6[5] , \wRegOut_4_6[4] , \wRegOut_4_6[3] , \wRegOut_4_6[2] , 
        \wRegOut_4_6[1] , \wRegOut_4_6[0] }), .P_Out({\wRegInBot_4_6[31] , 
        \wRegInBot_4_6[30] , \wRegInBot_4_6[29] , \wRegInBot_4_6[28] , 
        \wRegInBot_4_6[27] , \wRegInBot_4_6[26] , \wRegInBot_4_6[25] , 
        \wRegInBot_4_6[24] , \wRegInBot_4_6[23] , \wRegInBot_4_6[22] , 
        \wRegInBot_4_6[21] , \wRegInBot_4_6[20] , \wRegInBot_4_6[19] , 
        \wRegInBot_4_6[18] , \wRegInBot_4_6[17] , \wRegInBot_4_6[16] , 
        \wRegInBot_4_6[15] , \wRegInBot_4_6[14] , \wRegInBot_4_6[13] , 
        \wRegInBot_4_6[12] , \wRegInBot_4_6[11] , \wRegInBot_4_6[10] , 
        \wRegInBot_4_6[9] , \wRegInBot_4_6[8] , \wRegInBot_4_6[7] , 
        \wRegInBot_4_6[6] , \wRegInBot_4_6[5] , \wRegInBot_4_6[4] , 
        \wRegInBot_4_6[3] , \wRegInBot_4_6[2] , \wRegInBot_4_6[1] , 
        \wRegInBot_4_6[0] }), .L_WR(\wRegEnTop_5_12[0] ), .L_In({
        \wRegOut_5_12[31] , \wRegOut_5_12[30] , \wRegOut_5_12[29] , 
        \wRegOut_5_12[28] , \wRegOut_5_12[27] , \wRegOut_5_12[26] , 
        \wRegOut_5_12[25] , \wRegOut_5_12[24] , \wRegOut_5_12[23] , 
        \wRegOut_5_12[22] , \wRegOut_5_12[21] , \wRegOut_5_12[20] , 
        \wRegOut_5_12[19] , \wRegOut_5_12[18] , \wRegOut_5_12[17] , 
        \wRegOut_5_12[16] , \wRegOut_5_12[15] , \wRegOut_5_12[14] , 
        \wRegOut_5_12[13] , \wRegOut_5_12[12] , \wRegOut_5_12[11] , 
        \wRegOut_5_12[10] , \wRegOut_5_12[9] , \wRegOut_5_12[8] , 
        \wRegOut_5_12[7] , \wRegOut_5_12[6] , \wRegOut_5_12[5] , 
        \wRegOut_5_12[4] , \wRegOut_5_12[3] , \wRegOut_5_12[2] , 
        \wRegOut_5_12[1] , \wRegOut_5_12[0] }), .L_Out({\wRegInTop_5_12[31] , 
        \wRegInTop_5_12[30] , \wRegInTop_5_12[29] , \wRegInTop_5_12[28] , 
        \wRegInTop_5_12[27] , \wRegInTop_5_12[26] , \wRegInTop_5_12[25] , 
        \wRegInTop_5_12[24] , \wRegInTop_5_12[23] , \wRegInTop_5_12[22] , 
        \wRegInTop_5_12[21] , \wRegInTop_5_12[20] , \wRegInTop_5_12[19] , 
        \wRegInTop_5_12[18] , \wRegInTop_5_12[17] , \wRegInTop_5_12[16] , 
        \wRegInTop_5_12[15] , \wRegInTop_5_12[14] , \wRegInTop_5_12[13] , 
        \wRegInTop_5_12[12] , \wRegInTop_5_12[11] , \wRegInTop_5_12[10] , 
        \wRegInTop_5_12[9] , \wRegInTop_5_12[8] , \wRegInTop_5_12[7] , 
        \wRegInTop_5_12[6] , \wRegInTop_5_12[5] , \wRegInTop_5_12[4] , 
        \wRegInTop_5_12[3] , \wRegInTop_5_12[2] , \wRegInTop_5_12[1] , 
        \wRegInTop_5_12[0] }), .R_WR(\wRegEnTop_5_13[0] ), .R_In({
        \wRegOut_5_13[31] , \wRegOut_5_13[30] , \wRegOut_5_13[29] , 
        \wRegOut_5_13[28] , \wRegOut_5_13[27] , \wRegOut_5_13[26] , 
        \wRegOut_5_13[25] , \wRegOut_5_13[24] , \wRegOut_5_13[23] , 
        \wRegOut_5_13[22] , \wRegOut_5_13[21] , \wRegOut_5_13[20] , 
        \wRegOut_5_13[19] , \wRegOut_5_13[18] , \wRegOut_5_13[17] , 
        \wRegOut_5_13[16] , \wRegOut_5_13[15] , \wRegOut_5_13[14] , 
        \wRegOut_5_13[13] , \wRegOut_5_13[12] , \wRegOut_5_13[11] , 
        \wRegOut_5_13[10] , \wRegOut_5_13[9] , \wRegOut_5_13[8] , 
        \wRegOut_5_13[7] , \wRegOut_5_13[6] , \wRegOut_5_13[5] , 
        \wRegOut_5_13[4] , \wRegOut_5_13[3] , \wRegOut_5_13[2] , 
        \wRegOut_5_13[1] , \wRegOut_5_13[0] }), .R_Out({\wRegInTop_5_13[31] , 
        \wRegInTop_5_13[30] , \wRegInTop_5_13[29] , \wRegInTop_5_13[28] , 
        \wRegInTop_5_13[27] , \wRegInTop_5_13[26] , \wRegInTop_5_13[25] , 
        \wRegInTop_5_13[24] , \wRegInTop_5_13[23] , \wRegInTop_5_13[22] , 
        \wRegInTop_5_13[21] , \wRegInTop_5_13[20] , \wRegInTop_5_13[19] , 
        \wRegInTop_5_13[18] , \wRegInTop_5_13[17] , \wRegInTop_5_13[16] , 
        \wRegInTop_5_13[15] , \wRegInTop_5_13[14] , \wRegInTop_5_13[13] , 
        \wRegInTop_5_13[12] , \wRegInTop_5_13[11] , \wRegInTop_5_13[10] , 
        \wRegInTop_5_13[9] , \wRegInTop_5_13[8] , \wRegInTop_5_13[7] , 
        \wRegInTop_5_13[6] , \wRegInTop_5_13[5] , \wRegInTop_5_13[4] , 
        \wRegInTop_5_13[3] , \wRegInTop_5_13[2] , \wRegInTop_5_13[1] , 
        \wRegInTop_5_13[0] }) );
endmodule

