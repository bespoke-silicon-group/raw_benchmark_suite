
module BubbleSort_Node_WIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n100, n112, n32, n29, n85, n47, n60, 
        n109, n40, n67, n82, n99, n27, n35, n49, n107, n90, n52, n75, n98, 
        n114, n34, n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, 
        n21, n46, n54, n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, n113, 
        n94, n23, n103, n16, n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, 
        n58, n104, n18, n24, n88, n37, n51, n93, n59, n76, n80, n42, n65, n19, 
        n50, n77, n89, n92, n25, n102, n105, n22, n39, n95, n45, n57, n70, n62, 
        n87, n17, n30, n79, n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_OR2 U54 ( .A(B[26]), .B(n96), .Z(n99) );
    VMW_INV U73 ( .A(B[27]), .Z(n105) );
    VMW_INV U96 ( .A(B[31]), .Z(n15) );
    VMW_INV U68 ( .A(A[30]), .Z(n113) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n66), .C(n62), .D(n57), .Z(n65) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U34 ( .A(B[16]), .B(n64), .Z(n67) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n75), .D(n70), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_NAND2 U61 ( .A(n110), .B(A[29]), .Z(n111) );
    VMW_INV U84 ( .A(B[15]), .Z(n66) );
    VMW_INV U101 ( .A(A[6]), .Z(n32) );
    VMW_INV U66 ( .A(B[7]), .Z(n41) );
    VMW_INV U83 ( .A(A[15]), .Z(n69) );
    VMW_INV U98 ( .A(B[13]), .Z(n60) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_NAND2 U48 ( .A(n90), .B(B[24]), .Z(n89) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n69), .C(n67), .D(n65), .Z(n68) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n98), .C(n94), .D(n89), .Z(n97) );
    VMW_INV U91 ( .A(B[11]), .Z(n54) );
    VMW_INV U74 ( .A(A[3]), .Z(n30) );
    VMW_INV U99 ( .A(A[26]), .Z(n96) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U40 ( .A(n78), .B(B[20]), .Z(n77) );
    VMW_INV U82 ( .A(B[29]), .Z(n110) );
    VMW_NAND2 U52 ( .A(n96), .B(B[26]), .Z(n95) );
    VMW_INV U67 ( .A(A[7]), .Z(n44) );
    VMW_INV U75 ( .A(B[3]), .Z(n27) );
    VMW_INV U90 ( .A(A[14]), .Z(n58) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n92), .C(n88), .D(n83), .Z(n91) );
    VMW_INV U69 ( .A(B[17]), .Z(n73) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n101), .C(n99), .D(n97), .Z(n100) );
    VMW_INV U72 ( .A(A[27]), .Z(n108) );
    VMW_INV U97 ( .A(A[16]), .Z(n64) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n110), .C(n107), .D(n102), .Z(n109) );
    VMW_INV U100 ( .A(B[23]), .Z(n92) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_INV U85 ( .A(A[4]), .Z(n25) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_NAND2 U32 ( .A(n64), .B(B[16]), .Z(n63) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n76), .C(n74), .D(n72), .Z(n75) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_INV U70 ( .A(A[17]), .Z(n76) );
    VMW_INV U95 ( .A(A[1]), .Z(n21) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_INV U79 ( .A(B[19]), .Z(n80) );
    VMW_INV U87 ( .A(A[8]), .Z(n39) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n77), .Z(n85) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n113), .C(n111), .D(n109), .Z(n112) );
    VMW_INV U65 ( .A(A[12]), .Z(n52) );
    VMW_INV U102 ( .A(A[2]), .Z(n18) );
    VMW_INV U80 ( .A(A[10]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n73), .C(n68), .D(n63), .Z(n72) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n108), .C(n106), .D(n104), .Z(n107) );
    VMW_INV U89 ( .A(A[18]), .Z(n71) );
    VMW_NAND2 U50 ( .A(n92), .B(A[23]), .Z(n93) );
    VMW_INV U77 ( .A(A[25]), .Z(n101) );
    VMW_INV U92 ( .A(A[28]), .Z(n103) );
    VMW_OR2 U58 ( .A(B[28]), .B(n103), .Z(n106) );
    VMW_NAND2 U36 ( .A(n71), .B(B[18]), .Z(n70) );
    VMW_INV U81 ( .A(B[9]), .Z(n48) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n78), .C(n81), .D(n79), .Z(n82) );
    VMW_AO22 U64 ( .A(n112), .B(n114), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n90), .C(n93), .D(n91), .Z(n94) );
    VMW_INV U76 ( .A(B[25]), .Z(n98) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_INV U88 ( .A(B[21]), .Z(n86) );
    VMW_INV U93 ( .A(A[5]), .Z(n37) );
    VMW_OR2 U38 ( .A(B[18]), .B(n71), .Z(n74) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n103), .B(B[28]), .Z(n102) );
    VMW_INV U94 ( .A(B[5]), .Z(n34) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_NAND2 U63 ( .A(n113), .B(B[30]), .Z(n114) );
    VMW_INV U86 ( .A(A[24]), .Z(n90) );
    VMW_INV U103 ( .A(A[0]), .Z(n20) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_INV U78 ( .A(A[20]), .Z(n78) );
endmodule


module BubbleSort_Node_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, 
    AIn, BIn, HiOut, LoOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
output [31:0] LoOut;
input  [31:0] AIn;
input  [31:0] BIn;
output [31:0] HiOut;
input  Clk, Reset, RD, WR;
    wire n159, a58;
    VMW_PULLDOWN U21 ( .Z(n159) );
    VMW_MUX2 U54 ( .A(BIn[9]), .B(AIn[9]), .S(a58), .Z(HiOut[9]) );
    VMW_MUX2 U73 ( .A(BIn[20]), .B(AIn[20]), .S(a58), .Z(HiOut[20]) );
    VMW_MUX2 U22 ( .A(AIn[9]), .B(BIn[9]), .S(a58), .Z(LoOut[9]) );
    VMW_MUX2 U26 ( .A(AIn[5]), .B(BIn[5]), .S(a58), .Z(LoOut[5]) );
    VMW_MUX2 U28 ( .A(AIn[3]), .B(BIn[3]), .S(a58), .Z(LoOut[3]) );
    VMW_MUX2 U33 ( .A(AIn[28]), .B(BIn[28]), .S(a58), .Z(LoOut[28]) );
    VMW_MUX2 U68 ( .A(BIn[25]), .B(AIn[25]), .S(a58), .Z(HiOut[25]) );
    VMW_MUX2 U34 ( .A(AIn[27]), .B(BIn[27]), .S(a58), .Z(LoOut[27]) );
    VMW_MUX2 U41 ( .A(AIn[20]), .B(BIn[20]), .S(a58), .Z(LoOut[20]) );
    VMW_MUX2 U46 ( .A(AIn[16]), .B(BIn[16]), .S(a58), .Z(LoOut[16]) );
    VMW_MUX2 U61 ( .A(BIn[31]), .B(AIn[31]), .S(a58), .Z(HiOut[31]) );
    VMW_MUX2 U84 ( .A(BIn[10]), .B(AIn[10]), .S(a58), .Z(HiOut[10]) );
    VMW_MUX2 U66 ( .A(BIn[27]), .B(AIn[27]), .S(a58), .Z(HiOut[27]) );
    VMW_MUX2 U83 ( .A(BIn[11]), .B(AIn[11]), .S(a58), .Z(HiOut[11]) );
    VMW_MUX2 U48 ( .A(AIn[14]), .B(BIn[14]), .S(a58), .Z(LoOut[14]) );
    VMW_MUX2 U27 ( .A(AIn[4]), .B(BIn[4]), .S(a58), .Z(LoOut[4]) );
    VMW_MUX2 U35 ( .A(AIn[26]), .B(BIn[26]), .S(a58), .Z(LoOut[26]) );
    VMW_MUX2 U53 ( .A(AIn[0]), .B(BIn[0]), .S(a58), .Z(LoOut[0]) );
    VMW_MUX2 U74 ( .A(BIn[1]), .B(AIn[1]), .S(a58), .Z(HiOut[1]) );
    VMW_MUX2 U40 ( .A(AIn[21]), .B(BIn[21]), .S(a58), .Z(LoOut[21]) );
    VMW_MUX2 U82 ( .A(BIn[12]), .B(AIn[12]), .S(a58), .Z(HiOut[12]) );
    VMW_MUX2 U52 ( .A(AIn[10]), .B(BIn[10]), .S(a58), .Z(LoOut[10]) );
    VMW_MUX2 U67 ( .A(BIn[26]), .B(AIn[26]), .S(a58), .Z(HiOut[26]) );
    VMW_MUX2 U75 ( .A(BIn[19]), .B(AIn[19]), .S(a58), .Z(HiOut[19]) );
    VMW_MUX2 U29 ( .A(AIn[31]), .B(BIn[31]), .S(a58), .Z(LoOut[31]) );
    VMW_MUX2 U47 ( .A(AIn[15]), .B(BIn[15]), .S(a58), .Z(LoOut[15]) );
    VMW_MUX2 U49 ( .A(AIn[13]), .B(BIn[13]), .S(a58), .Z(LoOut[13]) );
    VMW_MUX2 U55 ( .A(BIn[8]), .B(AIn[8]), .S(a58), .Z(HiOut[8]) );
    VMW_MUX2 U69 ( .A(BIn[24]), .B(AIn[24]), .S(a58), .Z(HiOut[24]) );
    VMW_MUX2 U72 ( .A(BIn[21]), .B(AIn[21]), .S(a58), .Z(HiOut[21]) );
    VMW_MUX2 U60 ( .A(BIn[3]), .B(AIn[3]), .S(a58), .Z(HiOut[3]) );
    VMW_MUX2 U32 ( .A(AIn[29]), .B(BIn[29]), .S(a58), .Z(LoOut[29]) );
    VMW_MUX2 U85 ( .A(BIn[0]), .B(AIn[0]), .S(a58), .Z(HiOut[0]) );
    VMW_MUX2 U39 ( .A(AIn[22]), .B(BIn[22]), .S(a58), .Z(LoOut[22]) );
    VMW_MUX2 U57 ( .A(BIn[6]), .B(AIn[6]), .S(a58), .Z(HiOut[6]) );
    VMW_MUX2 U70 ( .A(BIn[23]), .B(AIn[23]), .S(a58), .Z(HiOut[23]) );
    VMW_MUX2 U23 ( .A(AIn[8]), .B(BIn[8]), .S(a58), .Z(LoOut[8]) );
    VMW_MUX2 U24 ( .A(AIn[7]), .B(BIn[7]), .S(a58), .Z(LoOut[7]) );
    VMW_MUX2 U25 ( .A(AIn[6]), .B(BIn[6]), .S(a58), .Z(LoOut[6]) );
    VMW_MUX2 U30 ( .A(AIn[30]), .B(BIn[30]), .S(a58), .Z(LoOut[30]) );
    VMW_MUX2 U79 ( .A(BIn[15]), .B(AIn[15]), .S(a58), .Z(HiOut[15]) );
    BubbleSort_Node_WIDTH32_DW01_cmp2_32_0 gt_41 ( .A(BIn), .B(AIn), .LEQ(n159
        ), .TC(n159), .LT_LE(a58) );
    VMW_MUX2 U37 ( .A(AIn[24]), .B(BIn[24]), .S(a58), .Z(LoOut[24]) );
    VMW_MUX2 U42 ( .A(AIn[1]), .B(BIn[1]), .S(a58), .Z(LoOut[1]) );
    VMW_MUX2 U45 ( .A(AIn[17]), .B(BIn[17]), .S(a58), .Z(LoOut[17]) );
    VMW_MUX2 U62 ( .A(BIn[30]), .B(AIn[30]), .S(a58), .Z(HiOut[30]) );
    VMW_MUX2 U65 ( .A(BIn[28]), .B(AIn[28]), .S(a58), .Z(HiOut[28]) );
    VMW_MUX2 U80 ( .A(BIn[14]), .B(AIn[14]), .S(a58), .Z(HiOut[14]) );
    VMW_MUX2 U59 ( .A(BIn[4]), .B(AIn[4]), .S(a58), .Z(HiOut[4]) );
    VMW_MUX2 U36 ( .A(AIn[25]), .B(BIn[25]), .S(a58), .Z(LoOut[25]) );
    VMW_MUX2 U50 ( .A(AIn[12]), .B(BIn[12]), .S(a58), .Z(LoOut[12]) );
    VMW_MUX2 U77 ( .A(BIn[17]), .B(AIn[17]), .S(a58), .Z(HiOut[17]) );
    VMW_MUX2 U58 ( .A(BIn[5]), .B(AIn[5]), .S(a58), .Z(HiOut[5]) );
    VMW_MUX2 U43 ( .A(AIn[19]), .B(BIn[19]), .S(a58), .Z(LoOut[19]) );
    VMW_MUX2 U64 ( .A(BIn[29]), .B(AIn[29]), .S(a58), .Z(HiOut[29]) );
    VMW_MUX2 U81 ( .A(BIn[13]), .B(AIn[13]), .S(a58), .Z(HiOut[13]) );
    VMW_MUX2 U51 ( .A(AIn[11]), .B(BIn[11]), .S(a58), .Z(LoOut[11]) );
    VMW_MUX2 U76 ( .A(BIn[18]), .B(AIn[18]), .S(a58), .Z(HiOut[18]) );
    VMW_MUX2 U31 ( .A(AIn[2]), .B(BIn[2]), .S(a58), .Z(LoOut[2]) );
    VMW_MUX2 U38 ( .A(AIn[23]), .B(BIn[23]), .S(a58), .Z(LoOut[23]) );
    VMW_MUX2 U44 ( .A(AIn[18]), .B(BIn[18]), .S(a58), .Z(LoOut[18]) );
    VMW_MUX2 U56 ( .A(BIn[7]), .B(AIn[7]), .S(a58), .Z(HiOut[7]) );
    VMW_MUX2 U71 ( .A(BIn[22]), .B(AIn[22]), .S(a58), .Z(HiOut[22]) );
    VMW_MUX2 U63 ( .A(BIn[2]), .B(AIn[2]), .S(a58), .Z(HiOut[2]) );
    VMW_MUX2 U78 ( .A(BIn[16]), .B(AIn[16]), .S(a58), .Z(HiOut[16]) );
endmodule


module BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, In, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[31] , \ScanOut[5]1 , \ScanOut[4]1 , n245, n262, n217, n230, 
        n222, n199, n205, n257, n239, \ScanOut[23]1 , \ScanOut[8]1 , n202, 
        n250, n219, n225, n259, n210, n237, \ScanOut[10]1 , \ScanOut[22]1 , 
        \ScanOut[11]1 , n242, \ScanOut[9]1 , n197, n203, n224, n251, n206, 
        \ScanOut[19]1 , n196, n218, \ScanOut[26]1 , \ScanOut[18]1 , 
        \ScanOut[1]1 , \ScanOut[0]1 , n258, n243, \ScanOut[15]1 , n211, n236, 
        n216, n231, \ScanOut[27]1 , n244, \ScanOut[14]1 , n256, n238, n223, 
        n198, n204, n233, n228, n261, n246, n214, \ScanOut[28]1 , n221, 
        \ScanOut[3]1 , \ScanOut[30]1 , \ScanOut[29]1 , \ScanOut[2]1 , n254, 
        \ScanOut[25]1 , \ScanOut[24]1 , \ScanOut[17]1 , n253, n248, 
        \ScanOut[16]1 , n226, n201, n213, n234, n241, n194, n208, 
        \ScanOut[6]1 , n200, n227, n249, \ScanOut[7]1 , n252, n195, n209, n212, 
        n240, n235, n215, n260, n232, n247, \ScanOut[21]1 , n229, 
        \ScanOut[13]1 , \ScanOut[12]1 , n255, \ScanOut[20]1 , n207, n220;
    assign ScanOut[31] = \ScanOut[31] ;
    assign ScanOut[30] = \ScanOut[30]1 ;
    assign ScanOut[29] = \ScanOut[29]1 ;
    assign ScanOut[28] = \ScanOut[28]1 ;
    assign ScanOut[27] = \ScanOut[27]1 ;
    assign ScanOut[26] = \ScanOut[26]1 ;
    assign ScanOut[25] = \ScanOut[25]1 ;
    assign ScanOut[24] = \ScanOut[24]1 ;
    assign ScanOut[23] = \ScanOut[23]1 ;
    assign ScanOut[22] = \ScanOut[22]1 ;
    assign ScanOut[21] = \ScanOut[21]1 ;
    assign ScanOut[20] = \ScanOut[20]1 ;
    assign ScanOut[19] = \ScanOut[19]1 ;
    assign ScanOut[18] = \ScanOut[18]1 ;
    assign ScanOut[17] = \ScanOut[17]1 ;
    assign ScanOut[16] = \ScanOut[16]1 ;
    assign ScanOut[15] = \ScanOut[15]1 ;
    assign ScanOut[14] = \ScanOut[14]1 ;
    assign ScanOut[13] = \ScanOut[13]1 ;
    assign ScanOut[12] = \ScanOut[12]1 ;
    assign ScanOut[11] = \ScanOut[11]1 ;
    assign ScanOut[10] = \ScanOut[10]1 ;
    assign ScanOut[9] = \ScanOut[9]1 ;
    assign ScanOut[8] = \ScanOut[8]1 ;
    assign ScanOut[7] = \ScanOut[7]1 ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[31] = \ScanOut[31] ;
    assign Out[30] = \ScanOut[30]1 ;
    assign Out[29] = \ScanOut[29]1 ;
    assign Out[28] = \ScanOut[28]1 ;
    assign Out[27] = \ScanOut[27]1 ;
    assign Out[26] = \ScanOut[26]1 ;
    assign Out[25] = \ScanOut[25]1 ;
    assign Out[24] = \ScanOut[24]1 ;
    assign Out[23] = \ScanOut[23]1 ;
    assign Out[22] = \ScanOut[22]1 ;
    assign Out[21] = \ScanOut[21]1 ;
    assign Out[20] = \ScanOut[20]1 ;
    assign Out[19] = \ScanOut[19]1 ;
    assign Out[18] = \ScanOut[18]1 ;
    assign Out[17] = \ScanOut[17]1 ;
    assign Out[16] = \ScanOut[16]1 ;
    assign Out[15] = \ScanOut[15]1 ;
    assign Out[14] = \ScanOut[14]1 ;
    assign Out[13] = \ScanOut[13]1 ;
    assign Out[12] = \ScanOut[12]1 ;
    assign Out[11] = \ScanOut[11]1 ;
    assign Out[10] = \ScanOut[10]1 ;
    assign Out[9] = \ScanOut[9]1 ;
    assign Out[8] = \ScanOut[8]1 ;
    assign Out[7] = \ScanOut[7]1 ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO21 U54 ( .A(\ScanOut[25]1 ), .B(n194), .C(n220), .Z(n237) );
    VMW_AO22 U73 ( .A(ScanIn[30]), .B(n230), .C(In[30]), .D(n228), .Z(n225) );
    VMW_AO22 U68 ( .A(ScanIn[6]), .B(n230), .C(In[6]), .D(n228), .Z(n201) );
    VMW_AO22 U96 ( .A(ScanIn[0]), .B(n230), .C(In[0]), .D(n228), .Z(n195) );
    VMW_AO21 U33 ( .A(\ScanOut[4]1 ), .B(n194), .C(n199), .Z(n258) );
    VMW_AO21 U34 ( .A(\ScanOut[5]1 ), .B(n194), .C(n200), .Z(n257) );
    VMW_AO21 U41 ( .A(\ScanOut[12]1 ), .B(n194), .C(n207), .Z(n250) );
    VMW_AO21 U46 ( .A(\ScanOut[17]1 ), .B(n194), .C(n212), .Z(n245) );
    VMW_NOR2 U61 ( .A(Reset), .B(n194), .Z(n227) );
    VMW_AO22 U84 ( .A(ScanIn[20]), .B(n230), .C(In[20]), .D(n228), .Z(n215) );
    VMW_AO22 U66 ( .A(ScanIn[8]), .B(n230), .C(In[8]), .D(n228), .Z(n203) );
    VMW_AO22 U83 ( .A(ScanIn[21]), .B(n230), .C(In[21]), .D(n228), .Z(n216) );
    VMW_AO21 U35 ( .A(\ScanOut[6]1 ), .B(n194), .C(n201), .Z(n256) );
    VMW_AO21 U48 ( .A(\ScanOut[19]1 ), .B(n194), .C(n214), .Z(n243) );
    VMW_AO21 U53 ( .A(\ScanOut[24]1 ), .B(n194), .C(n219), .Z(n238) );
    VMW_AO22 U91 ( .A(ScanIn[14]), .B(n230), .C(In[14]), .D(n228), .Z(n209) );
    VMW_AO22 U74 ( .A(ScanIn[2]), .B(n230), .C(In[2]), .D(n228), .Z(n197) );
    VMW_FD \Out_reg[25]  ( .D(n237), .CP(Clk), .Q(\ScanOut[25]1 ) );
    VMW_FD \Out_reg[16]  ( .D(n246), .CP(Clk), .Q(\ScanOut[16]1 ) );
    VMW_AO21 U29 ( .A(\ScanOut[0]1 ), .B(n194), .C(n195), .Z(n262) );
    VMW_AO21 U40 ( .A(\ScanOut[11]1 ), .B(n194), .C(n206), .Z(n251) );
    VMW_AO22 U82 ( .A(ScanIn[22]), .B(n230), .C(In[22]), .D(n228), .Z(n217) );
    VMW_FD \Out_reg[5]  ( .D(n257), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO21 U47 ( .A(\ScanOut[18]1 ), .B(n194), .C(n213), .Z(n244) );
    VMW_AO21 U49 ( .A(\ScanOut[20]1 ), .B(n194), .C(n215), .Z(n242) );
    VMW_AO21 U52 ( .A(\ScanOut[23]1 ), .B(n194), .C(n218), .Z(n239) );
    VMW_AO22 U67 ( .A(ScanIn[7]), .B(n230), .C(In[7]), .D(n228), .Z(n202) );
    VMW_AO22 U75 ( .A(ScanIn[29]), .B(n230), .C(In[29]), .D(n228), .Z(n224) );
    VMW_FD \Out_reg[12]  ( .D(n250), .CP(Clk), .Q(\ScanOut[12]1 ) );
    VMW_AO22 U90 ( .A(ScanIn[15]), .B(n230), .C(In[15]), .D(n228), .Z(n210) );
    VMW_FD \Out_reg[21]  ( .D(n241), .CP(Clk), .Q(\ScanOut[21]1 ) );
    VMW_FD \Out_reg[31]  ( .D(n231), .CP(Clk), .Q(\ScanOut[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n234), .CP(Clk), .Q(\ScanOut[28]1 ) );
    VMW_FD \Out_reg[8]  ( .D(n254), .CP(Clk), .Q(\ScanOut[8]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n261), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_AO21 U55 ( .A(\ScanOut[26]1 ), .B(n194), .C(n221), .Z(n236) );
    VMW_AO22 U69 ( .A(ScanIn[5]), .B(n230), .C(In[5]), .D(n228), .Z(n200) );
    VMW_FD \Out_reg[19]  ( .D(n243), .CP(Clk), .Q(\ScanOut[19]1 ) );
    VMW_AO22 U72 ( .A(ScanIn[31]), .B(n230), .C(In[31]), .D(n228), .Z(n226) );
    VMW_INV U97 ( .A(n227), .Z(n229) );
    VMW_FD \Out_reg[3]  ( .D(n259), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_FD \Out_reg[23]  ( .D(n239), .CP(Clk), .Q(\ScanOut[23]1 ) );
    VMW_FD \Out_reg[10]  ( .D(n252), .CP(Clk), .Q(\ScanOut[10]1 ) );
    VMW_AO21 U60 ( .A(\ScanOut[31] ), .B(n194), .C(n226), .Z(n231) );
    VMW_FD \Out_reg[7]  ( .D(n255), .CP(Clk), .Q(\ScanOut[7]1 ) );
    VMW_AO21 U32 ( .A(\ScanOut[3]1 ), .B(n194), .C(n198), .Z(n259) );
    VMW_AO22 U85 ( .A(ScanIn[1]), .B(n230), .C(In[1]), .D(n228), .Z(n196) );
    VMW_FD \Out_reg[27]  ( .D(n235), .CP(Clk), .Q(\ScanOut[27]1 ) );
    VMW_FD \Out_reg[14]  ( .D(n248), .CP(Clk), .Q(\ScanOut[14]1 ) );
    VMW_AO21 U30 ( .A(\ScanOut[1]1 ), .B(n194), .C(n196), .Z(n261) );
    VMW_AO21 U39 ( .A(\ScanOut[10]1 ), .B(n194), .C(n205), .Z(n252) );
    VMW_AO21 U57 ( .A(\ScanOut[28]1 ), .B(n194), .C(n223), .Z(n234) );
    VMW_FD \Out_reg[6]  ( .D(n256), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U70 ( .A(ScanIn[4]), .B(n230), .C(In[4]), .D(n228), .Z(n199) );
    VMW_AO22 U79 ( .A(ScanIn[25]), .B(n230), .C(In[25]), .D(n228), .Z(n220) );
    VMW_AO22 U95 ( .A(ScanIn[10]), .B(n230), .C(In[10]), .D(n228), .Z(n205) );
    VMW_FD \Out_reg[26]  ( .D(n236), .CP(Clk), .Q(\ScanOut[26]1 ) );
    VMW_FD \Out_reg[15]  ( .D(n247), .CP(Clk), .Q(\ScanOut[15]1 ) );
    VMW_FD \Out_reg[18]  ( .D(n244), .CP(Clk), .Q(\ScanOut[18]1 ) );
    VMW_AO21 U31 ( .A(\ScanOut[2]1 ), .B(n194), .C(n197), .Z(n260) );
    VMW_AO21 U36 ( .A(\ScanOut[7]1 ), .B(n194), .C(n202), .Z(n255) );
    VMW_AO21 U37 ( .A(\ScanOut[8]1 ), .B(n194), .C(n203), .Z(n254) );
    VMW_AO21 U42 ( .A(\ScanOut[13]1 ), .B(n194), .C(n208), .Z(n249) );
    VMW_AO21 U45 ( .A(\ScanOut[16]1 ), .B(n194), .C(n211), .Z(n246) );
    VMW_AO22 U87 ( .A(ScanIn[18]), .B(n230), .C(In[18]), .D(n228), .Z(n213) );
    VMW_FD \Out_reg[2]  ( .D(n260), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_FD \Out_reg[11]  ( .D(n251), .CP(Clk), .Q(\ScanOut[11]1 ) );
    VMW_NOR2 U62 ( .A(n229), .B(ScanEnable), .Z(n228) );
    VMW_FD \Out_reg[22]  ( .D(n240), .CP(Clk), .Q(\ScanOut[22]1 ) );
    VMW_AO22 U65 ( .A(ScanIn[9]), .B(n230), .C(In[9]), .D(n228), .Z(n204) );
    VMW_FD \Out_reg[20]  ( .D(n242), .CP(Clk), .Q(\ScanOut[20]1 ) );
    VMW_FD \Out_reg[13]  ( .D(n249), .CP(Clk), .Q(\ScanOut[13]1 ) );
    VMW_AO22 U80 ( .A(ScanIn[24]), .B(n230), .C(In[24]), .D(n228), .Z(n219) );
    VMW_FD \Out_reg[9]  ( .D(n253), .CP(Clk), .Q(\ScanOut[9]1 ) );
    VMW_AO21 U50 ( .A(\ScanOut[21]1 ), .B(n194), .C(n216), .Z(n241) );
    VMW_AO21 U59 ( .A(\ScanOut[30]1 ), .B(n194), .C(n225), .Z(n232) );
    VMW_FD \Out_reg[30]  ( .D(n232), .CP(Clk), .Q(\ScanOut[30]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n262), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_FD \Out_reg[29]  ( .D(n233), .CP(Clk), .Q(\ScanOut[29]1 ) );
    VMW_AO22 U77 ( .A(ScanIn[27]), .B(n230), .C(In[27]), .D(n228), .Z(n222) );
    VMW_AO22 U89 ( .A(ScanIn[16]), .B(n230), .C(In[16]), .D(n228), .Z(n211) );
    VMW_AO22 U92 ( .A(ScanIn[13]), .B(n230), .C(In[13]), .D(n228), .Z(n208) );
    VMW_FD \Out_reg[24]  ( .D(n238), .CP(Clk), .Q(\ScanOut[24]1 ) );
    VMW_FD \Out_reg[17]  ( .D(n245), .CP(Clk), .Q(\ScanOut[17]1 ) );
    VMW_FD \Out_reg[4]  ( .D(n258), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_AO21 U58 ( .A(\ScanOut[29]1 ), .B(n194), .C(n224), .Z(n233) );
    VMW_AO21 U38 ( .A(\ScanOut[9]1 ), .B(n194), .C(n204), .Z(n253) );
    VMW_AO21 U43 ( .A(\ScanOut[14]1 ), .B(n194), .C(n209), .Z(n248) );
    VMW_NOR3 U64 ( .A(ScanEnable), .B(Reset), .C(Enable), .Z(n194) );
    VMW_AO22 U81 ( .A(ScanIn[23]), .B(n230), .C(In[23]), .D(n228), .Z(n218) );
    VMW_AO21 U51 ( .A(\ScanOut[22]1 ), .B(n194), .C(n217), .Z(n240) );
    VMW_AO22 U76 ( .A(ScanIn[28]), .B(n230), .C(In[28]), .D(n228), .Z(n223) );
    VMW_AO22 U88 ( .A(ScanIn[17]), .B(n230), .C(In[17]), .D(n228), .Z(n212) );
    VMW_AO22 U93 ( .A(ScanIn[12]), .B(n230), .C(In[12]), .D(n228), .Z(n207) );
    VMW_AO21 U44 ( .A(\ScanOut[15]1 ), .B(n194), .C(n210), .Z(n247) );
    VMW_AO21 U56 ( .A(\ScanOut[27]1 ), .B(n194), .C(n222), .Z(n235) );
    VMW_AO22 U94 ( .A(ScanIn[11]), .B(n230), .C(In[11]), .D(n228), .Z(n206) );
    VMW_AO22 U71 ( .A(ScanIn[3]), .B(n230), .C(In[3]), .D(n228), .Z(n198) );
    VMW_AND2 U63 ( .A(ScanEnable), .B(n227), .Z(n230) );
    VMW_AO22 U86 ( .A(ScanIn[19]), .B(n230), .C(In[19]), .D(n228), .Z(n214) );
    VMW_AO22 U78 ( .A(ScanIn[26]), .B(n230), .C(In[26]), .D(n228), .Z(n221) );
endmodule


module BubbleSort_Control_CWIDTH2_IDWIDTH1_WIDTH32_SCAN1 ( Clk, Reset, RD, WR, 
    Addr, DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire n330, n317, n345, n339, n357, n322, n325, n350, n319, n342, 
        \count[0] , n359, n356, n337, n318, n351, \ScanReg[15] , \ScanReg[26] , 
        \ScanReg[2] , n324, \ScanReg[18] , n336, n358, n343, \ScanReg[22] , 
        \ScanReg[11] , \ScanReg[6] , \ScanReg[20] , \ScanReg[13] , 
        \ScanReg[4] , n344, \ScanReg[29] , n316, \ScanReg[30] , n331, n323, 
        \ScanReg[17] , \ScanReg[24] , \ScanReg[0] , \ScanReg[9] , n338, n314, 
        n333, \ScanReg[16] , \ScanReg[25] , \ScanReg[8] , n346, \ScanReg[1] , 
        \ScanReg[7] , n328, \ScanReg[5] , n354, \ScanReg[21] , \ScanReg[12] , 
        \ScanReg[28] , \ScanReg[31] , n321, n348, \ScanReg[19] , n326, n353, 
        \ScanReg[10] , \ScanReg[23] , n341, \ScanReg[14] , \ScanReg[27] , n313, 
        \ScanReg[3] , n334, \count[1] , n352, n349, n327, n335, n347, n340, 
        n329, n332, n315, n320, n355;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U54 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U73 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_AND2 U113 ( .A(\ScanReg[19] ), .B(n315), .Z(n325) );
    VMW_BUFIZ U134 ( .A(n327), .E(n330), .Z(\arr[23] ) );
    VMW_AND2 U68 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_AND2 U96 ( .A(\ScanReg[30] ), .B(n315), .Z(n343) );
    VMW_AND2 U108 ( .A(\ScanReg[4] ), .B(n315), .Z(n331) );
    VMW_BUFIZ U141 ( .A(n335), .E(n330), .Z(\arr[16] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AND2 U53 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U61 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_AND2 U84 ( .A(\ScanReg[11] ), .B(n315), .Z(n355) );
    VMW_BUFIZ U148 ( .A(n342), .E(n330), .Z(\arr[13] ) );
    VMW_BUFIZ U153 ( .A(n347), .E(n330), .Z(\arr[24] ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U66 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AND2 U101 ( .A(\ScanReg[31] ), .B(n315), .Z(n338) );
    VMW_AND2 U106 ( .A(\ScanReg[14] ), .B(n315), .Z(n333) );
    VMW_NAND3 U121 ( .A(n316), .B(n320), .C(ScanOut[1]), .Z(n314) );
    VMW_XNOR2 U126 ( .A(Addr[0]), .B(ScanId), .Z(n318) );
    VMW_AND2 U83 ( .A(\ScanReg[8] ), .B(n315), .Z(n357) );
    VMW_FD \count_reg[0]  ( .D(n359), .CP(Clk), .Q(\count[0] ) );
    VMW_AND2 U91 ( .A(\ScanReg[17] ), .B(n315), .Z(n348) );
    VMW_AND2 U98 ( .A(\ScanReg[2] ), .B(n315), .Z(n341) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_INV U128 ( .A(n319), .Z(n324) );
    VMW_BUFIZ U154 ( .A(n348), .E(n330), .Z(\arr[17] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U146 ( .A(n340), .E(n330), .Z(\arr[28] ) );
    VMW_BUFIZ U161 ( .A(n355), .E(n330), .Z(\arr[11] ) );
    VMW_AND2 U74 ( .A(DataIn[9]), .B(WR), .Z(ScanOut[9]) );
    VMW_XNOR2 U114 ( .A(Addr[0]), .B(Id), .Z(n316) );
    VMW_BUFIZ U133 ( .A(n326), .E(n330), .Z(\arr[0] ) );
    VMW_AND2 U99 ( .A(\ScanReg[28] ), .B(n315), .Z(n340) );
    VMW_BUFIZ U155 ( .A(n349), .E(n330), .Z(\arr[7] ) );
    VMW_AND2 U52 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U67 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_NAND2 U82 ( .A(n313), .B(n314), .Z(n358) );
    VMW_AND2 U107 ( .A(\ScanReg[27] ), .B(n315), .Z(n332) );
    VMW_NAND2 U120 ( .A(WR), .B(n316), .Z(n319) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U55 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U69 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U75 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U115 ( .A(WR), .B(DataIn[1]), .Z(ScanOut[1]) );
    VMW_BUFIZ U132 ( .A(n325), .E(n330), .Z(\arr[19] ) );
    VMW_AND2 U90 ( .A(\ScanReg[7] ), .B(n315), .Z(n349) );
    VMW_AND2 U109 ( .A(\ScanReg[9] ), .B(n315), .Z(n329) );
    VMW_INV U129 ( .A(n323), .Z(n359) );
    VMW_BUFIZ U147 ( .A(n341), .E(n330), .Z(\arr[2] ) );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_BUFIZ U160 ( .A(n354), .E(n330), .Z(\arr[22] ) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_AND2 U72 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_AND2 U97 ( .A(\ScanReg[13] ), .B(n315), .Z(n342) );
    VMW_BUFIZ U140 ( .A(n334), .E(n330), .Z(\arr[25] ) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_AO21 U112 ( .A(RD), .B(ScanEnable), .C(n316), .Z(n330) );
    VMW_BUFIZ U135 ( .A(n328), .E(n330), .Z(\arr[10] ) );
    VMW_AND2 U60 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U85 ( .A(\ScanReg[22] ), .B(n315), .Z(n354) );
    VMW_AND2 U100 ( .A(\ScanReg[21] ), .B(n315), .Z(n339) );
    VMW_INV U127 ( .A(\count[0] ), .Z(n322) );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_BUFIZ U149 ( .A(n343), .E(n330), .Z(\arr[30] ) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_BUFIZ U152 ( .A(n346), .E(n330), .Z(\arr[3] ) );
    VMW_OR2 U51 ( .A(\count[0] ), .B(\count[1] ), .Z(Enable) );
    VMW_AND2 U57 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_BUFIZ U137 ( .A(n331), .E(n330), .Z(\arr[4] ) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_AND2 U58 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U59 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_AND2 U62 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_AND2 U70 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AND2 U79 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AND2 U95 ( .A(\ScanReg[29] ), .B(n315), .Z(n344) );
    VMW_AND2 U110 ( .A(\ScanReg[10] ), .B(n315), .Z(n328) );
    VMW_BUFIZ U159 ( .A(n353), .E(n330), .Z(\arr[18] ) );
    VMW_AO22 U119 ( .A(\ScanReg[0] ), .B(n315), .C(\count[0] ), .D(n316), .Z(
        n326) );
    VMW_BUFIZ U142 ( .A(n336), .E(n330), .Z(\arr[12] ) );
    VMW_AND2 U87 ( .A(\ScanReg[15] ), .B(n315), .Z(n352) );
    VMW_BUFIZ U150 ( .A(n344), .E(n330), .Z(\arr[29] ) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_INV U125 ( .A(n316), .Z(n315) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U65 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AND2 U102 ( .A(\ScanReg[6] ), .B(n315), .Z(n337) );
    VMW_AND2 U105 ( .A(\ScanReg[25] ), .B(n315), .Z(n334) );
    VMW_AND2 U80 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_NAND4 U122 ( .A(\count[0] ), .B(\count[1] ), .C(n320), .D(n319), .Z(
        n313) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_BUFIZ U139 ( .A(n333), .E(n330), .Z(\arr[14] ) );
    VMW_BUFIZ U157 ( .A(n351), .E(n330), .Z(\arr[26] ) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AND2 U77 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_AND2 U89 ( .A(\ScanReg[5] ), .B(n315), .Z(n350) );
    VMW_AND2 U92 ( .A(\ScanReg[24] ), .B(n315), .Z(n347) );
    VMW_BUFIZ U145 ( .A(n339), .E(n330), .Z(\arr[21] ) );
    VMW_BUFIZ U162 ( .A(n356), .E(n330), .Z(\arr[1] ) );
    VMW_OAI21 U117 ( .A(RD), .B(WR), .C(n318), .Z(n317) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_INV U130 ( .A(Reset), .Z(n320) );
    VMW_BUFIZ U138 ( .A(n332), .E(n330), .Z(\arr[27] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AND2 U64 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AND2 U81 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_BUFIZ U156 ( .A(n350), .E(n330), .Z(\arr[5] ) );
    VMW_AND2 U104 ( .A(\ScanReg[16] ), .B(n315), .Z(n335) );
    VMW_AND2 U76 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_AND2 U116 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_AO22 U123 ( .A(ScanOut[0]), .B(n316), .C(n319), .D(n322), .Z(n321) );
    VMW_AND2 U56 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U88 ( .A(\ScanReg[26] ), .B(n315), .Z(n351) );
    VMW_AND2 U93 ( .A(\ScanReg[3] ), .B(n315), .Z(n346) );
    VMW_INV U131 ( .A(n317), .Z(ScanEnable) );
    VMW_FD \count_reg[1]  ( .D(n358), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(\ScanReg[20] ), .B(n315), .Z(n345) );
    VMW_BUFIZ U143 ( .A(n337), .E(n330), .Z(\arr[6] ) );
    VMW_BUFIZ U144 ( .A(n338), .E(n330), .Z(\arr[31] ) );
    VMW_BUFIZ U163 ( .A(n357), .E(n330), .Z(\arr[8] ) );
    VMW_BUFIZ U158 ( .A(n352), .E(n330), .Z(\arr[15] ) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_BUFIZ U136 ( .A(n329), .E(n330), .Z(\arr[9] ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AND2 U63 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U71 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_AND2 U111 ( .A(\ScanReg[23] ), .B(n315), .Z(n327) );
    VMW_OAI211 U124 ( .A(Enable), .B(n324), .C(n320), .D(n321), .Z(n323) );
    VMW_AND2 U78 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_AND2 U86 ( .A(\ScanReg[18] ), .B(n315), .Z(n353) );
    VMW_AND2 U103 ( .A(\ScanReg[12] ), .B(n315), .Z(n336) );
    VMW_AO22 U118 ( .A(\ScanReg[1] ), .B(n315), .C(\count[1] ), .D(n316), .Z(
        n356) );
    VMW_BUFIZ U151 ( .A(n345), .E(n330), .Z(\arr[20] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \wRegInA0[9] , \wAIn1[3] , \ScanLink0[13] , \wBIn0[27] , \wBIn0[9] , 
        \wRegInA0[26] , \wRegInA0[15] , \ScanLink4[11] , \ScanLink0[20] , 
        \wRegInB1[8] , \ScanLink4[22] , \wBIn0[14] , \ScanLink1[19] , 
        \wBIn0[0] , \wRegInA1[16] , \ScanLink4[3] , \wRegInA0[0] , \wBIn1[24] , 
        \wRegInB1[1] , \wRegInA1[25] , \wEnable[0] , \ScanLink2[4] , 
        \ScanLink1[10] , \ScanLink1[23] , \ScanLink1[7] , \ScanLink0[30] , 
        \ScanLink0[29] , \wBIn1[17] , \ScanLink4[18] , \wAMid0[4] , 
        \wBIn0[23] , \ScanLink4[7] , \wBIn0[10] , \wRegInA0[22] , 
        \wRegInA0[11] , \wRegInA1[31] , \wRegInA1[28] , \ScanLink2[9] , 
        \ScanLink4[26] , \ScanLink4[15] , \wAMid0[9] , \ScanEnable[0] , 
        \wAIn1[7] , \ScanLink0[17] , \wBIn1[30] , \wBIn1[29] , \ScanLink0[24] , 
        \wRegInA0[18] , \wAMid0[0] , \wBIn1[20] , \wBIn0[19] , \wRegInA0[4] , 
        \wBIn1[13] , \ScanLink2[0] , \ScanLink1[3] , \ScanLink1[27] , 
        \ScanLink1[14] , \wBIn0[31] , \wBIn0[28] , \wBIn0[4] , \wRegInB1[5] , 
        \wRegInA1[21] , \wRegInA1[12] , \ScanLink2[2] , \ScanLink1[16] , 
        \ScanLink1[1] , \wBIn0[6] , \wRegInB1[7] , \ScanLink1[25] , 
        \wRegInA1[10] , \wRegInA0[30] , \wAMid0[2] , \wRegInA1[23] , 
        \wRegInA0[29] , \wRegInA0[6] , \wBIn1[22] , \wRegInA0[20] , 
        \wRegInA0[13] , \wBIn1[11] , \ScanLink4[17] , \ScanLink4[24] , 
        \wAIn1[5] , \wBIn1[18] , \ScanLink0[15] , \ScanLink0[26] , \wBIn0[21] , 
        \ScanLink4[5] , \wBIn0[12] , \wRegInA0[2] , \wAIn1[8] , \wBIn1[26] , 
        \wRegInA1[19] , \ScanLink1[8] , \wBIn1[15] , \ScanLink0[18] , 
        \ScanLink4[30] , \ScanLink4[29] , \wBIn0[25] , \wBIn0[2] , \wAMid0[6] , 
        \wRegInB1[3] , \wRegInA1[27] , \wRegInA1[14] , \ScanLink4[8] , 
        \ScanLink2[6] , \ScanLink1[5] , \ScanLink1[31] , \ScanLink1[28] , 
        \ScanLink1[21] , \ScanLink1[12] , \wBIn0[16] , \wAIn1[1] , 
        \ScanLink4[1] , \ScanLink0[11] , \ScanLink0[22] , \wRegInA0[24] , 
        \wRegInA0[17] , \ScanLink4[20] , \ScanLink4[13] , \wAIn1[25] , 
        \wBMid0[31] , \wBMid0[28] , \wBMid0[5] , \wRegInB0[25] , 
        \wRegInB0[16] , \ScanLink2[24] , \ScanLink2[17] , \wAIn1[16] , 
        \wRegInA1[6] , \ScanLink3[2] , \ScanLink0[1] , \wRegInB0[7] , 
        \wAIn0[26] , \wAMid0[30] , \wAMid0[29] , \wBIn1[6] , \ScanLink0[8] , 
        \wAIn0[15] , \wAMid0[20] , \wAMid0[13] , \wRegInB1[26] , 
        \ScanLink3[27] , \wAIn0[5] , \wBMid0[21] , \wRegInB1[15] , 
        \ScanLink3[14] , \wBMid0[12] , \wBIn1[2] , \wRegInB1[18] , 
        \ScanLink3[19] , \wRegInB0[3] , \wAIn0[18] , \ScanLink3[6] , 
        \ScanLink0[5] , \wAIn0[8] , \wAIn1[21] , \wRegInA1[2] , \wAIn0[1] , 
        \wAIn1[31] , \wAIn1[12] , \wBMid0[1] , \wRegInB0[21] , \ScanLink2[20] , 
        \wRegInB0[12] , \ScanLink2[13] , \wAIn1[28] , \wBMid0[25] , 
        \wBMid0[8] , \ScanLink2[30] , \ScanLink2[29] , \wRegInB0[31] , 
        \wRegInB0[28] , \wBMid0[16] , \wRegInB1[22] , \wRegInB1[11] , 
        \ScanLink3[23] , \ScanLink3[10] , \wAMid0[24] , \wAMid0[17] , 
        \wAIn0[22] , \wAIn0[11] , \wRegInB1[20] , \ScanLink3[21] , 
        \wRegInB0[8] , \wAIn0[20] , \wAMid0[26] , \wBIn1[9] , \wRegInB1[13] , 
        \ScanLink3[12] , \wAMid0[15] , \wAIn0[13] , \wAIn0[3] , \wAIn1[19] , 
        \wRegInA1[9] , \wBMid0[27] , \wRegInB0[19] , \ScanLink2[18] , 
        \wBMid0[14] , \wAIn1[23] , \wAIn1[10] , \wRegInA1[0] , \wBIn1[0] , 
        \wBMid0[3] , \wRegInB0[23] , \wRegInB0[10] , \ScanLink2[22] , 
        \ScanLink2[11] , \wRegInB0[1] , \wAIn0[30] , \wAIn0[29] , 
        \wRegInB1[30] , \wRegInB1[29] , \ScanLink3[31] , \ScanLink3[28] , 
        \ScanLink0[7] , \wAIn0[24] , \wAIn0[7] , \wBMid0[23] , \ScanLink3[4] , 
        \wBMid0[10] , \ScanLink3[9] , \wAIn0[17] , \wAMid0[22] , \wAMid0[11] , 
        \wRegInB1[24] , \wRegInB1[17] , \ScanLink3[25] , \ScanLink3[16] , 
        \ScanLink3[0] , \ScanLink0[3] , \wRegInB0[5] , \wAMid0[18] , 
        \wAIn1[27] , \wBIn1[4] , \wBMid0[19] , \wBMid0[7] , \wRegInB0[27] , 
        \ScanLink2[26] , \wRegInB0[14] , \ScanLink2[15] , \wRegInA1[4] , 
        \wAIn1[14] , \wAIn0[25] , \wAIn0[6] , \wBMid0[22] , \wBMid0[11] , 
        \ScanLink3[8] , \wAIn0[16] , \wRegInB1[25] , \ScanLink3[24] , 
        \ScanLink3[17] , \wAMid0[23] , \wRegInB1[16] , \wAMid0[19] , 
        \wAMid0[10] , \ScanLink3[1] , \ScanLink0[2] , \wBIn1[5] , 
        \wRegInB0[4] , \wBMid0[18] , \wBMid0[6] , \ScanLink2[27] , 
        \wRegInB0[26] , \wRegInB0[15] , \ScanLink2[14] , \wAMid0[27] , 
        \wAIn1[26] , \wAIn1[15] , \wRegInA1[5] , \wAMid0[14] , \wBIn1[8] , 
        \wRegInB1[21] , \ScanLink3[20] , \wRegInB1[12] , \wAIn0[21] , 
        \wRegInB0[9] , \ScanLink3[13] , \wAIn0[12] , \wAIn0[2] , \wAIn1[18] , 
        \wRegInA1[8] , \wAIn1[22] , \wBMid0[26] , \wBMid0[15] , \wRegInB0[18] , 
        \ScanLink2[19] , \wRegInA1[1] , \wAIn1[11] , \wBMid0[2] , 
        \wRegInB0[22] , \wRegInB0[11] , \ScanLink2[23] , \ScanLink2[10] , 
        \wRegInB0[0] , \wRegInB1[31] , \ScanLink3[30] , \ScanLink3[29] , 
        \wRegInB1[28] , \wAIn0[31] , \wBIn1[1] , \wAIn0[28] , \wRegInB0[2] , 
        \ScanLink3[5] , \ScanLink0[6] , \wRegInB1[19] , \ScanLink3[18] , 
        \wAIn0[19] , \wBIn1[3] , \wAIn0[9] , \wAIn1[20] , \ScanLink3[7] , 
        \ScanLink0[4] , \wAIn1[13] , \wRegInA1[3] , \wAIn0[0] , \wAIn1[30] , 
        \wAIn1[29] , \wBMid0[0] , \ScanLink2[21] , \wRegInB0[20] , 
        \wRegInB0[13] , \ScanLink2[12] , \wAMid0[25] , \wBMid0[24] , 
        \wBMid0[17] , \wBMid0[9] , \wRegInB0[30] , \wRegInB0[29] , 
        \ScanLink2[31] , \ScanLink2[28] , \wAMid0[16] , \wRegInB1[23] , 
        \ScanLink3[22] , \ScanLink3[11] , \wAIn0[23] , \wRegInB1[10] , 
        \wAIn0[10] , \wBMid0[30] , \wBMid0[29] , \wBMid0[4] , \wRegInB0[24] , 
        \wRegInB0[17] , \ScanLink2[25] , \ScanLink2[16] , \wAMid0[31] , 
        \wAIn1[24] , \wRegInA1[7] , \wAIn1[17] , \wBIn1[7] , \ScanLink3[3] , 
        \ScanLink0[0] , \wAMid0[28] , \wRegInB0[6] , \wAIn0[27] , \wAIn0[14] , 
        \ScanLink0[9] , \wRegInB1[27] , \ScanLink3[26] , \wRegInB1[14] , 
        \wAIn0[4] , \wAMid0[21] , \ScanLink3[15] , \wAMid0[12] , \wBMid0[20] , 
        \wBMid0[13] , \wRegInA0[3] , \wBIn1[27] , \wAMid0[7] , \wAIn1[9] , 
        \ScanLink0[19] , \wBIn1[14] , \ScanLink4[31] , \ScanLink4[28] , 
        \wBIn0[3] , \wRegInB1[2] , \wRegInA1[26] , \wRegInA1[15] , 
        \ScanLink4[9] , \ScanLink2[7] , \ScanLink1[20] , \ScanLink1[13] , 
        \ScanLink1[4] , \ScanLink4[0] , \wBIn0[24] , \ScanLink1[30] , 
        \ScanLink1[29] , \wBIn0[17] , \wAIn1[0] , \ScanLink0[10] , \wBIn0[30] , 
        \wRegInA0[25] , \wRegInA0[16] , \ScanLink0[23] , \ScanLink4[21] , 
        \ScanLink4[12] , \ScanLink2[3] , \ScanLink1[17] , \ScanLink1[0] , 
        \wBIn0[29] , \wBIn0[7] , \wRegInA1[11] , \ScanLink1[24] , 
        \wRegInA0[31] , \wRegInA0[28] , \wRegInB1[6] , \wRegInA1[22] , 
        \wAMid0[3] , \wBIn1[23] , \wBIn1[10] , \wRegInA0[21] , \wRegInA0[12] , 
        \wRegInA0[7] , \ScanLink4[16] , \wAIn1[4] , \ScanLink4[25] , 
        \wBIn1[19] , \ScanLink0[14] , \ScanLink0[27] , \wBIn0[20] , 
        \wBIn0[13] , \ScanLink1[9] , \ScanLink4[4] , \wBIn0[22] , 
        \wRegInA1[18] , \wBIn0[11] , \ScanLink2[8] , \ScanLink4[6] , 
        \wRegInA0[23] , \wRegInA0[10] , \wAMid0[8] , \wRegInA1[30] , 
        \wRegInA1[29] , \ScanLink4[27] , \ScanLink4[14] , \wAIn1[6] , 
        \ScanLink0[16] , \wRegInA0[19] , \wBIn1[31] , \wBIn1[28] , 
        \ScanLink0[25] , \wAMid0[1] , \wRegInA0[5] , \wBIn1[21] , \wBIn1[12] , 
        \wBIn0[18] , \wBIn0[5] , \ScanLink2[1] , \ScanLink1[26] , 
        \ScanLink1[15] , \ScanLink1[2] , \wAIn1[2] , \wRegInB1[4] , 
        \wRegInA1[20] , \wRegInA1[13] , \ScanLink0[12] , \wRegInA0[8] , 
        \ScanLink0[21] , \wBIn0[8] , \wRegInA0[27] , \wRegInA0[14] , 
        \ScanLink4[10] , \ScanLink4[23] , \wRegInB1[9] , \ScanLink4[2] , 
        \wBIn0[26] , \wBIn0[15] , \ScanLink1[18] , \wBIn0[1] , \wRegInB1[0] , 
        \wRegInA1[17] , \wRegInA0[1] , \wBIn1[25] , \wRegInA1[24] , 
        \ScanLink2[5] , \ScanLink1[11] , \ScanLink1[6] , \ScanLink1[22] , 
        \ScanLink0[31] , \ScanLink0[28] , \wBIn1[16] , \wAMid0[5] , 
        \ScanLink4[19] ;
    BubbleSort_Node_WIDTH32 BSN1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn0[31] , 
        \wAIn0[30] , \wAIn0[29] , \wAIn0[28] , \wAIn0[27] , \wAIn0[26] , 
        \wAIn0[25] , \wAIn0[24] , \wAIn0[23] , \wAIn0[22] , \wAIn0[21] , 
        \wAIn0[20] , \wAIn0[19] , \wAIn0[18] , \wAIn0[17] , \wAIn0[16] , 
        \wAIn0[15] , \wAIn0[14] , \wAIn0[13] , \wAIn0[12] , \wAIn0[11] , 
        \wAIn0[10] , \wAIn0[9] , \wAIn0[8] , \wAIn0[7] , \wAIn0[6] , 
        \wAIn0[5] , \wAIn0[4] , \wAIn0[3] , \wAIn0[2] , \wAIn0[1] , \wAIn0[0] 
        }), .BIn({\wBIn0[31] , \wBIn0[30] , \wBIn0[29] , \wBIn0[28] , 
        \wBIn0[27] , \wBIn0[26] , \wBIn0[25] , \wBIn0[24] , \wBIn0[23] , 
        \wBIn0[22] , \wBIn0[21] , \wBIn0[20] , \wBIn0[19] , \wBIn0[18] , 
        \wBIn0[17] , \wBIn0[16] , \wBIn0[15] , \wBIn0[14] , \wBIn0[13] , 
        \wBIn0[12] , \wBIn0[11] , \wBIn0[10] , \wBIn0[9] , \wBIn0[8] , 
        \wBIn0[7] , \wBIn0[6] , \wBIn0[5] , \wBIn0[4] , \wBIn0[3] , \wBIn0[2] , 
        \wBIn0[1] , \wBIn0[0] }), .HiOut({\wRegInA0[31] , \wRegInA0[30] , 
        \wRegInA0[29] , \wRegInA0[28] , \wRegInA0[27] , \wRegInA0[26] , 
        \wRegInA0[25] , \wRegInA0[24] , \wRegInA0[23] , \wRegInA0[22] , 
        \wRegInA0[21] , \wRegInA0[20] , \wRegInA0[19] , \wRegInA0[18] , 
        \wRegInA0[17] , \wRegInA0[16] , \wRegInA0[15] , \wRegInA0[14] , 
        \wRegInA0[13] , \wRegInA0[12] , \wRegInA0[11] , \wRegInA0[10] , 
        \wRegInA0[9] , \wRegInA0[8] , \wRegInA0[7] , \wRegInA0[6] , 
        \wRegInA0[5] , \wRegInA0[4] , \wRegInA0[3] , \wRegInA0[2] , 
        \wRegInA0[1] , \wRegInA0[0] }), .LoOut({\wAMid0[31] , \wAMid0[30] , 
        \wAMid0[29] , \wAMid0[28] , \wAMid0[27] , \wAMid0[26] , \wAMid0[25] , 
        \wAMid0[24] , \wAMid0[23] , \wAMid0[22] , \wAMid0[21] , \wAMid0[20] , 
        \wAMid0[19] , \wAMid0[18] , \wAMid0[17] , \wAMid0[16] , \wAMid0[15] , 
        \wAMid0[14] , \wAMid0[13] , \wAMid0[12] , \wAMid0[11] , \wAMid0[10] , 
        \wAMid0[9] , \wAMid0[8] , \wAMid0[7] , \wAMid0[6] , \wAMid0[5] , 
        \wAMid0[4] , \wAMid0[3] , \wAMid0[2] , \wAMid0[1] , \wAMid0[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid0[31] , 
        \wAMid0[30] , \wAMid0[29] , \wAMid0[28] , \wAMid0[27] , \wAMid0[26] , 
        \wAMid0[25] , \wAMid0[24] , \wAMid0[23] , \wAMid0[22] , \wAMid0[21] , 
        \wAMid0[20] , \wAMid0[19] , \wAMid0[18] , \wAMid0[17] , \wAMid0[16] , 
        \wAMid0[15] , \wAMid0[14] , \wAMid0[13] , \wAMid0[12] , \wAMid0[11] , 
        \wAMid0[10] , \wAMid0[9] , \wAMid0[8] , \wAMid0[7] , \wAMid0[6] , 
        \wAMid0[5] , \wAMid0[4] , \wAMid0[3] , \wAMid0[2] , \wAMid0[1] , 
        \wAMid0[0] }), .BIn({\wBMid0[31] , \wBMid0[30] , \wBMid0[29] , 
        \wBMid0[28] , \wBMid0[27] , \wBMid0[26] , \wBMid0[25] , \wBMid0[24] , 
        \wBMid0[23] , \wBMid0[22] , \wBMid0[21] , \wBMid0[20] , \wBMid0[19] , 
        \wBMid0[18] , \wBMid0[17] , \wBMid0[16] , \wBMid0[15] , \wBMid0[14] , 
        \wBMid0[13] , \wBMid0[12] , \wBMid0[11] , \wBMid0[10] , \wBMid0[9] , 
        \wBMid0[8] , \wBMid0[7] , \wBMid0[6] , \wBMid0[5] , \wBMid0[4] , 
        \wBMid0[3] , \wBMid0[2] , \wBMid0[1] , \wBMid0[0] }), .HiOut({
        \wRegInB0[31] , \wRegInB0[30] , \wRegInB0[29] , \wRegInB0[28] , 
        \wRegInB0[27] , \wRegInB0[26] , \wRegInB0[25] , \wRegInB0[24] , 
        \wRegInB0[23] , \wRegInB0[22] , \wRegInB0[21] , \wRegInB0[20] , 
        \wRegInB0[19] , \wRegInB0[18] , \wRegInB0[17] , \wRegInB0[16] , 
        \wRegInB0[15] , \wRegInB0[14] , \wRegInB0[13] , \wRegInB0[12] , 
        \wRegInB0[11] , \wRegInB0[10] , \wRegInB0[9] , \wRegInB0[8] , 
        \wRegInB0[7] , \wRegInB0[6] , \wRegInB0[5] , \wRegInB0[4] , 
        \wRegInB0[3] , \wRegInB0[2] , \wRegInB0[1] , \wRegInB0[0] }), .LoOut({
        \wRegInA1[31] , \wRegInA1[30] , \wRegInA1[29] , \wRegInA1[28] , 
        \wRegInA1[27] , \wRegInA1[26] , \wRegInA1[25] , \wRegInA1[24] , 
        \wRegInA1[23] , \wRegInA1[22] , \wRegInA1[21] , \wRegInA1[20] , 
        \wRegInA1[19] , \wRegInA1[18] , \wRegInA1[17] , \wRegInA1[16] , 
        \wRegInA1[15] , \wRegInA1[14] , \wRegInA1[13] , \wRegInA1[12] , 
        \wRegInA1[11] , \wRegInA1[10] , \wRegInA1[9] , \wRegInA1[8] , 
        \wRegInA1[7] , \wRegInA1[6] , \wRegInA1[5] , \wRegInA1[4] , 
        \wRegInA1[3] , \wRegInA1[2] , \wRegInA1[1] , \wRegInA1[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_3 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink4[31] , \ScanLink4[30] , \ScanLink4[29] , 
        \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , \ScanLink4[25] , 
        \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , \ScanLink4[21] , 
        \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , \ScanLink4[17] , 
        \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , \ScanLink4[13] , 
        \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , \ScanLink4[9] , 
        \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , \ScanLink4[5] , 
        \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , \ScanLink4[1] , 
        \ScanLink4[0] }), .ScanOut({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA0[31] , \wRegInA0[30] , 
        \wRegInA0[29] , \wRegInA0[28] , \wRegInA0[27] , \wRegInA0[26] , 
        \wRegInA0[25] , \wRegInA0[24] , \wRegInA0[23] , \wRegInA0[22] , 
        \wRegInA0[21] , \wRegInA0[20] , \wRegInA0[19] , \wRegInA0[18] , 
        \wRegInA0[17] , \wRegInA0[16] , \wRegInA0[15] , \wRegInA0[14] , 
        \wRegInA0[13] , \wRegInA0[12] , \wRegInA0[11] , \wRegInA0[10] , 
        \wRegInA0[9] , \wRegInA0[8] , \wRegInA0[7] , \wRegInA0[6] , 
        \wRegInA0[5] , \wRegInA0[4] , \wRegInA0[3] , \wRegInA0[2] , 
        \wRegInA0[1] , \wRegInA0[0] }), .Out({\wAIn0[31] , \wAIn0[30] , 
        \wAIn0[29] , \wAIn0[28] , \wAIn0[27] , \wAIn0[26] , \wAIn0[25] , 
        \wAIn0[24] , \wAIn0[23] , \wAIn0[22] , \wAIn0[21] , \wAIn0[20] , 
        \wAIn0[19] , \wAIn0[18] , \wAIn0[17] , \wAIn0[16] , \wAIn0[15] , 
        \wAIn0[14] , \wAIn0[13] , \wAIn0[12] , \wAIn0[11] , \wAIn0[10] , 
        \wAIn0[9] , \wAIn0[8] , \wAIn0[7] , \wAIn0[6] , \wAIn0[5] , \wAIn0[4] , 
        \wAIn0[3] , \wAIn0[2] , \wAIn0[1] , \wAIn0[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_2 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink3[31] , \ScanLink3[30] , \ScanLink3[29] , 
        \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , \ScanLink3[25] , 
        \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , \ScanLink3[21] , 
        \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , \ScanLink3[17] , 
        \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , \ScanLink3[13] , 
        \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , \ScanLink3[9] , 
        \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , \ScanLink3[5] , 
        \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , \ScanLink3[1] , 
        \ScanLink3[0] }), .ScanOut({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB0[31] , \wRegInB0[30] , 
        \wRegInB0[29] , \wRegInB0[28] , \wRegInB0[27] , \wRegInB0[26] , 
        \wRegInB0[25] , \wRegInB0[24] , \wRegInB0[23] , \wRegInB0[22] , 
        \wRegInB0[21] , \wRegInB0[20] , \wRegInB0[19] , \wRegInB0[18] , 
        \wRegInB0[17] , \wRegInB0[16] , \wRegInB0[15] , \wRegInB0[14] , 
        \wRegInB0[13] , \wRegInB0[12] , \wRegInB0[11] , \wRegInB0[10] , 
        \wRegInB0[9] , \wRegInB0[8] , \wRegInB0[7] , \wRegInB0[6] , 
        \wRegInB0[5] , \wRegInB0[4] , \wRegInB0[3] , \wRegInB0[2] , 
        \wRegInB0[1] , \wRegInB0[0] }), .Out({\wBIn0[31] , \wBIn0[30] , 
        \wBIn0[29] , \wBIn0[28] , \wBIn0[27] , \wBIn0[26] , \wBIn0[25] , 
        \wBIn0[24] , \wBIn0[23] , \wBIn0[22] , \wBIn0[21] , \wBIn0[20] , 
        \wBIn0[19] , \wBIn0[18] , \wBIn0[17] , \wBIn0[16] , \wBIn0[15] , 
        \wBIn0[14] , \wBIn0[13] , \wBIn0[12] , \wBIn0[11] , \wBIn0[10] , 
        \wBIn0[9] , \wBIn0[8] , \wBIn0[7] , \wBIn0[6] , \wBIn0[5] , \wBIn0[4] , 
        \wBIn0[3] , \wBIn0[2] , \wBIn0[1] , \wBIn0[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_0 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink1[31] , \ScanLink1[30] , \ScanLink1[29] , 
        \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , \ScanLink1[25] , 
        \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , \ScanLink1[21] , 
        \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , \ScanLink1[17] , 
        \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , \ScanLink1[13] , 
        \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , \ScanLink1[9] , 
        \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , \ScanLink1[5] , 
        \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , \ScanLink1[1] , 
        \ScanLink1[0] }), .ScanOut({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB1[31] , \wRegInB1[30] , 
        \wRegInB1[29] , \wRegInB1[28] , \wRegInB1[27] , \wRegInB1[26] , 
        \wRegInB1[25] , \wRegInB1[24] , \wRegInB1[23] , \wRegInB1[22] , 
        \wRegInB1[21] , \wRegInB1[20] , \wRegInB1[19] , \wRegInB1[18] , 
        \wRegInB1[17] , \wRegInB1[16] , \wRegInB1[15] , \wRegInB1[14] , 
        \wRegInB1[13] , \wRegInB1[12] , \wRegInB1[11] , \wRegInB1[10] , 
        \wRegInB1[9] , \wRegInB1[8] , \wRegInB1[7] , \wRegInB1[6] , 
        \wRegInB1[5] , \wRegInB1[4] , \wRegInB1[3] , \wRegInB1[2] , 
        \wRegInB1[1] , \wRegInB1[0] }), .Out({\wBIn1[31] , \wBIn1[30] , 
        \wBIn1[29] , \wBIn1[28] , \wBIn1[27] , \wBIn1[26] , \wBIn1[25] , 
        \wBIn1[24] , \wBIn1[23] , \wBIn1[22] , \wBIn1[21] , \wBIn1[20] , 
        \wBIn1[19] , \wBIn1[18] , \wBIn1[17] , \wBIn1[16] , \wBIn1[15] , 
        \wBIn1[14] , \wBIn1[13] , \wBIn1[12] , \wBIn1[11] , \wBIn1[10] , 
        \wBIn1[9] , \wBIn1[8] , \wBIn1[7] , \wBIn1[6] , \wBIn1[5] , \wBIn1[4] , 
        \wBIn1[3] , \wBIn1[2] , \wBIn1[1] , \wBIn1[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn1[31] , 
        \wAIn1[30] , \wAIn1[29] , \wAIn1[28] , \wAIn1[27] , \wAIn1[26] , 
        \wAIn1[25] , \wAIn1[24] , \wAIn1[23] , \wAIn1[22] , \wAIn1[21] , 
        \wAIn1[20] , \wAIn1[19] , \wAIn1[18] , \wAIn1[17] , \wAIn1[16] , 
        \wAIn1[15] , \wAIn1[14] , \wAIn1[13] , \wAIn1[12] , \wAIn1[11] , 
        \wAIn1[10] , \wAIn1[9] , \wAIn1[8] , \wAIn1[7] , \wAIn1[6] , 
        \wAIn1[5] , \wAIn1[4] , \wAIn1[3] , \wAIn1[2] , \wAIn1[1] , \wAIn1[0] 
        }), .BIn({\wBIn1[31] , \wBIn1[30] , \wBIn1[29] , \wBIn1[28] , 
        \wBIn1[27] , \wBIn1[26] , \wBIn1[25] , \wBIn1[24] , \wBIn1[23] , 
        \wBIn1[22] , \wBIn1[21] , \wBIn1[20] , \wBIn1[19] , \wBIn1[18] , 
        \wBIn1[17] , \wBIn1[16] , \wBIn1[15] , \wBIn1[14] , \wBIn1[13] , 
        \wBIn1[12] , \wBIn1[11] , \wBIn1[10] , \wBIn1[9] , \wBIn1[8] , 
        \wBIn1[7] , \wBIn1[6] , \wBIn1[5] , \wBIn1[4] , \wBIn1[3] , \wBIn1[2] , 
        \wBIn1[1] , \wBIn1[0] }), .HiOut({\wBMid0[31] , \wBMid0[30] , 
        \wBMid0[29] , \wBMid0[28] , \wBMid0[27] , \wBMid0[26] , \wBMid0[25] , 
        \wBMid0[24] , \wBMid0[23] , \wBMid0[22] , \wBMid0[21] , \wBMid0[20] , 
        \wBMid0[19] , \wBMid0[18] , \wBMid0[17] , \wBMid0[16] , \wBMid0[15] , 
        \wBMid0[14] , \wBMid0[13] , \wBMid0[12] , \wBMid0[11] , \wBMid0[10] , 
        \wBMid0[9] , \wBMid0[8] , \wBMid0[7] , \wBMid0[6] , \wBMid0[5] , 
        \wBMid0[4] , \wBMid0[3] , \wBMid0[2] , \wBMid0[1] , \wBMid0[0] }), 
        .LoOut({\wRegInB1[31] , \wRegInB1[30] , \wRegInB1[29] , \wRegInB1[28] , 
        \wRegInB1[27] , \wRegInB1[26] , \wRegInB1[25] , \wRegInB1[24] , 
        \wRegInB1[23] , \wRegInB1[22] , \wRegInB1[21] , \wRegInB1[20] , 
        \wRegInB1[19] , \wRegInB1[18] , \wRegInB1[17] , \wRegInB1[16] , 
        \wRegInB1[15] , \wRegInB1[14] , \wRegInB1[13] , \wRegInB1[12] , 
        \wRegInB1[11] , \wRegInB1[10] , \wRegInB1[9] , \wRegInB1[8] , 
        \wRegInB1[7] , \wRegInB1[6] , \wRegInB1[5] , \wRegInB1[4] , 
        \wRegInB1[3] , \wRegInB1[2] , \wRegInB1[1] , \wRegInB1[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_1 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink2[31] , \ScanLink2[30] , \ScanLink2[29] , 
        \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , \ScanLink2[25] , 
        \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , \ScanLink2[21] , 
        \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , \ScanLink2[17] , 
        \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , \ScanLink2[13] , 
        \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , \ScanLink2[9] , 
        \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , \ScanLink2[5] , 
        \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , \ScanLink2[1] , 
        \ScanLink2[0] }), .ScanOut({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA1[31] , \wRegInA1[30] , 
        \wRegInA1[29] , \wRegInA1[28] , \wRegInA1[27] , \wRegInA1[26] , 
        \wRegInA1[25] , \wRegInA1[24] , \wRegInA1[23] , \wRegInA1[22] , 
        \wRegInA1[21] , \wRegInA1[20] , \wRegInA1[19] , \wRegInA1[18] , 
        \wRegInA1[17] , \wRegInA1[16] , \wRegInA1[15] , \wRegInA1[14] , 
        \wRegInA1[13] , \wRegInA1[12] , \wRegInA1[11] , \wRegInA1[10] , 
        \wRegInA1[9] , \wRegInA1[8] , \wRegInA1[7] , \wRegInA1[6] , 
        \wRegInA1[5] , \wRegInA1[4] , \wRegInA1[3] , \wRegInA1[2] , 
        \wRegInA1[1] , \wRegInA1[0] }), .Out({\wAIn1[31] , \wAIn1[30] , 
        \wAIn1[29] , \wAIn1[28] , \wAIn1[27] , \wAIn1[26] , \wAIn1[25] , 
        \wAIn1[24] , \wAIn1[23] , \wAIn1[22] , \wAIn1[21] , \wAIn1[20] , 
        \wAIn1[19] , \wAIn1[18] , \wAIn1[17] , \wAIn1[16] , \wAIn1[15] , 
        \wAIn1[14] , \wAIn1[13] , \wAIn1[12] , \wAIn1[11] , \wAIn1[10] , 
        \wAIn1[9] , \wAIn1[8] , \wAIn1[7] , \wAIn1[6] , \wAIn1[5] , \wAIn1[4] , 
        \wAIn1[3] , \wAIn1[2] , \wAIn1[1] , \wAIn1[0] }) );
    BubbleSort_Control_CWIDTH2_IDWIDTH1_WIDTH32_SCAN1 U_BSC ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanOut({\ScanLink4[31] , 
        \ScanLink4[30] , \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , 
        \ScanLink4[26] , \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , 
        \ScanLink4[22] , \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , 
        \ScanLink4[18] , \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , 
        \ScanLink4[14] , \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , 
        \ScanLink4[10] , \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , 
        \ScanLink4[6] , \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , 
        \ScanLink4[2] , \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(
        \ScanEnable[0] ), .ScanId(1'b0), .Id(1'b1), .Enable(\wEnable[0] ) );
endmodule

