
module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_15 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15;
    VMW_AOI21 U3 ( .A(A[3]), .B(n15), .C(A[4]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[2]), .B(A[1]), .C(A[0]), .Z(n15) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_14 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR3 U3 ( .A(A[2]), .B(A[4]), .C(A[3]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_13 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n16;
    VMW_NOR2 U3 ( .A(A[4]), .B(n16), .Z(LT_LE) );
    VMW_AND3 U4 ( .A(A[3]), .B(A[2]), .C(A[1]), .Z(n16) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_12 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n17;
    VMW_NOR3 U3 ( .A(n17), .B(A[4]), .C(A[3]), .Z(LT_LE) );
    VMW_AND3 U4 ( .A(A[1]), .B(A[2]), .C(A[0]), .Z(n17) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_11 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n18, n19;
    VMW_NOR2 U3 ( .A(n18), .B(A[4]), .Z(LT_LE) );
    VMW_INV U5 ( .A(n19), .Z(n18) );
    VMW_OAI211 U4 ( .A(A[1]), .B(A[0]), .C(A[2]), .D(A[3]), .Z(n19) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_10 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR2 U3 ( .A(A[4]), .B(A[3]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_9 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n20;
    VMW_NOR3 U3 ( .A(n20), .B(A[4]), .C(A[3]), .Z(LT_LE) );
    VMW_AO21 U4 ( .A(A[0]), .B(A[1]), .C(A[2]), .Z(n20) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_7 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n21;
    VMW_AOI21 U3 ( .A(A[3]), .B(n21), .C(A[4]), .Z(LT_LE) );
    VMW_AO21 U4 ( .A(A[0]), .B(A[1]), .C(A[2]), .Z(n21) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_6 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n22;
    VMW_AOI211 U3 ( .A(A[2]), .B(n22), .C(A[3]), .D(A[4]), .Z(LT_LE) );
    VMW_OR2 U4 ( .A(A[1]), .B(A[0]), .Z(n22) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_5 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n23;
    VMW_AOI21 U3 ( .A(A[3]), .B(n23), .C(A[4]), .Z(LT_LE) );
    VMW_OR2 U4 ( .A(A[2]), .B(A[1]), .Z(n23) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_4 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_AOI21 U3 ( .A(A[2]), .B(A[3]), .C(A[4]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_3 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR4 U3 ( .A(A[4]), .B(A[3]), .C(A[2]), .D(A[1]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_2 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n24;
    VMW_NOR2 U3 ( .A(A[4]), .B(n24), .Z(LT_LE) );
    VMW_AND4 U4 ( .A(A[0]), .B(A[3]), .C(A[1]), .D(A[2]), .Z(n24) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_1 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_AOI211 U3 ( .A(A[1]), .B(A[2]), .C(A[4]), .D(A[3]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_0 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [4:0] A;
input  [4:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR5 U3 ( .A(A[1]), .B(A[0]), .C(A[2]), .D(A[4]), .E(A[3]), .Z(LT_LE)
         );
endmodule


module NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, CallIn, ReturnIn, ColIn, PDiagIn, 
    NDiagIn, CallOut, ReturnOut, ColOut, PDiagOut, NDiagOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [4:0] Id;
input  [15:0] ColIn;
output [15:0] ColOut;
input  [4:0] ScanIn;
output [4:0] ScanOut;
input  [15:0] NDiagIn;
output [15:0] PDiagOut;
output [15:0] NDiagOut;
input  [15:0] PDiagIn;
input  Clk, Reset, RD, WR, ScanEnable, CallIn, ReturnIn;
output CallOut, ReturnOut;
    wire \NDiagOut[0] , n2010, n2037, n1996, n2059, n2065, n468, n2042, n2137, 
        n2080, n2110, n596, n2125, n2019, Logic11, \n768[3] , ReturnOut723, 
        n2092, n2102, n2077, n2050, n2002, n2089, n484, n2119, n2005, n2025, 
        n2022, n1998, \n768[1] , n2057, n2070, n2039, n2095, n2105, n2122, 
        n2087, n2117, n2130, n2045, n2062, n1991, n2079, n548, n2030, n2104, 
        n2017, n2038, n2094, n1999, n2123, n2056, n2071, n2138, n1990, n2004, 
        n2023, n388, n2031, n2016, n500, n2044, n2078, n452, n2063, n2131, 
        n2086, n2116, n2136, n2043, n2064, n2081, n420, n2111, n1997, n2011, 
        n2058, n2036, n2088, n2118, n1985, n2003, n532, n2024, n2051, n2076, 
        n2124, n2018, n2093, n2103, n2098, n612, n2108, n2126, n2134, n1995, 
        n2013, n2034, n2041, n2008, n2066, n2083, n2113, n2091, n2101, n2053, 
        n2074, n1987, n2001, n2048, n2026, n2006, n2021, n2054, n2068, n2073, 
        n2128, n2133, n2028, n2121, n2096, n2106, n580, n1989, n2084, n2114, 
        n1992, n2061, n2046, n2014, n2033, n2120, n2097, n2107, n436, n2055, 
        n2072, n564, n2007, n2069, n2020, n2129, \n768[4] , CallOut730, n2015, 
        n2032, n1993, n1988, \n768[0] , n2060, n2029, n2047, n2132, n2009, 
        n2085, n404, n2115, n2135, n2082, n2112, \n768[2] , n2040, n2067, 
        n1994, n2000, n2012, n2035, n2099, n2109, n2027, n1986, n516, n2049, 
        n2052, n2075, n2127, n2090, n2100;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 ;
    assign PDiagOut[15] = \NDiagOut[0] ;
    assign NDiagOut[0] = \NDiagOut[0] ;
    VMW_PULLDOWN U460 ( .Z(n2125) );
    VMW_OR3 U529 ( .A(n2024), .B(n2025), .C(n2026), .Z(n2123) );
    VMW_OR2 U585 ( .A(n2086), .B(n2085), .Z(n1994) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_7 gt_104_4 ( .A({\n768[4] , 
        \n768[3] , \n768[2] , \n768[1] , \n768[0] }), .B({\NDiagOut[0] , 
        Logic11, \NDiagOut[0] , Logic11, Logic11}), .LEQ(n2131), .TC(n2131), 
        .LT_LE(n452) );
    VMW_AND2 U547 ( .A(n2064), .B(n2062), .Z(n2053) );
    VMW_NAND2 U560 ( .A(ScanOut[1]), .B(ScanOut[2]), .Z(n2086) );
    VMW_NAND4 U619 ( .A(n2111), .B(n2016), .C(n2006), .D(n1993), .Z(n2060) );
    VMW_INV U650 ( .A(CallIn), .Z(n2073) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_6 gt_104_10 ( .A({
        \n768[4] , \n768[3] , \n768[2] , \n768[1] , \n768[0] }), .B({
        \NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11}), .LEQ(
        n2130), .TC(n2130), .LT_LE(n548) );
    VMW_NAND2 U485 ( .A(n1995), .B(n1996), .Z(ColOut[6]) );
    VMW_OR2 U515 ( .A(NDiagIn[11]), .B(n1989), .Z(NDiagOut[12]) );
    VMW_OR3 U532 ( .A(n2024), .B(n2031), .C(n2032), .Z(n2120) );
    VMW_OR4 U602 ( .A(n2102), .B(NDiagIn[10]), .C(PDiagIn[10]), .D(ColIn[10]), 
        .Z(n2069) );
    VMW_OAI211 U625 ( .A(n2098), .B(n2097), .C(n2068), .D(n2069), .Z(n2036) );
    VMW_PULLDOWN U467 ( .Z(n2132) );
    VMW_PULLDOWN U469 ( .Z(n2134) );
    VMW_PULLDOWN U472 ( .Z(n2137) );
    VMW_OR2 U497 ( .A(PDiagIn[10]), .B(n1990), .Z(PDiagOut[9]) );
    VMW_OR2 U507 ( .A(CallIn), .B(n2011), .Z(\n768[4] ) );
    VMW_NAND2 U520 ( .A(n1996), .B(n2017), .Z(NDiagOut[7]) );
    VMW_NAND4 U610 ( .A(n2106), .B(n2018), .C(n2008), .D(n1997), .Z(n2042) );
    VMW_INV U637 ( .A(PDiagIn[5]), .Z(n2008) );
    VMW_MUX2I U569 ( .A(n2082), .B(n2095), .S(ScanEnable), .Z(n2014) );
    VMW_INV U659 ( .A(n2052), .Z(n2054) );
    VMW_PULLDOWN U475 ( .Z(\NDiagOut[0] ) );
    VMW_NOR2 U549 ( .A(n2049), .B(n2056), .Z(n2052) );
    VMW_AO21 U552 ( .A(n2072), .B(n2073), .C(Reset), .Z(n2023) );
    VMW_NAND2 U555 ( .A(ScanOut[1]), .B(n2079), .Z(n2078) );
    VMW_OAI22 U572 ( .A(n2084), .B(n2090), .C(n2092), .D(n2089), .Z(n2051) );
    VMW_INV U642 ( .A(ScanOut[2]), .Z(n2079) );
    VMW_NOR2 U590 ( .A(n2078), .B(n2087), .Z(n2002) );
    VMW_NOR2 U597 ( .A(CallIn), .B(n420), .Z(n2100) );
    VMW_INV U665 ( .A(n2045), .Z(n2058) );
    VMW_INV U662 ( .A(n2101), .Z(n2097) );
    VMW_AO21 U575 ( .A(n2059), .B(n2062), .C(n2047), .Z(n2037) );
    VMW_INV U645 ( .A(NDiagIn[7]), .Z(n2016) );
    VMW_OR2 U482 ( .A(n1991), .B(ColIn[9]), .Z(ColOut[9]) );
    VMW_NAND2 U490 ( .A(n2003), .B(n2004), .Z(ColOut[1]) );
    VMW_AND2 U527 ( .A(n2021), .B(n2022), .Z(ReturnOut723) );
    VMW_AND4 U617 ( .A(n2109), .B(n2017), .C(n2007), .D(n1995), .Z(n2110) );
    VMW_INV U630 ( .A(ColIn[7]), .Z(n1993) );
    VMW_NAND2 U500 ( .A(n1994), .B(n2006), .Z(PDiagOut[6]) );
    VMW_OR2 U512 ( .A(NDiagIn[14]), .B(n1986), .Z(NDiagOut[15]) );
    VMW_NOR4 U535 ( .A(n2040), .B(NDiagIn[14]), .C(PDiagIn[14]), .D(ColIn[14]), 
        .Z(n2039) );
    VMW_NOR2 U605 ( .A(CallIn), .B(n484), .Z(n2104) );
    VMW_NOR4 U622 ( .A(PDiagIn[0]), .B(n2073), .C(ColIn[0]), .D(NDiagIn[0]), 
        .Z(n2056) );
    VMW_NOR2 U599 ( .A(CallIn), .B(n404), .Z(n2040) );
    VMW_PULLUP U474 ( .Z(Logic11) );
    VMW_OR2 U491 ( .A(ColIn[0]), .B(n2005), .Z(ColOut[0]) );
    VMW_OR2 U499 ( .A(PDiagIn[8]), .B(n1992), .Z(PDiagOut[7]) );
    VMW_OR2 U509 ( .A(CallIn), .B(n2013), .Z(\n768[2] ) );
    VMW_NOR3 U540 ( .A(n2054), .B(n2055), .C(n2023), .Z(n2029) );
    VMW_MUX2I U567 ( .A(n2075), .B(n2093), .S(ScanEnable), .Z(n2012) );
    VMW_NOR2 U582 ( .A(n2076), .B(n2078), .Z(n1990) );
    VMW_INV U657 ( .A(n2044), .Z(n2063) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_4 gt_104_3 ( .A({\n768[4] , 
        \n768[3] , \n768[2] , UNCONNECTED_1, UNCONNECTED_2}), .B({
        \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , \NDiagOut[0] }), .LEQ(
        n2128), .TC(n2128), .LT_LE(n436) );
    VMW_NAND2 U501 ( .A(n1996), .B(n2007), .Z(PDiagOut[5]) );
    VMW_OR2 U526 ( .A(NDiagIn[0]), .B(n2005), .Z(NDiagOut[1]) );
    VMW_INV U639 ( .A(PDiagIn[1]), .Z(n2010) );
    VMW_OR2 U616 ( .A(CallIn), .B(n532), .Z(n2109) );
    VMW_INV U631 ( .A(ColIn[6]), .Z(n1995) );
    VMW_AND3 U548 ( .A(n2065), .B(n2066), .C(n2053), .Z(n2035) );
    VMW_PULLDOWN U461 ( .Z(n2126) );
    VMW_PULLDOWN U466 ( .Z(n2131) );
    VMW_OR2 U498 ( .A(PDiagIn[9]), .B(n1991), .Z(PDiagOut[8]) );
    VMW_NOR2 U553 ( .A(ScanOut[4]), .B(n2075), .Z(n2074) );
    VMW_INV U663 ( .A(n2069), .Z(n2116) );
    VMW_OAI22 U574 ( .A(n2079), .B(n2090), .C(n2094), .D(n2089), .Z(n2030) );
    VMW_NOR2 U583 ( .A(n2080), .B(n2081), .Z(n1991) );
    VMW_OR2 U591 ( .A(n2085), .B(n2081), .Z(n2004) );
    VMW_INV U644 ( .A(ScanOut[0]), .Z(n2077) );
    VMW_FD CallOut_reg ( .D(CallOut730), .CP(Clk), .Q(CallOut) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_11 gt_104_2 ( .A({
        \n768[4] , \n768[3] , \n768[2] , \n768[1] , \n768[0] }), .B({
        \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , Logic11}), .LEQ(n2134), 
        .TC(n2134), .LT_LE(n420) );
    VMW_OR2 U508 ( .A(CallIn), .B(n2012), .Z(\n768[3] ) );
    VMW_NOR3 U541 ( .A(n2023), .B(n2034), .C(n2054), .Z(n2027) );
    VMW_INV U638 ( .A(PDiagIn[3]), .Z(n2009) );
    VMW_MUX2I U566 ( .A(n2084), .B(n2092), .S(ScanEnable), .Z(n2011) );
    VMW_INV U656 ( .A(ReturnIn), .Z(n2072) );
    VMW_OR2 U483 ( .A(n1992), .B(ColIn[8]), .Z(ColOut[8]) );
    VMW_AOI211 U534 ( .A(n2035), .B(n2036), .C(n2037), .D(n2038), .Z(n2034) );
    VMW_FD \MyColumn_reg[1]  ( .D(n2122), .CP(Clk), .Q(ScanOut[1]) );
    VMW_OR4 U604 ( .A(n2103), .B(NDiagIn[11]), .C(PDiagIn[11]), .D(ColIn[11]), 
        .Z(n2068) );
    VMW_NOR2 U623 ( .A(n2044), .B(n2057), .Z(n2113) );
    VMW_NAND2 U484 ( .A(n1993), .B(n1994), .Z(ColOut[7]) );
    VMW_OR2 U513 ( .A(NDiagIn[13]), .B(n1987), .Z(NDiagOut[14]) );
    VMW_OR2 U514 ( .A(NDiagIn[12]), .B(n1988), .Z(NDiagOut[13]) );
    VMW_OR4 U598 ( .A(n2100), .B(NDiagIn[13]), .C(PDiagIn[13]), .D(ColIn[13]), 
        .Z(n2101) );
    VMW_NOR2 U533 ( .A(CallIn), .B(n388), .Z(n2033) );
    VMW_NOR2 U603 ( .A(CallIn), .B(n452), .Z(n2103) );
    VMW_AOI211 U624 ( .A(n2059), .B(n2062), .C(n2113), .D(n2067), .Z(n2055) );
    VMW_PULLDOWN U468 ( .Z(n2133) );
    VMW_NOR2 U528 ( .A(n2023), .B(n2021), .Z(CallOut730) );
    VMW_AND2 U546 ( .A(n2057), .B(n2063), .Z(n2062) );
    VMW_OR2 U561 ( .A(ScanOut[0]), .B(n2083), .Z(n2087) );
    VMW_INV U651 ( .A(ScanIn[4]), .Z(n2092) );
    VMW_FD \MyColumn_reg[3]  ( .D(n2120), .CP(Clk), .Q(ScanOut[3]) );
    VMW_NOR2 U584 ( .A(n2076), .B(n2081), .Z(n1992) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_5 gt_104_5 ( .A({\n768[4] , 
        \n768[3] , \n768[2] , \n768[1] , UNCONNECTED_3}), .B({\NDiagOut[0] , 
        Logic11, \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n2129), .TC(
        n2129), .LT_LE(n468) );
    VMW_NOR4 U596 ( .A(n2099), .B(NDiagIn[12]), .C(PDiagIn[12]), .D(ColIn[12]), 
        .Z(n2098) );
    VMW_OR2 U618 ( .A(CallIn), .B(n516), .Z(n2111) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_14 gt_104_11 ( .A({
        \n768[4] , \n768[3] , \n768[2] , UNCONNECTED_4, UNCONNECTED_5}), .B({
        \NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] }), 
        .LEQ(n2137), .TC(n2137), .LT_LE(n564) );
    VMW_PULLDOWN U473 ( .Z(n2138) );
    VMW_NAND2 U554 ( .A(n2074), .B(n2077), .Z(n2076) );
    VMW_OAI22 U573 ( .A(n2075), .B(n2090), .C(n2093), .D(n2089), .Z(n2032) );
    VMW_INV U643 ( .A(ScanOut[1]), .Z(n2082) );
    VMW_MUX2I U568 ( .A(n2079), .B(n2094), .S(ScanEnable), .Z(n2013) );
    VMW_INV U664 ( .A(n2065), .Z(n2118) );
    VMW_INV U658 ( .A(n2059), .Z(n2064) );
    VMW_PULLDOWN U459 ( .Z(n2124) );
    VMW_PULLDOWN U463 ( .Z(n2128) );
    VMW_OR2 U478 ( .A(n1987), .B(ColIn[13]), .Z(ColOut[13]) );
    VMW_OR2 U496 ( .A(PDiagIn[11]), .B(n1989), .Z(PDiagOut[10]) );
    VMW_NAND2 U506 ( .A(n2004), .B(n2010), .Z(PDiagOut[0]) );
    VMW_NAND2 U521 ( .A(n1998), .B(n2018), .Z(NDiagOut[6]) );
    VMW_NOR2 U611 ( .A(CallIn), .B(n564), .Z(n2107) );
    VMW_INV U636 ( .A(PDiagIn[6]), .Z(n2007) );
    VMW_OR2 U586 ( .A(n2087), .B(n2086), .Z(n1996) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_3 gt_104_13 ( .A({
        \n768[4] , \n768[3] , \n768[2] , \n768[1] , UNCONNECTED_6}), .B({
        \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] }), 
        .LEQ(n2127), .TC(n2127), .LT_LE(n596) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_10 gt_104_7 ( .A({
        \n768[4] , \n768[3] , UNCONNECTED_7, UNCONNECTED_8, UNCONNECTED_9}), 
        .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] }), .LEQ(n2133), .TC(n2133), .LT_LE(n500) );
    VMW_OR2 U544 ( .A(n2047), .B(n2038), .Z(n2044) );
    VMW_NAND2 U563 ( .A(n2090), .B(n2023), .Z(n2089) );
    VMW_INV U653 ( .A(ScanIn[2]), .Z(n2094) );
    VMW_NOR2 U578 ( .A(n2076), .B(n2086), .Z(n1986) );
    VMW_INV U648 ( .A(NDiagIn[3]), .Z(n2019) );
    VMW_PULLDOWN U464 ( .Z(n2129) );
    VMW_PULLDOWN U471 ( .Z(n2136) );
    VMW_NAND2 U486 ( .A(n1997), .B(n1998), .Z(ColOut[5]) );
    VMW_OR2 U516 ( .A(NDiagIn[10]), .B(n1990), .Z(NDiagOut[11]) );
    VMW_OR3 U531 ( .A(n2024), .B(n2029), .C(n2030), .Z(n2121) );
    VMW_NOR2 U601 ( .A(CallIn), .B(n468), .Z(n2102) );
    VMW_OR2 U494 ( .A(PDiagIn[13]), .B(n1987), .Z(PDiagOut[12]) );
    VMW_NAND2 U523 ( .A(n2001), .B(n2019), .Z(NDiagOut[4]) );
    VMW_OR2 U613 ( .A(CallIn), .B(n580), .Z(n2091) );
    VMW_AO21 U626 ( .A(n2039), .B(n2101), .C(n2098), .Z(n2114) );
    VMW_NAND2 U504 ( .A(n2001), .B(n2009), .Z(PDiagOut[2]) );
    VMW_INV U634 ( .A(ColIn[1]), .Z(n2003) );
    VMW_OR2 U476 ( .A(n1985), .B(ColIn[15]), .Z(ColOut[15]) );
    VMW_NAND2 U488 ( .A(n2000), .B(n2001), .Z(ColOut[3]) );
    VMW_OR2 U518 ( .A(NDiagIn[8]), .B(n1992), .Z(NDiagOut[9]) );
    VMW_AOI211 U538 ( .A(n2022), .B(n2021), .C(n2051), .D(n2024), .Z(n2050) );
    VMW_NAND2 U556 ( .A(n2074), .B(ScanOut[0]), .Z(n2080) );
    VMW_FD \MyColumn_reg[2]  ( .D(n2121), .CP(Clk), .Q(ScanOut[2]) );
    VMW_NOR3 U571 ( .A(n2097), .B(n2098), .C(n2039), .Z(n2071) );
    VMW_INV U641 ( .A(ScanOut[3]), .Z(n2075) );
    VMW_INV U666 ( .A(n2048), .Z(n2038) );
    VMW_NOR2 U594 ( .A(n2087), .B(n2081), .Z(n2005) );
    VMW_NOR2 U593 ( .A(n2080), .B(n2086), .Z(n1985) );
    VMW_OR4 U608 ( .A(n2105), .B(NDiagIn[8]), .C(PDiagIn[8]), .D(ColIn[8]), 
        .Z(n2065) );
    VMW_AND4 U551 ( .A(n2052), .B(n2070), .C(n2067), .D(n2071), .Z(n2021) );
    VMW_OAI22 U576 ( .A(n2082), .B(n2090), .C(n2095), .D(n2089), .Z(n2028) );
    VMW_AO21 U628 ( .A(n2066), .B(n2115), .C(n2118), .Z(n2117) );
    VMW_INV U646 ( .A(NDiagIn[6]), .Z(n2017) );
    VMW_INV U661 ( .A(n2023), .Z(n2022) );
    VMW_OR2 U481 ( .A(n1990), .B(ColIn[10]), .Z(ColOut[10]) );
    VMW_OR2 U493 ( .A(PDiagIn[14]), .B(n1986), .Z(PDiagOut[13]) );
    VMW_OR2 U503 ( .A(PDiagIn[4]), .B(n1999), .Z(PDiagOut[3]) );
    VMW_INV U633 ( .A(ColIn[3]), .Z(n2000) );
    VMW_FD \MyColumn_reg[0]  ( .D(n2123), .CP(Clk), .Q(ScanOut[0]) );
    VMW_OR2 U524 ( .A(NDiagIn[2]), .B(n2002), .Z(NDiagOut[3]) );
    VMW_NOR2 U588 ( .A(n2087), .B(n2088), .Z(n1999) );
    VMW_NOR2 U614 ( .A(CallIn), .B(n596), .Z(n2108) );
    VMW_AND4 U621 ( .A(n2112), .B(n2020), .C(n2010), .D(n2003), .Z(n2049) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_1 gt_104_9 ( .A({\n768[4] , 
        \n768[3] , \n768[2] , \n768[1] , UNCONNECTED_10}), .B({\NDiagOut[0] , 
        \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] }), .LEQ(n2125), .TC(
        n2125), .LT_LE(n532) );
    VMW_OR2 U511 ( .A(CallIn), .B(n2015), .Z(\n768[0] ) );
    VMW_AOI211 U536 ( .A(n2042), .B(n2043), .C(n2044), .D(n2045), .Z(n2041) );
    VMW_NAND2 U558 ( .A(n2084), .B(n2075), .Z(n2083) );
    VMW_OR4 U606 ( .A(n2104), .B(NDiagIn[9]), .C(PDiagIn[9]), .D(ColIn[9]), 
        .Z(n2066) );
    VMW_OR2 U477 ( .A(n1986), .B(ColIn[14]), .Z(ColOut[14]) );
    VMW_OR2 U492 ( .A(n1985), .B(PDiagIn[15]), .Z(PDiagOut[14]) );
    VMW_AND2 U543 ( .A(n2042), .B(n2058), .Z(n2057) );
    VMW_OR3 U564 ( .A(CallIn), .B(ScanEnable), .C(n2022), .Z(n2090) );
    VMW_INV U654 ( .A(ScanIn[1]), .Z(n2095) );
    VMW_NOR2 U581 ( .A(n2078), .B(n2080), .Z(n1989) );
    VMW_FD \MyColumn_reg[4]  ( .D(n2119), .CP(Clk), .Q(ScanOut[4]) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_0 gt_104_14 ( .A({
        \n768[4] , \n768[3] , \n768[2] , \n768[1] , \n768[0] }), .B({
        \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11}), 
        .LEQ(n2124), .TC(n2124), .LT_LE(n612) );
    VMW_INV U632 ( .A(ColIn[5]), .Z(n1997) );
    VMW_NAND2 U502 ( .A(n1998), .B(n2008), .Z(PDiagOut[4]) );
    VMW_NAND2 U525 ( .A(n2004), .B(n2020), .Z(NDiagOut[2]) );
    VMW_OR2 U589 ( .A(n2078), .B(n2085), .Z(n2001) );
    VMW_OR4 U615 ( .A(n2108), .B(NDiagIn[2]), .C(PDiagIn[2]), .D(ColIn[2]), 
        .Z(n2048) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_12 gt_104_8 ( .A({
        \n768[4] , \n768[3] , \n768[2] , \n768[1] , \n768[0] }), .B({
        \NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, Logic11}), .LEQ(n2135), 
        .TC(n2135), .LT_LE(n516) );
    VMW_OR2 U489 ( .A(n2002), .B(ColIn[2]), .Z(ColOut[2]) );
    VMW_AND3 U550 ( .A(n2068), .B(n2069), .C(n2035), .Z(n2067) );
    VMW_OAI22 U577 ( .A(n2077), .B(n2090), .C(n2096), .D(n2089), .Z(n2026) );
    VMW_INV U647 ( .A(NDiagIn[5]), .Z(n2018) );
    VMW_INV U660 ( .A(n2050), .Z(n2119) );
    VMW_NOR2 U592 ( .A(n2089), .B(n2073), .Z(n2024) );
    VMW_NAND2 U519 ( .A(n1994), .B(n2016), .Z(NDiagOut[8]) );
    VMW_NOR2 U580 ( .A(n2076), .B(n2088), .Z(n1988) );
    VMW_AO21 U629 ( .A(n2060), .B(n2117), .C(n2110), .Z(n2043) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_13 gt_104_1 ( .A({
        \n768[4] , \n768[3] , \n768[2] , \n768[1] , UNCONNECTED_11}), .B({
        \NDiagOut[0] , Logic11, Logic11, Logic11, \NDiagOut[0] }), .LEQ(n2136), 
        .TC(n2136), .LT_LE(n404) );
    VMW_PULLDOWN U462 ( .Z(n2127) );
    VMW_PULLDOWN U465 ( .Z(n2130) );
    VMW_NOR3 U542 ( .A(n2023), .B(n2056), .C(n2046), .Z(n2025) );
    VMW_AND4 U565 ( .A(n2091), .B(n2019), .C(n2009), .D(n2000), .Z(n2047) );
    VMW_INV U655 ( .A(ScanIn[0]), .Z(n2096) );
    VMW_OR2 U559 ( .A(n2083), .B(n2077), .Z(n2085) );
    VMW_OR2 U480 ( .A(n1989), .B(ColIn[11]), .Z(ColOut[11]) );
    VMW_OR2 U510 ( .A(CallIn), .B(n2014), .Z(\n768[1] ) );
    VMW_OR2 U620 ( .A(CallIn), .B(n612), .Z(n2112) );
    VMW_OR2 U487 ( .A(n1999), .B(ColIn[4]), .Z(ColOut[4]) );
    VMW_OR3 U530 ( .A(n2024), .B(n2027), .C(n2028), .Z(n2122) );
    VMW_AOI211 U537 ( .A(n2047), .B(n2048), .C(n2049), .D(n2041), .Z(n2046) );
    VMW_OR4 U600 ( .A(NDiagIn[15]), .B(n2033), .C(ColIn[15]), .D(PDiagIn[15]), 
        .Z(n2070) );
    VMW_NOR2 U607 ( .A(CallIn), .B(n500), .Z(n2105) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_2 gt_104 ( .A({\n768[4] , 
        \n768[3] , \n768[2] , \n768[1] , \n768[0] }), .B({\NDiagOut[0] , 
        Logic11, Logic11, Logic11, Logic11}), .LEQ(n2126), .TC(n2126), .LT_LE(
        n388) );
    VMW_OR2 U517 ( .A(NDiagIn[9]), .B(n1991), .Z(NDiagOut[10]) );
    VMW_NOR2 U579 ( .A(n2080), .B(n2088), .Z(n1987) );
    VMW_AO21 U627 ( .A(n2068), .B(n2114), .C(n2116), .Z(n2115) );
    VMW_INV U649 ( .A(NDiagIn[1]), .Z(n2020) );
    VMW_PULLDOWN U470 ( .Z(n2135) );
    VMW_OR2 U479 ( .A(n1988), .B(ColIn[12]), .Z(ColOut[12]) );
    VMW_FD ReturnOut_reg ( .D(ReturnOut723), .CP(Clk), .Q(ReturnOut) );
    VMW_AND3 U539 ( .A(n2052), .B(n2053), .C(n2022), .Z(n2031) );
    VMW_NAND2 U545 ( .A(n2060), .B(n2061), .Z(n2059) );
    VMW_NAND2 U562 ( .A(ScanOut[2]), .B(n2082), .Z(n2088) );
    VMW_INV U652 ( .A(ScanIn[3]), .Z(n2093) );
    VMW_OR2 U587 ( .A(n2085), .B(n2088), .Z(n1998) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_9 gt_104_12 ( .A({
        \n768[4] , \n768[3] , \n768[2] , \n768[1] , \n768[0] }), .B({
        \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11}), .LEQ(
        n2132), .TC(n2132), .LT_LE(n580) );
    VMW_NOR2 U595 ( .A(CallIn), .B(n436), .Z(n2099) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1_DW01_cmp2_5_15 gt_104_6 ( .A({
        \n768[4] , \n768[3] , \n768[2] , \n768[1] , \n768[0] }), .B({
        \NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(
        n2138), .TC(n2138), .LT_LE(n484) );
    VMW_NAND2 U557 ( .A(n2079), .B(n2082), .Z(n2081) );
    VMW_OR2 U609 ( .A(CallIn), .B(n548), .Z(n2106) );
    VMW_MUX2I U570 ( .A(n2077), .B(n2096), .S(ScanEnable), .Z(n2015) );
    VMW_INV U640 ( .A(ScanOut[4]), .Z(n2084) );
    VMW_INV U667 ( .A(n2110), .Z(n2061) );
    VMW_OR2 U495 ( .A(PDiagIn[12]), .B(n1988), .Z(PDiagOut[11]) );
    VMW_OR2 U505 ( .A(PDiagIn[2]), .B(n2002), .Z(PDiagOut[1]) );
    VMW_OR2 U522 ( .A(NDiagIn[4]), .B(n1999), .Z(NDiagOut[5]) );
    VMW_NOR4 U612 ( .A(n2107), .B(NDiagIn[4]), .C(PDiagIn[4]), .D(ColIn[4]), 
        .Z(n2045) );
    VMW_INV U635 ( .A(PDiagIn[7]), .Z(n2006) );
endmodule


module NQueens_Control_IDWIDTH5_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, ScanId, CallIn, ReturnIn, 
    CallOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [4:0] Id;
input  [4:0] ScanIn;
output [4:0] ScanOut;
input  [4:0] ScanId;
input  Clk, Reset, RD, WR, CallIn, ReturnIn;
output ScanEnable, CallOut;
    wire n421, n387, n406, n433, n414, n395, n446, n428, n389, n408, n441, 
        n413, n434, n392, n448, n401, n426, n412, n393, n435, \status[4] , 
        n440, \ScanReg[2] , n388, n409, n449, \status[0] , n427, n400, n420, 
        \ScanReg[4] , n386, n407, \status[2] , n429, n447, \ScanReg[0] , n432, 
        n415, n394, n439, \status[6] , \ScanReg[1] , \status[7] , n422, n405, 
        n417, n430, n396, \status[3] , n445, \status[1] , n442, n410, n437, 
        n391, n425, n402, \status[5] , n450, n419, n398, \ScanReg[3] , n436, 
        n390, n411, n443, n418, n399, n424, n403, n423, n385, n404, Logic01, 
        n438, n444, n431, n397, n416;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    assign ScanOut[4] = Logic01;
    assign ScanOut[3] = Logic01;
    assign ScanOut[2] = Logic01;
    assign ScanOut[1] = Logic01;
    assign ScanOut[0] = Logic01;
    VMW_PULLDOWN U96 ( .Z(n435) );
    VMW_OAI21 U113 ( .A(n392), .B(n393), .C(n394), .Z(n449) );
    VMW_XNOR2 U134 ( .A(Addr[1]), .B(Id[1]), .Z(n397) );
    VMW_AND2 U108 ( .A(\status[5] ), .B(n387), .Z(n437) );
    VMW_INV U141 ( .A(\status[0] ), .Z(n395) );
    VMW_BUFIZ U166 ( .A(n431), .E(n415), .Z(\arr[24] ) );
    VMW_PULLDOWN U83 ( .Z(n419) );
    VMW_PULLDOWN U84 ( .Z(n420) );
    VMW_BUFIZ U148 ( .A(n412), .E(n415), .Z(\arr[23] ) );
    VMW_BUFIZ U153 ( .A(n418), .E(n415), .Z(\arr[14] ) );
    VMW_BUFIZ U174 ( .A(n439), .E(n415), .Z(\arr[18] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_PULLDOWN U101 ( .Z(Logic01) );
    VMW_AND2 U106 ( .A(\status[6] ), .B(n386), .Z(n444) );
    VMW_AO22 U121 ( .A(\ScanReg[4] ), .B(n385), .C(\status[4] ), .D(n387), .Z(
        n416) );
    VMW_AND2 U126 ( .A(n404), .B(n405), .Z(CallOut) );
    VMW_BUFIZ U168 ( .A(n433), .E(n415), .Z(\arr[3] ) );
    VMW_PULLDOWN U91 ( .Z(n429) );
    VMW_PULLDOWN U98 ( .Z(n439) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AND2 U128 ( .A(n403), .B(CallIn), .Z(n407) );
    VMW_BUFIZ U154 ( .A(n419), .E(n415), .Z(\arr[25] ) );
    VMW_BUFIZ U173 ( .A(n438), .E(n415), .Z(\arr[22] ) );
    VMW_BUFIZ U146 ( .A(n410), .E(n415), .Z(\arr[19] ) );
    VMW_BUFIZ U161 ( .A(n426), .E(n415), .Z(\arr[2] ) );
    VMW_PULLDOWN U99 ( .Z(n440) );
    VMW_OAI21 U114 ( .A(n395), .B(n393), .C(n396), .Z(n450) );
    VMW_XNOR2 U133 ( .A(Addr[3]), .B(Id[3]), .Z(n398) );
    VMW_FD \status_reg[7]  ( .D(n443), .CP(Clk), .Q(\status[7] ) );
    VMW_BUFIZ U155 ( .A(n420), .E(n415), .Z(\arr[16] ) );
    VMW_BUFIZ U172 ( .A(n437), .E(n415), .Z(\arr[5] ) );
    VMW_PULLDOWN U82 ( .Z(n418) );
    VMW_BUFIZ U169 ( .A(n434), .E(n415), .Z(\arr[26] ) );
    VMW_PULLDOWN U85 ( .Z(n421) );
    VMW_PULLDOWN U90 ( .Z(n428) );
    VMW_AND2 U107 ( .A(\status[7] ), .B(n386), .Z(n443) );
    VMW_NAND4 U120 ( .A(n406), .B(n408), .C(n390), .D(n391), .Z(n393) );
    VMW_AND5 U115 ( .A(n397), .B(n398), .C(n399), .D(n400), .E(n401), .Z(n387)
         );
    VMW_OAI21 U132 ( .A(n407), .B(n409), .C(n390), .Z(n396) );
    VMW_FD \status_reg[3]  ( .D(n447), .CP(Clk), .Q(\status[3] ) );
    VMW_PULLDOWN U97 ( .Z(n438) );
    VMW_AND2 U109 ( .A(\status[7] ), .B(n387), .Z(n436) );
    VMW_NAND2 U129 ( .A(ReturnIn), .B(n403), .Z(n408) );
    VMW_BUFIZ U147 ( .A(n411), .E(n415), .Z(\arr[0] ) );
    VMW_BUFIZ U160 ( .A(n425), .E(n415), .Z(\arr[28] ) );
    VMW_INV U140 ( .A(\status[1] ), .Z(n392) );
    VMW_BUFIZ U167 ( .A(n432), .E(n415), .Z(\arr[17] ) );
    VMW_PULLDOWN U100 ( .Z(n442) );
    VMW_AND4 U112 ( .A(n388), .B(n389), .C(n390), .D(n391), .Z(n448) );
    VMW_XNOR2 U135 ( .A(Addr[4]), .B(Id[4]), .Z(n399) );
    VMW_FD \status_reg[1]  ( .D(n449), .CP(Clk), .Q(\status[1] ) );
    VMW_AND2 U127 ( .A(n387), .B(WR), .Z(n409) );
    VMW_BUFIZ U149 ( .A(n413), .E(n415), .Z(\arr[10] ) );
    VMW_BUFIZ U152 ( .A(n417), .E(n415), .Z(\arr[27] ) );
    VMW_BUFIZ U175 ( .A(n440), .E(n415), .Z(\arr[11] ) );
    VMW_FD \status_reg[5]  ( .D(n445), .CP(Clk), .Q(\status[5] ) );
    VMW_PULLDOWN U77 ( .Z(n410) );
    VMW_PULLDOWN U79 ( .Z(n413) );
    VMW_PULLDOWN U95 ( .Z(n434) );
    VMW_AND2 U110 ( .A(\status[6] ), .B(n387), .Z(n422) );
    VMW_XNOR2 U137 ( .A(Addr[0]), .B(Id[0]), .Z(n400) );
    VMW_BUFIZ U159 ( .A(n424), .E(n415), .Z(\arr[21] ) );
    VMW_NOR2 U119 ( .A(n407), .B(CallOut), .Z(n406) );
    VMW_INV U142 ( .A(Reset), .Z(n390) );
    VMW_FD \status_reg[4]  ( .D(n446), .CP(Clk), .Q(\status[4] ) );
    VMW_BUFIZ U165 ( .A(n430), .E(n415), .Z(\arr[20] ) );
    VMW_PULLDOWN U80 ( .Z(n414) );
    VMW_PULLDOWN U87 ( .Z(n424) );
    VMW_BUFIZ U150 ( .A(n414), .E(n415), .Z(\arr[9] ) );
    VMW_BUFIZ U177 ( .A(n442), .E(n415), .Z(\arr[8] ) );
    VMW_AND2 U102 ( .A(RD), .B(n385), .Z(ScanEnable) );
    VMW_AO22 U125 ( .A(\ScanReg[0] ), .B(n385), .C(\status[0] ), .D(n387), .Z(
        n411) );
    VMW_AND2 U105 ( .A(\status[5] ), .B(n386), .Z(n445) );
    VMW_FD \status_reg[0]  ( .D(n450), .CP(Clk), .Q(\status[0] ) );
    VMW_AO22 U122 ( .A(\ScanReg[3] ), .B(n385), .C(\status[3] ), .D(n387), .Z(
        n433) );
    VMW_FD \status_reg[2]  ( .D(n448), .CP(Clk), .Q(\status[2] ) );
    VMW_PULLDOWN U89 ( .Z(n427) );
    VMW_INV U139 ( .A(\status[2] ), .Z(n404) );
    VMW_BUFIZ U157 ( .A(n422), .E(n415), .Z(\arr[6] ) );
    VMW_BUFIZ U170 ( .A(n435), .E(n415), .Z(\arr[15] ) );
    VMW_PULLDOWN U92 ( .Z(n430) );
    VMW_INV U145 ( .A(n407), .Z(n389) );
    VMW_BUFIZ U162 ( .A(n427), .E(n415), .Z(\arr[13] ) );
    VMW_FD \status_reg[6]  ( .D(n444), .CP(Clk), .Q(\status[6] ) );
    VMW_AND4 U117 ( .A(\status[1] ), .B(n402), .C(n395), .D(n404), .Z(n403) );
    VMW_PULLDOWN U78 ( .Z(n412) );
    VMW_PULLDOWN U81 ( .Z(n417) );
    VMW_OAI21 U130 ( .A(n405), .B(n386), .C(n404), .Z(n388) );
    VMW_INV U138 ( .A(n387), .Z(n385) );
    VMW_BUFIZ U156 ( .A(n421), .E(n415), .Z(\arr[12] ) );
    VMW_BUFIZ U171 ( .A(n436), .E(n415), .Z(\arr[7] ) );
    VMW_PULLDOWN U86 ( .Z(n423) );
    VMW_PULLDOWN U88 ( .Z(n425) );
    VMW_PULLDOWN U93 ( .Z(n431) );
    VMW_AND2 U104 ( .A(\status[4] ), .B(n386), .Z(n446) );
    VMW_NOR5 U116 ( .A(\status[6] ), .B(\status[7] ), .C(\status[5] ), .D(
        \status[3] ), .E(\status[4] ), .Z(n402) );
    VMW_AO22 U123 ( .A(\ScanReg[2] ), .B(n385), .C(\status[2] ), .D(n387), .Z(
        n426) );
    VMW_OR3 U131 ( .A(Reset), .B(n409), .C(n406), .Z(n394) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_PULLDOWN U94 ( .Z(n432) );
    VMW_INV U143 ( .A(n393), .Z(n386) );
    VMW_INV U144 ( .A(n409), .Z(n391) );
    VMW_BUFIZ U163 ( .A(n428), .E(n415), .Z(\arr[30] ) );
    VMW_BUFIZ U158 ( .A(n423), .E(n415), .Z(\arr[31] ) );
    VMW_BUFIZ U164 ( .A(n429), .E(n415), .Z(\arr[29] ) );
    VMW_AND2 U103 ( .A(\status[3] ), .B(n386), .Z(n447) );
    VMW_OR2 U111 ( .A(n387), .B(RD), .Z(n415) );
    VMW_XNOR2 U136 ( .A(Addr[2]), .B(Id[2]), .Z(n401) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AO22 U124 ( .A(\ScanReg[1] ), .B(n385), .C(\status[1] ), .D(n387), .Z(
        n441) );
    VMW_AND3 U118 ( .A(n402), .B(n392), .C(\status[0] ), .Z(n405) );
    VMW_BUFIZ U151 ( .A(n416), .E(n415), .Z(\arr[4] ) );
    VMW_BUFIZ U176 ( .A(n441), .E(n415), .Z(\arr[1] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \wPDiag_8[4] , \wPDiag_1[12] , \wColumn_3[4] , \wPDiag_5[10] , 
        \wColumn_13[14] , \wColumn_9[15] , \wNDiag_10[11] , \wColumn_12[8] , 
        \wNDiag_15[4] , \wNDiag_14[13] , \wColumn_3[13] , \wNDiag_4[12] , 
        \wColumn_6[9] , \wColumn_14[6] , \wNDiag_4[1] , \wNDiag_9[4] , 
        \wNDiag_10[9] , \wReturn_13[0] , \wNDiag_7[2] , \wPDiag_5[1] , 
        \wPDiag_6[2] , \wColumn_7[11] , \wPDiag_13[12] , \wPDiag_10[1] , 
        \wPDiag_13[2] , \wNDiag_1[13] , \wNDiag_1[5] , \wNDiag_2[6] , 
        \wNDiag_4[8] , \wColumn_8[6] , \wCall_11[0] , \wNDiag_5[11] , 
        \wNDiag_15[10] , \wPDiag_3[6] , \wPDiag_4[13] , \wScan_5[2] , 
        \wPDiag_10[8] , \wScan_6[1] , \wNDiag_11[12] , \wScan_11[1] , 
        \wScan_12[2] , \wColumn_5[3] , \wPDiag_5[8] , \wPDiag_15[5] , 
        \wCall_6[0] , \wColumn_6[12] , \wColumn_6[0] , \wPDiag_12[11] , 
        \wNDiag_13[3] , \wNDiag_10[0] , \wColumn_2[10] , \wPDiag_10[5] , 
        \wColumn_11[2] , \wColumn_12[1] , \wPDiag_13[6] , \wScan_0[2] , 
        \wScan_14[1] , \wPDiag_5[5] , \wPDiag_15[8] , \wNDiag_1[8] , 
        \wScan_3[1] , \wNDiag_4[5] , \wPDiag_6[6] , \wColumn_7[15] , 
        \wNDiag_7[6] , \wCall_3[0] , \wColumn_3[0] , \wNDiag_9[0] , 
        \wColumn_14[2] , \wColumn_9[11] , \wNDiag_15[0] , \wPDiag_5[14] , 
        \wNDiag_10[15] , \wColumn_13[10] , \wColumn_2[14] , \wColumn_3[9] , 
        \wPDiag_8[0] , \wColumn_5[7] , \wColumn_11[6] , \wColumn_12[5] , 
        \wNDiag_15[9] , \wColumn_6[4] , \wNDiag_9[9] , \wNDiag_10[4] , 
        \wNDiag_13[7] , \wScan_8[3] , \wPDiag_8[9] , \wPDiag_12[15] , 
        \wColumn_12[13] , \wCall_14[0] , \wPDiag_15[1] , \wNDiag_1[15] , 
        \wNDiag_1[1] , \wPDiag_3[2] , \wNDiag_2[2] , \wNDiag_5[15] , 
        \wColumn_8[12] , \wNDiag_15[14] , \wColumn_8[2] , \wScan_12[4] , 
        \wNDiag_1[3] , \wNDiag_2[0] , \wPDiag_3[0] , \wPDiag_4[15] , 
        \wScan_5[4] , \wColumn_12[11] , \wPDiag_15[3] , \wNDiag_11[14] , 
        \wColumn_8[10] , \wColumn_5[5] , \wColumn_6[6] , \wCall_8[0] , 
        \wColumn_8[0] , \wColumn_11[4] , \wColumn_12[7] , \wNDiag_13[5] , 
        \wNDiag_10[6] , \wColumn_14[9] , \wReturn_0[0] , \wPDiag_1[14] , 
        \wNDiag_4[14] , \wColumn_6[14] , \wScan_8[1] , \wColumn_14[0] , 
        \wColumn_9[13] , \wNDiag_9[2] , \wNDiag_15[2] , \wNDiag_14[15] , 
        \wColumn_3[2] , \wPDiag_3[9] , \wPDiag_8[2] , \wPDiag_10[7] , 
        \wColumn_13[12] , \wPDiag_13[4] , \wScan_0[0] , \wScan_3[3] , 
        \wPDiag_6[4] , \wScan_14[3] , \wColumn_2[12] , \wNDiag_2[9] , 
        \wColumn_3[15] , \wNDiag_4[7] , \wPDiag_5[7] , \wColumn_8[9] , 
        \wPDiag_13[14] , \wNDiag_7[4] , \wReturn_5[0] , \wColumn_5[1] , 
        \wColumn_6[10] , \wPDiag_12[13] , \wColumn_6[2] , \wNDiag_10[2] , 
        \wNDiag_13[1] , \wScan_0[4] , \wNDiag_1[11] , \wNDiag_1[7] , 
        \wNDiag_5[13] , \wNDiag_7[9] , \wColumn_11[0] , \wColumn_12[3] , 
        \wColumn_8[4] , \wNDiag_2[4] , \wColumn_8[14] , \wPDiag_3[4] , 
        \wNDiag_15[12] , \wPDiag_4[11] , \wScan_5[0] , \wScan_6[3] , 
        \wNDiag_11[10] , \wPDiag_13[9] , \wScan_11[3] , \wScan_12[0] , 
        \wColumn_12[15] , \wPDiag_15[7] , \wColumn_3[11] , \wNDiag_4[3] , 
        \wPDiag_6[9] , \wNDiag_7[0] , \wPDiag_5[3] , \wPDiag_6[0] , 
        \wColumn_7[13] , \wPDiag_10[3] , \wPDiag_13[10] , \wPDiag_13[0] , 
        \wPDiag_8[6] , \wColumn_1[8] , \wPDiag_1[10] , \wPDiag_5[12] , 
        \wNDiag_10[13] , \wNDiag_2[14] , \wColumn_3[6] , \wNDiag_4[10] , 
        \wColumn_5[8] , \wColumn_11[9] , \wNDiag_14[11] , \wNDiag_15[6] , 
        \wNDiag_9[6] , \wNDiag_13[8] , \wColumn_14[4] , \wColumn_10[4] , 
        \wColumn_11[10] , \wColumn_4[5] , \wPDiag_7[14] , \wNDiag_12[15] , 
        \wColumn_13[7] , \wNDiag_11[6] , \wColumn_7[6] , \wNDiag_12[5] , 
        \wScan_9[1] , \wColumn_15[12] , \wColumn_15[9] , \wPDiag_1[3] , 
        \wPDiag_2[0] , \wScan_13[4] , \wPDiag_14[3] , \wPDiag_15[14] , 
        \wScan_4[4] , \wPDiag_9[10] , \wNDiag_3[0] , \wColumn_5[15] , 
        \wScan_1[0] , \wPDiag_2[15] , \wPDiag_2[9] , \wNDiag_7[15] , 
        \wNDiag_8[12] , \wCall_9[0] , \wColumn_9[0] , \wScan_16[0] , 
        \wPDiag_12[4] , \wColumn_14[11] , \wScan_15[3] , \wPDiag_11[7] , 
        \wScan_2[3] , \wPDiag_4[7] , \wPDiag_7[4] , \wNDiag_5[7] , 
        \wNDiag_6[4] , \wColumn_9[9] , \wColumn_10[13] , \wReturn_1[0] , 
        \wColumn_1[1] , \wColumn_2[2] , \wNDiag_3[9] , \wNDiag_8[2] , 
        \wNDiag_9[11] , \wColumn_15[0] , \wPDiag_10[15] , \wNDiag_14[2] , 
        \wNDiag_3[4] , \wNDiag_6[9] , \wPDiag_8[13] , \wColumn_9[4] , 
        \wPDiag_9[2] , \wColumn_5[11] , \wPDiag_11[12] , \wColumn_1[13] , 
        \wPDiag_1[7] , \wScan_4[0] , \wPDiag_9[14] , \wPDiag_2[4] , 
        \wNDiag_6[12] , \wScan_7[3] , \wPDiag_15[10] , \wPDiag_7[9] , 
        \wPDiag_12[9] , \wScan_10[3] , \wScan_13[0] , \wPDiag_14[7] , 
        \wColumn_1[5] , \wNDiag_2[10] , \wPDiag_3[12] , \wReturn_4[0] , 
        \wColumn_4[1] , \wColumn_7[2] , \wPDiag_7[10] , \wNDiag_12[11] , 
        \wNDiag_12[1] , \wColumn_11[14] , \wNDiag_11[2] , \wColumn_4[12] , 
        \wPDiag_9[6] , \wColumn_10[0] , \wColumn_13[3] , \wPDiag_14[13] , 
        \wNDiag_14[6] , \wColumn_2[6] , \wPDiag_10[11] , \wNDiag_3[13] , 
        \wColumn_4[8] , \wNDiag_9[15] , \wColumn_10[9] , \wNDiag_12[8] , 
        \wColumn_15[4] , \wNDiag_8[6] , \wPDiag_2[11] , \wNDiag_5[3] , 
        \wPDiag_6[13] , \wNDiag_13[12] , \wNDiag_6[0] , \wScan_1[4] , 
        \wPDiag_4[3] , \wPDiag_7[0] , \wNDiag_3[11] , \wNDiag_7[11] , 
        \wColumn_14[15] , \wColumn_10[15] , \wPDiag_11[3] , \wScan_16[4] , 
        \wPDiag_12[0] , \wReturn_12[0] , \wPDiag_2[13] , \wNDiag_5[1] , 
        \wPDiag_6[11] , \wNDiag_6[2] , \wNDiag_13[10] , \wPDiag_4[1] , 
        \wPDiag_7[2] , \wNDiag_7[13] , \wPDiag_8[15] , \wPDiag_9[4] , 
        \wCall_10[0] , \wPDiag_11[1] , \wPDiag_12[2] , \wColumn_1[7] , 
        \wColumn_2[4] , \wPDiag_10[13] , \wPDiag_14[11] , \wColumn_4[10] , 
        \wNDiag_6[10] , \wColumn_7[9] , \wNDiag_8[4] , \wColumn_13[8] , 
        \wNDiag_14[4] , \wNDiag_11[9] , \wColumn_15[14] , \wColumn_15[6] , 
        \wPDiag_3[10] , \wScanEnable[0] , \wNDiag_2[12] , \wColumn_4[3] , 
        \wPDiag_7[12] , \wNDiag_12[13] , \wNDiag_11[0] , \wCall_7[0] , 
        \wColumn_7[0] , \wNDiag_12[3] , \wNDiag_5[8] , \wNDiag_8[14] , 
        \wColumn_10[2] , \wColumn_13[1] , \wColumn_9[6] , \wNDiag_3[6] , 
        \wColumn_5[13] , \wPDiag_11[10] , \wScan_1[2] , \wColumn_1[11] , 
        \wPDiag_2[6] , \wScan_7[1] , \wPDiag_15[12] , \wColumn_1[3] , 
        \wPDiag_1[5] , \wCall_2[0] , \wScan_4[2] , \wPDiag_11[8] , 
        \wPDiag_4[8] , \wPDiag_14[5] , \wNDiag_8[0] , \wNDiag_9[13] , 
        \wScan_10[1] , \wScan_13[2] , \wColumn_15[2] , \wNDiag_14[0] , 
        \wPDiag_1[8] , \wColumn_2[0] , \wColumn_4[14] , \wPDiag_8[11] , 
        \wPDiag_14[15] , \wPDiag_9[0] , \wPDiag_11[5] , \wColumn_14[13] , 
        \wScan_15[1] , \wScan_16[2] , \wScan_2[1] , \wPDiag_12[6] , 
        \wPDiag_4[5] , \wPDiag_7[6] , \wPDiag_14[8] , \wNDiag_3[15] , 
        \wNDiag_5[5] , \wPDiag_6[15] , \wNDiag_13[14] , \wNDiag_6[6] , 
        \wColumn_10[11] , \wColumn_1[15] , \wPDiag_1[1] , \wPDiag_9[12] , 
        \wPDiag_14[1] , \wCall_15[0] , \wPDiag_2[2] , \wNDiag_3[2] , 
        \wPDiag_11[14] , \wColumn_2[9] , \wNDiag_8[10] , \wColumn_9[2] , 
        \wColumn_11[12] , \wColumn_13[5] , \wNDiag_14[9] , \wPDiag_3[14] , 
        \wColumn_4[7] , \wColumn_7[4] , \wColumn_10[6] , \wNDiag_12[7] , 
        \wNDiag_8[9] , \wNDiag_11[4] , \wNDiag_6[14] , \wPDiag_9[9] , 
        \wScan_9[3] , \wColumn_15[10] , \wScan_1[3] , \wColumn_1[2] , 
        \wColumn_2[1] , \wReturn_2[0] , \wColumn_4[15] , \wPDiag_8[10] , 
        \wNDiag_8[1] , \wNDiag_14[1] , \wPDiag_9[1] , \wNDiag_9[12] , 
        \wColumn_15[3] , \wPDiag_4[4] , \wPDiag_14[14] , \wPDiag_1[9] , 
        \wScan_2[0] , \wPDiag_14[9] , \wPDiag_7[7] , \wPDiag_11[4] , 
        \wPDiag_12[7] , \wColumn_14[12] , \wScan_15[0] , \wScan_16[3] , 
        \wNDiag_3[14] , \wColumn_10[10] , \wColumn_1[14] , \wPDiag_2[3] , 
        \wNDiag_5[4] , \wPDiag_6[14] , \wNDiag_13[15] , \wNDiag_6[7] , 
        \wScan_7[4] , \wPDiag_9[13] , \wPDiag_1[0] , \wNDiag_8[11] , 
        \wColumn_9[3] , \wScan_10[4] , \wPDiag_14[0] , \wNDiag_3[3] , 
        \wPDiag_11[15] , \wColumn_2[8] , \wColumn_4[6] , \wNDiag_11[5] , 
        \wColumn_7[5] , \wNDiag_8[8] , \wNDiag_12[6] , \wColumn_11[13] , 
        \wNDiag_6[15] , \wColumn_10[7] , \wColumn_13[4] , \wNDiag_14[8] , 
        \wColumn_15[11] , \wPDiag_3[15] , \wScan_9[2] , \wNDiag_3[10] , 
        \wNDiag_5[0] , \wPDiag_6[10] , \wPDiag_9[8] , \wNDiag_13[11] , 
        \wNDiag_6[3] , \wColumn_10[14] , \wScan_2[4] , \wPDiag_2[12] , 
        \wNDiag_7[12] , \wScan_15[4] , \wPDiag_11[0] , \wPDiag_12[3] , 
        \wPDiag_7[3] , \wPDiag_4[0] , \wPDiag_8[14] , \wPDiag_14[10] , 
        \wColumn_1[6] , \wColumn_7[8] , \wPDiag_9[5] , \wNDiag_8[5] , 
        \wNDiag_11[8] , \wColumn_15[7] , \wNDiag_14[5] , \wColumn_2[5] , 
        \wColumn_4[11] , \wColumn_13[9] , \wPDiag_3[11] , \wPDiag_10[12] , 
        \wNDiag_6[11] , \wReturn_7[0] , \wColumn_15[15] , \wNDiag_2[13] , 
        \wNDiag_3[7] , \wColumn_4[2] , \wColumn_7[1] , \wPDiag_7[13] , 
        \wColumn_10[3] , \wColumn_13[0] , \wNDiag_12[12] , \wNDiag_12[2] , 
        \wPDiag_11[11] , \wNDiag_11[1] , \wColumn_5[12] , \wColumn_1[10] , 
        \wPDiag_1[4] , \wPDiag_4[9] , \wNDiag_5[9] , \wNDiag_8[15] , 
        \wColumn_9[7] , \wPDiag_14[4] , \wScan_10[0] , \wScan_13[3] , 
        \wPDiag_2[7] , \wScan_4[3] , \wScan_7[0] , \wPDiag_11[9] , 
        \wColumn_5[10] , \wPDiag_15[13] , \wNDiag_3[5] , \wPDiag_11[13] , 
        \wColumn_1[12] , \wPDiag_2[5] , \wNDiag_6[8] , \wPDiag_7[8] , 
        \wColumn_9[5] , \wPDiag_14[6] , \wScan_10[2] , \wScan_13[1] , 
        \wPDiag_15[11] , \wScan_4[1] , \wScan_7[2] , \wPDiag_12[8] , 
        \wPDiag_9[15] , \wPDiag_1[6] , \wPDiag_3[13] , \wNDiag_6[13] , 
        \wScan_9[4] , \wColumn_1[4] , \wColumn_2[7] , \wNDiag_2[11] , 
        \wCall_4[0] , \wColumn_4[0] , \wPDiag_7[11] , \wColumn_10[1] , 
        \wColumn_11[15] , \wColumn_13[2] , \wNDiag_11[3] , \wNDiag_12[10] , 
        \wColumn_7[3] , \wNDiag_12[0] , \wColumn_4[9] , \wPDiag_9[7] , 
        \wPDiag_14[12] , \wNDiag_8[7] , \wNDiag_9[14] , \wNDiag_12[9] , 
        \wColumn_15[5] , \wColumn_4[13] , \wColumn_10[8] , \wPDiag_10[10] , 
        \wPDiag_6[12] , \wNDiag_13[13] , \wNDiag_14[7] , \wNDiag_3[12] , 
        \wNDiag_5[2] , \wNDiag_6[1] , \wReturn_11[0] , \wColumn_1[9] , 
        \wPDiag_2[10] , \wNDiag_7[10] , \wPDiag_11[2] , \wPDiag_12[1] , 
        \wCall_13[0] , \wColumn_14[14] , \wNDiag_2[15] , \wColumn_4[4] , 
        \wPDiag_4[2] , \wColumn_7[7] , \wPDiag_7[15] , \wPDiag_7[1] , 
        \wNDiag_12[14] , \wNDiag_12[4] , \wColumn_15[8] , \wColumn_11[11] , 
        \wNDiag_11[7] , \wColumn_10[5] , \wColumn_13[6] , \wColumn_15[13] , 
        \wPDiag_1[2] , \wScan_9[0] , \wPDiag_2[1] , \wPDiag_9[11] , 
        \wNDiag_3[1] , \wNDiag_8[13] , \wReturn_9[0] , \wPDiag_14[2] , 
        \wPDiag_15[15] , \wCall_16[0] , \wColumn_9[1] , \wReturn_14[0] , 
        \wColumn_5[14] , \wScan_1[1] , \wScan_2[2] , \wPDiag_2[14] , 
        \wPDiag_7[5] , \wPDiag_2[8] , \wPDiag_4[6] , \wNDiag_7[14] , 
        \wColumn_14[10] , \wScan_15[2] , \wScan_16[1] , \wPDiag_11[6] , 
        \wPDiag_12[5] , \wColumn_10[12] , \wCall_1[0] , \wColumn_1[0] , 
        \wNDiag_3[8] , \wNDiag_5[6] , \wColumn_9[8] , \wNDiag_6[5] , 
        \wNDiag_14[3] , \wPDiag_10[14] , \wColumn_2[3] , \wCall_5[0] , 
        \wColumn_6[11] , \wPDiag_8[12] , \wNDiag_8[3] , \wNDiag_9[10] , 
        \wColumn_15[1] , \wPDiag_9[3] , \wScan_8[4] , \wPDiag_12[12] , 
        \wColumn_11[1] , \wColumn_12[2] , \wNDiag_13[0] , \wColumn_5[0] , 
        \wColumn_6[3] , \wNDiag_10[3] , \wNDiag_1[10] , \wNDiag_1[6] , 
        \wColumn_2[13] , \wNDiag_2[5] , \wColumn_8[15] , \wNDiag_15[13] , 
        \wNDiag_5[12] , \wColumn_8[5] , \wNDiag_7[8] , \wScan_11[2] , 
        \wScan_12[1] , \wColumn_3[10] , \wPDiag_3[5] , \wPDiag_4[10] , 
        \wScan_5[1] , \wPDiag_6[8] , \wColumn_12[14] , \wPDiag_15[6] , 
        \wNDiag_4[2] , \wScan_6[2] , \wPDiag_13[8] , \wNDiag_11[11] , 
        \wNDiag_7[1] , \wReturn_10[0] , \wPDiag_10[2] , \wPDiag_13[1] , 
        \wPDiag_5[13] , \wPDiag_5[2] , \wPDiag_6[1] , \wCall_12[0] , 
        \wColumn_7[12] , \wPDiag_13[11] , \wNDiag_10[12] , \wPDiag_1[11] , 
        \wNDiag_4[11] , \wPDiag_8[7] , \wColumn_14[5] , \wColumn_5[9] , 
        \wNDiag_13[9] , \wNDiag_9[7] , \wNDiag_15[7] , \wNDiag_1[14] , 
        \wColumn_3[7] , \wPDiag_3[1] , \wColumn_11[8] , \wNDiag_11[15] , 
        \wNDiag_14[10] , \wPDiag_4[14] , \wReturn_8[0] , \wColumn_12[10] , 
        \wPDiag_15[2] , \wNDiag_1[2] , \wColumn_8[1] , \wReturn_15[0] , 
        \wNDiag_2[1] , \wColumn_8[11] , \wColumn_5[4] , \wColumn_6[7] , 
        \wNDiag_10[7] , \wNDiag_13[4] , \wColumn_14[8] , \wScan_8[0] , 
        \wColumn_11[5] , \wColumn_12[6] , \wCall_0[0] , \wPDiag_1[15] , 
        \wColumn_6[15] , \wColumn_9[12] , \wNDiag_14[14] , \wColumn_3[3] , 
        \wNDiag_4[15] , \wNDiag_9[3] , \wNDiag_15[3] , \wColumn_14[1] , 
        \wPDiag_8[3] , \wColumn_13[13] , \wScan_0[1] , \wScan_3[2] , 
        \wPDiag_5[6] , \wPDiag_6[5] , \wPDiag_3[8] , \wPDiag_13[15] , 
        \wPDiag_13[5] , \wPDiag_10[6] , \wScan_14[2] , \wScan_0[3] , 
        \wNDiag_2[8] , \wScan_3[0] , \wColumn_3[14] , \wNDiag_4[6] , 
        \wNDiag_7[5] , \wColumn_8[8] , \wPDiag_5[4] , \wPDiag_6[7] , 
        \wColumn_7[14] , \wPDiag_15[9] , \wPDiag_10[4] , \wPDiag_13[7] , 
        \wScan_14[0] , \wNDiag_1[9] , \wColumn_3[1] , \wNDiag_4[4] , 
        \wNDiag_7[7] , \wNDiag_15[1] , \wColumn_9[10] , \wNDiag_9[1] , 
        \wColumn_14[3] , \wPDiag_8[1] , \wColumn_2[15] , \wReturn_3[0] , 
        \wNDiag_10[14] , \wColumn_13[11] , \wColumn_5[6] , \wPDiag_5[15] , 
        \wColumn_6[5] , \wNDiag_13[6] , \wNDiag_10[5] , \wNDiag_9[8] , 
        \wColumn_3[8] , \wColumn_12[4] , \wNDiag_15[8] , \wScan_8[2] , 
        \wColumn_11[7] , \wPDiag_8[8] , \wPDiag_12[14] , \wNDiag_1[0] , 
        \wNDiag_2[3] , \wPDiag_3[3] , \wNDiag_5[14] , \wScan_6[4] , 
        \wColumn_8[3] , \wScan_11[4] , \wColumn_12[12] , \wPDiag_15[0] , 
        \wNDiag_15[15] , \wColumn_8[13] , \wPDiag_5[11] , \wNDiag_10[10] , 
        \wColumn_13[15] , \wPDiag_1[13] , \wColumn_3[5] , \wNDiag_4[13] , 
        \wColumn_6[8] , \wPDiag_8[5] , \wNDiag_9[5] , \wNDiag_10[8] , 
        \wColumn_9[14] , \wColumn_14[7] , \wNDiag_14[12] , \wColumn_3[12] , 
        \wNDiag_4[0] , \wNDiag_7[3] , \wColumn_12[9] , \wNDiag_15[5] , 
        \wPDiag_10[0] , \wPDiag_13[3] , \wNDiag_1[12] , \wNDiag_1[4] , 
        \wScan_3[4] , \wPDiag_5[0] , \wScan_14[4] , \wPDiag_6[3] , 
        \wColumn_7[10] , \wPDiag_13[13] , \wNDiag_2[7] , \wNDiag_4[9] , 
        \wNDiag_5[10] , \wNDiag_15[11] , \wColumn_8[7] , \wPDiag_5[9] , 
        \wScan_11[0] , \wScan_12[3] , \wPDiag_15[4] , \wColumn_2[11] , 
        \wPDiag_3[7] , \wScan_6[0] , \wNDiag_11[13] , \wPDiag_4[12] , 
        \wScan_5[3] , \wColumn_5[2] , \wReturn_6[0] , \wPDiag_10[9] , 
        \wColumn_6[13] , \wPDiag_12[10] , \wColumn_11[3] , \wColumn_12[0] , 
        \wColumn_6[1] , \wNDiag_10[1] , \wNDiag_13[2] ;
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_12 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_13[4] , \wScan_13[3] , \wScan_13[2] , 
        \wScan_13[1] , \wScan_13[0] }), .ScanOut({\wScan_12[4] , \wScan_12[3] , 
        \wScan_12[2] , \wScan_12[1] , \wScan_12[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_12[0] ), .ReturnIn(\wReturn_13[0] ), .ColIn({\wColumn_12[15] , 
        \wColumn_12[14] , \wColumn_12[13] , \wColumn_12[12] , \wColumn_12[11] , 
        \wColumn_12[10] , \wColumn_12[9] , \wColumn_12[8] , \wColumn_12[7] , 
        \wColumn_12[6] , \wColumn_12[5] , \wColumn_12[4] , \wColumn_12[3] , 
        \wColumn_12[2] , \wColumn_12[1] , \wColumn_12[0] }), .PDiagIn({
        \wPDiag_12[15] , \wPDiag_12[14] , \wPDiag_12[13] , \wPDiag_12[12] , 
        \wPDiag_12[11] , \wPDiag_12[10] , \wPDiag_12[9] , \wPDiag_12[8] , 
        \wPDiag_12[7] , \wPDiag_12[6] , \wPDiag_12[5] , \wPDiag_12[4] , 
        \wPDiag_12[3] , \wPDiag_12[2] , \wPDiag_12[1] , \wPDiag_12[0] }), 
        .NDiagIn({\wNDiag_12[15] , \wNDiag_12[14] , \wNDiag_12[13] , 
        \wNDiag_12[12] , \wNDiag_12[11] , \wNDiag_12[10] , \wNDiag_12[9] , 
        \wNDiag_12[8] , \wNDiag_12[7] , \wNDiag_12[6] , \wNDiag_12[5] , 
        \wNDiag_12[4] , \wNDiag_12[3] , \wNDiag_12[2] , \wNDiag_12[1] , 
        \wNDiag_12[0] }), .CallOut(\wCall_13[0] ), .ReturnOut(\wReturn_12[0] ), 
        .ColOut({\wColumn_13[15] , \wColumn_13[14] , \wColumn_13[13] , 
        \wColumn_13[12] , \wColumn_13[11] , \wColumn_13[10] , \wColumn_13[9] , 
        \wColumn_13[8] , \wColumn_13[7] , \wColumn_13[6] , \wColumn_13[5] , 
        \wColumn_13[4] , \wColumn_13[3] , \wColumn_13[2] , \wColumn_13[1] , 
        \wColumn_13[0] }), .PDiagOut({\wPDiag_13[15] , \wPDiag_13[14] , 
        \wPDiag_13[13] , \wPDiag_13[12] , \wPDiag_13[11] , \wPDiag_13[10] , 
        \wPDiag_13[9] , \wPDiag_13[8] , \wPDiag_13[7] , \wPDiag_13[6] , 
        \wPDiag_13[5] , \wPDiag_13[4] , \wPDiag_13[3] , \wPDiag_13[2] , 
        \wPDiag_13[1] , \wPDiag_13[0] }), .NDiagOut({\wNDiag_13[15] , 
        \wNDiag_13[14] , \wNDiag_13[13] , \wNDiag_13[12] , \wNDiag_13[11] , 
        \wNDiag_13[10] , \wNDiag_13[9] , \wNDiag_13[8] , \wNDiag_13[7] , 
        \wNDiag_13[6] , \wNDiag_13[5] , \wNDiag_13[4] , \wNDiag_13[3] , 
        \wNDiag_13[2] , \wNDiag_13[1] , \wNDiag_13[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_0 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_1[4] , \wScan_1[3] , \wScan_1[2] , 
        \wScan_1[1] , \wScan_1[0] }), .ScanOut({\wScan_0[4] , \wScan_0[3] , 
        \wScan_0[2] , \wScan_0[1] , \wScan_0[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_0[0] ), .ReturnIn(\wReturn_1[0] ), .ColIn({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .PDiagIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .NDiagIn({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CallOut(\wCall_1[0] ), .ReturnOut(\wReturn_0[0] ), .ColOut({
        \wColumn_1[15] , \wColumn_1[14] , \wColumn_1[13] , \wColumn_1[12] , 
        \wColumn_1[11] , \wColumn_1[10] , \wColumn_1[9] , \wColumn_1[8] , 
        \wColumn_1[7] , \wColumn_1[6] , \wColumn_1[5] , \wColumn_1[4] , 
        \wColumn_1[3] , \wColumn_1[2] , \wColumn_1[1] , \wColumn_1[0] }), 
        .PDiagOut({\wPDiag_1[15] , \wPDiag_1[14] , \wPDiag_1[13] , 
        \wPDiag_1[12] , \wPDiag_1[11] , \wPDiag_1[10] , \wPDiag_1[9] , 
        \wPDiag_1[8] , \wPDiag_1[7] , \wPDiag_1[6] , \wPDiag_1[5] , 
        \wPDiag_1[4] , \wPDiag_1[3] , \wPDiag_1[2] , \wPDiag_1[1] , 
        \wPDiag_1[0] }), .NDiagOut({\wNDiag_1[15] , \wNDiag_1[14] , 
        \wNDiag_1[13] , \wNDiag_1[12] , \wNDiag_1[11] , \wNDiag_1[10] , 
        \wNDiag_1[9] , \wNDiag_1[8] , \wNDiag_1[7] , \wNDiag_1[6] , 
        \wNDiag_1[5] , \wNDiag_1[4] , \wNDiag_1[3] , \wNDiag_1[2] , 
        \wNDiag_1[1] , \wNDiag_1[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_2 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_3[4] , \wScan_3[3] , \wScan_3[2] , 
        \wScan_3[1] , \wScan_3[0] }), .ScanOut({\wScan_2[4] , \wScan_2[3] , 
        \wScan_2[2] , \wScan_2[1] , \wScan_2[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_2[0] ), .ReturnIn(\wReturn_3[0] ), .ColIn({\wColumn_2[15] , 
        \wColumn_2[14] , \wColumn_2[13] , \wColumn_2[12] , \wColumn_2[11] , 
        \wColumn_2[10] , \wColumn_2[9] , \wColumn_2[8] , \wColumn_2[7] , 
        \wColumn_2[6] , \wColumn_2[5] , \wColumn_2[4] , \wColumn_2[3] , 
        \wColumn_2[2] , \wColumn_2[1] , \wColumn_2[0] }), .PDiagIn({
        \wPDiag_2[15] , \wPDiag_2[14] , \wPDiag_2[13] , \wPDiag_2[12] , 
        \wPDiag_2[11] , \wPDiag_2[10] , \wPDiag_2[9] , \wPDiag_2[8] , 
        \wPDiag_2[7] , \wPDiag_2[6] , \wPDiag_2[5] , \wPDiag_2[4] , 
        \wPDiag_2[3] , \wPDiag_2[2] , \wPDiag_2[1] , \wPDiag_2[0] }), 
        .NDiagIn({\wNDiag_2[15] , \wNDiag_2[14] , \wNDiag_2[13] , 
        \wNDiag_2[12] , \wNDiag_2[11] , \wNDiag_2[10] , \wNDiag_2[9] , 
        \wNDiag_2[8] , \wNDiag_2[7] , \wNDiag_2[6] , \wNDiag_2[5] , 
        \wNDiag_2[4] , \wNDiag_2[3] , \wNDiag_2[2] , \wNDiag_2[1] , 
        \wNDiag_2[0] }), .CallOut(\wCall_3[0] ), .ReturnOut(\wReturn_2[0] ), 
        .ColOut({\wColumn_3[15] , \wColumn_3[14] , \wColumn_3[13] , 
        \wColumn_3[12] , \wColumn_3[11] , \wColumn_3[10] , \wColumn_3[9] , 
        \wColumn_3[8] , \wColumn_3[7] , \wColumn_3[6] , \wColumn_3[5] , 
        \wColumn_3[4] , \wColumn_3[3] , \wColumn_3[2] , \wColumn_3[1] , 
        \wColumn_3[0] }), .PDiagOut({\wPDiag_3[15] , \wPDiag_3[14] , 
        \wPDiag_3[13] , \wPDiag_3[12] , \wPDiag_3[11] , \wPDiag_3[10] , 
        \wPDiag_3[9] , \wPDiag_3[8] , \wPDiag_3[7] , \wPDiag_3[6] , 
        \wPDiag_3[5] , \wPDiag_3[4] , \wPDiag_3[3] , \wPDiag_3[2] , 
        \wPDiag_3[1] , \wPDiag_3[0] }), .NDiagOut({\wNDiag_3[15] , 
        \wNDiag_3[14] , \wNDiag_3[13] , \wNDiag_3[12] , \wNDiag_3[11] , 
        \wNDiag_3[10] , \wNDiag_3[9] , \wNDiag_3[8] , \wNDiag_3[7] , 
        \wNDiag_3[6] , \wNDiag_3[5] , \wNDiag_3[4] , \wNDiag_3[3] , 
        \wNDiag_3[2] , \wNDiag_3[1] , \wNDiag_3[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_3 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_4[4] , \wScan_4[3] , \wScan_4[2] , 
        \wScan_4[1] , \wScan_4[0] }), .ScanOut({\wScan_3[4] , \wScan_3[3] , 
        \wScan_3[2] , \wScan_3[1] , \wScan_3[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_3[0] ), .ReturnIn(\wReturn_4[0] ), .ColIn({\wColumn_3[15] , 
        \wColumn_3[14] , \wColumn_3[13] , \wColumn_3[12] , \wColumn_3[11] , 
        \wColumn_3[10] , \wColumn_3[9] , \wColumn_3[8] , \wColumn_3[7] , 
        \wColumn_3[6] , \wColumn_3[5] , \wColumn_3[4] , \wColumn_3[3] , 
        \wColumn_3[2] , \wColumn_3[1] , \wColumn_3[0] }), .PDiagIn({
        \wPDiag_3[15] , \wPDiag_3[14] , \wPDiag_3[13] , \wPDiag_3[12] , 
        \wPDiag_3[11] , \wPDiag_3[10] , \wPDiag_3[9] , \wPDiag_3[8] , 
        \wPDiag_3[7] , \wPDiag_3[6] , \wPDiag_3[5] , \wPDiag_3[4] , 
        \wPDiag_3[3] , \wPDiag_3[2] , \wPDiag_3[1] , \wPDiag_3[0] }), 
        .NDiagIn({\wNDiag_3[15] , \wNDiag_3[14] , \wNDiag_3[13] , 
        \wNDiag_3[12] , \wNDiag_3[11] , \wNDiag_3[10] , \wNDiag_3[9] , 
        \wNDiag_3[8] , \wNDiag_3[7] , \wNDiag_3[6] , \wNDiag_3[5] , 
        \wNDiag_3[4] , \wNDiag_3[3] , \wNDiag_3[2] , \wNDiag_3[1] , 
        \wNDiag_3[0] }), .CallOut(\wCall_4[0] ), .ReturnOut(\wReturn_3[0] ), 
        .ColOut({\wColumn_4[15] , \wColumn_4[14] , \wColumn_4[13] , 
        \wColumn_4[12] , \wColumn_4[11] , \wColumn_4[10] , \wColumn_4[9] , 
        \wColumn_4[8] , \wColumn_4[7] , \wColumn_4[6] , \wColumn_4[5] , 
        \wColumn_4[4] , \wColumn_4[3] , \wColumn_4[2] , \wColumn_4[1] , 
        \wColumn_4[0] }), .PDiagOut({\wPDiag_4[15] , \wPDiag_4[14] , 
        \wPDiag_4[13] , \wPDiag_4[12] , \wPDiag_4[11] , \wPDiag_4[10] , 
        \wPDiag_4[9] , \wPDiag_4[8] , \wPDiag_4[7] , \wPDiag_4[6] , 
        \wPDiag_4[5] , \wPDiag_4[4] , \wPDiag_4[3] , \wPDiag_4[2] , 
        \wPDiag_4[1] , \wPDiag_4[0] }), .NDiagOut({\wNDiag_4[15] , 
        \wNDiag_4[14] , \wNDiag_4[13] , \wNDiag_4[12] , \wNDiag_4[11] , 
        \wNDiag_4[10] , \wNDiag_4[9] , \wNDiag_4[8] , \wNDiag_4[7] , 
        \wNDiag_4[6] , \wNDiag_4[5] , \wNDiag_4[4] , \wNDiag_4[3] , 
        \wNDiag_4[2] , \wNDiag_4[1] , \wNDiag_4[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_4 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_5[4] , \wScan_5[3] , \wScan_5[2] , 
        \wScan_5[1] , \wScan_5[0] }), .ScanOut({\wScan_4[4] , \wScan_4[3] , 
        \wScan_4[2] , \wScan_4[1] , \wScan_4[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_4[0] ), .ReturnIn(\wReturn_5[0] ), .ColIn({\wColumn_4[15] , 
        \wColumn_4[14] , \wColumn_4[13] , \wColumn_4[12] , \wColumn_4[11] , 
        \wColumn_4[10] , \wColumn_4[9] , \wColumn_4[8] , \wColumn_4[7] , 
        \wColumn_4[6] , \wColumn_4[5] , \wColumn_4[4] , \wColumn_4[3] , 
        \wColumn_4[2] , \wColumn_4[1] , \wColumn_4[0] }), .PDiagIn({
        \wPDiag_4[15] , \wPDiag_4[14] , \wPDiag_4[13] , \wPDiag_4[12] , 
        \wPDiag_4[11] , \wPDiag_4[10] , \wPDiag_4[9] , \wPDiag_4[8] , 
        \wPDiag_4[7] , \wPDiag_4[6] , \wPDiag_4[5] , \wPDiag_4[4] , 
        \wPDiag_4[3] , \wPDiag_4[2] , \wPDiag_4[1] , \wPDiag_4[0] }), 
        .NDiagIn({\wNDiag_4[15] , \wNDiag_4[14] , \wNDiag_4[13] , 
        \wNDiag_4[12] , \wNDiag_4[11] , \wNDiag_4[10] , \wNDiag_4[9] , 
        \wNDiag_4[8] , \wNDiag_4[7] , \wNDiag_4[6] , \wNDiag_4[5] , 
        \wNDiag_4[4] , \wNDiag_4[3] , \wNDiag_4[2] , \wNDiag_4[1] , 
        \wNDiag_4[0] }), .CallOut(\wCall_5[0] ), .ReturnOut(\wReturn_4[0] ), 
        .ColOut({\wColumn_5[15] , \wColumn_5[14] , \wColumn_5[13] , 
        \wColumn_5[12] , \wColumn_5[11] , \wColumn_5[10] , \wColumn_5[9] , 
        \wColumn_5[8] , \wColumn_5[7] , \wColumn_5[6] , \wColumn_5[5] , 
        \wColumn_5[4] , \wColumn_5[3] , \wColumn_5[2] , \wColumn_5[1] , 
        \wColumn_5[0] }), .PDiagOut({\wPDiag_5[15] , \wPDiag_5[14] , 
        \wPDiag_5[13] , \wPDiag_5[12] , \wPDiag_5[11] , \wPDiag_5[10] , 
        \wPDiag_5[9] , \wPDiag_5[8] , \wPDiag_5[7] , \wPDiag_5[6] , 
        \wPDiag_5[5] , \wPDiag_5[4] , \wPDiag_5[3] , \wPDiag_5[2] , 
        \wPDiag_5[1] , \wPDiag_5[0] }), .NDiagOut({\wNDiag_5[15] , 
        \wNDiag_5[14] , \wNDiag_5[13] , \wNDiag_5[12] , \wNDiag_5[11] , 
        \wNDiag_5[10] , \wNDiag_5[9] , \wNDiag_5[8] , \wNDiag_5[7] , 
        \wNDiag_5[6] , \wNDiag_5[5] , \wNDiag_5[4] , \wNDiag_5[3] , 
        \wNDiag_5[2] , \wNDiag_5[1] , \wNDiag_5[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_5 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_6[4] , \wScan_6[3] , \wScan_6[2] , 
        \wScan_6[1] , \wScan_6[0] }), .ScanOut({\wScan_5[4] , \wScan_5[3] , 
        \wScan_5[2] , \wScan_5[1] , \wScan_5[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_5[0] ), .ReturnIn(\wReturn_6[0] ), .ColIn({\wColumn_5[15] , 
        \wColumn_5[14] , \wColumn_5[13] , \wColumn_5[12] , \wColumn_5[11] , 
        \wColumn_5[10] , \wColumn_5[9] , \wColumn_5[8] , \wColumn_5[7] , 
        \wColumn_5[6] , \wColumn_5[5] , \wColumn_5[4] , \wColumn_5[3] , 
        \wColumn_5[2] , \wColumn_5[1] , \wColumn_5[0] }), .PDiagIn({
        \wPDiag_5[15] , \wPDiag_5[14] , \wPDiag_5[13] , \wPDiag_5[12] , 
        \wPDiag_5[11] , \wPDiag_5[10] , \wPDiag_5[9] , \wPDiag_5[8] , 
        \wPDiag_5[7] , \wPDiag_5[6] , \wPDiag_5[5] , \wPDiag_5[4] , 
        \wPDiag_5[3] , \wPDiag_5[2] , \wPDiag_5[1] , \wPDiag_5[0] }), 
        .NDiagIn({\wNDiag_5[15] , \wNDiag_5[14] , \wNDiag_5[13] , 
        \wNDiag_5[12] , \wNDiag_5[11] , \wNDiag_5[10] , \wNDiag_5[9] , 
        \wNDiag_5[8] , \wNDiag_5[7] , \wNDiag_5[6] , \wNDiag_5[5] , 
        \wNDiag_5[4] , \wNDiag_5[3] , \wNDiag_5[2] , \wNDiag_5[1] , 
        \wNDiag_5[0] }), .CallOut(\wCall_6[0] ), .ReturnOut(\wReturn_5[0] ), 
        .ColOut({\wColumn_6[15] , \wColumn_6[14] , \wColumn_6[13] , 
        \wColumn_6[12] , \wColumn_6[11] , \wColumn_6[10] , \wColumn_6[9] , 
        \wColumn_6[8] , \wColumn_6[7] , \wColumn_6[6] , \wColumn_6[5] , 
        \wColumn_6[4] , \wColumn_6[3] , \wColumn_6[2] , \wColumn_6[1] , 
        \wColumn_6[0] }), .PDiagOut({\wPDiag_6[15] , \wPDiag_6[14] , 
        \wPDiag_6[13] , \wPDiag_6[12] , \wPDiag_6[11] , \wPDiag_6[10] , 
        \wPDiag_6[9] , \wPDiag_6[8] , \wPDiag_6[7] , \wPDiag_6[6] , 
        \wPDiag_6[5] , \wPDiag_6[4] , \wPDiag_6[3] , \wPDiag_6[2] , 
        \wPDiag_6[1] , \wPDiag_6[0] }), .NDiagOut({\wNDiag_6[15] , 
        \wNDiag_6[14] , \wNDiag_6[13] , \wNDiag_6[12] , \wNDiag_6[11] , 
        \wNDiag_6[10] , \wNDiag_6[9] , \wNDiag_6[8] , \wNDiag_6[7] , 
        \wNDiag_6[6] , \wNDiag_6[5] , \wNDiag_6[4] , \wNDiag_6[3] , 
        \wNDiag_6[2] , \wNDiag_6[1] , \wNDiag_6[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_15 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_16[4] , \wScan_16[3] , \wScan_16[2] , 
        \wScan_16[1] , \wScan_16[0] }), .ScanOut({\wScan_15[4] , \wScan_15[3] , 
        \wScan_15[2] , \wScan_15[1] , \wScan_15[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_15[0] ), .ReturnIn(1'b0), .ColIn({\wColumn_15[15] , 
        \wColumn_15[14] , \wColumn_15[13] , \wColumn_15[12] , \wColumn_15[11] , 
        \wColumn_15[10] , \wColumn_15[9] , \wColumn_15[8] , \wColumn_15[7] , 
        \wColumn_15[6] , \wColumn_15[5] , \wColumn_15[4] , \wColumn_15[3] , 
        \wColumn_15[2] , \wColumn_15[1] , \wColumn_15[0] }), .PDiagIn({
        \wPDiag_15[15] , \wPDiag_15[14] , \wPDiag_15[13] , \wPDiag_15[12] , 
        \wPDiag_15[11] , \wPDiag_15[10] , \wPDiag_15[9] , \wPDiag_15[8] , 
        \wPDiag_15[7] , \wPDiag_15[6] , \wPDiag_15[5] , \wPDiag_15[4] , 
        \wPDiag_15[3] , \wPDiag_15[2] , \wPDiag_15[1] , \wPDiag_15[0] }), 
        .NDiagIn({\wNDiag_15[15] , \wNDiag_15[14] , \wNDiag_15[13] , 
        \wNDiag_15[12] , \wNDiag_15[11] , \wNDiag_15[10] , \wNDiag_15[9] , 
        \wNDiag_15[8] , \wNDiag_15[7] , \wNDiag_15[6] , \wNDiag_15[5] , 
        \wNDiag_15[4] , \wNDiag_15[3] , \wNDiag_15[2] , \wNDiag_15[1] , 
        \wNDiag_15[0] }), .CallOut(\wCall_16[0] ), .ReturnOut(\wReturn_15[0] )
         );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_13 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_14[4] , \wScan_14[3] , \wScan_14[2] , 
        \wScan_14[1] , \wScan_14[0] }), .ScanOut({\wScan_13[4] , \wScan_13[3] , 
        \wScan_13[2] , \wScan_13[1] , \wScan_13[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_13[0] ), .ReturnIn(\wReturn_14[0] ), .ColIn({\wColumn_13[15] , 
        \wColumn_13[14] , \wColumn_13[13] , \wColumn_13[12] , \wColumn_13[11] , 
        \wColumn_13[10] , \wColumn_13[9] , \wColumn_13[8] , \wColumn_13[7] , 
        \wColumn_13[6] , \wColumn_13[5] , \wColumn_13[4] , \wColumn_13[3] , 
        \wColumn_13[2] , \wColumn_13[1] , \wColumn_13[0] }), .PDiagIn({
        \wPDiag_13[15] , \wPDiag_13[14] , \wPDiag_13[13] , \wPDiag_13[12] , 
        \wPDiag_13[11] , \wPDiag_13[10] , \wPDiag_13[9] , \wPDiag_13[8] , 
        \wPDiag_13[7] , \wPDiag_13[6] , \wPDiag_13[5] , \wPDiag_13[4] , 
        \wPDiag_13[3] , \wPDiag_13[2] , \wPDiag_13[1] , \wPDiag_13[0] }), 
        .NDiagIn({\wNDiag_13[15] , \wNDiag_13[14] , \wNDiag_13[13] , 
        \wNDiag_13[12] , \wNDiag_13[11] , \wNDiag_13[10] , \wNDiag_13[9] , 
        \wNDiag_13[8] , \wNDiag_13[7] , \wNDiag_13[6] , \wNDiag_13[5] , 
        \wNDiag_13[4] , \wNDiag_13[3] , \wNDiag_13[2] , \wNDiag_13[1] , 
        \wNDiag_13[0] }), .CallOut(\wCall_14[0] ), .ReturnOut(\wReturn_13[0] ), 
        .ColOut({\wColumn_14[15] , \wColumn_14[14] , \wColumn_14[13] , 
        \wColumn_14[12] , \wColumn_14[11] , \wColumn_14[10] , \wColumn_14[9] , 
        \wColumn_14[8] , \wColumn_14[7] , \wColumn_14[6] , \wColumn_14[5] , 
        \wColumn_14[4] , \wColumn_14[3] , \wColumn_14[2] , \wColumn_14[1] , 
        \wColumn_14[0] }), .PDiagOut({\wPDiag_14[15] , \wPDiag_14[14] , 
        \wPDiag_14[13] , \wPDiag_14[12] , \wPDiag_14[11] , \wPDiag_14[10] , 
        \wPDiag_14[9] , \wPDiag_14[8] , \wPDiag_14[7] , \wPDiag_14[6] , 
        \wPDiag_14[5] , \wPDiag_14[4] , \wPDiag_14[3] , \wPDiag_14[2] , 
        \wPDiag_14[1] , \wPDiag_14[0] }), .NDiagOut({\wNDiag_14[15] , 
        \wNDiag_14[14] , \wNDiag_14[13] , \wNDiag_14[12] , \wNDiag_14[11] , 
        \wNDiag_14[10] , \wNDiag_14[9] , \wNDiag_14[8] , \wNDiag_14[7] , 
        \wNDiag_14[6] , \wNDiag_14[5] , \wNDiag_14[4] , \wNDiag_14[3] , 
        \wNDiag_14[2] , \wNDiag_14[1] , \wNDiag_14[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_14 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_15[4] , \wScan_15[3] , \wScan_15[2] , 
        \wScan_15[1] , \wScan_15[0] }), .ScanOut({\wScan_14[4] , \wScan_14[3] , 
        \wScan_14[2] , \wScan_14[1] , \wScan_14[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_14[0] ), .ReturnIn(\wReturn_15[0] ), .ColIn({\wColumn_14[15] , 
        \wColumn_14[14] , \wColumn_14[13] , \wColumn_14[12] , \wColumn_14[11] , 
        \wColumn_14[10] , \wColumn_14[9] , \wColumn_14[8] , \wColumn_14[7] , 
        \wColumn_14[6] , \wColumn_14[5] , \wColumn_14[4] , \wColumn_14[3] , 
        \wColumn_14[2] , \wColumn_14[1] , \wColumn_14[0] }), .PDiagIn({
        \wPDiag_14[15] , \wPDiag_14[14] , \wPDiag_14[13] , \wPDiag_14[12] , 
        \wPDiag_14[11] , \wPDiag_14[10] , \wPDiag_14[9] , \wPDiag_14[8] , 
        \wPDiag_14[7] , \wPDiag_14[6] , \wPDiag_14[5] , \wPDiag_14[4] , 
        \wPDiag_14[3] , \wPDiag_14[2] , \wPDiag_14[1] , \wPDiag_14[0] }), 
        .NDiagIn({\wNDiag_14[15] , \wNDiag_14[14] , \wNDiag_14[13] , 
        \wNDiag_14[12] , \wNDiag_14[11] , \wNDiag_14[10] , \wNDiag_14[9] , 
        \wNDiag_14[8] , \wNDiag_14[7] , \wNDiag_14[6] , \wNDiag_14[5] , 
        \wNDiag_14[4] , \wNDiag_14[3] , \wNDiag_14[2] , \wNDiag_14[1] , 
        \wNDiag_14[0] }), .CallOut(\wCall_15[0] ), .ReturnOut(\wReturn_14[0] ), 
        .ColOut({\wColumn_15[15] , \wColumn_15[14] , \wColumn_15[13] , 
        \wColumn_15[12] , \wColumn_15[11] , \wColumn_15[10] , \wColumn_15[9] , 
        \wColumn_15[8] , \wColumn_15[7] , \wColumn_15[6] , \wColumn_15[5] , 
        \wColumn_15[4] , \wColumn_15[3] , \wColumn_15[2] , \wColumn_15[1] , 
        \wColumn_15[0] }), .PDiagOut({\wPDiag_15[15] , \wPDiag_15[14] , 
        \wPDiag_15[13] , \wPDiag_15[12] , \wPDiag_15[11] , \wPDiag_15[10] , 
        \wPDiag_15[9] , \wPDiag_15[8] , \wPDiag_15[7] , \wPDiag_15[6] , 
        \wPDiag_15[5] , \wPDiag_15[4] , \wPDiag_15[3] , \wPDiag_15[2] , 
        \wPDiag_15[1] , \wPDiag_15[0] }), .NDiagOut({\wNDiag_15[15] , 
        \wNDiag_15[14] , \wNDiag_15[13] , \wNDiag_15[12] , \wNDiag_15[11] , 
        \wNDiag_15[10] , \wNDiag_15[9] , \wNDiag_15[8] , \wNDiag_15[7] , 
        \wNDiag_15[6] , \wNDiag_15[5] , \wNDiag_15[4] , \wNDiag_15[3] , 
        \wNDiag_15[2] , \wNDiag_15[1] , \wNDiag_15[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_9 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_10[4] , \wScan_10[3] , \wScan_10[2] , 
        \wScan_10[1] , \wScan_10[0] }), .ScanOut({\wScan_9[4] , \wScan_9[3] , 
        \wScan_9[2] , \wScan_9[1] , \wScan_9[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_9[0] ), .ReturnIn(\wReturn_10[0] ), .ColIn({\wColumn_9[15] , 
        \wColumn_9[14] , \wColumn_9[13] , \wColumn_9[12] , \wColumn_9[11] , 
        \wColumn_9[10] , \wColumn_9[9] , \wColumn_9[8] , \wColumn_9[7] , 
        \wColumn_9[6] , \wColumn_9[5] , \wColumn_9[4] , \wColumn_9[3] , 
        \wColumn_9[2] , \wColumn_9[1] , \wColumn_9[0] }), .PDiagIn({
        \wPDiag_9[15] , \wPDiag_9[14] , \wPDiag_9[13] , \wPDiag_9[12] , 
        \wPDiag_9[11] , \wPDiag_9[10] , \wPDiag_9[9] , \wPDiag_9[8] , 
        \wPDiag_9[7] , \wPDiag_9[6] , \wPDiag_9[5] , \wPDiag_9[4] , 
        \wPDiag_9[3] , \wPDiag_9[2] , \wPDiag_9[1] , \wPDiag_9[0] }), 
        .NDiagIn({\wNDiag_9[15] , \wNDiag_9[14] , \wNDiag_9[13] , 
        \wNDiag_9[12] , \wNDiag_9[11] , \wNDiag_9[10] , \wNDiag_9[9] , 
        \wNDiag_9[8] , \wNDiag_9[7] , \wNDiag_9[6] , \wNDiag_9[5] , 
        \wNDiag_9[4] , \wNDiag_9[3] , \wNDiag_9[2] , \wNDiag_9[1] , 
        \wNDiag_9[0] }), .CallOut(\wCall_10[0] ), .ReturnOut(\wReturn_9[0] ), 
        .ColOut({\wColumn_10[15] , \wColumn_10[14] , \wColumn_10[13] , 
        \wColumn_10[12] , \wColumn_10[11] , \wColumn_10[10] , \wColumn_10[9] , 
        \wColumn_10[8] , \wColumn_10[7] , \wColumn_10[6] , \wColumn_10[5] , 
        \wColumn_10[4] , \wColumn_10[3] , \wColumn_10[2] , \wColumn_10[1] , 
        \wColumn_10[0] }), .PDiagOut({\wPDiag_10[15] , \wPDiag_10[14] , 
        \wPDiag_10[13] , \wPDiag_10[12] , \wPDiag_10[11] , \wPDiag_10[10] , 
        \wPDiag_10[9] , \wPDiag_10[8] , \wPDiag_10[7] , \wPDiag_10[6] , 
        \wPDiag_10[5] , \wPDiag_10[4] , \wPDiag_10[3] , \wPDiag_10[2] , 
        \wPDiag_10[1] , \wPDiag_10[0] }), .NDiagOut({\wNDiag_10[15] , 
        \wNDiag_10[14] , \wNDiag_10[13] , \wNDiag_10[12] , \wNDiag_10[11] , 
        \wNDiag_10[10] , \wNDiag_10[9] , \wNDiag_10[8] , \wNDiag_10[7] , 
        \wNDiag_10[6] , \wNDiag_10[5] , \wNDiag_10[4] , \wNDiag_10[3] , 
        \wNDiag_10[2] , \wNDiag_10[1] , \wNDiag_10[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_11 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_12[4] , \wScan_12[3] , \wScan_12[2] , 
        \wScan_12[1] , \wScan_12[0] }), .ScanOut({\wScan_11[4] , \wScan_11[3] , 
        \wScan_11[2] , \wScan_11[1] , \wScan_11[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_11[0] ), .ReturnIn(\wReturn_12[0] ), .ColIn({\wColumn_11[15] , 
        \wColumn_11[14] , \wColumn_11[13] , \wColumn_11[12] , \wColumn_11[11] , 
        \wColumn_11[10] , \wColumn_11[9] , \wColumn_11[8] , \wColumn_11[7] , 
        \wColumn_11[6] , \wColumn_11[5] , \wColumn_11[4] , \wColumn_11[3] , 
        \wColumn_11[2] , \wColumn_11[1] , \wColumn_11[0] }), .PDiagIn({
        \wPDiag_11[15] , \wPDiag_11[14] , \wPDiag_11[13] , \wPDiag_11[12] , 
        \wPDiag_11[11] , \wPDiag_11[10] , \wPDiag_11[9] , \wPDiag_11[8] , 
        \wPDiag_11[7] , \wPDiag_11[6] , \wPDiag_11[5] , \wPDiag_11[4] , 
        \wPDiag_11[3] , \wPDiag_11[2] , \wPDiag_11[1] , \wPDiag_11[0] }), 
        .NDiagIn({\wNDiag_11[15] , \wNDiag_11[14] , \wNDiag_11[13] , 
        \wNDiag_11[12] , \wNDiag_11[11] , \wNDiag_11[10] , \wNDiag_11[9] , 
        \wNDiag_11[8] , \wNDiag_11[7] , \wNDiag_11[6] , \wNDiag_11[5] , 
        \wNDiag_11[4] , \wNDiag_11[3] , \wNDiag_11[2] , \wNDiag_11[1] , 
        \wNDiag_11[0] }), .CallOut(\wCall_12[0] ), .ReturnOut(\wReturn_11[0] ), 
        .ColOut({\wColumn_12[15] , \wColumn_12[14] , \wColumn_12[13] , 
        \wColumn_12[12] , \wColumn_12[11] , \wColumn_12[10] , \wColumn_12[9] , 
        \wColumn_12[8] , \wColumn_12[7] , \wColumn_12[6] , \wColumn_12[5] , 
        \wColumn_12[4] , \wColumn_12[3] , \wColumn_12[2] , \wColumn_12[1] , 
        \wColumn_12[0] }), .PDiagOut({\wPDiag_12[15] , \wPDiag_12[14] , 
        \wPDiag_12[13] , \wPDiag_12[12] , \wPDiag_12[11] , \wPDiag_12[10] , 
        \wPDiag_12[9] , \wPDiag_12[8] , \wPDiag_12[7] , \wPDiag_12[6] , 
        \wPDiag_12[5] , \wPDiag_12[4] , \wPDiag_12[3] , \wPDiag_12[2] , 
        \wPDiag_12[1] , \wPDiag_12[0] }), .NDiagOut({\wNDiag_12[15] , 
        \wNDiag_12[14] , \wNDiag_12[13] , \wNDiag_12[12] , \wNDiag_12[11] , 
        \wNDiag_12[10] , \wNDiag_12[9] , \wNDiag_12[8] , \wNDiag_12[7] , 
        \wNDiag_12[6] , \wNDiag_12[5] , \wNDiag_12[4] , \wNDiag_12[3] , 
        \wNDiag_12[2] , \wNDiag_12[1] , \wNDiag_12[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_1 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_2[4] , \wScan_2[3] , \wScan_2[2] , 
        \wScan_2[1] , \wScan_2[0] }), .ScanOut({\wScan_1[4] , \wScan_1[3] , 
        \wScan_1[2] , \wScan_1[1] , \wScan_1[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_1[0] ), .ReturnIn(\wReturn_2[0] ), .ColIn({\wColumn_1[15] , 
        \wColumn_1[14] , \wColumn_1[13] , \wColumn_1[12] , \wColumn_1[11] , 
        \wColumn_1[10] , \wColumn_1[9] , \wColumn_1[8] , \wColumn_1[7] , 
        \wColumn_1[6] , \wColumn_1[5] , \wColumn_1[4] , \wColumn_1[3] , 
        \wColumn_1[2] , \wColumn_1[1] , \wColumn_1[0] }), .PDiagIn({
        \wPDiag_1[15] , \wPDiag_1[14] , \wPDiag_1[13] , \wPDiag_1[12] , 
        \wPDiag_1[11] , \wPDiag_1[10] , \wPDiag_1[9] , \wPDiag_1[8] , 
        \wPDiag_1[7] , \wPDiag_1[6] , \wPDiag_1[5] , \wPDiag_1[4] , 
        \wPDiag_1[3] , \wPDiag_1[2] , \wPDiag_1[1] , \wPDiag_1[0] }), 
        .NDiagIn({\wNDiag_1[15] , \wNDiag_1[14] , \wNDiag_1[13] , 
        \wNDiag_1[12] , \wNDiag_1[11] , \wNDiag_1[10] , \wNDiag_1[9] , 
        \wNDiag_1[8] , \wNDiag_1[7] , \wNDiag_1[6] , \wNDiag_1[5] , 
        \wNDiag_1[4] , \wNDiag_1[3] , \wNDiag_1[2] , \wNDiag_1[1] , 
        \wNDiag_1[0] }), .CallOut(\wCall_2[0] ), .ReturnOut(\wReturn_1[0] ), 
        .ColOut({\wColumn_2[15] , \wColumn_2[14] , \wColumn_2[13] , 
        \wColumn_2[12] , \wColumn_2[11] , \wColumn_2[10] , \wColumn_2[9] , 
        \wColumn_2[8] , \wColumn_2[7] , \wColumn_2[6] , \wColumn_2[5] , 
        \wColumn_2[4] , \wColumn_2[3] , \wColumn_2[2] , \wColumn_2[1] , 
        \wColumn_2[0] }), .PDiagOut({\wPDiag_2[15] , \wPDiag_2[14] , 
        \wPDiag_2[13] , \wPDiag_2[12] , \wPDiag_2[11] , \wPDiag_2[10] , 
        \wPDiag_2[9] , \wPDiag_2[8] , \wPDiag_2[7] , \wPDiag_2[6] , 
        \wPDiag_2[5] , \wPDiag_2[4] , \wPDiag_2[3] , \wPDiag_2[2] , 
        \wPDiag_2[1] , \wPDiag_2[0] }), .NDiagOut({\wNDiag_2[15] , 
        \wNDiag_2[14] , \wNDiag_2[13] , \wNDiag_2[12] , \wNDiag_2[11] , 
        \wNDiag_2[10] , \wNDiag_2[9] , \wNDiag_2[8] , \wNDiag_2[7] , 
        \wNDiag_2[6] , \wNDiag_2[5] , \wNDiag_2[4] , \wNDiag_2[3] , 
        \wNDiag_2[2] , \wNDiag_2[1] , \wNDiag_2[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_6 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_7[4] , \wScan_7[3] , \wScan_7[2] , 
        \wScan_7[1] , \wScan_7[0] }), .ScanOut({\wScan_6[4] , \wScan_6[3] , 
        \wScan_6[2] , \wScan_6[1] , \wScan_6[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_6[0] ), .ReturnIn(\wReturn_7[0] ), .ColIn({\wColumn_6[15] , 
        \wColumn_6[14] , \wColumn_6[13] , \wColumn_6[12] , \wColumn_6[11] , 
        \wColumn_6[10] , \wColumn_6[9] , \wColumn_6[8] , \wColumn_6[7] , 
        \wColumn_6[6] , \wColumn_6[5] , \wColumn_6[4] , \wColumn_6[3] , 
        \wColumn_6[2] , \wColumn_6[1] , \wColumn_6[0] }), .PDiagIn({
        \wPDiag_6[15] , \wPDiag_6[14] , \wPDiag_6[13] , \wPDiag_6[12] , 
        \wPDiag_6[11] , \wPDiag_6[10] , \wPDiag_6[9] , \wPDiag_6[8] , 
        \wPDiag_6[7] , \wPDiag_6[6] , \wPDiag_6[5] , \wPDiag_6[4] , 
        \wPDiag_6[3] , \wPDiag_6[2] , \wPDiag_6[1] , \wPDiag_6[0] }), 
        .NDiagIn({\wNDiag_6[15] , \wNDiag_6[14] , \wNDiag_6[13] , 
        \wNDiag_6[12] , \wNDiag_6[11] , \wNDiag_6[10] , \wNDiag_6[9] , 
        \wNDiag_6[8] , \wNDiag_6[7] , \wNDiag_6[6] , \wNDiag_6[5] , 
        \wNDiag_6[4] , \wNDiag_6[3] , \wNDiag_6[2] , \wNDiag_6[1] , 
        \wNDiag_6[0] }), .CallOut(\wCall_7[0] ), .ReturnOut(\wReturn_6[0] ), 
        .ColOut({\wColumn_7[15] , \wColumn_7[14] , \wColumn_7[13] , 
        \wColumn_7[12] , \wColumn_7[11] , \wColumn_7[10] , \wColumn_7[9] , 
        \wColumn_7[8] , \wColumn_7[7] , \wColumn_7[6] , \wColumn_7[5] , 
        \wColumn_7[4] , \wColumn_7[3] , \wColumn_7[2] , \wColumn_7[1] , 
        \wColumn_7[0] }), .PDiagOut({\wPDiag_7[15] , \wPDiag_7[14] , 
        \wPDiag_7[13] , \wPDiag_7[12] , \wPDiag_7[11] , \wPDiag_7[10] , 
        \wPDiag_7[9] , \wPDiag_7[8] , \wPDiag_7[7] , \wPDiag_7[6] , 
        \wPDiag_7[5] , \wPDiag_7[4] , \wPDiag_7[3] , \wPDiag_7[2] , 
        \wPDiag_7[1] , \wPDiag_7[0] }), .NDiagOut({\wNDiag_7[15] , 
        \wNDiag_7[14] , \wNDiag_7[13] , \wNDiag_7[12] , \wNDiag_7[11] , 
        \wNDiag_7[10] , \wNDiag_7[9] , \wNDiag_7[8] , \wNDiag_7[7] , 
        \wNDiag_7[6] , \wNDiag_7[5] , \wNDiag_7[4] , \wNDiag_7[3] , 
        \wNDiag_7[2] , \wNDiag_7[1] , \wNDiag_7[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_7 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_8[4] , \wScan_8[3] , \wScan_8[2] , 
        \wScan_8[1] , \wScan_8[0] }), .ScanOut({\wScan_7[4] , \wScan_7[3] , 
        \wScan_7[2] , \wScan_7[1] , \wScan_7[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_7[0] ), .ReturnIn(\wReturn_8[0] ), .ColIn({\wColumn_7[15] , 
        \wColumn_7[14] , \wColumn_7[13] , \wColumn_7[12] , \wColumn_7[11] , 
        \wColumn_7[10] , \wColumn_7[9] , \wColumn_7[8] , \wColumn_7[7] , 
        \wColumn_7[6] , \wColumn_7[5] , \wColumn_7[4] , \wColumn_7[3] , 
        \wColumn_7[2] , \wColumn_7[1] , \wColumn_7[0] }), .PDiagIn({
        \wPDiag_7[15] , \wPDiag_7[14] , \wPDiag_7[13] , \wPDiag_7[12] , 
        \wPDiag_7[11] , \wPDiag_7[10] , \wPDiag_7[9] , \wPDiag_7[8] , 
        \wPDiag_7[7] , \wPDiag_7[6] , \wPDiag_7[5] , \wPDiag_7[4] , 
        \wPDiag_7[3] , \wPDiag_7[2] , \wPDiag_7[1] , \wPDiag_7[0] }), 
        .NDiagIn({\wNDiag_7[15] , \wNDiag_7[14] , \wNDiag_7[13] , 
        \wNDiag_7[12] , \wNDiag_7[11] , \wNDiag_7[10] , \wNDiag_7[9] , 
        \wNDiag_7[8] , \wNDiag_7[7] , \wNDiag_7[6] , \wNDiag_7[5] , 
        \wNDiag_7[4] , \wNDiag_7[3] , \wNDiag_7[2] , \wNDiag_7[1] , 
        \wNDiag_7[0] }), .CallOut(\wCall_8[0] ), .ReturnOut(\wReturn_7[0] ), 
        .ColOut({\wColumn_8[15] , \wColumn_8[14] , \wColumn_8[13] , 
        \wColumn_8[12] , \wColumn_8[11] , \wColumn_8[10] , \wColumn_8[9] , 
        \wColumn_8[8] , \wColumn_8[7] , \wColumn_8[6] , \wColumn_8[5] , 
        \wColumn_8[4] , \wColumn_8[3] , \wColumn_8[2] , \wColumn_8[1] , 
        \wColumn_8[0] }), .PDiagOut({\wPDiag_8[15] , \wPDiag_8[14] , 
        \wPDiag_8[13] , \wPDiag_8[12] , \wPDiag_8[11] , \wPDiag_8[10] , 
        \wPDiag_8[9] , \wPDiag_8[8] , \wPDiag_8[7] , \wPDiag_8[6] , 
        \wPDiag_8[5] , \wPDiag_8[4] , \wPDiag_8[3] , \wPDiag_8[2] , 
        \wPDiag_8[1] , \wPDiag_8[0] }), .NDiagOut({\wNDiag_8[15] , 
        \wNDiag_8[14] , \wNDiag_8[13] , \wNDiag_8[12] , \wNDiag_8[11] , 
        \wNDiag_8[10] , \wNDiag_8[9] , \wNDiag_8[8] , \wNDiag_8[7] , 
        \wNDiag_8[6] , \wNDiag_8[5] , \wNDiag_8[4] , \wNDiag_8[3] , 
        \wNDiag_8[2] , \wNDiag_8[1] , \wNDiag_8[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_8 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_9[4] , \wScan_9[3] , \wScan_9[2] , 
        \wScan_9[1] , \wScan_9[0] }), .ScanOut({\wScan_8[4] , \wScan_8[3] , 
        \wScan_8[2] , \wScan_8[1] , \wScan_8[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_8[0] ), .ReturnIn(\wReturn_9[0] ), .ColIn({\wColumn_8[15] , 
        \wColumn_8[14] , \wColumn_8[13] , \wColumn_8[12] , \wColumn_8[11] , 
        \wColumn_8[10] , \wColumn_8[9] , \wColumn_8[8] , \wColumn_8[7] , 
        \wColumn_8[6] , \wColumn_8[5] , \wColumn_8[4] , \wColumn_8[3] , 
        \wColumn_8[2] , \wColumn_8[1] , \wColumn_8[0] }), .PDiagIn({
        \wPDiag_8[15] , \wPDiag_8[14] , \wPDiag_8[13] , \wPDiag_8[12] , 
        \wPDiag_8[11] , \wPDiag_8[10] , \wPDiag_8[9] , \wPDiag_8[8] , 
        \wPDiag_8[7] , \wPDiag_8[6] , \wPDiag_8[5] , \wPDiag_8[4] , 
        \wPDiag_8[3] , \wPDiag_8[2] , \wPDiag_8[1] , \wPDiag_8[0] }), 
        .NDiagIn({\wNDiag_8[15] , \wNDiag_8[14] , \wNDiag_8[13] , 
        \wNDiag_8[12] , \wNDiag_8[11] , \wNDiag_8[10] , \wNDiag_8[9] , 
        \wNDiag_8[8] , \wNDiag_8[7] , \wNDiag_8[6] , \wNDiag_8[5] , 
        \wNDiag_8[4] , \wNDiag_8[3] , \wNDiag_8[2] , \wNDiag_8[1] , 
        \wNDiag_8[0] }), .CallOut(\wCall_9[0] ), .ReturnOut(\wReturn_8[0] ), 
        .ColOut({\wColumn_9[15] , \wColumn_9[14] , \wColumn_9[13] , 
        \wColumn_9[12] , \wColumn_9[11] , \wColumn_9[10] , \wColumn_9[9] , 
        \wColumn_9[8] , \wColumn_9[7] , \wColumn_9[6] , \wColumn_9[5] , 
        \wColumn_9[4] , \wColumn_9[3] , \wColumn_9[2] , \wColumn_9[1] , 
        \wColumn_9[0] }), .PDiagOut({\wPDiag_9[15] , \wPDiag_9[14] , 
        \wPDiag_9[13] , \wPDiag_9[12] , \wPDiag_9[11] , \wPDiag_9[10] , 
        \wPDiag_9[9] , \wPDiag_9[8] , \wPDiag_9[7] , \wPDiag_9[6] , 
        \wPDiag_9[5] , \wPDiag_9[4] , \wPDiag_9[3] , \wPDiag_9[2] , 
        \wPDiag_9[1] , \wPDiag_9[0] }), .NDiagOut({\wNDiag_9[15] , 
        \wNDiag_9[14] , \wNDiag_9[13] , \wNDiag_9[12] , \wNDiag_9[11] , 
        \wNDiag_9[10] , \wNDiag_9[9] , \wNDiag_9[8] , \wNDiag_9[7] , 
        \wNDiag_9[6] , \wNDiag_9[5] , \wNDiag_9[4] , \wNDiag_9[3] , 
        \wNDiag_9[2] , \wNDiag_9[1] , \wNDiag_9[0] }) );
    NQueens_Node_WIDTH16_IDWIDTH5_SCAN1 U_NQueens_Node_10 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_11[4] , \wScan_11[3] , \wScan_11[2] , 
        \wScan_11[1] , \wScan_11[0] }), .ScanOut({\wScan_10[4] , \wScan_10[3] , 
        \wScan_10[2] , \wScan_10[1] , \wScan_10[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_10[0] ), .ReturnIn(\wReturn_11[0] ), .ColIn({\wColumn_10[15] , 
        \wColumn_10[14] , \wColumn_10[13] , \wColumn_10[12] , \wColumn_10[11] , 
        \wColumn_10[10] , \wColumn_10[9] , \wColumn_10[8] , \wColumn_10[7] , 
        \wColumn_10[6] , \wColumn_10[5] , \wColumn_10[4] , \wColumn_10[3] , 
        \wColumn_10[2] , \wColumn_10[1] , \wColumn_10[0] }), .PDiagIn({
        \wPDiag_10[15] , \wPDiag_10[14] , \wPDiag_10[13] , \wPDiag_10[12] , 
        \wPDiag_10[11] , \wPDiag_10[10] , \wPDiag_10[9] , \wPDiag_10[8] , 
        \wPDiag_10[7] , \wPDiag_10[6] , \wPDiag_10[5] , \wPDiag_10[4] , 
        \wPDiag_10[3] , \wPDiag_10[2] , \wPDiag_10[1] , \wPDiag_10[0] }), 
        .NDiagIn({\wNDiag_10[15] , \wNDiag_10[14] , \wNDiag_10[13] , 
        \wNDiag_10[12] , \wNDiag_10[11] , \wNDiag_10[10] , \wNDiag_10[9] , 
        \wNDiag_10[8] , \wNDiag_10[7] , \wNDiag_10[6] , \wNDiag_10[5] , 
        \wNDiag_10[4] , \wNDiag_10[3] , \wNDiag_10[2] , \wNDiag_10[1] , 
        \wNDiag_10[0] }), .CallOut(\wCall_11[0] ), .ReturnOut(\wReturn_10[0] ), 
        .ColOut({\wColumn_11[15] , \wColumn_11[14] , \wColumn_11[13] , 
        \wColumn_11[12] , \wColumn_11[11] , \wColumn_11[10] , \wColumn_11[9] , 
        \wColumn_11[8] , \wColumn_11[7] , \wColumn_11[6] , \wColumn_11[5] , 
        \wColumn_11[4] , \wColumn_11[3] , \wColumn_11[2] , \wColumn_11[1] , 
        \wColumn_11[0] }), .PDiagOut({\wPDiag_11[15] , \wPDiag_11[14] , 
        \wPDiag_11[13] , \wPDiag_11[12] , \wPDiag_11[11] , \wPDiag_11[10] , 
        \wPDiag_11[9] , \wPDiag_11[8] , \wPDiag_11[7] , \wPDiag_11[6] , 
        \wPDiag_11[5] , \wPDiag_11[4] , \wPDiag_11[3] , \wPDiag_11[2] , 
        \wPDiag_11[1] , \wPDiag_11[0] }), .NDiagOut({\wNDiag_11[15] , 
        \wNDiag_11[14] , \wNDiag_11[13] , \wNDiag_11[12] , \wNDiag_11[11] , 
        \wNDiag_11[10] , \wNDiag_11[9] , \wNDiag_11[8] , \wNDiag_11[7] , 
        \wNDiag_11[6] , \wNDiag_11[5] , \wNDiag_11[4] , \wNDiag_11[3] , 
        \wNDiag_11[2] , \wNDiag_11[1] , \wNDiag_11[0] }) );
    NQueens_Control_IDWIDTH5_SCAN1 U_NQueens_Control ( .Clk(Clk), .Reset(Reset
        ), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\wScan_0[4] , \wScan_0[3] , \wScan_0[2] , \wScan_0[1] , 
        \wScan_0[0] }), .ScanOut({\wScan_16[4] , \wScan_16[3] , \wScan_16[2] , 
        \wScan_16[1] , \wScan_16[0] }), .ScanEnable(\wScanEnable[0] ), .Id({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .ScanId({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}
        ), .CallIn(\wCall_16[0] ), .ReturnIn(\wReturn_0[0] ), .CallOut(
        \wCall_0[0] ) );
endmodule

