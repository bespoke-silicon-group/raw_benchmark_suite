
module NORMALIZE_SIZE16_DW01_dec_16_0 ( A, SUM );
input  [15:0] A;
output [15:0] SUM;
    wire n5, n20, n15, n9, n7, n12, n13, n6, n21, n8, n14, n23, n16, n11, n24, 
        n18, n10, n19, n25, n22, n17;
    VMW_AO21 U3 ( .A(n5), .B(A[9]), .C(n6), .Z(SUM[9]) );
    VMW_OAI21 U5 ( .A(n7), .B(n8), .C(n9), .Z(SUM[6]) );
    VMW_AO21 U6 ( .A(A[0]), .B(A[1]), .C(n10), .Z(SUM[1]) );
    VMW_OAI21 U14 ( .A(n20), .B(n21), .C(n16), .Z(SUM[12]) );
    VMW_NAND2 U21 ( .A(n13), .B(n14), .Z(n15) );
    VMW_NOR2 U28 ( .A(n23), .B(A[11]), .Z(n20) );
    VMW_INV U33 ( .A(n25), .Z(n17) );
    VMW_OAI21 U7 ( .A(n10), .B(n11), .C(n12), .Z(SUM[2]) );
    VMW_OAI21 U8 ( .A(n13), .B(n14), .C(n15), .Z(SUM[4]) );
    VMW_AO21 U13 ( .A(n12), .B(A[3]), .C(n13), .Z(SUM[3]) );
    VMW_INV U34 ( .A(A[6]), .Z(n8) );
    VMW_NOR2 U26 ( .A(n5), .B(A[9]), .Z(n6) );
    VMW_AO21 U9 ( .A(n15), .B(A[5]), .C(n7), .Z(SUM[5]) );
    VMW_AO21 U12 ( .A(n9), .B(A[7]), .C(n18), .Z(SUM[7]) );
    VMW_INV U35 ( .A(A[2]), .Z(n11) );
    VMW_NAND2 U27 ( .A(n22), .B(n6), .Z(n23) );
    VMW_NOR2 U20 ( .A(n12), .B(A[3]), .Z(n13) );
    VMW_NAND2 U29 ( .A(n21), .B(n20), .Z(n16) );
    VMW_OAI21 U15 ( .A(n6), .B(n22), .C(n23), .Z(SUM[10]) );
    VMW_NOR2 U17 ( .A(A[14]), .B(n25), .Z(n24) );
    VMW_NOR2 U22 ( .A(n15), .B(A[5]), .Z(n7) );
    VMW_MUX2I U32 ( .A(n25), .B(n17), .S(A[14]), .Z(SUM[14]) );
    VMW_INV U39 ( .A(A[10]), .Z(n22) );
    VMW_OR2 U30 ( .A(n16), .B(A[13]), .Z(n25) );
    VMW_AO21 U10 ( .A(n16), .B(A[13]), .C(n17), .Z(SUM[13]) );
    VMW_OAI21 U11 ( .A(n18), .B(n19), .C(n5), .Z(SUM[8]) );
    VMW_NAND2 U19 ( .A(n10), .B(n11), .Z(n12) );
    VMW_NAND2 U25 ( .A(n18), .B(n19), .Z(n5) );
    VMW_INV U37 ( .A(A[8]), .Z(n19) );
    VMW_INV U36 ( .A(A[4]), .Z(n14) );
    VMW_INV U4 ( .A(A[0]), .Z(SUM[0]) );
    VMW_NOR2 U18 ( .A(A[1]), .B(A[0]), .Z(n10) );
    VMW_NAND2 U23 ( .A(n7), .B(n8), .Z(n9) );
    VMW_NOR2 U24 ( .A(A[7]), .B(n9), .Z(n18) );
    VMW_INV U38 ( .A(A[12]), .Z(n21) );
    VMW_AO21 U16 ( .A(n23), .B(A[11]), .C(n20), .Z(SUM[11]) );
    VMW_XOR2 U31 ( .A(A[15]), .B(n24), .Z(SUM[15]) );
endmodule


module NORMALIZE_SIZE16 ( a, b );
input  [16:0] a;
output [16:0] b;
    wire \b99[9] , n175, \b99[4] , \b99[6] , n169, n172, \b99[2] , n168, n173, 
        \b99[15] , \b99[11] , n174, \b99[13] , \b99[16] , \b99[10] , \b99[12] , 
        n171, \b99[14] , \b99[3] , n170, \b99[7] , \b99[5] , \b99[8] , 
        \b99[1] ;
    VMW_AND2 U22 ( .A(a[16]), .B(n168), .Z(b[16]) );
    VMW_AO22 U26 ( .A(a[7]), .B(n173), .C(\b99[8] ), .D(n174), .Z(b[7]) );
    VMW_AO22 U28 ( .A(a[5]), .B(n173), .C(\b99[6] ), .D(n174), .Z(b[5]) );
    VMW_AO22 U33 ( .A(a[15]), .B(n173), .C(\b99[16] ), .D(n174), .Z(b[15]) );
    VMW_AO22 U34 ( .A(a[14]), .B(n173), .C(\b99[15] ), .D(n174), .Z(b[14]) );
    VMW_NOR4 U41 ( .A(a[8]), .B(a[9]), .C(a[10]), .D(a[11]), .Z(n171) );
    VMW_INV U46 ( .A(n168), .Z(n175) );
    VMW_AO22 U27 ( .A(a[6]), .B(n173), .C(\b99[7] ), .D(n174), .Z(b[6]) );
    VMW_AO22 U35 ( .A(a[13]), .B(n173), .C(\b99[14] ), .D(n174), .Z(b[13]) );
    VMW_NOR4 U40 ( .A(a[12]), .B(a[13]), .C(a[14]), .D(a[15]), .Z(n172) );
    NORMALIZE_SIZE16_DW01_dec_16_0 sub_217 ( .A(a[15:0]), .SUM({\b99[16] , 
        \b99[15] , \b99[14] , \b99[13] , \b99[12] , \b99[11] , \b99[10] , 
        \b99[9] , \b99[8] , \b99[7] , \b99[6] , \b99[5] , \b99[4] , \b99[3] , 
        \b99[2] , \b99[1] }) );
    VMW_AO22 U29 ( .A(a[4]), .B(n173), .C(\b99[5] ), .D(n174), .Z(b[4]) );
    VMW_AO22 U32 ( .A(a[1]), .B(n173), .C(\b99[2] ), .D(n174), .Z(b[1]) );
    VMW_AO22 U39 ( .A(a[0]), .B(n173), .C(\b99[1] ), .D(n174), .Z(b[0]) );
    VMW_AND4 U23 ( .A(n169), .B(n170), .C(n171), .D(n172), .Z(n168) );
    VMW_AO22 U24 ( .A(a[9]), .B(n173), .C(\b99[10] ), .D(n174), .Z(b[9]) );
    VMW_AO22 U25 ( .A(a[8]), .B(n173), .C(\b99[9] ), .D(n174), .Z(b[8]) );
    VMW_AO22 U30 ( .A(a[3]), .B(n173), .C(\b99[4] ), .D(n174), .Z(b[3]) );
    VMW_AO22 U37 ( .A(a[11]), .B(n173), .C(\b99[12] ), .D(n174), .Z(b[11]) );
    VMW_NOR4 U42 ( .A(a[4]), .B(a[5]), .C(a[6]), .D(a[7]), .Z(n170) );
    VMW_INV U45 ( .A(n173), .Z(n174) );
    VMW_AO22 U36 ( .A(a[12]), .B(n173), .C(\b99[13] ), .D(n174), .Z(b[12]) );
    VMW_NOR4 U43 ( .A(a[0]), .B(a[1]), .C(a[2]), .D(a[3]), .Z(n169) );
    VMW_AO22 U31 ( .A(a[2]), .B(n173), .C(\b99[3] ), .D(n174), .Z(b[2]) );
    VMW_AO22 U38 ( .A(a[10]), .B(n173), .C(\b99[11] ), .D(n174), .Z(b[10]) );
    VMW_NAND2 U44 ( .A(a[16]), .B(n175), .Z(n173) );
endmodule


module ADD_NN_SIZE16_DW01_add_16_0 ( A, B, CI, SUM, CO );
input  [15:0] A;
input  [15:0] B;
output [15:0] SUM;
input  CI;
output CO;
    wire \carry[9] , \carry[4] , \carry[2] , \carry[6] , \carry[13] , 
        \carry[15] , \carry[11] , \carry[10] , \carry[14] , \carry[12] , 
        \carry[7] , \carry[3] , \carry[8] , \carry[1] , \carry[5] ;
    VMW_AND2 U1 ( .A(A[0]), .B(B[0]), .Z(\carry[1] ) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_8 ( .CI(\carry[8] ), .A(A[8]), .B(B[8]), .S(SUM[8]), .CO(
        \carry[9] ) );
    VMW_FADD U1_11 ( .CI(\carry[11] ), .A(A[11]), .B(B[11]), .S(SUM[11]), .CO(
        \carry[12] ) );
    VMW_XOR2 U2 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]), .CO(
        \carry[8] ) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_9 ( .CI(\carry[9] ), .A(A[9]), .B(B[9]), .S(SUM[9]), .CO(
        \carry[10] ) );
    VMW_FADD U1_10 ( .CI(\carry[10] ), .A(A[10]), .B(B[10]), .S(SUM[10]), .CO(
        \carry[11] ) );
    VMW_FADD U1_12 ( .CI(\carry[12] ), .A(A[12]), .B(B[12]), .S(SUM[12]), .CO(
        \carry[13] ) );
    VMW_FADD U1_15 ( .CI(\carry[15] ), .A(A[15]), .B(B[15]), .S(SUM[15]) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
    VMW_FADD U1_14 ( .CI(\carry[14] ), .A(A[14]), .B(B[14]), .S(SUM[14]), .CO(
        \carry[15] ) );
    VMW_FADD U1_13 ( .CI(\carry[13] ), .A(A[13]), .B(B[13]), .S(SUM[13]), .CO(
        \carry[14] ) );
endmodule


module ADD_NN_SIZE16 ( a, b, c );
input  [16:0] a;
input  [16:0] b;
output [16:0] c;
    wire \arr[16] , \arr[15] , \arr[11] , \arr[13] , \arr[12] , \arr[9] , 
        \arr[8] , \arr[7] , \arr[3] , \arr[5] , \arr[1] , \arr[6] , \arr[4] , 
        \arr[0] , n56, \arr[2] , n58, n59, \arr[14] , \arr[10] , n57;
    NORMALIZE_SIZE16 norm ( .a({\arr[16] , \arr[15] , \arr[14] , \arr[13] , 
        \arr[12] , \arr[11] , \arr[10] , \arr[9] , \arr[8] , \arr[7] , 
        \arr[6] , \arr[5] , \arr[4] , \arr[3] , \arr[2] , \arr[1] , \arr[0] }), 
        .b(c) );
    VMW_INV U6 ( .A(n58), .Z(n57) );
    ADD_NN_SIZE16_DW01_add_16_0 add_234 ( .A(a[15:0]), .B(b[15:0]), .CI(n59), 
        .SUM({\arr[15] , \arr[14] , \arr[13] , \arr[12] , \arr[11] , \arr[10] , 
        \arr[9] , \arr[8] , \arr[7] , \arr[6] , \arr[5] , \arr[4] , \arr[3] , 
        \arr[2] , \arr[1] , \arr[0] }) );
    VMW_PULLDOWN U2 ( .Z(n59) );
    VMW_INV U5 ( .A(\arr[15] ), .Z(n56) );
    VMW_AO21 U3 ( .A(n56), .B(b[15]), .C(n57), .Z(\arr[16] ) );
    VMW_OAI21 U4 ( .A(b[15]), .B(n56), .C(a[15]), .Z(n58) );
endmodule


module ADD_MINUS_1_SIZE16_DW01_dec_16_0 ( A, SUM );
input  [15:0] A;
output [15:0] SUM;
    wire n5, n20, n15, n9, n7, n12, n13, n6, n21, n8, n14, n23, n16, n11, n24, 
        n18, n10, n19, n25, n22, n17;
    VMW_AO21 U3 ( .A(n5), .B(A[9]), .C(n6), .Z(SUM[9]) );
    VMW_OAI21 U5 ( .A(n7), .B(n8), .C(n9), .Z(SUM[6]) );
    VMW_AO21 U6 ( .A(A[0]), .B(A[1]), .C(n10), .Z(SUM[1]) );
    VMW_OAI21 U14 ( .A(n20), .B(n21), .C(n16), .Z(SUM[12]) );
    VMW_NAND2 U21 ( .A(n13), .B(n14), .Z(n15) );
    VMW_NOR2 U28 ( .A(n23), .B(A[11]), .Z(n20) );
    VMW_INV U33 ( .A(n25), .Z(n17) );
    VMW_OAI21 U7 ( .A(n10), .B(n11), .C(n12), .Z(SUM[2]) );
    VMW_OAI21 U8 ( .A(n13), .B(n14), .C(n15), .Z(SUM[4]) );
    VMW_AO21 U13 ( .A(n12), .B(A[3]), .C(n13), .Z(SUM[3]) );
    VMW_INV U34 ( .A(A[6]), .Z(n8) );
    VMW_NOR2 U26 ( .A(n5), .B(A[9]), .Z(n6) );
    VMW_AO21 U9 ( .A(n15), .B(A[5]), .C(n7), .Z(SUM[5]) );
    VMW_AO21 U12 ( .A(n9), .B(A[7]), .C(n18), .Z(SUM[7]) );
    VMW_INV U35 ( .A(A[2]), .Z(n11) );
    VMW_NAND2 U27 ( .A(n22), .B(n6), .Z(n23) );
    VMW_NOR2 U20 ( .A(n12), .B(A[3]), .Z(n13) );
    VMW_NAND2 U29 ( .A(n21), .B(n20), .Z(n16) );
    VMW_OAI21 U15 ( .A(n6), .B(n22), .C(n23), .Z(SUM[10]) );
    VMW_NOR2 U17 ( .A(A[14]), .B(n25), .Z(n24) );
    VMW_NOR2 U22 ( .A(n15), .B(A[5]), .Z(n7) );
    VMW_MUX2I U32 ( .A(n25), .B(n17), .S(A[14]), .Z(SUM[14]) );
    VMW_INV U39 ( .A(A[10]), .Z(n22) );
    VMW_OR2 U30 ( .A(n16), .B(A[13]), .Z(n25) );
    VMW_AO21 U10 ( .A(n16), .B(A[13]), .C(n17), .Z(SUM[13]) );
    VMW_OAI21 U11 ( .A(n18), .B(n19), .C(n5), .Z(SUM[8]) );
    VMW_NAND2 U19 ( .A(n10), .B(n11), .Z(n12) );
    VMW_NAND2 U25 ( .A(n18), .B(n19), .Z(n5) );
    VMW_INV U37 ( .A(A[8]), .Z(n19) );
    VMW_INV U36 ( .A(A[4]), .Z(n14) );
    VMW_INV U4 ( .A(A[0]), .Z(SUM[0]) );
    VMW_NOR2 U18 ( .A(A[1]), .B(A[0]), .Z(n10) );
    VMW_NAND2 U23 ( .A(n7), .B(n8), .Z(n9) );
    VMW_NOR2 U24 ( .A(A[7]), .B(n9), .Z(n18) );
    VMW_INV U38 ( .A(A[12]), .Z(n21) );
    VMW_AO21 U16 ( .A(n23), .B(A[11]), .C(n20), .Z(SUM[11]) );
    VMW_XOR2 U31 ( .A(A[15]), .B(n24), .Z(SUM[15]) );
endmodule


module ADD_MINUS_1_SIZE16 ( a, b );
input  [16:0] a;
output [16:0] b;
    wire n150, n151, n152, n153, \c82[7] , \c82[3] , \c82[1] , \c82[8] , 
        \c82[5] , \c82[12] , \c82[16] , \c82[14] , \c82[10] , \c82[15] , 
        \c82[11] , \c82[13] , \c82[4] , \c82[9] , \c82[2] , \c82[6] ;
    VMW_AND4 U20 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(b[16]) );
    VMW_OR2 U21 ( .A(\c82[16] ), .B(a[16]), .Z(b[15]) );
    VMW_OR2 U26 ( .A(\c82[11] ), .B(a[16]), .Z(b[10]) );
    VMW_OR2 U28 ( .A(\c82[9] ), .B(a[16]), .Z(b[8]) );
    VMW_OR2 U33 ( .A(\c82[4] ), .B(a[16]), .Z(b[3]) );
    VMW_OR2 U34 ( .A(\c82[3] ), .B(a[16]), .Z(b[2]) );
    VMW_OR2 U27 ( .A(\c82[10] ), .B(a[16]), .Z(b[9]) );
    VMW_OR2 U35 ( .A(\c82[2] ), .B(a[16]), .Z(b[1]) );
    VMW_NOR4 U40 ( .A(a[3]), .B(a[2]), .C(a[1]), .D(a[0]), .Z(n150) );
    ADD_MINUS_1_SIZE16_DW01_dec_16_0 sub_199 ( .A(a[15:0]), .SUM({\c82[16] , 
        \c82[15] , \c82[14] , \c82[13] , \c82[12] , \c82[11] , \c82[10] , 
        \c82[9] , \c82[8] , \c82[7] , \c82[6] , \c82[5] , \c82[4] , \c82[3] , 
        \c82[2] , \c82[1] }) );
    VMW_OR2 U22 ( .A(\c82[15] ), .B(a[16]), .Z(b[14]) );
    VMW_OR2 U29 ( .A(\c82[8] ), .B(a[16]), .Z(b[7]) );
    VMW_OR2 U32 ( .A(\c82[5] ), .B(a[16]), .Z(b[4]) );
    VMW_NOR4 U39 ( .A(a[7]), .B(a[6]), .C(a[5]), .D(a[4]), .Z(n151) );
    VMW_OR2 U23 ( .A(\c82[14] ), .B(a[16]), .Z(b[13]) );
    VMW_OR2 U24 ( .A(\c82[13] ), .B(a[16]), .Z(b[12]) );
    VMW_OR2 U25 ( .A(\c82[12] ), .B(a[16]), .Z(b[11]) );
    VMW_OR2 U30 ( .A(\c82[7] ), .B(a[16]), .Z(b[6]) );
    VMW_NOR5 U37 ( .A(a[13]), .B(a[12]), .C(a[14]), .D(a[16]), .E(a[15]), .Z(
        n153) );
    VMW_OR2 U36 ( .A(\c82[1] ), .B(a[16]), .Z(b[0]) );
    VMW_OR2 U31 ( .A(\c82[6] ), .B(a[16]), .Z(b[5]) );
    VMW_NOR4 U38 ( .A(a[11]), .B(a[10]), .C(a[9]), .D(a[8]), .Z(n152) );
endmodule


module ADD_SIZE16 ( a, b, c );
input  [16:0] a;
input  [16:0] b;
output [16:0] c;
    wire \sum1[6] , n97, \sum2[5] , \sum3[13] , \sum2[14] , n100, \sum2[8] , 
        \sum2[10] , \sum1[2] , \sum2[1] , \sum1[0] , \sum2[12] , \sum2[3] , 
        n99, \sum1[9] , \sum3[11] , \sum1[4] , \sum2[16] , \sum2[7] , n107, 
        \sum3[15] , n90, \sum1[13] , n98, \sum3[3] , \sum3[7] , n91, n106, 
        \sum1[15] , \sum3[5] , n96, n101, \sum1[11] , \sum3[8] , \sum3[1] , 
        \sum1[16] , \sum1[14] , \sum1[10] , \sum3[9] , n94, \sum3[4] , 
        \sum3[0] , n103, \sum3[6] , \sum1[12] , n104, \sum3[2] , n93, 
        \sum1[5] , \sum3[14] , \sum2[6] , \sum1[1] , \sum2[2] , \sum2[13] , 
        n92, n89, \sum1[8] , \sum3[10] , n105, \sum3[12] , n102, \sum2[9] , 
        \sum2[11] , n95, \sum1[3] , \sum2[0] , \sum1[7] , \sum3[16] , 
        \sum2[4] , \sum2[15] ;
    ADD_NN_SIZE16 add_nn ( .a(a), .b(b), .c({\sum1[16] , \sum1[15] , 
        \sum1[14] , \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , 
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    ADD_MINUS_1_SIZE16 am2 ( .a(b), .b({\sum3[16] , \sum3[15] , \sum3[14] , 
        \sum3[13] , \sum3[12] , \sum3[11] , \sum3[10] , \sum3[9] , \sum3[8] , 
        \sum3[7] , \sum3[6] , \sum3[5] , \sum3[4] , \sum3[3] , \sum3[2] , 
        \sum3[1] , \sum3[0] }) );
    VMW_AO21 U20 ( .A(\sum1[13] ), .B(n89), .C(n93), .Z(c[13]) );
    VMW_AO21 U21 ( .A(\sum1[12] ), .B(n89), .C(n94), .Z(c[12]) );
    VMW_AO21 U26 ( .A(\sum1[7] ), .B(n89), .C(n99), .Z(c[7]) );
    VMW_AO21 U28 ( .A(\sum1[5] ), .B(n89), .C(n101), .Z(c[5]) );
    VMW_AO21 U33 ( .A(\sum1[0] ), .B(n89), .C(n106), .Z(c[0]) );
    VMW_NOR2 U34 ( .A(n89), .B(a[16]), .Z(n107) );
    VMW_AO22 U41 ( .A(\sum3[4] ), .B(a[16]), .C(\sum2[4] ), .D(n107), .Z(n102)
         );
    VMW_AO22 U46 ( .A(\sum3[15] ), .B(a[16]), .C(\sum2[15] ), .D(n107), .Z(n91
        ) );
    VMW_AO22 U48 ( .A(\sum3[13] ), .B(a[16]), .C(\sum2[13] ), .D(n107), .Z(n93
        ) );
    VMW_AO21 U27 ( .A(\sum1[6] ), .B(n89), .C(n100), .Z(c[6]) );
    VMW_NOR2 U35 ( .A(a[16]), .B(b[16]), .Z(n89) );
    VMW_AO22 U40 ( .A(\sum3[5] ), .B(a[16]), .C(\sum2[5] ), .D(n107), .Z(n101)
         );
    VMW_AO22 U52 ( .A(\sum3[0] ), .B(a[16]), .C(\sum2[0] ), .D(n107), .Z(n106)
         );
    VMW_AO22 U49 ( .A(\sum3[12] ), .B(a[16]), .C(\sum2[12] ), .D(n107), .Z(n94
        ) );
    VMW_AO21 U29 ( .A(\sum1[4] ), .B(n89), .C(n102), .Z(c[4]) );
    VMW_AO22 U47 ( .A(\sum3[14] ), .B(a[16]), .C(\sum2[14] ), .D(n107), .Z(n92
        ) );
    VMW_AO21 U17 ( .A(\sum1[16] ), .B(n89), .C(n90), .Z(c[16]) );
    VMW_AO21 U22 ( .A(\sum1[11] ), .B(n89), .C(n95), .Z(c[11]) );
    VMW_AO21 U32 ( .A(\sum1[1] ), .B(n89), .C(n105), .Z(c[1]) );
    VMW_AO22 U39 ( .A(\sum3[6] ), .B(a[16]), .C(\sum2[6] ), .D(n107), .Z(n100)
         );
    VMW_AO21 U30 ( .A(\sum1[3] ), .B(n89), .C(n103), .Z(c[3]) );
    VMW_AO21 U18 ( .A(\sum1[15] ), .B(n89), .C(n91), .Z(c[15]) );
    VMW_AO21 U19 ( .A(\sum1[14] ), .B(n89), .C(n92), .Z(c[14]) );
    VMW_AO21 U25 ( .A(\sum1[8] ), .B(n89), .C(n98), .Z(c[8]) );
    VMW_AO22 U37 ( .A(\sum3[8] ), .B(a[16]), .C(\sum2[8] ), .D(n107), .Z(n98)
         );
    VMW_AO22 U42 ( .A(\sum3[3] ), .B(a[16]), .C(\sum2[3] ), .D(n107), .Z(n103)
         );
    VMW_AO22 U45 ( .A(\sum3[16] ), .B(a[16]), .C(\sum2[16] ), .D(n107), .Z(n90
        ) );
    VMW_AO22 U36 ( .A(\sum3[9] ), .B(a[16]), .C(\sum2[9] ), .D(n107), .Z(n97)
         );
    VMW_AO22 U50 ( .A(\sum3[11] ), .B(a[16]), .C(\sum2[11] ), .D(n107), .Z(n95
        ) );
    VMW_AO22 U43 ( .A(\sum3[2] ), .B(a[16]), .C(\sum2[2] ), .D(n107), .Z(n104)
         );
    VMW_AO22 U51 ( .A(\sum3[10] ), .B(a[16]), .C(\sum2[10] ), .D(n107), .Z(n96
        ) );
    VMW_AO21 U23 ( .A(\sum1[10] ), .B(n89), .C(n96), .Z(c[10]) );
    VMW_AO21 U24 ( .A(n89), .B(\sum1[9] ), .C(n97), .Z(c[9]) );
    VMW_AO22 U38 ( .A(\sum3[7] ), .B(a[16]), .C(\sum2[7] ), .D(n107), .Z(n99)
         );
    ADD_MINUS_1_SIZE16 am1 ( .a(a), .b({\sum2[16] , \sum2[15] , \sum2[14] , 
        \sum2[13] , \sum2[12] , \sum2[11] , \sum2[10] , \sum2[9] , \sum2[8] , 
        \sum2[7] , \sum2[6] , \sum2[5] , \sum2[4] , \sum2[3] , \sum2[2] , 
        \sum2[1] , \sum2[0] }) );
    VMW_AO21 U31 ( .A(\sum1[2] ), .B(n89), .C(n104), .Z(c[2]) );
    VMW_AO22 U44 ( .A(\sum3[1] ), .B(a[16]), .C(\sum2[1] ), .D(n107), .Z(n105)
         );
endmodule


module NEGATE_SIZE16_DW01_sub_17_0 ( A, B, CI, DIFF, CO );
input  [16:0] A;
input  [16:0] B;
output [16:0] DIFF;
input  CI;
output CO;
    wire \carry[16] , \B_not[16] , \B_not[14] , \B_not[12] , \carry[9] , 
        \carry[4] , \B_not[3] , \B_not[10] , \B_not[7] , \B_not[5] , 
        \carry[2] , \B_not[8] , \carry[6] , \carry[13] , \carry[15] , 
        \carry[11] , \carry[14] , \carry[10] , \carry[12] , \B_not[15] , 
        \B_not[9] , \carry[7] , \B_not[13] , \B_not[11] , \B_not[4] , 
        \carry[3] , \carry[8] , \B_not[6] , \carry[5] , \B_not[2] ;
    VMW_XNOR2 U3 ( .A(\carry[16] ), .B(\B_not[16] ), .Z(DIFF[16]) );
    VMW_XOR2 U5 ( .A(\carry[15] ), .B(\B_not[15] ), .Z(DIFF[15]) );
    VMW_AND2 U6 ( .A(\carry[14] ), .B(\B_not[14] ), .Z(\carry[15] ) );
    VMW_AND2 U14 ( .A(\carry[10] ), .B(\B_not[10] ), .Z(\carry[11] ) );
    VMW_XOR2 U21 ( .A(\carry[7] ), .B(\B_not[7] ), .Z(DIFF[7]) );
    VMW_AND2 U28 ( .A(\carry[3] ), .B(\B_not[3] ), .Z(\carry[4] ) );
    VMW_INV U33 ( .A(B[13]), .Z(\B_not[13] ) );
    VMW_XOR2 U7 ( .A(\carry[14] ), .B(\B_not[14] ), .Z(DIFF[14]) );
    VMW_AND2 U8 ( .A(\carry[13] ), .B(\B_not[13] ), .Z(\carry[14] ) );
    VMW_XOR2 U13 ( .A(\carry[11] ), .B(\B_not[11] ), .Z(DIFF[11]) );
    VMW_INV U34 ( .A(B[14]), .Z(\B_not[14] ) );
    VMW_INV U41 ( .A(B[9]), .Z(\B_not[9] ) );
    VMW_INV U46 ( .A(B[16]), .Z(\B_not[16] ) );
    VMW_AND2 U26 ( .A(\carry[4] ), .B(\B_not[4] ), .Z(\carry[5] ) );
    VMW_INV U48 ( .A(B[8]), .Z(\B_not[8] ) );
    VMW_XOR2 U9 ( .A(\carry[13] ), .B(\B_not[13] ), .Z(DIFF[13]) );
    VMW_AND2 U12 ( .A(\carry[11] ), .B(\B_not[11] ), .Z(\carry[12] ) );
    VMW_INV U35 ( .A(B[4]), .Z(\B_not[4] ) );
    VMW_XOR2 U27 ( .A(\carry[4] ), .B(\B_not[4] ), .Z(DIFF[4]) );
    VMW_INV U40 ( .A(B[10]), .Z(\B_not[10] ) );
    VMW_AND2 U20 ( .A(\carry[7] ), .B(\B_not[7] ), .Z(\carry[8] ) );
    VMW_INV U49 ( .A(B[1]), .Z(\carry[2] ) );
    VMW_XOR2 U29 ( .A(\carry[3] ), .B(\B_not[3] ), .Z(DIFF[3]) );
    VMW_INV U47 ( .A(B[11]), .Z(\B_not[11] ) );
    VMW_XOR2 U15 ( .A(\carry[10] ), .B(\B_not[10] ), .Z(DIFF[10]) );
    VMW_XOR2 U17 ( .A(\carry[9] ), .B(\B_not[9] ), .Z(DIFF[9]) );
    VMW_AND2 U22 ( .A(\carry[6] ), .B(\B_not[6] ), .Z(\carry[7] ) );
    VMW_INV U32 ( .A(\carry[2] ), .Z(DIFF[1]) );
    VMW_INV U39 ( .A(B[12]), .Z(\B_not[12] ) );
    VMW_AND2 U30 ( .A(\carry[2] ), .B(\B_not[2] ), .Z(\carry[3] ) );
    VMW_AND2 U10 ( .A(\carry[12] ), .B(\B_not[12] ), .Z(\carry[13] ) );
    VMW_INV U42 ( .A(B[2]), .Z(\B_not[2] ) );
    VMW_INV U45 ( .A(B[0]), .Z(DIFF[0]) );
    VMW_XOR2 U11 ( .A(\carry[12] ), .B(\B_not[12] ), .Z(DIFF[12]) );
    VMW_XOR2 U19 ( .A(\carry[8] ), .B(\B_not[8] ), .Z(DIFF[8]) );
    VMW_XOR2 U25 ( .A(\carry[5] ), .B(\B_not[5] ), .Z(DIFF[5]) );
    VMW_INV U37 ( .A(B[5]), .Z(\B_not[5] ) );
    VMW_INV U36 ( .A(B[3]), .Z(\B_not[3] ) );
    VMW_AND2 U4 ( .A(\carry[15] ), .B(\B_not[15] ), .Z(\carry[16] ) );
    VMW_AND2 U18 ( .A(\carry[8] ), .B(\B_not[8] ), .Z(\carry[9] ) );
    VMW_INV U43 ( .A(B[7]), .Z(\B_not[7] ) );
    VMW_XOR2 U23 ( .A(\carry[6] ), .B(\B_not[6] ), .Z(DIFF[6]) );
    VMW_AND2 U24 ( .A(\carry[5] ), .B(\B_not[5] ), .Z(\carry[6] ) );
    VMW_INV U38 ( .A(B[15]), .Z(\B_not[15] ) );
    VMW_INV U44 ( .A(B[6]), .Z(\B_not[6] ) );
    VMW_AND2 U16 ( .A(\carry[9] ), .B(\B_not[9] ), .Z(\carry[10] ) );
    VMW_XOR2 U31 ( .A(\carry[2] ), .B(\B_not[2] ), .Z(DIFF[2]) );
endmodule


module NEGATE_SIZE16 ( a, b );
input  [16:0] a;
output [16:0] b;
    wire n330, \c260[9] , \ozzo[1] , \ozzo[0] , n322, \c260[4] , n323, n325, 
        \c260[6] , \c260[2] , \c260[16] , \c260[12] , n324, \c260[10] , 
        \c260[14] , \c260[17] , \c260[15] , \c260[13] , \c260[11] , n328, n326, 
        \c260[3] , n327, \c260[7] , n329, \c260[5] , \c260[8] , \c260[1] ;
    VMW_PULLDOWN U83 ( .Z(n330) );
    VMW_PULLDOWN U84 ( .Z(\ozzo[1] ) );
    VMW_AND2 U96 ( .A(\c260[7] ), .B(n322), .Z(b[6]) );
    VMW_NOR3 U108 ( .A(a[1]), .B(a[3]), .C(a[2]), .Z(n325) );
    NEGATE_SIZE16_DW01_sub_17_0 sub_276 ( .A({\ozzo[0] , \ozzo[1] , \ozzo[1] , 
        \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[1] , 
        \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[1] , 
        \ozzo[1] , \ozzo[0] }), .B(a), .CI(n330), .DIFF({\c260[17] , 
        \c260[16] , \c260[15] , \c260[14] , \c260[13] , \c260[12] , \c260[11] , 
        \c260[10] , \c260[9] , \c260[8] , \c260[7] , \c260[6] , \c260[5] , 
        \c260[4] , \c260[3] , \c260[2] , \c260[1] }) );
    VMW_AND2 U101 ( .A(\c260[2] ), .B(n322), .Z(b[1]) );
    VMW_NOR4 U106 ( .A(a[9]), .B(a[10]), .C(a[11]), .D(a[12]), .Z(n327) );
    VMW_PULLUP U85 ( .Z(\ozzo[0] ) );
    VMW_AND2 U90 ( .A(\c260[13] ), .B(n322), .Z(b[12]) );
    VMW_AND2 U91 ( .A(\c260[12] ), .B(n322), .Z(b[11]) );
    VMW_AND2 U98 ( .A(\c260[5] ), .B(n322), .Z(b[4]) );
    VMW_AND2 U99 ( .A(\c260[4] ), .B(n322), .Z(b[3]) );
    VMW_NOR4 U107 ( .A(a[13]), .B(a[15]), .C(a[14]), .D(a[4]), .Z(n326) );
    VMW_AND2 U97 ( .A(\c260[6] ), .B(n322), .Z(b[5]) );
    VMW_NOR2 U109 ( .A(a[16]), .B(n324), .Z(n323) );
    VMW_AND2 U100 ( .A(\c260[3] ), .B(n322), .Z(b[2]) );
    VMW_AO22 U86 ( .A(\c260[17] ), .B(n322), .C(n323), .D(a[0]), .Z(b[16]) );
    VMW_AND2 U87 ( .A(\c260[16] ), .B(n322), .Z(b[15]) );
    VMW_AND2 U95 ( .A(\c260[8] ), .B(n322), .Z(b[7]) );
    VMW_INV U110 ( .A(n324), .Z(n329) );
    VMW_AND2 U88 ( .A(\c260[15] ), .B(n322), .Z(b[14]) );
    VMW_AND2 U89 ( .A(\c260[14] ), .B(n322), .Z(b[13]) );
    VMW_AO21 U102 ( .A(\c260[1] ), .B(n324), .C(a[16]), .Z(b[0]) );
    VMW_NOR4 U105 ( .A(a[5]), .B(a[6]), .C(a[7]), .D(a[8]), .Z(n328) );
    VMW_AND2 U92 ( .A(\c260[11] ), .B(n322), .Z(b[10]) );
    VMW_AND2 U93 ( .A(\c260[10] ), .B(n322), .Z(b[9]) );
    VMW_NOR2 U104 ( .A(a[16]), .B(n329), .Z(n322) );
    VMW_AND2 U94 ( .A(\c260[9] ), .B(n322), .Z(b[8]) );
    VMW_NAND4 U103 ( .A(n325), .B(n326), .C(n327), .D(n328), .Z(n324) );
endmodule


module SHIFT_UP_SIZE16_s33 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , \nb2[1] , \sum1[0] , 
        \nb2[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \sum1[14] , 
        \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , \sum1[5] , \nb2[6] , 
        \sum1[1] , \nb2[15] , \nb2[11] , \nb2[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \nb2[4] , \nb2[0] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), 
        .c({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , \sum1[12] , 
        \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , \sum1[6] , 
        \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U9 ( .Z(Logic0) );
endmodule


module COMBINATIONAL_SIZE16_s33 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \a[1]1 , \a[2]1 , \t1[2] , \t1[15] , \t2[5] , \t1[6] , \b[4] , 
        \t2[1] , \t1[13] , \b[0] , \b[9] , \t2[8] , \t1[11] , \t1[9] , \b[2] , 
        \b[6] , \a[3]1 , \t2[3] , \t1[0] , \a[16]1 , \t2[7] , \t1[4] , 
        \t2[12] , \b[10] , \a[13]1 , \a[12]1 , \a[6]1 , \b[14] , \t2[16] , 
        \b[16] , \a[7]1 , \t2[14] , \b[12] , \t2[10] , \a[11]1 , \a[10]1 , 
        \a[9]1 , \a[8]1 , \b[13] , \t2[11] , \a[4]1 , \t2[15] , \a[5]1 , 
        \b[15] , \b[11] , \t2[13] , \b[7] , \t1[16] , \t2[6] , \t1[5] , 
        \t2[0] , \b[3] , \t1[8] , \t1[12] , \t2[2] , \t1[1] , \t1[3] , 
        \t1[10] , \b[8] , \b[1] , \t2[9] , \b[5] , \a[15]1 , \t2[4] , \t1[7] , 
        \a[14]1 , \a[0]1 , \t1[14] ;
    assign \a[16]1  = a[16];
    assign \a[15]1  = a[15];
    assign \a[14]1  = a[14];
    assign \a[13]1  = a[13];
    assign \a[12]1  = a[12];
    assign \a[11]1  = a[11];
    assign \a[10]1  = a[10];
    assign \a[9]1  = a[9];
    assign \a[8]1  = a[8];
    assign \a[7]1  = a[7];
    assign \a[6]1  = a[6];
    assign \a[5]1  = a[5];
    assign \a[4]1  = a[4];
    assign \a[3]1  = a[3];
    assign \a[2]1  = a[2];
    assign \a[1]1  = a[1];
    assign \a[0]1  = a[0];
    assign \b[16]  = b[16];
    assign \b[15]  = b[15];
    assign \b[14]  = b[14];
    assign \b[13]  = b[13];
    assign \b[12]  = b[12];
    assign \b[11]  = b[11];
    assign \b[10]  = b[10];
    assign \b[9]  = b[9];
    assign \b[8]  = b[8];
    assign \b[7]  = b[7];
    assign \b[6]  = b[6];
    assign \b[5]  = b[5];
    assign \b[4]  = b[4];
    assign \b[3]  = b[3];
    assign \b[2]  = b[2];
    assign \b[1]  = b[1];
    assign \b[0]  = b[0];
    assign x[16] = \a[16]1 ;
    assign x[15] = \a[15]1 ;
    assign x[14] = \a[14]1 ;
    assign x[13] = \a[13]1 ;
    assign x[12] = \a[12]1 ;
    assign x[11] = \a[11]1 ;
    assign x[10] = \a[10]1 ;
    assign x[9] = \a[9]1 ;
    assign x[8] = \a[8]1 ;
    assign x[7] = \a[7]1 ;
    assign x[6] = \a[6]1 ;
    assign x[5] = \a[5]1 ;
    assign x[4] = \a[4]1 ;
    assign x[3] = \a[3]1 ;
    assign x[2] = \a[2]1 ;
    assign x[1] = \a[1]1 ;
    assign x[0] = \a[0]1 ;
    assign y[16] = \b[16] ;
    assign y[15] = \b[15] ;
    assign y[14] = \b[14] ;
    assign y[13] = \b[13] ;
    assign y[12] = \b[12] ;
    assign y[11] = \b[11] ;
    assign y[10] = \b[10] ;
    assign y[9] = \b[9] ;
    assign y[8] = \b[8] ;
    assign y[7] = \b[7] ;
    assign y[6] = \b[6] ;
    assign y[5] = \b[5] ;
    assign y[4] = \b[4] ;
    assign y[3] = \b[3] ;
    assign y[2] = \b[2] ;
    assign y[1] = \b[1] ;
    assign y[0] = \b[0] ;
    ADD_SIZE16 add2 ( .a({\a[16]1 , \a[15]1 , \a[14]1 , \a[13]1 , \a[12]1 , 
        \a[11]1 , \a[10]1 , \a[9]1 , \a[8]1 , \a[7]1 , \a[6]1 , \a[5]1 , 
        \a[4]1 , \a[3]1 , \a[2]1 , \a[1]1 , \a[0]1 }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    ADD_SIZE16 add1 ( .a({\a[16]1 , \a[15]1 , \a[14]1 , \a[13]1 , \a[12]1 , 
        \a[11]1 , \a[10]1 , \a[9]1 , \a[8]1 , \a[7]1 , \a[6]1 , \a[5]1 , 
        \a[4]1 , \a[3]1 , \a[2]1 , \a[1]1 , \a[0]1 }), .b({\t1[16] , \t1[15] , 
        \t1[14] , \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , 
        \t1[7] , \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] 
        }) );
    SHIFT_UP_SIZE16_s33 shift ( .a({\b[16] , \b[15] , \b[14] , \b[13] , 
        \b[12] , \b[11] , \b[10] , \b[9] , \b[8] , \b[7] , \b[6] , \b[5] , 
        \b[4] , \b[3] , \b[2] , \b[1] , \b[0] }), .c({\t1[16] , \t1[15] , 
        \t1[14] , \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , 
        \t1[7] , \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] 
        }) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s33 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s0 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \a[16] , \a[15] , \a[13] , \a[7] , \sum1[6] , \nb2[16] , \b1[16] , 
        \b1[5] , \nb2[5] , \nb2[12] , \nb2[8] , \b1[12] , \b1[1] , \a[11] , 
        \a[3] , \b1[8] , \a[1] , \sum1[2] , \nb2[1] , \sum1[0] , \nb2[3] , 
        \b1[10] , \b1[3] , \a[8] , \a[5] , \sum1[9] , \nb2[10] , \nb2[7] , 
        \sum1[4] , \nb2[14] , \b1[14] , \a[14] , \a[4] , \b1[7] , \sum1[13] , 
        \sum1[15] , \sum1[11] , \sum1[10] , \sum1[14] , \sum1[16] , \sum1[12] , 
        \sum1[5] , \nb2[6] , \nb2[15] , \b1[15] , \b1[6] , \a[12] , \a[10] , 
        \a[0] , \sum1[1] , \nb2[2] , \b1[11] , \a[9] , \b1[2] , \sum1[8] , 
        \nb2[11] , \nb2[13] , \nb2[9] , \b1[13] , \a[2] , Logic01, \b1[9] , 
        \b1[0] , n150, \nb2[0] , \sum1[3] , \b1[4] , \a[6] , \nb2[4] , 
        \sum1[7] ;
    assign \a[16]  = a[16];
    assign \a[15]  = a[15];
    assign \a[14]  = a[14];
    assign \a[13]  = a[13];
    assign \a[12]  = a[12];
    assign \a[11]  = a[11];
    assign \a[10]  = a[10];
    assign \a[9]  = a[9];
    assign \a[8]  = a[8];
    assign \a[7]  = a[7];
    assign \a[6]  = a[6];
    assign \a[5]  = a[5];
    assign \a[4]  = a[4];
    assign \a[3]  = a[3];
    assign \a[2]  = a[2];
    assign \a[1]  = a[1];
    assign \a[0]  = a[0];
    assign c[16] = \a[16] ;
    assign c[15] = \a[15] ;
    assign c[14] = \a[14] ;
    assign c[13] = \a[13] ;
    assign c[12] = \a[12] ;
    assign c[11] = \a[11] ;
    assign c[10] = \a[10] ;
    assign c[9] = \a[9] ;
    assign c[8] = \a[8] ;
    assign c[7] = \a[7] ;
    assign c[6] = \a[6] ;
    assign c[5] = \a[5] ;
    assign c[4] = \a[4] ;
    assign c[3] = \a[3] ;
    assign c[2] = \a[2] ;
    assign c[1] = \a[1] ;
    assign c[0] = \a[0] ;
    VMW_AND2 U21 ( .A(\a[9] ), .B(n150), .Z(\b1[9] ) );
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, 
        Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, 
        Logic01, Logic01, Logic01}) );
    VMW_PULLDOWN U13 ( .Z(Logic01) );
    VMW_PULLDOWN U14 ( .Z(\b1[16] ) );
    VMW_AND2 U28 ( .A(\a[2] ), .B(n150), .Z(\b1[2] ) );
    VMW_AND2 U26 ( .A(\a[4] ), .B(n150), .Z(\b1[4] ) );
    VMW_AND2 U15 ( .A(\a[15] ), .B(n150), .Z(\b1[15] ) );
    VMW_AND2 U20 ( .A(\a[10] ), .B(n150), .Z(\b1[10] ) );
    VMW_AND2 U27 ( .A(\a[3] ), .B(n150), .Z(\b1[3] ) );
    VMW_AND2 U29 ( .A(\a[1] ), .B(n150), .Z(\b1[1] ) );
    NEGATE_SIZE16 negate ( .a({Logic01, Logic01, Logic01, Logic01, Logic01, 
        Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, 
        Logic01, Logic01, Logic01, Logic01}), .b({\nb2[16] , \nb2[15] , 
        \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , 
        \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , 
        \nb2[1] , \nb2[0] }) );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_AND2 U17 ( .A(\a[13] ), .B(n150), .Z(\b1[13] ) );
    VMW_AND2 U22 ( .A(\a[8] ), .B(n150), .Z(\b1[8] ) );
    VMW_AND2 U30 ( .A(\a[0] ), .B(n150), .Z(\b1[0] ) );
    VMW_AND2 U25 ( .A(\a[5] ), .B(n150), .Z(\b1[5] ) );
    VMW_AND2 U16 ( .A(\a[14] ), .B(n150), .Z(\b1[14] ) );
    VMW_AND2 U18 ( .A(\a[12] ), .B(n150), .Z(\b1[12] ) );
    VMW_AND2 U19 ( .A(\a[11] ), .B(n150), .Z(\b1[11] ) );
    VMW_AND2 U23 ( .A(\a[7] ), .B(n150), .Z(\b1[7] ) );
    VMW_AND2 U24 ( .A(\a[6] ), .B(n150), .Z(\b1[6] ) );
    VMW_INV U31 ( .A(\a[16] ), .Z(n150) );
endmodule


module COMBINATIONAL_SIZE16_s0 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s0 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, n509, 
        n468, \comleft[4] , \comright[11] , n454, n473, n483, \outleft[11] , 
        \comleft[0] , \comright[15] , \comright[3] , n528, \comleft[12] , 
        \comleft[9] , n461, n533, n514, n484, n534, n513, \outleft[13] , 
        \comright[8] , n466, \comleft[10] , \comright[1] , n541, \comleft[2] , 
        n508, n498, \outleft[9] , \comleft[6] , n474, \comleft[14] , 
        \comright[13] , \comright[5] , n453, n526, n491, n501, n499, n540, 
        \outleft[6] , \outleft[4] , \outleft[0] , n467, \ScanReg[2] , 
        \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, \ScanReg[4] , 
        \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, \outleft[2] , 
        n455, n472, n507, n497, n520, n532, n515, n485, n460, \ScanReg[9] , 
        \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , \outleft[7] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s0 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s8 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , n158, \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[5] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n158), .Z(\b1[10] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n158), .Z(\b1[12] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U20 ( .Z(Logic0) );
    VMW_AND2 U27 ( .A(a[3]), .B(n158), .Z(\b1[11] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n158), .Z(\b1[9] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[7] ) );
    VMW_PULLDOWN U22 ( .Z(\b1[16] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n158), .Z(\b1[8] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n158), .Z(\b1[13] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[3] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[1] ) );
    VMW_AND2 U23 ( .A(a[7]), .B(n158), .Z(\b1[15] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n158), .Z(\b1[14] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n158) );
endmodule


module COMBINATIONAL_SIZE16_s8 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s8 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, n516, n486, \comleft[5] , n463, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s8 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s4 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        n154, \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[2] ) );
    VMW_AND2 U21 ( .A(a[9]), .B(n154), .Z(\b1[13] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n154), .Z(\b1[6] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n154), .Z(\b1[8] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[3] ) );
    VMW_AND2 U20 ( .A(a[10]), .B(n154), .Z(\b1[14] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n154), .Z(\b1[7] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n154), .Z(\b1[5] ) );
    VMW_PULLDOWN U17 ( .Z(Logic0) );
    VMW_AND2 U22 ( .A(a[8]), .B(n154), .Z(\b1[12] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n154), .Z(\b1[4] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n154), .Z(\b1[9] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[1] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[16] ) );
    VMW_AND2 U19 ( .A(a[11]), .B(n154), .Z(\b1[15] ) );
    VMW_AND2 U23 ( .A(a[7]), .B(n154), .Z(\b1[11] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n154), .Z(\b1[10] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n154) );
endmodule


module COMBINATIONAL_SIZE16_s4 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s4 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s4_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s4 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s12 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , \sum1[5] , 
        \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , n162, \nb2[11] , 
        \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , \nb2[13] , \nb2[9] , 
        \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[9] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[3] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n162), .Z(\b1[14] ) );
    VMW_PULLDOWN U26 ( .Z(\b1[16] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[10] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n162), .Z(\b1[15] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n162), .Z(\b1[13] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[11] ) );
    VMW_PULLDOWN U22 ( .Z(\b1[8] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n162), .Z(\b1[12] ) );
    VMW_PULLDOWN U25 ( .Z(\b1[5] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[7] ) );
    VMW_PULLDOWN U23 ( .Z(\b1[1] ) );
    VMW_PULLDOWN U24 ( .Z(Logic0) );
    VMW_INV U31 ( .A(a[16]), .Z(n162) );
endmodule


module COMBINATIONAL_SIZE16_s12 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s12 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s12_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , n461, \comleft[9] , n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s12 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s2 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , n152, \sum1[2] , Logic0, \nb2[5] , \nb2[12] , 
        \nb2[8] , \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , 
        \b1[10] , \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , 
        \b1[7] , \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[1] ) );
    VMW_AND2 U21 ( .A(a[9]), .B(n152), .Z(\b1[11] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n152), .Z(\b1[4] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n152), .Z(\b1[6] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(Logic0) );
    VMW_AND2 U20 ( .A(a[10]), .B(n152), .Z(\b1[12] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n152), .Z(\b1[5] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n152), .Z(\b1[3] ) );
    VMW_AND2 U17 ( .A(a[13]), .B(n152), .Z(\b1[15] ) );
    VMW_AND2 U22 ( .A(a[8]), .B(n152), .Z(\b1[10] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n152), .Z(\b1[2] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n152), .Z(\b1[7] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[16] ) );
    VMW_AND2 U18 ( .A(a[12]), .B(n152), .Z(\b1[14] ) );
    VMW_AND2 U19 ( .A(a[11]), .B(n152), .Z(\b1[13] ) );
    VMW_AND2 U23 ( .A(a[7]), .B(n152), .Z(\b1[9] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n152), .Z(\b1[8] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n152) );
endmodule


module COMBINATIONAL_SIZE16_s2 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s2 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s2_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[4] , \outleft[0] , n467, \ScanReg[2] , 
        \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, \outleft[6] , 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s2 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s6 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , \sum1[5] , 
        \nb2[6] , n156, \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , \nb2[11] , 
        \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , \nb2[13] , \nb2[9] , 
        \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_AND2 U21 ( .A(a[9]), .B(n156), .Z(\b1[15] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n156), .Z(\b1[8] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n156), .Z(\b1[10] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[16] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n156), .Z(\b1[9] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n156), .Z(\b1[7] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[1] ) );
    VMW_AND2 U22 ( .A(a[8]), .B(n156), .Z(\b1[14] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n156), .Z(\b1[6] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n156), .Z(\b1[11] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[3] ) );
    VMW_PULLDOWN U18 ( .Z(Logic0) );
    VMW_PULLDOWN U19 ( .Z(\b1[5] ) );
    VMW_AND2 U23 ( .A(a[7]), .B(n156), .Z(\b1[13] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n156), .Z(\b1[12] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n156) );
endmodule


module COMBINATIONAL_SIZE16_s6 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s6 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s6_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s6 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s10 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , n160, \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , 
        \b1[7] , \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[9] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[1] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n160), .Z(\b1[12] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n160), .Z(\b1[14] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[8] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n160), .Z(\b1[13] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n160), .Z(\b1[11] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U22 ( .Z(Logic0) );
    VMW_AND2 U30 ( .A(a[0]), .B(n160), .Z(\b1[10] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n160), .Z(\b1[15] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[7] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[3] ) );
    VMW_PULLDOWN U23 ( .Z(\b1[5] ) );
    VMW_PULLDOWN U24 ( .Z(\b1[16] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n160) );
endmodule


module COMBINATIONAL_SIZE16_s10 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s10 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s10_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[0] , n467, \ScanReg[2] , \ScanReg[15] , n535, 
        n512, n482, n527, n500, n490, n475, \outleft[6] , \outleft[4] , 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s10 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s14 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , n164, \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[9] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[10] ) );
    VMW_PULLDOWN U28 ( .Z(\b1[16] ) );
    VMW_PULLDOWN U26 ( .Z(Logic0) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[7] ) );
    VMW_PULLDOWN U27 ( .Z(\b1[5] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n164), .Z(\b1[15] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U22 ( .Z(\b1[3] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n164), .Z(\b1[14] ) );
    VMW_PULLDOWN U25 ( .Z(\b1[1] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[13] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[11] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U23 ( .Z(\b1[8] ) );
    VMW_PULLDOWN U24 ( .Z(\b1[12] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n164) );
endmodule


module COMBINATIONAL_SIZE16_s14 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s14 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s14_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s14 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s1 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , n151, \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U14 ( .Z(Logic0) );
    VMW_AND2 U21 ( .A(a[9]), .B(n151), .Z(\b1[10] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n151), .Z(\b1[3] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n151), .Z(\b1[5] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[16] ) );
    VMW_AND2 U20 ( .A(a[10]), .B(n151), .Z(\b1[11] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n151), .Z(\b1[4] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n151), .Z(\b1[2] ) );
    VMW_AND2 U17 ( .A(a[13]), .B(n151), .Z(\b1[14] ) );
    VMW_AND2 U22 ( .A(a[8]), .B(n151), .Z(\b1[9] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n151), .Z(\b1[1] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n151), .Z(\b1[6] ) );
    VMW_AND2 U16 ( .A(a[14]), .B(n151), .Z(\b1[15] ) );
    VMW_AND2 U18 ( .A(a[12]), .B(n151), .Z(\b1[13] ) );
    VMW_AND2 U19 ( .A(a[11]), .B(n151), .Z(\b1[12] ) );
    VMW_AND2 U23 ( .A(a[7]), .B(n151), .Z(\b1[8] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n151), .Z(\b1[7] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n151) );
endmodule


module COMBINATIONAL_SIZE16_s1 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s1 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , n519, n489, \outleft[1] , 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s1 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s3 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        n153, \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[2] ) );
    VMW_AND2 U21 ( .A(a[9]), .B(n153), .Z(\b1[12] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n153), .Z(\b1[5] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n153), .Z(\b1[7] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[1] ) );
    VMW_AND2 U20 ( .A(a[10]), .B(n153), .Z(\b1[13] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n153), .Z(\b1[6] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n153), .Z(\b1[4] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[16] ) );
    VMW_AND2 U22 ( .A(a[8]), .B(n153), .Z(\b1[11] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n153), .Z(\b1[3] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n153), .Z(\b1[8] ) );
    VMW_PULLDOWN U16 ( .Z(Logic0) );
    VMW_AND2 U18 ( .A(a[12]), .B(n153), .Z(\b1[15] ) );
    VMW_AND2 U19 ( .A(a[11]), .B(n153), .Z(\b1[14] ) );
    VMW_AND2 U23 ( .A(a[7]), .B(n153), .Z(\b1[10] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n153), .Z(\b1[9] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n153) );
endmodule


module COMBINATIONAL_SIZE16_s3 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s3 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s3_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s3 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s5 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , n155, 
        \b1[7] , \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_AND2 U21 ( .A(a[9]), .B(n155), .Z(\b1[14] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n155), .Z(\b1[7] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n155), .Z(\b1[9] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[2] ) );
    VMW_AND2 U20 ( .A(a[10]), .B(n155), .Z(\b1[15] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n155), .Z(\b1[8] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n155), .Z(\b1[6] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[1] ) );
    VMW_AND2 U22 ( .A(a[8]), .B(n155), .Z(\b1[13] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n155), .Z(\b1[5] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n155), .Z(\b1[10] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[3] ) );
    VMW_PULLDOWN U18 ( .Z(Logic0) );
    VMW_PULLDOWN U19 ( .Z(\b1[16] ) );
    VMW_AND2 U23 ( .A(a[7]), .B(n155), .Z(\b1[12] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n155), .Z(\b1[11] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n155) );
endmodule


module COMBINATIONAL_SIZE16_s5 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s5 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s5_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s5 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s7 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , \sum1[5] , 
        \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , \nb2[11] , \nb2[2] , 
        \b1[11] , n157, \b1[2] , \sum1[7] , \sum1[3] , \nb2[13] , \nb2[9] , 
        \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[16] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n157), .Z(\b1[9] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n157), .Z(\b1[11] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[5] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n157), .Z(\b1[10] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n157), .Z(\b1[8] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[3] ) );
    VMW_AND2 U22 ( .A(a[8]), .B(n157), .Z(\b1[15] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n157), .Z(\b1[7] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n157), .Z(\b1[12] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[1] ) );
    VMW_PULLDOWN U19 ( .Z(Logic0) );
    VMW_AND2 U23 ( .A(a[7]), .B(n157), .Z(\b1[14] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n157), .Z(\b1[13] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n157) );
endmodule


module COMBINATIONAL_SIZE16_s7 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s7 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s7_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s7 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s9 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , \sum1[5] , 
        \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , \nb2[11] , \nb2[2] , 
        \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , \nb2[13] , \nb2[9] , \b1[13] , 
        \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , \b1[4] , n159;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U21 ( .Z(Logic0) );
    VMW_AND2 U28 ( .A(a[2]), .B(n159), .Z(\b1[11] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n159), .Z(\b1[13] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[1] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n159), .Z(\b1[12] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n159), .Z(\b1[10] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[7] ) );
    VMW_PULLDOWN U22 ( .Z(\b1[5] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n159), .Z(\b1[9] ) );
    VMW_AND2 U25 ( .A(a[5]), .B(n159), .Z(\b1[14] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[3] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[8] ) );
    VMW_PULLDOWN U23 ( .Z(\b1[16] ) );
    VMW_AND2 U24 ( .A(a[6]), .B(n159), .Z(\b1[15] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n159) );
endmodule


module COMBINATIONAL_SIZE16_s9 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s9 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s9_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, \comleft[4] , \comright[11] , n454, n468, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s9 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s11 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        n161, \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[9] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[8] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n161), .Z(\b1[13] ) );
    VMW_AND2 U26 ( .A(a[4]), .B(n161), .Z(\b1[15] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[3] ) );
    VMW_AND2 U27 ( .A(a[3]), .B(n161), .Z(\b1[14] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n161), .Z(\b1[12] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U22 ( .Z(\b1[1] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n161), .Z(\b1[11] ) );
    VMW_PULLDOWN U25 ( .Z(\b1[16] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[7] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[10] ) );
    VMW_PULLDOWN U23 ( .Z(Logic0) );
    VMW_PULLDOWN U24 ( .Z(\b1[5] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n161) );
endmodule


module COMBINATIONAL_SIZE16_s11 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s11 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s11_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[4] , \outleft[0] , n467, \ScanReg[2] , 
        \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, \ScanReg[4] , 
        \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, \outleft[6] , n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s11 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s13 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , n163, \sum1[8] , 
        \sum1[5] , \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , 
        \nb2[11] , \nb2[2] , \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , 
        \nb2[13] , \nb2[9] , \b1[13] , \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , 
        \b1[4] ;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[9] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[3] ) );
    VMW_AND2 U28 ( .A(a[2]), .B(n163), .Z(\b1[15] ) );
    VMW_PULLDOWN U26 ( .Z(\b1[5] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[10] ) );
    VMW_PULLDOWN U27 ( .Z(\b1[16] ) );
    VMW_AND2 U29 ( .A(a[1]), .B(n163), .Z(\b1[14] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[11] ) );
    VMW_PULLDOWN U22 ( .Z(\b1[8] ) );
    VMW_AND2 U30 ( .A(a[0]), .B(n163), .Z(\b1[13] ) );
    VMW_PULLDOWN U25 ( .Z(Logic0) );
    VMW_PULLDOWN U16 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[7] ) );
    VMW_PULLDOWN U23 ( .Z(\b1[12] ) );
    VMW_PULLDOWN U24 ( .Z(\b1[1] ) );
    VMW_INV U31 ( .A(a[16]), .Z(n163) );
endmodule


module COMBINATIONAL_SIZE16_s13 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s13 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s13_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \comright[8] , n466, \outleft[13] , \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, \outleft[6] , \outleft[4] , \outleft[0] , n467, 
        \ScanReg[2] , \ScanReg[15] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s13 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE16_s15 ( a, c );
input  [16:0] a;
output [16:0] c;
    wire \sum1[16] , \sum1[15] , \sum1[13] , \sum1[9] , \sum1[6] , \nb2[16] , 
        \b1[16] , \b1[5] , \sum1[2] , Logic0, \nb2[5] , \nb2[12] , \nb2[8] , 
        \nb2[1] , \b1[12] , \b1[1] , \b1[8] , \sum1[0] , \nb2[3] , \b1[10] , 
        \b1[3] , \sum1[4] , \nb2[10] , \nb2[14] , \nb2[7] , \b1[14] , \b1[7] , 
        \sum1[14] , \sum1[11] , \sum1[10] , \sum1[12] , \sum1[8] , \sum1[5] , 
        \nb2[6] , \sum1[1] , \nb2[15] , \b1[15] , \b1[6] , \nb2[11] , \nb2[2] , 
        \b1[11] , \b1[2] , \sum1[7] , \sum1[3] , \nb2[13] , \nb2[9] , \b1[13] , 
        \b1[9] , \b1[0] , \nb2[4] , \nb2[0] , \b1[4] , n165;
    ADD_SIZE16 add2 ( .a({\sum1[16] , \sum1[15] , \sum1[14] , \sum1[13] , 
        \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , \sum1[7] , 
        \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , 
        \sum1[0] }), .b({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[14] ) );
    VMW_PULLDOWN U28 ( .Z(\b1[5] ) );
    VMW_PULLDOWN U26 ( .Z(\b1[1] ) );
    NEGATE_SIZE16 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0}), .b({\nb2[16] , \nb2[15] , \nb2[14] , \nb2[13] , 
        \nb2[12] , \nb2[11] , \nb2[10] , \nb2[9] , \nb2[8] , \nb2[7] , 
        \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] })
         );
    ADD_SIZE16 add1 ( .a({\b1[16] , \b1[15] , \b1[14] , \b1[13] , \b1[12] , 
        \b1[11] , \b1[10] , \b1[9] , \b1[8] , \b1[7] , \b1[6] , \b1[5] , 
        \b1[4] , \b1[3] , \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[16] , 
        \nb2[15] , \nb2[14] , \nb2[13] , \nb2[12] , \nb2[11] , \nb2[10] , 
        \nb2[9] , \nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , \nb2[4] , \nb2[3] , 
        \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[16] , \sum1[15] , \sum1[14] , 
        \sum1[13] , \sum1[12] , \sum1[11] , \sum1[10] , \sum1[9] , \sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[9] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[7] ) );
    VMW_PULLDOWN U27 ( .Z(Logic0) );
    VMW_PULLDOWN U29 ( .Z(\b1[16] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U22 ( .Z(\b1[10] ) );
    VMW_NOR2 U30 ( .A(n165), .B(a[16]), .Z(\b1[15] ) );
    VMW_PULLDOWN U25 ( .Z(\b1[12] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[13] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[11] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U23 ( .Z(\b1[3] ) );
    VMW_PULLDOWN U24 ( .Z(\b1[8] ) );
    VMW_INV U31 ( .A(a[0]), .Z(n165) );
endmodule


module COMBINATIONAL_SIZE16_s15 ( a, b, x, y );
input  [16:0] a;
output [16:0] y;
input  [16:0] b;
output [16:0] x;
    wire \t2[5] , \t4[14] , \t1[6] , \t4[2] , \t1[15] , \t2[1] , \t4[10] , 
        \t1[2] , \t2[8] , \t4[6] , \t1[11] , \t4[4] , \t1[9] , \t1[13] , 
        \t2[3] , \t1[0] , \t4[12] , \t2[7] , \t4[9] , \t4[0] , \t1[4] , 
        \t2[16] , \t2[12] , \t3[3] , \t3[11] , \t2[15] , \t2[14] , \t3[15] , 
        \t3[7] , \t3[5] , \t2[11] , \t2[10] , \t3[13] , \t3[1] , \t3[12] , 
        \t3[8] , \t3[0] , \t3[9] , \t3[4] , \t2[13] , \t3[14] , \t3[6] , 
        \t3[10] , \t3[2] , n138, \t2[6] , \t4[1] , \t1[16] , \t1[5] , \t4[8] , 
        \t4[5] , \t1[8] , \t1[12] , \t2[2] , \t4[13] , \t2[0] , \t4[11] , 
        \t1[1] , \t1[3] , \t1[10] , \t2[9] , \t4[7] , \t2[4] , \t4[15] , 
        \t1[7] , \t4[3] , \t1[14] , n137;
    ADD_SIZE16 add2 ( .a(a), .b({\t2[16] , \t2[15] , \t2[14] , \t2[13] , 
        \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[16], 
        \t4[15] , \t4[14] , \t4[13] , \t4[12] , \t4[11] , \t4[10] , \t4[9] , 
        \t4[8] , \t4[7] , \t4[6] , \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , 
        \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[14] ), .B(n137), .Z(x[14]) );
    VMW_AND2 U26 ( .A(\t3[9] ), .B(n137), .Z(x[9]) );
    VMW_AND2 U28 ( .A(\t3[7] ), .B(n137), .Z(x[7]) );
    VMW_AND2 U33 ( .A(\t3[2] ), .B(n137), .Z(x[2]) );
    VMW_AND2 U34 ( .A(\t3[1] ), .B(n137), .Z(x[1]) );
    VMW_AND2 U41 ( .A(\t4[10] ), .B(n138), .Z(y[10]) );
    VMW_AND2 U46 ( .A(\t4[5] ), .B(n138), .Z(y[5]) );
    VMW_AND2 U48 ( .A(\t4[3] ), .B(n138), .Z(y[3]) );
    ADD_SIZE16 add1 ( .a(a), .b({\t1[16] , \t1[15] , \t1[14] , \t1[13] , 
        \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[16], 
        \t3[15] , \t3[14] , \t3[13] , \t3[12] , \t3[11] , \t3[10] , \t3[9] , 
        \t3[8] , \t3[7] , \t3[6] , \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , 
        \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[15] ), .B(n137), .Z(x[15]) );
    VMW_AND2 U27 ( .A(\t3[8] ), .B(n137), .Z(x[8]) );
    VMW_AND2 U35 ( .A(\t3[0] ), .B(n137), .Z(x[0]) );
    VMW_INV U53 ( .A(x[16]), .Z(n137) );
    VMW_AND2 U40 ( .A(\t4[11] ), .B(n138), .Z(y[11]) );
    VMW_INV U52 ( .A(y[16]), .Z(n138) );
    VMW_AND2 U49 ( .A(\t4[2] ), .B(n138), .Z(y[2]) );
    VMW_AND2 U22 ( .A(\t3[13] ), .B(n137), .Z(x[13]) );
    VMW_AND2 U29 ( .A(\t3[6] ), .B(n137), .Z(x[6]) );
    VMW_AND2 U47 ( .A(\t4[4] ), .B(n138), .Z(y[4]) );
    VMW_AND2 U32 ( .A(\t3[3] ), .B(n137), .Z(x[3]) );
    VMW_AND2 U39 ( .A(\t4[12] ), .B(n138), .Z(y[12]) );
    VMW_AND2 U30 ( .A(\t3[5] ), .B(n137), .Z(x[5]) );
    VMW_AND2 U37 ( .A(\t4[14] ), .B(n138), .Z(y[14]) );
    VMW_AND2 U42 ( .A(\t4[9] ), .B(n138), .Z(y[9]) );
    VMW_AND2 U45 ( .A(\t4[6] ), .B(n138), .Z(y[6]) );
    SHIFT_UP_SIZE16_s15 shift ( .a(b), .c({\t1[16] , \t1[15] , \t1[14] , 
        \t1[13] , \t1[12] , \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , 
        \t1[6] , \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[10] ), .B(n137), .Z(x[10]) );
    VMW_AND2 U36 ( .A(\t4[15] ), .B(n138), .Z(y[15]) );
    VMW_AND2 U50 ( .A(\t4[1] ), .B(n138), .Z(y[1]) );
    NEGATE_SIZE16 neg ( .a({\t1[16] , \t1[15] , \t1[14] , \t1[13] , \t1[12] , 
        \t1[11] , \t1[10] , \t1[9] , \t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[16] , \t2[15] , 
        \t2[14] , \t2[13] , \t2[12] , \t2[11] , \t2[10] , \t2[9] , \t2[8] , 
        \t2[7] , \t2[6] , \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] 
        }) );
    VMW_AND2 U23 ( .A(\t3[12] ), .B(n137), .Z(x[12]) );
    VMW_AND2 U24 ( .A(\t3[11] ), .B(n137), .Z(x[11]) );
    VMW_AND2 U43 ( .A(\t4[8] ), .B(n138), .Z(y[8]) );
    VMW_AND2 U51 ( .A(\t4[0] ), .B(n138), .Z(y[0]) );
    VMW_AND2 U31 ( .A(\t3[4] ), .B(n137), .Z(x[4]) );
    VMW_AND2 U38 ( .A(\t4[13] ), .B(n138), .Z(y[13]) );
    VMW_AND2 U44 ( .A(\t4[7] ), .B(n138), .Z(y[7]) );
endmodule


module FFT_Node_SIZE16_IDWIDTH1_s15_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [16:0] outleft;
input  [15:0] ScanIn;
input  [0:0] Idr;
input  [16:0] inleft;
input  [16:0] inright;
output [15:0] ScanOut;
output [16:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[15] , \comleft[16] , \comright[7] , n506, n496, n521, 
        \outleft[7] , n509, n468, \comleft[4] , \comright[11] , n454, n473, 
        n483, \outleft[11] , \comleft[0] , \comright[15] , \comright[3] , n528, 
        \comleft[12] , \comleft[9] , n461, n533, n514, n484, n534, n513, 
        \outleft[13] , \comright[8] , n466, \comleft[10] , \comright[1] , n541, 
        \comleft[2] , n508, n498, \outleft[9] , \comleft[6] , n474, 
        \comleft[14] , \comright[13] , \comright[5] , n453, n526, n491, n501, 
        n499, n540, n467, \ScanReg[15] , \outleft[6] , \outleft[4] , 
        \outleft[0] , \ScanReg[2] , n535, n512, n482, n527, n500, n490, n475, 
        \ScanReg[4] , \ScanReg[6] , \ScanReg[11] , \ScanReg[13] , n469, n529, 
        \outleft[2] , n455, n472, n507, n497, n520, n532, n515, n485, n460, 
        \ScanReg[9] , \outleft[3] , n522, n505, n495, n457, n470, \ScanReg[8] , 
        \ScanReg[5] , n539, \ScanReg[12] , n479, \outleft[8] , \outleft[5] , 
        n537, n462, n530, n517, n487, n480, n510, n465, n459, n542, 
        \ScanReg[7] , \ScanReg[10] , \comright[14] , \outleft[1] , n519, n489, 
        \ScanReg[3] , \ScanReg[14] , n477, n502, n492, n525, n458, n503, 
        \comleft[7] , n464, \comright[12] , \comleft[15] , \comright[4] , n511, 
        n481, n536, n493, \outleft[12] , \comright[9] , n524, \comright[0] , 
        n476, \comleft[11] , \comleft[3] , \comright[16] , n518, n488, 
        \comleft[1] , n523, \outleft[10] , \comleft[13] , \comright[2] , n538, 
        n471, n456, \outleft[14] , \comleft[8] , n504, \comright[6] , n531, 
        n494, \comleft[5] , n463, n516, n486, \comright[10] , n478;
    assign ScanOut[15] = \outleft[15] ;
    assign ScanOut[14] = \outleft[14] ;
    assign ScanOut[13] = \outleft[13] ;
    assign ScanOut[12] = \outleft[12] ;
    assign ScanOut[11] = \outleft[11] ;
    assign ScanOut[10] = \outleft[10] ;
    assign ScanOut[9] = \outleft[9] ;
    assign ScanOut[8] = \outleft[8] ;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[15] = \outleft[15] ;
    assign outleft[14] = \outleft[14] ;
    assign outleft[13] = \outleft[13] ;
    assign outleft[12] = \outleft[12] ;
    assign outleft[11] = \outleft[11] ;
    assign outleft[10] = \outleft[10] ;
    assign outleft[9] = \outleft[9] ;
    assign outleft[8] = \outleft[8] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n453), .C(\ScanReg[3] ), .D(n454), .Z(
        n541) );
    VMW_AO21 U73 ( .A(outright[6]), .B(n455), .C(n462), .Z(n522) );
    VMW_AO22 U113 ( .A(\ScanReg[3] ), .B(n494), .C(\comright[3] ), .D(n492), 
        .Z(n459) );
    VMW_AO22 U134 ( .A(outright[15]), .B(n494), .C(\comleft[15] ), .D(n492), 
        .Z(n488) );
    VMW_AO21 U68 ( .A(outright[1]), .B(n455), .C(n457), .Z(n527) );
    VMW_AO21 U96 ( .A(\outleft[12] ), .B(n455), .C(n485), .Z(n499) );
    VMW_FD \outright_reg[0]  ( .D(n528), .CP(Clk), .Q(outright[0]) );
    VMW_AO22 U108 ( .A(\ScanReg[8] ), .B(n494), .C(\comright[8] ), .D(n492), 
        .Z(n464) );
    VMW_INV U141 ( .A(ScanEnable), .Z(n493) );
    VMW_FD \outleft_reg[4]  ( .D(n507), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n539), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \outright_reg[9]  ( .D(n519), .CP(Clk), .Q(outright[9]) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n453), .C(\ScanReg[2] ), .D(n454), .Z(
        n542) );
    VMW_AO22 U61 ( .A(ScanIn[10]), .B(n453), .C(\ScanReg[10] ), .D(n454), .Z(
        n534) );
    VMW_AO21 U84 ( .A(\outleft[0] ), .B(n455), .C(n473), .Z(n511) );
    VMW_FD \outleft_reg[9]  ( .D(n502), .CP(Clk), .Q(\outleft[9] ) );
    VMW_FD \outright_reg[4]  ( .D(n524), .CP(Clk), .Q(outright[4]) );
    VMW_FD \ScanReg_reg[8]  ( .D(n536), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \outleft_reg[0]  ( .D(n511), .CP(Clk), .Q(\outleft[0] ) );
    VMW_AO22 U66 ( .A(ScanIn[15]), .B(n453), .C(\ScanReg[15] ), .D(n454), .Z(
        n529) );
    VMW_OR2 U101 ( .A(ScanEnable), .B(Reset), .Z(n490) );
    VMW_NOR2 U106 ( .A(n493), .B(Reset), .Z(n453) );
    VMW_AO22 U121 ( .A(\ScanReg[11] ), .B(n494), .C(\comright[11] ), .D(n492), 
        .Z(n467) );
    VMW_AO22 U126 ( .A(outright[7]), .B(n494), .C(\comleft[7] ), .D(n492), .Z(
        n480) );
    VMW_AO21 U83 ( .A(outright[16]), .B(n455), .C(n472), .Z(n512) );
    VMW_AO21 U91 ( .A(\outleft[7] ), .B(n455), .C(n480), .Z(n504) );
    VMW_AO21 U98 ( .A(\outleft[14] ), .B(n455), .C(n487), .Z(n497) );
    VMW_FD \outleft_reg[2]  ( .D(n509), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n522), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n541), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(outright[5]), .B(n494), .C(\comleft[5] ), .D(n492), .Z(
        n478) );
    VMW_FD \outleft_reg[6]  ( .D(n505), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n537), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(outright[7]), .B(n455), .C(n463), .Z(n521) );
    VMW_AO22 U114 ( .A(\ScanReg[2] ), .B(n494), .C(\comright[2] ), .D(n492), 
        .Z(n458) );
    VMW_AO22 U133 ( .A(ScanIn[0]), .B(n494), .C(\comleft[16] ), .D(n492), .Z(
        n489) );
    VMW_AO21 U99 ( .A(\outleft[15] ), .B(n455), .C(n488), .Z(n496) );
    VMW_FD \outright_reg[2]  ( .D(n526), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n453), .C(\ScanReg[4] ), .D(n454), .Z(
        n540) );
    VMW_AO21 U67 ( .A(outright[0]), .B(n455), .C(n456), .Z(n528) );
    VMW_AO21 U82 ( .A(outright[15]), .B(n455), .C(n471), .Z(n513) );
    VMW_AO22 U107 ( .A(\ScanReg[9] ), .B(n494), .C(\comright[9] ), .D(n492), 
        .Z(n465) );
    VMW_AO22 U120 ( .A(\ScanReg[12] ), .B(n494), .C(\comright[12] ), .D(n492), 
        .Z(n468) );
    VMW_FD \outleft_reg[11]  ( .D(n500), .CP(Clk), .Q(\outleft[11] ) );
    VMW_AO21 U69 ( .A(outright[2]), .B(n455), .C(n458), .Z(n526) );
    VMW_AO21 U75 ( .A(outright[8]), .B(n455), .C(n464), .Z(n520) );
    VMW_AO22 U115 ( .A(outright[16]), .B(n494), .C(\comright[1] ), .D(n492), 
        .Z(n457) );
    VMW_AO22 U132 ( .A(outright[1]), .B(n494), .C(\comleft[1] ), .D(n492), .Z(
        n474) );
    VMW_FD \ScanReg_reg[14]  ( .D(n530), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO21 U90 ( .A(\outleft[6] ), .B(n455), .C(n479), .Z(n505) );
    VMW_AO22 U109 ( .A(\ScanReg[7] ), .B(n494), .C(\comright[7] ), .D(n492), 
        .Z(n463) );
    VMW_AO22 U129 ( .A(outright[4]), .B(n494), .C(\comleft[4] ), .D(n492), .Z(
        n477) );
    VMW_FD \outleft_reg[15]  ( .D(n496), .CP(Clk), .Q(\outleft[15] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(n534), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_FD \outright_reg[13]  ( .D(n515), .CP(Clk), .Q(outright[13]) );
    VMW_FD \outright_reg[11]  ( .D(n517), .CP(Clk), .Q(outright[11]) );
    VMW_AO21 U72 ( .A(outright[5]), .B(n455), .C(n461), .Z(n523) );
    VMW_AO21 U97 ( .A(\outleft[13] ), .B(n455), .C(n486), .Z(n498) );
    VMW_AO22 U140 ( .A(outright[0]), .B(n494), .C(\comleft[0] ), .D(n492), .Z(
        n473) );
    VMW_FD \ScanReg_reg[12]  ( .D(n532), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_AO22 U112 ( .A(\ScanReg[4] ), .B(n494), .C(\comright[4] ), .D(n492), 
        .Z(n460) );
    VMW_AO22 U135 ( .A(outright[14]), .B(n494), .C(\comleft[14] ), .D(n492), 
        .Z(n487) );
    VMW_AO22 U60 ( .A(ScanIn[9]), .B(n453), .C(\ScanReg[9] ), .D(n454), .Z(
        n535) );
    VMW_AO21 U85 ( .A(\outleft[1] ), .B(n455), .C(n474), .Z(n510) );
    VMW_AO21 U100 ( .A(outleft[16]), .B(n455), .C(n489), .Z(n495) );
    VMW_AO22 U127 ( .A(outright[6]), .B(n494), .C(\comleft[6] ), .D(n492), .Z(
        n479) );
    VMW_FD \outleft_reg[13]  ( .D(n498), .CP(Clk), .Q(\outleft[13] ) );
    VMW_FD \outright_reg[15]  ( .D(n513), .CP(Clk), .Q(outright[15]) );
    COMBINATIONAL_SIZE16_s15 com ( .a(inleft), .b(inright), .x({\comleft[16] , 
        \comleft[15] , \comleft[14] , \comleft[13] , \comleft[12] , 
        \comleft[11] , \comleft[10] , \comleft[9] , \comleft[8] , \comleft[7] , 
        \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , \comleft[2] , 
        \comleft[1] , \comleft[0] }), .y({\comright[16] , \comright[15] , 
        \comright[14] , \comright[13] , \comright[12] , \comright[11] , 
        \comright[10] , \comright[9] , \comright[8] , \comright[7] , 
        \comright[6] , \comright[5] , \comright[4] , \comright[3] , 
        \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n453), .C(\ScanReg[6] ), .D(n454), .Z(
        n538) );
    VMW_AO22 U137 ( .A(outright[12]), .B(n494), .C(\comleft[12] ), .D(n492), 
        .Z(n485) );
    VMW_AO22 U62 ( .A(ScanIn[11]), .B(n453), .C(\ScanReg[11] ), .D(n454), .Z(
        n533) );
    VMW_AO21 U70 ( .A(outright[3]), .B(n455), .C(n459), .Z(n525) );
    VMW_AO21 U79 ( .A(outright[12]), .B(n455), .C(n468), .Z(n516) );
    VMW_AO21 U95 ( .A(\outleft[11] ), .B(n455), .C(n484), .Z(n500) );
    VMW_AO22 U110 ( .A(\ScanReg[6] ), .B(n494), .C(\comright[6] ), .D(n492), 
        .Z(n462) );
    VMW_FD \outleft_reg[12]  ( .D(n499), .CP(Clk), .Q(\outleft[12] ) );
    VMW_FD \outright_reg[14]  ( .D(n514), .CP(Clk), .Q(outright[14]) );
    VMW_AO22 U119 ( .A(\ScanReg[13] ), .B(n494), .C(\comright[13] ), .D(n492), 
        .Z(n469) );
    VMW_INV U142 ( .A(n490), .Z(n454) );
    VMW_FD \outright_reg[10]  ( .D(n518), .CP(Clk), .Q(outright[10]) );
    VMW_AO21 U87 ( .A(\outleft[3] ), .B(n455), .C(n476), .Z(n508) );
    VMW_FD \outleft_reg[16]  ( .D(n495), .CP(Clk), .Q(outleft[16]) );
    VMW_FD \ScanReg_reg[13]  ( .D(n531), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(outright[8]), .B(n494), .C(\comleft[8] ), .D(n492), .Z(
        n481) );
    VMW_AO22 U65 ( .A(ScanIn[14]), .B(n453), .C(\ScanReg[14] ), .D(n454), .Z(
        n530) );
    VMW_NOR2 U102 ( .A(Reset), .B(n455), .Z(n491) );
    VMW_NOR2 U105 ( .A(Enable), .B(n490), .Z(n455) );
    VMW_AO22 U122 ( .A(\ScanReg[10] ), .B(n494), .C(\comright[10] ), .D(n492), 
        .Z(n466) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n453), .C(\ScanReg[5] ), .D(n454), .Z(
        n539) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n453), .C(\ScanReg[7] ), .D(n454), .Z(
        n537) );
    VMW_AO22 U59 ( .A(ScanIn[8]), .B(n453), .C(\ScanReg[8] ), .D(n454), .Z(
        n536) );
    VMW_AO21 U80 ( .A(outright[13]), .B(n455), .C(n469), .Z(n515) );
    VMW_AO22 U139 ( .A(outright[10]), .B(n494), .C(\comleft[10] ), .D(n492), 
        .Z(n483) );
    VMW_FD \outleft_reg[14]  ( .D(n497), .CP(Clk), .Q(\outleft[14] ) );
    VMW_FD \outright_reg[12]  ( .D(n516), .CP(Clk), .Q(outright[12]) );
    VMW_FD \ScanReg_reg[11]  ( .D(n533), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO21 U77 ( .A(outright[10]), .B(n455), .C(n466), .Z(n518) );
    VMW_AO21 U89 ( .A(\outleft[5] ), .B(n455), .C(n478), .Z(n506) );
    VMW_AO21 U92 ( .A(\outleft[8] ), .B(n455), .C(n481), .Z(n503) );
    VMW_FD \outright_reg[16]  ( .D(n512), .CP(Clk), .Q(outright[16]) );
    VMW_AO22 U117 ( .A(\ScanReg[15] ), .B(n494), .C(\comright[15] ), .D(n492), 
        .Z(n471) );
    VMW_FD \ScanReg_reg[15]  ( .D(n529), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(outright[3]), .B(n494), .C(\comleft[3] ), .D(n492), .Z(
        n476) );
    VMW_FD \outleft_reg[10]  ( .D(n501), .CP(Clk), .Q(\outleft[10] ) );
    VMW_AO22 U138 ( .A(outright[11]), .B(n494), .C(\comleft[11] ), .D(n492), 
        .Z(n484) );
    VMW_FD \outleft_reg[7]  ( .D(n504), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n538), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO22 U64 ( .A(ScanIn[13]), .B(n453), .C(\ScanReg[13] ), .D(n454), .Z(
        n531) );
    VMW_AO21 U81 ( .A(outright[14]), .B(n455), .C(n470), .Z(n514) );
    VMW_AND2 U104 ( .A(n491), .B(ScanEnable), .Z(n494) );
    VMW_AO21 U76 ( .A(outright[9]), .B(n455), .C(n465), .Z(n519) );
    VMW_AO22 U116 ( .A(ScanIn[1]), .B(n494), .C(\comright[16] ), .D(n492), .Z(
        n472) );
    VMW_AO22 U123 ( .A(outleft[16]), .B(n494), .C(\comright[0] ), .D(n492), 
        .Z(n456) );
    VMW_FD \outright_reg[3]  ( .D(n525), .CP(Clk), .Q(outright[3]) );
    VMW_AO21 U88 ( .A(\outleft[4] ), .B(n455), .C(n477), .Z(n507) );
    VMW_AO21 U93 ( .A(\outleft[9] ), .B(n455), .C(n482), .Z(n502) );
    VMW_AO22 U131 ( .A(outright[2]), .B(n494), .C(\comleft[2] ), .D(n492), .Z(
        n475) );
    VMW_FD \ScanReg_reg[2]  ( .D(n542), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n508), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO21 U94 ( .A(\outleft[10] ), .B(n455), .C(n483), .Z(n501) );
    VMW_FD \outleft_reg[8]  ( .D(n503), .CP(Clk), .Q(\outleft[8] ) );
    VMW_FD \outright_reg[7]  ( .D(n521), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n523), .CP(Clk), .Q(outright[5]) );
    VMW_FD \ScanReg_reg[9]  ( .D(n535), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(outright[13]), .B(n494), .C(\comleft[13] ), .D(n492), 
        .Z(n486) );
    VMW_FD \outleft_reg[1]  ( .D(n510), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO22 U63 ( .A(ScanIn[12]), .B(n453), .C(\ScanReg[12] ), .D(n454), .Z(
        n532) );
    VMW_AO21 U71 ( .A(outright[4]), .B(n455), .C(n460), .Z(n524) );
    VMW_AO22 U111 ( .A(\ScanReg[5] ), .B(n494), .C(\comright[5] ), .D(n492), 
        .Z(n461) );
    VMW_AO22 U124 ( .A(outright[9]), .B(n494), .C(\comleft[9] ), .D(n492), .Z(
        n482) );
    VMW_AO21 U78 ( .A(outright[11]), .B(n455), .C(n467), .Z(n517) );
    VMW_AO21 U86 ( .A(\outleft[2] ), .B(n455), .C(n475), .Z(n509) );
    VMW_AND2 U103 ( .A(n493), .B(n491), .Z(n492) );
    VMW_FD \outright_reg[1]  ( .D(n527), .CP(Clk), .Q(outright[1]) );
    VMW_AO22 U118 ( .A(\ScanReg[14] ), .B(n494), .C(\comright[14] ), .D(n492), 
        .Z(n470) );
    VMW_FD \outleft_reg[5]  ( .D(n506), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n540), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n520), .CP(Clk), .Q(outright[8]) );
endmodule


module FFT_Control_SIZE16_IDWIDTH1_SCAN1_DW01_dec_32_0 ( A, SUM );
input  [31:0] A;
output [31:0] SUM;
    wire n20, n15, n32, n29, n9, n47, n7, n12, n40, n35, n27, n49, n13, n34, 
        n41, n6, n26, n48, n21, n8, n46, n28, n33, n14, n38, n23, n16, n31, 
        n43, n44, n36, n11, n24, n18, n10, n37, n42, n5, n19, n25, n22, n39, 
        n45, n17, n30;
    VMW_INV U3 ( .A(A[0]), .Z(SUM[0]) );
    VMW_OAI21 U5 ( .A(n8), .B(n9), .C(n10), .Z(SUM[20]) );
    VMW_OAI21 U6 ( .A(n11), .B(n12), .C(n13), .Z(SUM[2]) );
    VMW_AO21 U14 ( .A(n25), .B(A[17]), .C(n14), .Z(SUM[17]) );
    VMW_AO21 U21 ( .A(n33), .B(A[29]), .C(n34), .Z(SUM[29]) );
    VMW_NOR2 U54 ( .A(n10), .B(A[21]), .Z(n41) );
    VMW_INV U73 ( .A(A[4]), .Z(n35) );
    VMW_INV U68 ( .A(A[2]), .Z(n12) );
    VMW_AO21 U28 ( .A(n36), .B(A[5]), .C(n43), .Z(SUM[5]) );
    VMW_NOR2 U33 ( .A(A[30]), .B(n49), .Z(n48) );
    VMW_OAI21 U7 ( .A(n14), .B(n15), .C(n16), .Z(SUM[18]) );
    VMW_AO21 U8 ( .A(n17), .B(A[25]), .C(n18), .Z(SUM[25]) );
    VMW_AO21 U13 ( .A(n13), .B(A[3]), .C(n24), .Z(SUM[3]) );
    VMW_NOR2 U34 ( .A(A[1]), .B(A[0]), .Z(n11) );
    VMW_NAND2 U41 ( .A(n39), .B(n46), .Z(n30) );
    VMW_NOR2 U46 ( .A(n7), .B(A[13]), .Z(n22) );
    VMW_NAND2 U61 ( .A(n47), .B(n45), .Z(n33) );
    VMW_INV U66 ( .A(A[12]), .Z(n6) );
    VMW_OAI21 U26 ( .A(n41), .B(n42), .C(n28), .Z(SUM[22]) );
    VMW_NOR2 U48 ( .A(n19), .B(A[15]), .Z(n20) );
    VMW_AO21 U9 ( .A(n19), .B(A[15]), .C(n20), .Z(SUM[15]) );
    VMW_AO21 U12 ( .A(A[0]), .B(A[1]), .C(n11), .Z(SUM[1]) );
    VMW_NAND2 U35 ( .A(n11), .B(n12), .Z(n13) );
    VMW_NAND2 U53 ( .A(n9), .B(n8), .Z(n10) );
    VMW_INV U74 ( .A(A[16]), .Z(n37) );
    VMW_AO21 U27 ( .A(n10), .B(A[21]), .C(n41), .Z(SUM[21]) );
    VMW_NOR2 U40 ( .A(A[7]), .B(n38), .Z(n39) );
    VMW_NOR2 U52 ( .A(n16), .B(A[19]), .Z(n8) );
    VMW_INV U67 ( .A(A[20]), .Z(n9) );
    VMW_INV U75 ( .A(A[10]), .Z(n40) );
    VMW_OAI21 U20 ( .A(n29), .B(n32), .C(n17), .Z(SUM[24]) );
    VMW_NAND2 U49 ( .A(n37), .B(n20), .Z(n25) );
    VMW_INV U69 ( .A(A[18]), .Z(n15) );
    VMW_OAI21 U29 ( .A(n43), .B(n44), .C(n38), .Z(SUM[6]) );
    VMW_NAND2 U47 ( .A(n23), .B(n22), .Z(n19) );
    VMW_NAND2 U55 ( .A(n42), .B(n41), .Z(n28) );
    VMW_INV U72 ( .A(A[24]), .Z(n32) );
    VMW_NOR2 U60 ( .A(n27), .B(A[27]), .Z(n45) );
    VMW_OAI21 U15 ( .A(n18), .B(n26), .C(n27), .Z(SUM[26]) );
    VMW_AO21 U17 ( .A(n28), .B(A[23]), .C(n29), .Z(SUM[23]) );
    VMW_OAI21 U22 ( .A(n24), .B(n35), .C(n36), .Z(SUM[4]) );
    VMW_OAI21 U32 ( .A(n45), .B(n47), .C(n33), .Z(SUM[28]) );
    VMW_NAND2 U39 ( .A(n43), .B(n44), .Z(n38) );
    VMW_NAND2 U57 ( .A(n32), .B(n29), .Z(n17) );
    VMW_INV U70 ( .A(A[14]), .Z(n23) );
    VMW_AO21 U30 ( .A(n27), .B(A[27]), .C(n45), .Z(SUM[27]) );
    VMW_INV U79 ( .A(A[28]), .Z(n47) );
    VMW_AO21 U10 ( .A(n21), .B(A[11]), .C(n5), .Z(SUM[11]) );
    VMW_NOR2 U42 ( .A(n30), .B(A[9]), .Z(n31) );
    VMW_NAND2 U45 ( .A(n6), .B(n5), .Z(n7) );
    VMW_OR2 U62 ( .A(n33), .B(A[29]), .Z(n49) );
    VMW_INV U65 ( .A(n49), .Z(n34) );
    VMW_OAI21 U11 ( .A(n22), .B(n23), .C(n19), .Z(SUM[14]) );
    VMW_AO21 U19 ( .A(n30), .B(A[9]), .C(n31), .Z(SUM[9]) );
    VMW_OAI21 U25 ( .A(n31), .B(n40), .C(n21), .Z(SUM[10]) );
    VMW_NAND2 U37 ( .A(n24), .B(n35), .Z(n36) );
    VMW_NAND2 U59 ( .A(n26), .B(n18), .Z(n27) );
    VMW_NOR2 U50 ( .A(n25), .B(A[17]), .Z(n14) );
    VMW_INV U77 ( .A(A[6]), .Z(n44) );
    VMW_NOR2 U58 ( .A(n17), .B(A[25]), .Z(n18) );
    VMW_NOR2 U36 ( .A(n13), .B(A[3]), .Z(n24) );
    VMW_OAI21 U4 ( .A(n5), .B(n6), .C(n7), .Z(SUM[12]) );
    VMW_AO21 U18 ( .A(n7), .B(A[13]), .C(n22), .Z(SUM[13]) );
    VMW_NAND2 U43 ( .A(n40), .B(n31), .Z(n21) );
    VMW_MUX2I U64 ( .A(n49), .B(n34), .S(A[30]), .Z(SUM[30]) );
    VMW_NAND2 U51 ( .A(n15), .B(n14), .Z(n16) );
    VMW_INV U76 ( .A(A[22]), .Z(n42) );
    VMW_OAI21 U23 ( .A(n20), .B(n37), .C(n25), .Z(SUM[16]) );
    VMW_AO21 U24 ( .A(n38), .B(A[7]), .C(n39), .Z(SUM[7]) );
    VMW_NOR2 U38 ( .A(n36), .B(A[5]), .Z(n43) );
    VMW_NOR2 U44 ( .A(n21), .B(A[11]), .Z(n5) );
    VMW_NOR2 U56 ( .A(n28), .B(A[23]), .Z(n29) );
    VMW_INV U71 ( .A(A[26]), .Z(n26) );
    VMW_XOR2 U63 ( .A(A[31]), .B(n48), .Z(SUM[31]) );
    VMW_AO21 U16 ( .A(n16), .B(A[19]), .C(n8), .Z(SUM[19]) );
    VMW_OAI21 U31 ( .A(n39), .B(n46), .C(n30), .Z(SUM[8]) );
    VMW_INV U78 ( .A(A[8]), .Z(n46) );
endmodule


module FFT_Control_SIZE16_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [15:0] ScanIn;
output [15:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire \DataIn[9] , \DataIn[4] , n317, \count241[28] , n330, \count[17] , 
        \count[24] , \count[2] , \DataIn[0] , n362, \count241[12] , 
        \count241[21] , n345, n370, n339, \count[20] , \count[6] , \count[13] , 
        n357, \count241[16] , \count241[25] , n295, n305, n322, \DataIn[6] , 
        \DataIn[2] , n302, n292, \count[29] , \count[30] , n325, 
        \count241[14] , \count241[27] , \count[18] , n350, \n239[1] , n359, 
        n365, n289, \count[4] , \count[11] , \count[22] , n319, \count241[10] , 
        \count241[23] , n342, \count[9] , \count[26] , \count[15] , \count[0] , 
        \count241[19] , n310, n337, n318, \count241[1] , n351, \DataIn[11] , 
        \ScanReg[2] , \ScanReg[15] , n293, n324, n303, \count241[8] , 
        \DataIn[15] , n311, n336, \count241[5] , n358, n364, n343, 
        \ScanReg[6] , \ScanReg[11] , \ScanReg[4] , \ScanReg[13] , n363, n344, 
        \count241[7] , n316, n294, n331, n323, n304, \ScanReg[0] , n356, 
        \DataIn[13] , \ScanReg[9] , n338, \count241[3] , n333, n314, n361, 
        n346, \ScanReg[1] , \ScanReg[8] , \DataIn[12] , \count241[2] , n328, 
        \ScanReg[5] , \ScanReg[12] , n354, n368, \count241[6] , n296, n321, 
        n306, \DataIn[14] , n291, n301, \count241[4] , n326, n348, 
        \ScanReg[7] , n353, \ScanReg[10] , \count241[0] , n366, n298, n308, 
        n341, \DataIn[10] , \ScanReg[14] , \DataIn[8] , \DataIn[7] , 
        \count241[9] , n334, n313, \ScanReg[3] , \count241[11] , 
        \count241[22] , \count[8] , n352, \count[1] , \count[14] , n349, 
        \count[27] , \DataIn[3] , n300, n290, \count241[18] , n312, n327, 
        \count241[15] , \count241[26] , n335, \count[19] , n340, n367, 
        \DataIn[1] , n299, \count[23] , \count[5] , \count[10] , n309, n360, 
        n347, n329, \count[7] , \count[12] , \count[21] , \count241[17] , 
        \count241[24] , \DataIn[5] , n332, \count[28] , n315, \count[31] , 
        n369, \count241[29] , n320, \count241[30] , n297, n307, \count[16] , 
        \count[3] , \count[25] , n355, \count241[20] , \count241[13] ;
    tri \DataOut[27]1 , \DataOut[14]1 , \DataOut[26]1 , \DataOut[15]1 , 
        \DataOut[31] , \DataOut[18]1 , \DataOut[0]1 , \DataOut[19]1 , 
        \DataOut[1]1 , \DataOut[23]1 , \DataOut[22]1 , \DataOut[11]1 , 
        \DataOut[10]1 , \DataOut[9]1 , \DataOut[8]1 , \DataOut[5]1 , 
        \DataOut[4]1 , \DataOut[21]1 , \DataOut[20]1 , \DataOut[13]1 , 
        \DataOut[12]1 , \DataOut[7]1 , \DataOut[6]1 , \DataOut[25]1 , 
        \DataOut[16]1 , \DataOut[24]1 , \DataOut[17]1 , \DataOut[29]1 , 
        \DataOut[30]1 , \DataOut[2]1 , \DataOut[28]1 , \DataOut[3]1 ;
    assign \DataIn[15]  = DataIn[15];
    assign \DataIn[14]  = DataIn[14];
    assign \DataIn[13]  = DataIn[13];
    assign \DataIn[12]  = DataIn[12];
    assign \DataIn[11]  = DataIn[11];
    assign \DataIn[10]  = DataIn[10];
    assign \DataIn[9]  = DataIn[9];
    assign \DataIn[8]  = DataIn[8];
    assign \DataIn[7]  = DataIn[7];
    assign \DataIn[6]  = DataIn[6];
    assign \DataIn[5]  = DataIn[5];
    assign \DataIn[4]  = DataIn[4];
    assign \DataIn[3]  = DataIn[3];
    assign \DataIn[2]  = DataIn[2];
    assign \DataIn[1]  = DataIn[1];
    assign \DataIn[0]  = DataIn[0];
    assign DataOut[31] = \DataOut[31] ;
    assign DataOut[30] = \DataOut[30]1 ;
    assign DataOut[29] = \DataOut[29]1 ;
    assign DataOut[28] = \DataOut[28]1 ;
    assign DataOut[27] = \DataOut[27]1 ;
    assign DataOut[26] = \DataOut[26]1 ;
    assign DataOut[25] = \DataOut[25]1 ;
    assign DataOut[24] = \DataOut[24]1 ;
    assign DataOut[23] = \DataOut[23]1 ;
    assign DataOut[22] = \DataOut[22]1 ;
    assign DataOut[21] = \DataOut[21]1 ;
    assign DataOut[20] = \DataOut[20]1 ;
    assign DataOut[19] = \DataOut[19]1 ;
    assign DataOut[18] = \DataOut[18]1 ;
    assign DataOut[17] = \DataOut[17]1 ;
    assign DataOut[16] = \DataOut[16]1 ;
    assign DataOut[15] = \DataOut[15]1 ;
    assign DataOut[14] = \DataOut[14]1 ;
    assign DataOut[13] = \DataOut[13]1 ;
    assign DataOut[12] = \DataOut[12]1 ;
    assign DataOut[11] = \DataOut[11]1 ;
    assign DataOut[10] = \DataOut[10]1 ;
    assign DataOut[9] = \DataOut[9]1 ;
    assign DataOut[8] = \DataOut[8]1 ;
    assign DataOut[7] = \DataOut[7]1 ;
    assign DataOut[6] = \DataOut[6]1 ;
    assign DataOut[5] = \DataOut[5]1 ;
    assign DataOut[4] = \DataOut[4]1 ;
    assign DataOut[3] = \DataOut[3]1 ;
    assign DataOut[2] = \DataOut[2]1 ;
    assign DataOut[1] = \DataOut[1]1 ;
    assign DataOut[0] = \DataOut[0]1 ;
    assign ScanOut[15] = \DataIn[15] ;
    assign ScanOut[14] = \DataIn[14] ;
    assign ScanOut[13] = \DataIn[13] ;
    assign ScanOut[12] = \DataIn[12] ;
    assign ScanOut[11] = \DataIn[11] ;
    assign ScanOut[10] = \DataIn[10] ;
    assign ScanOut[9] = \DataIn[9] ;
    assign ScanOut[8] = \DataIn[8] ;
    assign ScanOut[7] = \DataIn[7] ;
    assign ScanOut[6] = \DataIn[6] ;
    assign ScanOut[5] = \DataIn[5] ;
    assign ScanOut[4] = \DataIn[4] ;
    assign ScanOut[3] = \DataIn[3] ;
    assign ScanOut[2] = \DataIn[2] ;
    assign ScanOut[1] = \DataIn[1] ;
    assign ScanOut[0] = \DataIn[0] ;
    VMW_AO22 U54 ( .A(\DataIn[8] ), .B(n295), .C(\count241[8] ), .D(n296), .Z(
        n362) );
    VMW_AO22 U73 ( .A(DataIn[27]), .B(n295), .C(\count241[27] ), .D(n296), .Z(
        n343) );
    VMW_AO22 U113 ( .A(\ScanReg[11] ), .B(n298), .C(\count[11] ), .D(n297), 
        .Z(n336) );
    VMW_BUFIZ U134 ( .A(n312), .E(n311), .Z(\DataOut[4]1 ) );
    VMW_AO22 U68 ( .A(DataIn[22]), .B(n295), .C(\count241[22] ), .D(n296), .Z(
        n348) );
    VMW_AOI211 U96 ( .A(n297), .B(WR), .C(n289), .D(Reset), .Z(n296) );
    VMW_AO22 U108 ( .A(\ScanReg[1] ), .B(n298), .C(\count[1] ), .D(n297), .Z(
        n337) );
    VMW_BUFIZ U141 ( .A(n319), .E(n311), .Z(\DataOut[31] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \count_reg[6]  ( .D(n364), .CP(Clk), .Q(\count[6] ) );
    VMW_AO22 U46 ( .A(\DataIn[0] ), .B(n295), .C(\count241[0] ), .D(n296), .Z(
        n370) );
    VMW_AO22 U61 ( .A(\DataIn[15] ), .B(n295), .C(\count241[15] ), .D(n296), 
        .Z(n355) );
    VMW_AND2 U84 ( .A(n297), .B(\count[29] ), .Z(n325) );
    VMW_BUFIZ U148 ( .A(n326), .E(n311), .Z(\DataOut[20]1 ) );
    VMW_BUFIZ U153 ( .A(n331), .E(n311), .Z(\DataOut[5]1 ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \count_reg[2]  ( .D(n368), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AO22 U101 ( .A(\ScanReg[8] ), .B(n298), .C(\count[8] ), .D(n297), .Z(
        n338) );
    VMW_INV U126 ( .A(n289), .Z(Enable) );
    VMW_AO22 U48 ( .A(\DataIn[2] ), .B(n295), .C(\count241[2] ), .D(n296), .Z(
        n368) );
    VMW_AO22 U66 ( .A(DataIn[20]), .B(n295), .C(\count241[20] ), .D(n296), .Z(
        n350) );
    VMW_AO22 U106 ( .A(\ScanReg[3] ), .B(n298), .C(\count[3] ), .D(n297), .Z(
        n327) );
    VMW_NOR4 U121 ( .A(\count[12] ), .B(\count[13] ), .C(\count[14] ), .D(
        \count[15] ), .Z(n293) );
    VMW_AND2 U83 ( .A(n297), .B(\count[20] ), .Z(n326) );
    VMW_FD \count_reg[0]  ( .D(n370), .CP(Clk), .Q(\count[0] ) );
    VMW_OAI21 U98 ( .A(RD), .B(WR), .C(n301), .Z(n300) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_INV U128 ( .A(n300), .Z(ScanEnable) );
    VMW_BUFIZ U154 ( .A(n332), .E(n311), .Z(\DataOut[26]1 ) );
    VMW_FD \count_reg[9]  ( .D(n361), .CP(Clk), .Q(\count[9] ) );
    VMW_FD \count_reg[4]  ( .D(n366), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    FFT_Control_SIZE16_IDWIDTH1_SCAN1_DW01_dec_32_0 sub_183 ( .A({\count[31] , 
        \count[30] , \count[29] , \count[28] , \count[27] , \count[26] , 
        \count[25] , \count[24] , \count[23] , \count[22] , \count[21] , 
        \count[20] , \count[19] , \count[18] , \count[17] , \count[16] , 
        \count[15] , \count[14] , \count[13] , \count[12] , \count[11] , 
        \count[10] , \count[9] , \count[8] , \count[7] , \count[6] , 
        \count[5] , \count[4] , \count[3] , \count[2] , \count[1] , \count[0] 
        }), .SUM({\n239[1] , \count241[30] , \count241[29] , \count241[28] , 
        \count241[27] , \count241[26] , \count241[25] , \count241[24] , 
        \count241[23] , \count241[22] , \count241[21] , \count241[20] , 
        \count241[19] , \count241[18] , \count241[17] , \count241[16] , 
        \count241[15] , \count241[14] , \count241[13] , \count241[12] , 
        \count241[11] , \count241[10] , \count241[9] , \count241[8] , 
        \count241[7] , \count241[6] , \count241[5] , \count241[4] , 
        \count241[3] , \count241[2] , \count241[1] , \count241[0] }) );
    VMW_AO22 U53 ( .A(\DataIn[7] ), .B(n295), .C(\count241[7] ), .D(n296), .Z(
        n363) );
    VMW_AND2 U91 ( .A(n297), .B(\count[27] ), .Z(n313) );
    VMW_BUFIZ U146 ( .A(n324), .E(n311), .Z(\DataOut[30]1 ) );
    VMW_AO22 U74 ( .A(DataIn[28]), .B(n295), .C(\count241[28] ), .D(n296), .Z(
        n342) );
    VMW_AO22 U114 ( .A(\ScanReg[10] ), .B(n298), .C(\count[10] ), .D(n297), 
        .Z(n308) );
    VMW_BUFIZ U133 ( .A(n310), .E(n311), .Z(\DataOut[9]1 ) );
    VMW_XNOR2 U99 ( .A(Addr[0]), .B(ScanId), .Z(n301) );
    VMW_BUFIZ U155 ( .A(n333), .E(n311), .Z(\DataOut[15]1 ) );
    VMW_FD \count_reg[22]  ( .D(n348), .CP(Clk), .Q(\count[22] ) );
    VMW_FD \count_reg[11]  ( .D(n359), .CP(Clk), .Q(\count[11] ) );
    VMW_AO22 U47 ( .A(\DataIn[1] ), .B(n295), .C(\count241[1] ), .D(n296), .Z(
        n369) );
    VMW_AO22 U49 ( .A(\DataIn[3] ), .B(n295), .C(\count241[3] ), .D(n296), .Z(
        n367) );
    VMW_AO22 U52 ( .A(\DataIn[6] ), .B(n295), .C(\count241[6] ), .D(n296), .Z(
        n364) );
    VMW_AO22 U67 ( .A(DataIn[21]), .B(n295), .C(\count241[21] ), .D(n296), .Z(
        n349) );
    VMW_AND2 U82 ( .A(n297), .B(\count[24] ), .Z(n328) );
    VMW_FD \count_reg[18]  ( .D(n352), .CP(Clk), .Q(\count[18] ) );
    VMW_AO22 U107 ( .A(\ScanReg[2] ), .B(n298), .C(\count[2] ), .D(n297), .Z(
        n322) );
    VMW_AND4 U120 ( .A(n305), .B(n304), .C(n303), .D(n302), .Z(n294) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AO22 U75 ( .A(DataIn[29]), .B(n295), .C(\count241[29] ), .D(n296), .Z(
        n341) );
    VMW_AO22 U115 ( .A(\ScanReg[0] ), .B(n298), .C(\count[0] ), .D(n297), .Z(
        n309) );
    VMW_BUFIZ U132 ( .A(n309), .E(n311), .Z(\DataOut[0]1 ) );
    VMW_FD \count_reg[15]  ( .D(n355), .CP(Clk), .Q(\count[15] ) );
    VMW_FD \count_reg[26]  ( .D(n344), .CP(Clk), .Q(\count[26] ) );
    VMW_AND2 U90 ( .A(n297), .B(\count[25] ), .Z(n315) );
    VMW_BUFIZ U129 ( .A(n306), .E(n311), .Z(\DataOut[23]1 ) );
    VMW_BUFIZ U147 ( .A(n325), .E(n311), .Z(\DataOut[29]1 ) );
    VMW_BUFIZ U160 ( .A(n338), .E(n311), .Z(\DataOut[8]1 ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_AO22 U55 ( .A(\DataIn[9] ), .B(n295), .C(\count241[9] ), .D(n296), .Z(
        n361) );
    VMW_AO22 U69 ( .A(DataIn[23]), .B(n295), .C(\count241[23] ), .D(n296), .Z(
        n347) );
    VMW_AO22 U109 ( .A(\ScanReg[15] ), .B(n298), .C(\count[15] ), .D(n297), 
        .Z(n333) );
    VMW_AO22 U72 ( .A(DataIn[26]), .B(n295), .C(\count241[26] ), .D(n296), .Z(
        n344) );
    VMW_NOR3 U97 ( .A(n298), .B(Reset), .C(n299), .Z(n295) );
    VMW_BUFIZ U140 ( .A(n318), .E(n311), .Z(\DataOut[6]1 ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD \count_reg[17]  ( .D(n353), .CP(Clk), .Q(\count[17] ) );
    VMW_AO22 U112 ( .A(\ScanReg[12] ), .B(n298), .C(\count[12] ), .D(n297), 
        .Z(n317) );
    VMW_FD \count_reg[24]  ( .D(n346), .CP(Clk), .Q(\count[24] ) );
    VMW_BUFIZ U135 ( .A(n313), .E(n311), .Z(\DataOut[27]1 ) );
    VMW_AO22 U60 ( .A(\DataIn[14] ), .B(n295), .C(\count241[14] ), .D(n296), 
        .Z(n356) );
    VMW_AO22 U100 ( .A(\ScanReg[9] ), .B(n298), .C(\count[9] ), .D(n297), .Z(
        n310) );
    VMW_INV U127 ( .A(WR), .Z(n299) );
    VMW_AND2 U85 ( .A(n297), .B(\count[30] ), .Z(n324) );
    VMW_BUFIZ U149 ( .A(n327), .E(n311), .Z(\DataOut[3]1 ) );
    VMW_FD \count_reg[30]  ( .D(n340), .CP(Clk), .Q(\count[30] ) );
    VMW_FD \count_reg[29]  ( .D(n341), .CP(Clk), .Q(\count[29] ) );
    VMW_BUFIZ U152 ( .A(n330), .E(n311), .Z(\DataOut[7]1 ) );
    VMW_FD \count_reg[20]  ( .D(n350), .CP(Clk), .Q(\count[20] ) );
    VMW_FD \count_reg[13]  ( .D(n357), .CP(Clk), .Q(\count[13] ) );
    VMW_AND5 U45 ( .A(n290), .B(n291), .C(n292), .D(n293), .E(n294), .Z(n289)
         );
    VMW_AO22 U57 ( .A(\DataIn[11] ), .B(n295), .C(\count241[11] ), .D(n296), 
        .Z(n359) );
    VMW_BUFIZ U137 ( .A(n315), .E(n311), .Z(\DataOut[25]1 ) );
    VMW_AO22 U70 ( .A(DataIn[24]), .B(n295), .C(\count241[24] ), .D(n296), .Z(
        n346) );
    VMW_AND2 U79 ( .A(n297), .B(\count[18] ), .Z(n334) );
    VMW_XNOR2 U95 ( .A(Addr[0]), .B(Id), .Z(n297) );
    VMW_AO22 U110 ( .A(\ScanReg[14] ), .B(n298), .C(\count[14] ), .D(n297), 
        .Z(n314) );
    VMW_BUFIZ U159 ( .A(n337), .E(n311), .Z(\DataOut[1]1 ) );
    VMW_NOR4 U119 ( .A(\count[16] ), .B(\count[17] ), .C(\count[18] ), .D(
        \count[19] ), .Z(n305) );
    VMW_BUFIZ U142 ( .A(n320), .E(n311), .Z(\DataOut[21]1 ) );
    VMW_FD \count_reg[31]  ( .D(n339), .CP(Clk), .Q(\count[31] ) );
    VMW_FD \count_reg[28]  ( .D(n342), .CP(Clk), .Q(\count[28] ) );
    VMW_FD \count_reg[21]  ( .D(n349), .CP(Clk), .Q(\count[21] ) );
    VMW_FD \count_reg[12]  ( .D(n358), .CP(Clk), .Q(\count[12] ) );
    VMW_AND2 U87 ( .A(n297), .B(\count[21] ), .Z(n320) );
    VMW_BUFIZ U150 ( .A(n328), .E(n311), .Z(\DataOut[24]1 ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_INV U125 ( .A(n297), .Z(n298) );
    VMW_AO22 U50 ( .A(\DataIn[4] ), .B(n295), .C(\count241[4] ), .D(n296), .Z(
        n366) );
    VMW_AO22 U59 ( .A(\DataIn[13] ), .B(n295), .C(\count241[13] ), .D(n296), 
        .Z(n357) );
    VMW_AO22 U62 ( .A(DataIn[16]), .B(n295), .C(\count241[16] ), .D(n296), .Z(
        n354) );
    VMW_AO22 U65 ( .A(DataIn[19]), .B(n295), .C(\count241[19] ), .D(n296), .Z(
        n351) );
    VMW_AO22 U102 ( .A(\ScanReg[7] ), .B(n298), .C(\count[7] ), .D(n297), .Z(
        n330) );
    VMW_FD \count_reg[25]  ( .D(n345), .CP(Clk), .Q(\count[25] ) );
    VMW_FD \count_reg[16]  ( .D(n354), .CP(Clk), .Q(\count[16] ) );
    VMW_AO22 U105 ( .A(\ScanReg[4] ), .B(n298), .C(\count[4] ), .D(n297), .Z(
        n312) );
    VMW_AND2 U80 ( .A(n297), .B(\count[26] ), .Z(n332) );
    VMW_NOR4 U122 ( .A(\count[8] ), .B(\count[9] ), .C(\count[10] ), .D(
        \count[11] ), .Z(n292) );
    VMW_FD \count_reg[14]  ( .D(n356), .CP(Clk), .Q(\count[14] ) );
    VMW_FD \count_reg[27]  ( .D(n343), .CP(Clk), .Q(\count[27] ) );
    VMW_BUFIZ U139 ( .A(n317), .E(n311), .Z(\DataOut[12]1 ) );
    VMW_BUFIZ U157 ( .A(n335), .E(n311), .Z(\DataOut[22]1 ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO22 U77 ( .A(DataIn[31]), .B(n295), .C(\n239[1] ), .D(n296), .Z(n339)
         );
    VMW_AND2 U89 ( .A(n297), .B(\count[16] ), .Z(n316) );
    VMW_AO21 U92 ( .A(RD), .B(ScanEnable), .C(n297), .Z(n311) );
    VMW_BUFIZ U145 ( .A(n323), .E(n311), .Z(\DataOut[13]1 ) );
    VMW_FD \count_reg[23]  ( .D(n347), .CP(Clk), .Q(\count[23] ) );
    VMW_FD \count_reg[10]  ( .D(n360), .CP(Clk), .Q(\count[10] ) );
    VMW_NOR4 U117 ( .A(\count[24] ), .B(\count[25] ), .C(\count[26] ), .D(
        \count[27] ), .Z(n303) );
    VMW_FD \count_reg[19]  ( .D(n351), .CP(Clk), .Q(\count[19] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U51 ( .A(\DataIn[5] ), .B(n295), .C(\count241[5] ), .D(n296), .Z(
        n365) );
    VMW_AO22 U58 ( .A(\DataIn[12] ), .B(n295), .C(\count241[12] ), .D(n296), 
        .Z(n358) );
    VMW_BUFIZ U130 ( .A(n307), .E(n311), .Z(\DataOut[19]1 ) );
    VMW_BUFIZ U138 ( .A(n316), .E(n311), .Z(\DataOut[16]1 ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n365), .CP(Clk), .Q(\count[5] ) );
    VMW_AO22 U64 ( .A(DataIn[18]), .B(n295), .C(\count241[18] ), .D(n296), .Z(
        n352) );
    VMW_AND2 U81 ( .A(n297), .B(\count[17] ), .Z(n329) );
    VMW_BUFIZ U156 ( .A(n334), .E(n311), .Z(\DataOut[18]1 ) );
    VMW_AO22 U104 ( .A(\ScanReg[5] ), .B(n298), .C(\count[5] ), .D(n297), .Z(
        n331) );
    VMW_AO22 U76 ( .A(DataIn[30]), .B(n295), .C(\count241[30] ), .D(n296), .Z(
        n340) );
    VMW_NOR4 U116 ( .A(\count[28] ), .B(\count[29] ), .C(\count[30] ), .D(
        \count[31] ), .Z(n302) );
    VMW_NOR4 U123 ( .A(\count[4] ), .B(\count[5] ), .C(\count[6] ), .D(
        \count[7] ), .Z(n291) );
    VMW_AO22 U56 ( .A(\DataIn[10] ), .B(n295), .C(\count241[10] ), .D(n296), 
        .Z(n360) );
    VMW_AND2 U88 ( .A(n297), .B(\count[31] ), .Z(n319) );
    VMW_AND2 U93 ( .A(n297), .B(\count[19] ), .Z(n307) );
    VMW_BUFIZ U131 ( .A(n308), .E(n311), .Z(\DataOut[10]1 ) );
    VMW_FD \count_reg[1]  ( .D(n369), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(n297), .B(\count[23] ), .Z(n306) );
    VMW_BUFIZ U143 ( .A(n321), .E(n311), .Z(\DataOut[28]1 ) );
    VMW_BUFIZ U144 ( .A(n322), .E(n311), .Z(\DataOut[2]1 ) );
    VMW_FD \count_reg[8]  ( .D(n362), .CP(Clk), .Q(\count[8] ) );
    VMW_BUFIZ U158 ( .A(n336), .E(n311), .Z(\DataOut[11]1 ) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_FD \count_reg[3]  ( .D(n367), .CP(Clk), .Q(\count[3] ) );
    VMW_BUFIZ U136 ( .A(n314), .E(n311), .Z(\DataOut[14]1 ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AO22 U63 ( .A(DataIn[17]), .B(n295), .C(\count241[17] ), .D(n296), .Z(
        n353) );
    VMW_AO22 U71 ( .A(DataIn[25]), .B(n295), .C(\count241[25] ), .D(n296), .Z(
        n345) );
    VMW_AO22 U111 ( .A(\ScanReg[13] ), .B(n298), .C(\count[13] ), .D(n297), 
        .Z(n323) );
    VMW_NOR4 U124 ( .A(\count[0] ), .B(\count[1] ), .C(\count[2] ), .D(
        \count[3] ), .Z(n290) );
    VMW_AND2 U78 ( .A(n297), .B(\count[22] ), .Z(n335) );
    VMW_AND2 U86 ( .A(n297), .B(\count[28] ), .Z(n321) );
    VMW_AO22 U103 ( .A(\ScanReg[6] ), .B(n298), .C(\count[6] ), .D(n297), .Z(
        n318) );
    VMW_NOR4 U118 ( .A(\count[20] ), .B(\count[21] ), .C(\count[22] ), .D(
        \count[23] ), .Z(n304) );
    VMW_BUFIZ U151 ( .A(n329), .E(n311), .Z(\DataOut[17]1 ) );
    VMW_FD \count_reg[7]  ( .D(n363), .CP(Clk), .Q(\count[7] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \nLeftOut_7[13] , \nRightOut_86[5] , \ScanLink0[13] , 
        \nLeftOut_20[8] , \nRightOut_54[3] , \nRightOut_57[0] , 
        \nRightOut_30[7] , \nRightOut_85[6] , \nLeftOut_88[6] , 
        \nLeftOut_95[9] , \ScanLink29[3] , \nLeftOut_3[11] , \ScanLink4[11] , 
        \nLeftOut_8[6] , \nLeftOut_59[3] , \ScanLink9[6] , \nRightOut_10[16] , 
        \nLeftOut_25[5] , \nRightOut_33[4] , \nLeftOut_34[11] , 
        \nLeftOut_62[10] , \nLeftOut_54[15] , \nLeftOut_26[6] , 
        \nRightOut_70[12] , \nRightOut_26[13] , \nRightOut_9[12] , 
        \nRightOut_9[4] , \nLeftOut_17[13] , \nLeftOut_21[16] , 
        \nRightOut_36[9] , \nLeftOut_41[1] , \nRightOut_83[8] , 
        \ScanLink32[2] , \nLeftOut_93[7] , \nRightOut_28[5] , 
        \nLeftOut_41[12] , \nLeftOut_90[4] , \ScanLink19[11] , 
        \nRightOut_33[14] , \nLeftOut_42[2] , \nRightOut_42[15] , 
        \nRightOut_53[10] , \nRightOut_65[15] , \ScanLink31[1] , 
        \nLeftOut_13[11] , \nRightOut_14[14] , \ScanLink15[7] , 
        \nRightOut_22[11] , \nLeftOut_66[4] , \nRightOut_74[10] , 
        \ScanLink16[4] , \nLeftOut_65[7] , \nLeftOut_30[13] , 
        \nLeftOut_66[12] , \nLeftOut_78[8] , \nRightOut_37[16] , 
        \nRightOut_57[12] , \nRightOut_75[8] , \nRightOut_68[7] , 
        \nLeftOut_88[14] , \nLeftOut_25[14] , \nLeftOut_45[10] , 
        \nLeftOut_73[15] , \ScanLink13[9] , \nRightOut_17[2] , 
        \nRightOut_14[1] , \nLeftOut_63[9] , \nRightOut_3[14] , 
        \nLeftOut_11[9] , \nLeftOut_19[1] , \nRightOut_73[6] , 
        \nRightOut_66[1] , \nRightOut_70[5] , \nLeftOut_17[7] , 
        \nRightOut_65[2] , \nLeftOut_68[2] , \ScanLink18[2] , 
        \nRightOut_48[13] , \nRightOut_4[1] , \nLeftOut_5[3] , 
        \nLeftOut_14[4] , \nRightOut_19[4] , \nLeftOut_54[6] , 
        \nLeftOut_70[0] , \nLeftOut_73[3] , \nRightOut_90[10] , 
        \ScanLink17[15] , \nLeftOut_79[13] , \ScanLink21[10] , 
        \nLeftOut_82[12] , \ScanLink27[5] , \nLeftOut_6[0] , \nRightOut_7[16] , 
        \nLeftOut_49[9] , \nLeftOut_86[0] , \nLeftOut_57[5] , 
        \nRightOut_81[15] , \nLeftOut_85[3] , \ScanLink30[15] , 
        \nLeftOut_68[16] , \ScanLink24[6] , \nRightOut_25[0] , 
        \nLeftOut_30[2] , \nRightOut_39[12] , \nRightOut_59[16] , 
        \nLeftOut_33[1] , \nLeftOut_86[10] , \nRightOut_88[3] , 
        \nRightOut_44[9] , \ScanLink25[12] , \nLeftOut_52[8] , 
        \nRightOut_59[6] , \nRightOut_94[12] , \nRightOut_26[3] , 
        \ScanLink22[8] , \nRightOut_93[2] , \nLeftOut_0[7] , \nLeftOut_2[12] , 
        \ScanLink4[3] , \ScanLink7[0] , \nRightOut_41[4] , \nRightOut_7[2] , 
        \nLeftOut_28[0] , \nRightOut_42[7] , \nRightOut_90[1] , 
        \nLeftOut_3[4] , \nRightOut_4[8] , \ScanLink5[12] , \nLeftOut_70[9] , 
        \nRightOut_8[11] , \nRightOut_23[12] , \nLeftOut_31[10] , 
        \nRightOut_60[6] , \nRightOut_63[5] , \nLeftOut_51[14] , 
        \nLeftOut_67[11] , \nLeftOut_75[4] , \nLeftOut_76[7] , 
        \nRightOut_43[16] , \nRightOut_75[13] , \nLeftOut_11[0] , 
        \nRightOut_11[15] , \nLeftOut_12[12] , \nLeftOut_44[13] , 
        \nRightOut_66[8] , \nLeftOut_72[16] , \nLeftOut_12[3] , 
        \nRightOut_60[14] , \nRightOut_78[4] , \nRightOut_36[15] , 
        \nRightOut_56[11] , \nLeftOut_36[5] , \nRightOut_47[14] , 
        \ScanLink7[9] , \nRightOut_27[10] , \nRightOut_71[11] , 
        \nRightOut_25[9] , \nLeftOut_28[9] , \nLeftOut_35[12] , 
        \nLeftOut_35[6] , \nLeftOut_55[16] , \nRightOut_90[8] , 
        \nRightOut_52[13] , \nLeftOut_63[13] , \nLeftOut_52[1] , 
        \nRightOut_64[16] , \ScanLink21[2] , \nLeftOut_16[10] , 
        \nRightOut_38[6] , \nLeftOut_40[11] , \nLeftOut_80[7] , 
        \ScanLink18[12] , \nLeftOut_20[15] , \nLeftOut_76[14] , 
        \nLeftOut_83[4] , \nLeftOut_51[2] , \ScanLink22[1] , \ScanLink1[10] , 
        \nRightOut_95[5] , \ScanLink1[7] , \nRightOut_1[5] , \ScanLink2[4] , 
        \nRightOut_47[3] , \nRightOut_2[6] , \nLeftOut_33[8] , 
        \nRightOut_44[0] , \nLeftOut_6[10] , \nLeftOut_6[9] , 
        \nRightOut_20[4] , \nRightOut_23[7] , \nLeftOut_49[0] , 
        \nLeftOut_86[9] , \nRightOut_6[15] , \nRightOut_35[3] , 
        \nRightOut_36[0] , \nLeftOut_41[8] , \nLeftOut_38[3] , 
        \nRightOut_80[2] , \ScanLink31[8] , \nLeftOut_47[6] , 
        \nRightOut_51[7] , \nRightOut_52[4] , \nRightOut_83[1] , 
        \nLeftOut_69[15] , \nRightOut_80[16] , \nLeftOut_95[0] , 
        \ScanLink12[14] , \nLeftOut_44[5] , \nLeftOut_92[14] , 
        \nRightOut_49[5] , \nRightOut_95[11] , \nLeftOut_19[8] , 
        \nLeftOut_20[1] , \nLeftOut_23[2] , \nRightOut_57[9] , 
        \ScanLink24[11] , \nRightOut_38[11] , \nRightOut_58[15] , 
        \nLeftOut_87[13] , \nRightOut_29[14] , \nRightOut_49[10] , 
        \nLeftOut_60[3] , \nRightOut_84[14] , \nLeftOut_83[11] , 
        \nLeftOut_3[9] , \nLeftOut_8[14] , \ScanLink10[3] , \ScanLink13[0] , 
        \nLeftOut_63[0] , \nLeftOut_78[10] , \nRightOut_14[8] , 
        \nLeftOut_18[14] , \ScanLink20[13] , \nRightOut_75[1] , 
        \nRightOut_91[13] , \nRightOut_11[5] , \nRightOut_76[2] , 
        \nRightOut_12[6] , \nRightOut_25[4] , \nRightOut_26[7] , 
        \nLeftOut_78[1] , \nLeftOut_83[9] , \ScanLink7[4] , \nRightOut_7[6] , 
        \nLeftOut_28[4] , \nRightOut_90[5] , \nRightOut_42[3] , 
        \nRightOut_41[0] , \ScanLink4[7] , \nRightOut_4[5] , \nLeftOut_36[8] , 
        \nRightOut_93[6] , \ScanEnable[0] , \nRightOut_1[8] , \nLeftOut_5[7] , 
        \nLeftOut_6[4] , \nRightOut_20[9] , \nLeftOut_57[1] , \ScanLink30[11] , 
        \nLeftOut_68[12] , \ScanLink24[2] , \nRightOut_7[12] , 
        \nRightOut_81[11] , \nLeftOut_85[7] , \nLeftOut_54[2] , 
        \nLeftOut_86[4] , \nLeftOut_93[13] , \ScanLink27[1] , \ScanLink13[13] , 
        \nRightOut_59[2] , \nRightOut_94[16] , \nLeftOut_33[5] , 
        \ScanLink2[9] , \nLeftOut_30[6] , \nRightOut_88[7] , \nLeftOut_86[14] , 
        \nLeftOut_3[15] , \nRightOut_3[10] , \nLeftOut_14[0] , 
        \nRightOut_39[16] , \nRightOut_59[12] , \nRightOut_95[8] , 
        \nRightOut_28[13] , \nRightOut_63[8] , \nLeftOut_9[13] , 
        \nLeftOut_17[3] , \nRightOut_85[13] , \nLeftOut_19[13] , 
        \nLeftOut_70[4] , \nLeftOut_73[7] , \nLeftOut_82[16] , 
        \ScanLink21[14] , \nRightOut_19[0] , \nRightOut_90[14] , 
        \ScanLink17[11] , \nRightOut_65[6] , \nRightOut_78[9] , 
        \nRightOut_66[5] , \nLeftOut_68[6] , \nLeftOut_75[9] , \ScanLink18[6] , 
        \ScanLink4[15] , \nRightOut_14[5] , \nRightOut_17[6] , 
        \nRightOut_9[16] , \nRightOut_11[8] , \ScanLink15[3] , \ScanLink16[0] , 
        \nLeftOut_19[5] , \nRightOut_70[1] , \nLeftOut_50[13] , 
        \nLeftOut_66[16] , \nRightOut_73[2] , \nLeftOut_65[3] , 
        \nLeftOut_66[0] , \nRightOut_22[15] , \nRightOut_74[14] , 
        \nRightOut_14[10] , \nRightOut_42[11] , \ScanLink9[2] , 
        \nRightOut_9[0] , \nLeftOut_13[15] , \nLeftOut_25[10] , 
        \nLeftOut_73[11] , \nLeftOut_45[14] , \nRightOut_37[12] , 
        \nRightOut_61[13] , \nRightOut_68[3] , \nLeftOut_88[10] , 
        \nRightOut_57[16] , \nRightOut_10[12] , \nLeftOut_21[12] , 
        \nLeftOut_25[1] , \nLeftOut_26[2] , \nRightOut_46[13] , 
        \nRightOut_52[9] , \nRightOut_70[16] , \nRightOut_28[1] , 
        \nRightOut_33[10] , \nLeftOut_34[15] , \nLeftOut_54[11] , 
        \nLeftOut_42[6] , \nRightOut_53[14] , \nLeftOut_62[14] , 
        \nRightOut_65[11] , \ScanLink31[5] , \nLeftOut_41[16] , 
        \nLeftOut_90[0] , \nLeftOut_77[13] , \nLeftOut_93[3] , 
        \ScanLink19[15] , \nLeftOut_41[5] , \nRightOut_49[8] , 
        \nRightOut_54[7] , \nRightOut_57[4] , \nRightOut_85[2] , 
        \ScanLink32[6] , \nRightOut_86[1] , \nLeftOut_8[2] , \nRightOut_33[0] , 
        \nLeftOut_44[8] , \nLeftOut_59[7] , \nRightOut_2[13] , 
        \nLeftOut_8[10] , \nRightOut_30[3] , \ScanLink29[7] , 
        \nRightOut_76[6] , \nLeftOut_88[2] , \nRightOut_11[1] , 
        \nRightOut_12[2] , \nRightOut_75[5] , \nLeftOut_78[5] , 
        \ScanLink16[9] , \nRightOut_49[14] , \nLeftOut_66[9] , 
        \nRightOut_70[8] , \nRightOut_84[10] , \nRightOut_6[11] , 
        \ScanLink10[7] , \ScanLink16[12] , \nRightOut_29[10] , 
        \nLeftOut_18[10] , \nLeftOut_63[4] , \nLeftOut_78[14] , 
        \ScanLink13[4] , \nLeftOut_60[7] , \nLeftOut_83[15] , 
        \nRightOut_33[9] , \nLeftOut_44[1] , \nLeftOut_92[10] , 
        \nRightOut_80[12] , \ScanLink1[14] , \ScanLink1[3] , \nLeftOut_6[14] , 
        \nRightOut_9[9] , \ScanLink12[10] , \nLeftOut_20[5] , 
        \nRightOut_38[15] , \nLeftOut_47[2] , \nLeftOut_95[4] , 
        \ScanLink31[12] , \nLeftOut_69[11] , \nRightOut_58[11] , 
        \nLeftOut_23[6] , \ScanLink24[15] , \nRightOut_28[8] , 
        \nRightOut_35[7] , \nRightOut_49[1] , \nRightOut_86[8] , 
        \nRightOut_95[15] , \nLeftOut_90[9] , \nRightOut_36[4] , 
        \nLeftOut_25[8] , \nRightOut_51[3] , \nRightOut_83[5] , 
        \nLeftOut_38[7] , \nRightOut_52[0] , \nRightOut_80[6] , 
        \nRightOut_1[1] , \ScanLink2[0] , \nRightOut_2[2] , \nRightOut_44[4] , 
        \nRightOut_47[7] , \nRightOut_20[0] , \nLeftOut_57[8] , 
        \nRightOut_95[1] , \nRightOut_23[3] , \nLeftOut_49[4] , 
        \ScanLink27[8] , \nLeftOut_35[16] , \nLeftOut_35[2] , 
        \nLeftOut_55[12] , \nLeftOut_0[3] , \nRightOut_11[11] , 
        \nRightOut_27[14] , \nLeftOut_36[1] , \nRightOut_71[15] , 
        \nRightOut_41[9] , \nRightOut_47[10] , \nLeftOut_51[6] , 
        \ScanLink22[5] , \nLeftOut_0[1] , \ScanLink1[1] , \ScanLink2[2] , 
        \nLeftOut_2[16] , \nLeftOut_3[0] , \nLeftOut_16[14] , 
        \nLeftOut_20[11] , \nLeftOut_76[10] , \nLeftOut_83[0] , 
        \nRightOut_32[13] , \nRightOut_38[2] , \nLeftOut_40[15] , 
        \nLeftOut_80[3] , \nLeftOut_52[5] , \ScanLink21[6] , \nRightOut_8[15] , 
        \nRightOut_43[12] , \nRightOut_64[12] , \nLeftOut_11[4] , 
        \nLeftOut_12[16] , \nLeftOut_12[7] , \nRightOut_15[13] , 
        \nRightOut_23[16] , \nLeftOut_76[3] , \nLeftOut_31[14] , 
        \nLeftOut_51[10] , \nLeftOut_75[0] , \nLeftOut_67[15] , 
        \nRightOut_56[15] , \nRightOut_36[11] , \nRightOut_60[10] , 
        \nRightOut_78[0] , \nLeftOut_89[13] , \nLeftOut_24[13] , 
        \nLeftOut_72[12] , \nRightOut_19[9] , \nRightOut_2[0] , 
        \nLeftOut_14[9] , \nRightOut_63[1] , \nRightOut_47[5] , 
        \nRightOut_60[2] , \nRightOut_95[3] , \nRightOut_44[6] , 
        \nRightOut_1[3] , \nLeftOut_3[2] , \nLeftOut_6[16] , \nRightOut_59[9] , 
        \nRightOut_11[13] , \nRightOut_20[2] , \nRightOut_23[1] , 
        \nLeftOut_49[6] , \nLeftOut_54[9] , \nRightOut_47[12] , 
        \ScanLink24[9] , \nRightOut_27[16] , \nLeftOut_35[14] , 
        \nLeftOut_35[0] , \nLeftOut_36[3] , \nRightOut_42[8] , 
        \nLeftOut_55[10] , \nLeftOut_63[15] , \nRightOut_52[15] , 
        \nLeftOut_16[16] , \nRightOut_32[11] , \ScanLink21[4] , 
        \nRightOut_38[0] , \nLeftOut_52[7] , \nRightOut_64[10] , 
        \nLeftOut_80[1] , \nLeftOut_20[13] , \ScanLink18[14] , 
        \nLeftOut_76[12] , \nLeftOut_83[2] , \nLeftOut_2[14] , 
        \nLeftOut_11[6] , \nRightOut_15[11] , \nRightOut_23[14] , 
        \nLeftOut_31[16] , \nLeftOut_51[4] , \ScanLink22[7] , 
        \nLeftOut_51[12] , \nLeftOut_75[2] , \nRightOut_75[15] , 
        \nRightOut_43[10] , \nLeftOut_76[1] , \nLeftOut_12[14] , 
        \nLeftOut_24[11] , \nLeftOut_72[10] , \nLeftOut_12[5] , 
        \nRightOut_36[13] , \nLeftOut_44[15] , \nRightOut_78[2] , 
        \nLeftOut_89[11] , \nRightOut_60[12] , \nRightOut_2[11] , 
        \ScanLink5[14] , \nLeftOut_8[12] , \nLeftOut_17[8] , \nRightOut_60[0] , 
        \nRightOut_63[3] , \nRightOut_68[8] , \nRightOut_75[7] , 
        \nRightOut_11[3] , \ScanLink15[8] , \nRightOut_76[4] , 
        \nRightOut_12[0] , \nLeftOut_65[8] , \nRightOut_29[12] , 
        \nRightOut_73[9] , \nLeftOut_78[7] , \nRightOut_49[16] , 
        \nRightOut_6[13] , \ScanLink10[5] , \ScanLink13[6] , 
        \nRightOut_84[12] , \nLeftOut_60[5] , \ScanLink16[10] , 
        \nLeftOut_63[6] , \ScanLink20[15] , \nLeftOut_78[16] , 
        \nLeftOut_18[12] , \nRightOut_30[8] , \nRightOut_91[15] , 
        \nLeftOut_47[0] , \nLeftOut_69[13] , \nLeftOut_88[9] , 
        \ScanLink31[10] , \nRightOut_80[10] , \nLeftOut_95[6] , 
        \nLeftOut_8[9] , \nLeftOut_44[3] , \nRightOut_49[3] , 
        \nLeftOut_92[12] , \nLeftOut_7[15] , \ScanLink9[9] , \ScanLink12[12] , 
        \nLeftOut_20[7] , \nLeftOut_23[4] , \nLeftOut_87[15] , 
        \nLeftOut_26[9] , \nRightOut_35[5] , \nRightOut_36[6] , 
        \nRightOut_58[13] , \nRightOut_85[9] , \nLeftOut_93[8] , 
        \nLeftOut_38[5] , \nRightOut_80[4] , \nRightOut_51[1] , 
        \nRightOut_52[2] , \nRightOut_83[7] , \ScanLink9[0] , 
        \nRightOut_9[14] , \nRightOut_14[12] , \nRightOut_14[7] , 
        \nRightOut_17[4] , \nLeftOut_19[7] , \nRightOut_73[0] , 
        \nRightOut_70[3] , \nRightOut_42[13] , \nRightOut_9[2] , 
        \nRightOut_10[10] , \nRightOut_12[9] , \ScanLink15[1] , 
        \nLeftOut_66[2] , \nRightOut_74[16] , \ScanLink16[2] , 
        \nLeftOut_25[12] , \nLeftOut_30[15] , \nLeftOut_50[11] , 
        \nLeftOut_65[1] , \nRightOut_37[10] , \nRightOut_57[14] , 
        \nLeftOut_66[14] , \nRightOut_61[11] , \nLeftOut_45[16] , 
        \nRightOut_68[1] , \nLeftOut_88[12] , \nLeftOut_73[13] , 
        \nLeftOut_25[3] , \nLeftOut_54[13] , \nLeftOut_62[16] , 
        \nLeftOut_26[0] , \nRightOut_26[15] , \nRightOut_70[14] , 
        \nRightOut_46[11] , \nRightOut_51[8] , \nLeftOut_17[15] , 
        \nLeftOut_21[10] , \nLeftOut_41[7] , \ScanLink32[4] , 
        \nLeftOut_77[11] , \nLeftOut_93[1] , \nLeftOut_41[14] , 
        \nRightOut_28[3] , \nLeftOut_90[2] , \nRightOut_33[12] , 
        \nRightOut_65[13] , \ScanLink31[7] , \nLeftOut_42[4] , 
        \nRightOut_53[16] , \nRightOut_86[3] , \ScanLink0[15] , 
        \nRightOut_54[5] , \nRightOut_57[6] , \nRightOut_30[1] , 
        \nLeftOut_47[9] , \nRightOut_85[0] , \nLeftOut_88[0] , \nLeftOut_0[8] , 
        \nLeftOut_8[0] , \ScanLink29[5] , \nRightOut_25[6] , \nRightOut_33[2] , 
        \nLeftOut_59[5] , \nRightOut_38[9] , \nLeftOut_80[8] , 
        \nRightOut_26[5] , \nRightOut_93[4] , \ScanLink1[8] , \nRightOut_2[9] , 
        \ScanLink4[5] , \nRightOut_4[7] , \nLeftOut_5[5] , \ScanLink7[6] , 
        \nRightOut_7[4] , \nRightOut_41[2] , \nLeftOut_35[9] , 
        \nLeftOut_28[6] , \nRightOut_42[1] , \nRightOut_90[7] , 
        \nLeftOut_6[6] , \nRightOut_7[10] , \nRightOut_23[8] , 
        \nLeftOut_54[0] , \ScanLink27[3] , \nLeftOut_93[11] , \nLeftOut_86[6] , 
        \nLeftOut_68[10] , \nRightOut_81[13] , \nLeftOut_85[5] , 
        \nRightOut_39[14] , \nLeftOut_57[3] , \ScanLink24[0] , 
        \ScanLink30[13] , \nRightOut_59[10] , \nLeftOut_30[4] , 
        \nLeftOut_86[16] , \nRightOut_88[5] , \nRightOut_2[15] , 
        \nRightOut_3[12] , \ScanLink13[11] , \nLeftOut_33[7] , 
        \ScanLink25[14] , \nLeftOut_17[1] , \nRightOut_59[0] , 
        \nRightOut_94[14] , \nRightOut_60[9] , \nRightOut_48[15] , 
        \nRightOut_85[11] , \nLeftOut_9[11] , \nLeftOut_14[2] , 
        \nRightOut_28[11] , \nLeftOut_19[11] , \nRightOut_19[2] , 
        \nRightOut_90[16] , \nRightOut_66[7] , \nLeftOut_70[6] , 
        \nLeftOut_73[5] , \ScanLink17[13] , \nLeftOut_79[15] , 
        \nLeftOut_82[14] , \nLeftOut_20[3] , \nRightOut_35[1] , 
        \nLeftOut_42[9] , \nRightOut_65[4] , \nLeftOut_68[4] , 
        \nLeftOut_76[8] , \ScanLink18[4] , \nRightOut_36[2] , \ScanLink32[9] , 
        \nLeftOut_38[1] , \nRightOut_51[5] , \nRightOut_83[3] , 
        \nRightOut_52[6] , \nRightOut_38[13] , \nLeftOut_44[7] , 
        \nRightOut_80[0] , \nLeftOut_47[4] , \nLeftOut_59[8] , 
        \nLeftOut_92[16] , \nRightOut_80[14] , \nLeftOut_95[2] , 
        \ScanLink29[8] , \ScanLink31[14] , \nLeftOut_87[11] , \nLeftOut_23[0] , 
        \ScanLink24[13] , \nRightOut_49[12] , \nRightOut_49[7] , 
        \nRightOut_54[8] , \nRightOut_95[13] , \nRightOut_84[16] , 
        \ScanLink10[1] , \ScanLink16[14] , \nLeftOut_18[16] , 
        \nRightOut_29[16] , \nRightOut_91[11] , \ScanLink13[2] , 
        \nRightOut_17[9] , \nLeftOut_63[2] , \ScanLink20[11] , 
        \nLeftOut_78[12] , \nLeftOut_0[5] , \nLeftOut_2[10] , \ScanLink5[10] , 
        \nLeftOut_8[16] , \nLeftOut_60[1] , \nLeftOut_83[13] , 
        \nRightOut_76[0] , \nRightOut_11[7] , \nRightOut_12[4] , 
        \nRightOut_75[3] , \nLeftOut_78[3] , \nLeftOut_73[8] , \ScanLink4[8] , 
        \nRightOut_7[9] , \nRightOut_8[13] , \nRightOut_15[15] , 
        \nRightOut_60[4] , \nRightOut_63[7] , \ScanLink18[9] , 
        \nRightOut_43[14] , \nLeftOut_11[2] , \nLeftOut_12[10] , 
        \nLeftOut_12[1] , \nRightOut_23[10] , \nLeftOut_31[12] , 
        \nLeftOut_51[16] , \nLeftOut_75[6] , \nRightOut_75[11] , 
        \nLeftOut_76[5] , \nRightOut_56[13] , \nLeftOut_67[13] , 
        \nLeftOut_68[9] , \nRightOut_60[16] , \nRightOut_65[9] , 
        \nLeftOut_44[11] , \nRightOut_78[6] , \nLeftOut_89[15] , 
        \nLeftOut_24[15] , \nLeftOut_72[14] , \nLeftOut_35[10] , 
        \nLeftOut_55[14] , \nLeftOut_63[11] , \nRightOut_27[12] , 
        \nLeftOut_35[4] , \nLeftOut_36[7] , \nRightOut_71[13] , 
        \nRightOut_47[16] , \nRightOut_93[9] , \ScanLink1[12] , \ScanLink1[5] , 
        \nRightOut_1[7] , \nLeftOut_3[6] , \nLeftOut_16[12] , 
        \nRightOut_26[8] , \nLeftOut_51[0] , \ScanLink22[3] , 
        \nLeftOut_40[13] , \nLeftOut_76[16] , \nLeftOut_83[6] , 
        \ScanLink18[10] , \nRightOut_38[4] , \nLeftOut_80[5] , 
        \nRightOut_64[14] , \nLeftOut_6[12] , \nRightOut_32[15] , 
        \ScanLink21[0] , \nLeftOut_52[3] , \nRightOut_52[11] , \ScanLink2[6] , 
        \nRightOut_44[2] , \nRightOut_2[4] , \nLeftOut_30[9] , 
        \nRightOut_47[1] , \nRightOut_88[8] , \nRightOut_3[16] , 
        \nLeftOut_5[8] , \nRightOut_20[6] , \nRightOut_95[7] , 
        \nLeftOut_49[2] , \nLeftOut_85[8] , \nLeftOut_9[15] , \nLeftOut_12[8] , 
        \nRightOut_23[5] , \nRightOut_65[0] , \nLeftOut_14[6] , 
        \nRightOut_66[3] , \nLeftOut_68[0] , \ScanLink18[0] , 
        \nRightOut_28[15] , \nRightOut_48[11] , \nRightOut_4[3] , 
        \nLeftOut_5[1] , \nLeftOut_6[2] , \nLeftOut_17[5] , \nRightOut_85[15] , 
        \nLeftOut_19[15] , \nLeftOut_70[2] , \nLeftOut_82[10] , 
        \nLeftOut_73[1] , \ScanLink21[12] , \nLeftOut_79[11] , 
        \nRightOut_19[6] , \nRightOut_90[12] , \nLeftOut_68[14] , 
        \nRightOut_7[14] , \nLeftOut_57[7] , \ScanLink24[4] , \nLeftOut_85[1] , 
        \nLeftOut_86[2] , \ScanLink7[2] , \ScanLink13[15] , \nLeftOut_54[4] , 
        \ScanLink27[7] , \nRightOut_59[4] , \nLeftOut_93[15] , 
        \nRightOut_94[10] , \nRightOut_25[2] , \nRightOut_26[1] , 
        \nLeftOut_30[0] , \nLeftOut_33[3] , \ScanLink25[10] , 
        \nRightOut_47[8] , \nLeftOut_86[12] , \nRightOut_88[1] , 
        \nRightOut_39[10] , \nRightOut_59[14] , \nLeftOut_51[9] , 
        \nLeftOut_28[2] , \nRightOut_90[3] , \ScanLink21[9] , 
        \nRightOut_42[5] , \nRightOut_7[0] , \nRightOut_41[6] , 
        \ScanLink0[11] , \ScanLink4[1] , \nRightOut_85[4] , \nRightOut_93[0] , 
        \nLeftOut_23[9] , \nRightOut_54[1] , \nRightOut_57[2] , 
        \nRightOut_86[7] , \nLeftOut_7[11] , \nLeftOut_8[4] , 
        \nRightOut_33[6] , \nLeftOut_59[1] , \ScanLink29[1] , \nLeftOut_1[15] , 
        \nLeftOut_3[13] , \ScanLink9[4] , \nRightOut_30[5] , \nLeftOut_88[4] , 
        \nRightOut_9[10] , \nRightOut_9[6] , \nRightOut_10[14] , 
        \nRightOut_46[15] , \ScanLink15[5] , \ScanLink16[6] , 
        \nLeftOut_17[11] , \nLeftOut_25[7] , \nLeftOut_26[4] , 
        \nRightOut_26[11] , \nRightOut_70[10] , \nRightOut_28[7] , 
        \nRightOut_33[16] , \nLeftOut_34[13] , \nLeftOut_38[8] , 
        \nLeftOut_62[12] , \nRightOut_80[9] , \nRightOut_35[8] , 
        \nRightOut_53[12] , \ScanLink31[3] , \nLeftOut_42[0] , 
        \nLeftOut_90[6] , \nLeftOut_21[14] , \nLeftOut_41[10] , 
        \ScanLink19[13] , \nLeftOut_30[11] , \nLeftOut_41[3] , 
        \nLeftOut_77[15] , \nLeftOut_93[5] , \ScanLink32[0] , 
        \nLeftOut_66[10] , \nLeftOut_50[15] , \nLeftOut_65[5] , 
        \nRightOut_74[12] , \nRightOut_22[13] , \nLeftOut_66[6] , 
        \nLeftOut_13[13] , \nRightOut_14[16] , \nLeftOut_25[16] , 
        \nRightOut_76[9] , \nRightOut_37[14] , \nLeftOut_45[12] , 
        \nRightOut_68[5] , \nLeftOut_88[16] , \nRightOut_57[10] , 
        \nRightOut_61[15] , \ScanLink4[13] , \ScanLink10[8] , 
        \nRightOut_14[3] , \nRightOut_17[0] , \nLeftOut_60[8] , \ScanLink8[9] , 
        \nLeftOut_9[9] , \nRightOut_10[3] , \nRightOut_13[0] , 
        \nLeftOut_19[3] , \nRightOut_70[7] , \nLeftOut_64[8] , 
        \nRightOut_73[4] , \ScanLink14[8] , \nLeftOut_79[7] , \ScanLink11[5] , 
        \nRightOut_69[8] , \nRightOut_74[7] , \nRightOut_77[4] , 
        \nLeftOut_11[15] , \ScanLink12[6] , \nLeftOut_23[12] , 
        \nRightOut_31[10] , \nLeftOut_62[6] , \nRightOut_51[14] , 
        \nRightOut_67[11] , \nLeftOut_43[16] , \nLeftOut_75[13] , 
        \nRightOut_12[12] , \nRightOut_44[13] , \nLeftOut_61[5] , 
        \nRightOut_72[16] , \nLeftOut_21[7] , \nLeftOut_36[15] , 
        \nLeftOut_60[14] , \nRightOut_72[9] , \nLeftOut_56[11] , 
        \nLeftOut_22[4] , \nLeftOut_27[10] , \nLeftOut_47[14] , 
        \nRightOut_84[9] , \nRightOut_48[3] , \nLeftOut_71[11] , 
        \ScanLink29[12] , \nRightOut_55[16] , \nRightOut_35[12] , 
        \nLeftOut_52[13] , \nRightOut_63[13] , \nLeftOut_64[16] , 
        \nRightOut_16[10] , \nRightOut_40[11] , \nLeftOut_45[3] , 
        \nRightOut_20[15] , \nRightOut_31[8] , \nRightOut_76[14] , 
        \nLeftOut_27[9] , \nLeftOut_46[0] , \nRightOut_50[1] , 
        \nLeftOut_89[9] , \nLeftOut_94[6] , \nRightOut_82[7] , 
        \nLeftOut_39[5] , \nRightOut_81[4] , \nRightOut_53[2] , 
        \nRightOut_34[5] , \nRightOut_0[3] , \ScanLink0[1] , \ScanLink6[15] , 
        \nRightOut_37[6] , \nLeftOut_92[8] , \nRightOut_21[2] , 
        \nRightOut_22[1] , \ScanLink25[9] , \nRightOut_45[6] , 
        \nLeftOut_48[6] , \nLeftOut_55[9] , \nLeftOut_1[1] , \ScanLink3[2] , 
        \nRightOut_3[0] , \nRightOut_46[5] , \nRightOut_58[9] , 
        \nRightOut_94[3] , \nRightOut_69[15] , \nLeftOut_82[2] , 
        \nLeftOut_2[2] , \ScanLink15[11] , \nLeftOut_50[4] , \nLeftOut_80[16] , 
        \ScanLink23[7] , \ScanLink23[14] , \nLeftOut_34[0] , \nRightOut_39[0] , 
        \nLeftOut_53[7] , \ScanLink20[4] , \nRightOut_43[8] , \nLeftOut_81[1] , 
        \nRightOut_92[14] , \nLeftOut_95[11] , \nRightOut_1[10] , 
        \nLeftOut_37[3] , \nLeftOut_38[11] , \nLeftOut_58[15] , 
        \nRightOut_87[13] , \nRightOut_79[2] , \nLeftOut_10[6] , 
        \ScanLink11[13] , \nLeftOut_13[5] , \nLeftOut_29[14] , 
        \nLeftOut_49[10] , \nLeftOut_84[14] , \nLeftOut_77[1] , 
        \nRightOut_83[11] , \ScanLink32[11] , \nLeftOut_0[16] , 
        \nLeftOut_1[8] , \ScanLink5[5] , \nRightOut_5[12] , \nRightOut_18[14] , 
        \nRightOut_78[10] , \ScanLink6[6] , \nRightOut_6[4] , \ScanLink8[11] , 
        \nLeftOut_16[8] , \nRightOut_62[3] , \nLeftOut_74[2] , 
        \nLeftOut_91[13] , \nRightOut_61[0] , \nLeftOut_34[9] , 
        \nLeftOut_29[6] , \nRightOut_43[1] , \nRightOut_91[7] , 
        \nRightOut_92[4] , \nRightOut_5[7] , \nRightOut_40[2] , 
        \nRightOut_24[6] , \nRightOut_27[5] , \nLeftOut_81[8] , \ScanLink0[8] , 
        \nRightOut_39[9] , \nRightOut_62[10] , \nRightOut_3[9] , 
        \nLeftOut_10[16] , \nLeftOut_26[13] , \nLeftOut_32[7] , 
        \nRightOut_34[11] , \nRightOut_54[15] , \nRightOut_58[0] , 
        \nLeftOut_70[12] , \ScanLink28[11] , \nLeftOut_4[5] , \nLeftOut_7[6] , 
        \nLeftOut_31[4] , \nLeftOut_84[5] , \nRightOut_89[5] , 
        \nRightOut_17[13] , \nRightOut_21[16] , \ScanLink25[0] , 
        \nLeftOut_56[3] , \nRightOut_41[12] , \nRightOut_13[11] , 
        \nLeftOut_14[14] , \nRightOut_22[8] , \nLeftOut_55[0] , 
        \ScanLink26[3] , \nLeftOut_33[14] , \nLeftOut_42[15] , 
        \nLeftOut_53[10] , \nLeftOut_65[15] , \nLeftOut_87[6] , 
        \nLeftOut_71[6] , \nLeftOut_15[2] , \nRightOut_18[2] , 
        \nLeftOut_22[11] , \nLeftOut_74[10] , \nRightOut_30[13] , 
        \nRightOut_66[12] , \nLeftOut_72[5] , \nLeftOut_37[16] , 
        \nLeftOut_57[12] , \nRightOut_88[14] , \nLeftOut_16[1] , 
        \nRightOut_25[14] , \nRightOut_45[10] , \nRightOut_61[9] , 
        \nRightOut_73[15] , \nLeftOut_77[8] , \ScanLink19[4] , 
        \nLeftOut_4[14] , \nLeftOut_69[4] , \nRightOut_64[4] , 
        \nRightOut_0[13] , \ScanLink3[14] , \nRightOut_67[7] , 
        \nRightOut_4[11] , \ScanLink9[12] , \nRightOut_15[7] , 
        \nLeftOut_18[7] , \nRightOut_71[3] , \nRightOut_72[0] , 
        \ScanLink10[10] , \nRightOut_16[4] , \nRightOut_13[9] , 
        \nLeftOut_48[13] , \nRightOut_69[1] , \ScanLink26[15] , 
        \nLeftOut_64[1] , \nLeftOut_90[10] , \ScanLink17[2] , \ScanLink8[0] , 
        \nRightOut_8[2] , \ScanLink14[12] , \ScanLink14[1] , 
        \nRightOut_79[13] , \nRightOut_82[12] , \nRightOut_29[3] , 
        \nLeftOut_67[2] , \nLeftOut_91[2] , \nLeftOut_43[4] , \ScanLink30[7] , 
        \nLeftOut_27[0] , \nLeftOut_40[7] , \nLeftOut_81[15] , 
        \nRightOut_68[16] , \nLeftOut_92[1] , \nLeftOut_39[12] , 
        \nRightOut_50[8] , \nLeftOut_59[16] , \nRightOut_86[10] , 
        \ScanLink8[15] , \nLeftOut_9[0] , \nLeftOut_24[3] , \nLeftOut_94[12] , 
        \nRightOut_31[1] , \nRightOut_32[2] , \nLeftOut_58[5] , 
        \nLeftOut_46[9] , \nLeftOut_89[0] , \nRightOut_55[5] , 
        \nRightOut_56[6] , \ScanLink28[5] , \nRightOut_84[0] , 
        \nRightOut_87[3] , \nRightOut_61[4] , \nRightOut_62[7] , 
        \nLeftOut_72[8] , \nLeftOut_10[2] , \nLeftOut_84[10] , 
        \nLeftOut_13[1] , \nLeftOut_29[10] , \nLeftOut_49[14] , 
        \nRightOut_64[9] , \ScanLink27[12] , \nRightOut_5[16] , 
        \nLeftOut_74[6] , \nRightOut_79[6] , \nRightOut_18[10] , 
        \nLeftOut_69[9] , \nRightOut_78[14] , \ScanLink19[9] , 
        \nRightOut_0[7] , \nLeftOut_1[5] , \nLeftOut_2[6] , \nRightOut_39[4] , 
        \nLeftOut_77[5] , \nRightOut_83[15] , \nLeftOut_81[5] , 
        \nRightOut_92[10] , \ScanLink32[15] , \ScanLink23[10] , 
        \ScanLink15[15] , \nLeftOut_53[3] , \ScanLink20[0] , \nLeftOut_80[12] , 
        \nRightOut_1[14] , \ScanLink5[8] , \nRightOut_27[8] , \nLeftOut_50[0] , 
        \ScanLink23[3] , \nLeftOut_37[7] , \nRightOut_69[11] , 
        \nLeftOut_82[6] , \nLeftOut_38[15] , \nLeftOut_58[11] , 
        \nRightOut_92[9] , \ScanLink3[6] , \nLeftOut_4[8] , \nRightOut_6[9] , 
        \nLeftOut_34[4] , \nLeftOut_48[2] , \nLeftOut_95[15] , 
        \nRightOut_21[6] , \nRightOut_22[5] , \nLeftOut_84[8] , 
        \nRightOut_3[4] , \nLeftOut_31[9] , \nRightOut_46[1] , 
        \nRightOut_89[8] , \nRightOut_94[7] , \ScanLink0[5] , \ScanLink6[11] , 
        \nLeftOut_39[1] , \nRightOut_45[2] , \nRightOut_53[6] , 
        \nRightOut_50[5] , \nRightOut_81[0] , \nRightOut_82[3] , 
        \nRightOut_37[2] , \nLeftOut_1[11] , \nRightOut_34[1] , 
        \nLeftOut_43[9] , \ScanLink2[13] , \nLeftOut_5[13] , \nRightOut_10[7] , 
        \ScanLink11[1] , \nLeftOut_11[11] , \nLeftOut_22[0] , 
        \nLeftOut_27[14] , \nRightOut_35[16] , \nRightOut_48[7] , 
        \nRightOut_55[12] , \nRightOut_55[8] , \nLeftOut_71[15] , 
        \nLeftOut_47[10] , \ScanLink12[2] , \nRightOut_16[14] , 
        \nRightOut_20[11] , \nLeftOut_21[3] , \nLeftOut_94[2] , 
        \ScanLink28[8] , \nLeftOut_46[4] , \nRightOut_76[10] , 
        \nRightOut_16[9] , \nLeftOut_32[13] , \nRightOut_40[15] , 
        \nLeftOut_45[7] , \nLeftOut_58[8] , \nLeftOut_64[12] , 
        \nLeftOut_15[13] , \nLeftOut_43[12] , \nLeftOut_61[1] , 
        \nLeftOut_23[16] , \nRightOut_51[10] , \nRightOut_67[15] , 
        \nRightOut_12[16] , \nRightOut_31[14] , \nLeftOut_62[2] , 
        \nLeftOut_36[11] , \nLeftOut_56[15] , \nLeftOut_60[10] , 
        \nRightOut_89[13] , \nRightOut_24[13] , \nRightOut_72[12] , 
        \nRightOut_13[4] , \nLeftOut_79[3] , \nRightOut_74[3] , 
        \nRightOut_77[0] , \ScanLink3[10] , \nRightOut_4[15] , \ScanLink8[4] , 
        \nLeftOut_9[4] , \nRightOut_31[5] , \ScanLink28[1] , \nRightOut_32[6] , 
        \nLeftOut_89[4] , \nLeftOut_22[9] , \nRightOut_55[1] , 
        \nLeftOut_58[1] , \nLeftOut_24[7] , \nRightOut_29[7] , 
        \nRightOut_34[8] , \nLeftOut_40[3] , \nRightOut_56[2] , 
        \nRightOut_84[4] , \nRightOut_87[7] , \nRightOut_68[12] , 
        \nLeftOut_81[11] , \nLeftOut_92[5] , \nLeftOut_43[0] , 
        \ScanLink22[13] , \ScanLink30[3] , \nLeftOut_91[6] , 
        \nRightOut_93[13] , \nLeftOut_39[8] , \nRightOut_81[9] , 
        \nLeftOut_94[16] , \nRightOut_86[14] , \nRightOut_8[6] , 
        \ScanLink10[14] , \nLeftOut_27[4] , \nLeftOut_39[16] , 
        \nLeftOut_59[12] , \nLeftOut_28[13] , \nRightOut_69[5] , 
        \ScanLink26[11] , \ScanLink14[5] , \nRightOut_77[9] , 
        \nLeftOut_85[13] , \nRightOut_19[13] , \nLeftOut_67[6] , 
        \nRightOut_82[16] , \ScanLink11[8] , \nRightOut_16[0] , 
        \nLeftOut_18[3] , \nLeftOut_64[5] , \nLeftOut_90[14] , \ScanLink17[6] , 
        \nLeftOut_61[8] , \nRightOut_71[7] , \nRightOut_72[4] , 
        \nRightOut_15[3] , \nLeftOut_69[0] , \ScanLink19[0] , \nLeftOut_4[10] , 
        \nLeftOut_13[8] , \nRightOut_67[3] , \nRightOut_64[0] , 
        \nLeftOut_10[12] , \nRightOut_13[15] , \nLeftOut_14[10] , 
        \nRightOut_18[6] , \nRightOut_50[13] , \nRightOut_66[16] , 
        \nLeftOut_72[1] , \nLeftOut_22[15] , \nLeftOut_74[14] , 
        \nLeftOut_16[5] , \nRightOut_25[10] , \nLeftOut_42[11] , 
        \nLeftOut_71[2] , \nRightOut_73[11] , \nRightOut_45[14] , 
        \nLeftOut_15[6] , \nLeftOut_31[0] , \nLeftOut_37[12] , 
        \nLeftOut_61[13] , \nRightOut_88[10] , \nRightOut_46[8] , 
        \nLeftOut_57[16] , \nRightOut_89[1] , \nLeftOut_0[12] , 
        \nLeftOut_4[1] , \nLeftOut_32[3] , \nLeftOut_46[13] , 
        \nRightOut_54[11] , \nRightOut_58[4] , \nLeftOut_70[16] , 
        \ScanLink28[15] , \nLeftOut_33[10] , \nRightOut_34[15] , 
        \nLeftOut_53[14] , \nRightOut_62[14] , \nLeftOut_65[11] , 
        \nLeftOut_87[2] , \ScanLink5[1] , \nRightOut_5[3] , \nLeftOut_7[2] , 
        \nRightOut_41[16] , \nLeftOut_55[4] , \ScanLink26[7] , 
        \nRightOut_77[13] , \nRightOut_21[12] , \nRightOut_40[6] , 
        \nLeftOut_56[7] , \ScanLink25[4] , \nLeftOut_84[1] , \ScanLink6[2] , 
        \nLeftOut_29[2] , \nRightOut_91[3] , \nRightOut_92[0] , 
        \nRightOut_43[5] , \nRightOut_6[0] , \nLeftOut_4[12] , \ScanLink7[12] , 
        \nRightOut_24[2] , \nRightOut_27[1] , \ScanLink20[9] , 
        \nLeftOut_50[9] , \nLeftOut_69[2] , \ScanLink19[2] , \nRightOut_64[2] , 
        \nRightOut_67[1] , \nLeftOut_0[10] , \ScanLink3[12] , \nLeftOut_10[9] , 
        \nLeftOut_4[3] , \nLeftOut_7[0] , \nLeftOut_10[10] , \nLeftOut_14[12] , 
        \nLeftOut_71[0] , \nLeftOut_15[4] , \nRightOut_18[4] , 
        \nLeftOut_42[13] , \nLeftOut_74[16] , \nRightOut_30[15] , 
        \nRightOut_50[11] , \nLeftOut_37[10] , \nLeftOut_57[14] , 
        \nRightOut_66[14] , \nLeftOut_72[3] , \nLeftOut_61[11] , 
        \nLeftOut_16[7] , \nRightOut_45[16] , \nRightOut_88[12] , 
        \nRightOut_73[13] , \nRightOut_25[12] , \nLeftOut_26[15] , 
        \nLeftOut_32[1] , \nRightOut_45[9] , \nRightOut_62[16] , 
        \nRightOut_54[13] , \nRightOut_58[6] , \nLeftOut_70[14] , 
        \nRightOut_21[10] , \nLeftOut_31[2] , \nLeftOut_46[11] , 
        \nLeftOut_56[5] , \nRightOut_77[11] , \nLeftOut_84[3] , 
        \nRightOut_89[3] , \ScanLink25[6] , \nRightOut_17[15] , 
        \nRightOut_41[14] , \nLeftOut_55[6] , \ScanLink26[5] , \ScanLink5[3] , 
        \nRightOut_5[1] , \ScanLink6[0] , \nLeftOut_33[12] , \nLeftOut_48[9] , 
        \nLeftOut_87[0] , \nLeftOut_65[13] , \nLeftOut_53[16] , 
        \nRightOut_6[2] , \nLeftOut_29[0] , \nRightOut_43[7] , 
        \nRightOut_91[1] , \nRightOut_92[2] , \ScanLink7[10] , 
        \nRightOut_40[4] , \nRightOut_24[0] , \nRightOut_27[3] , 
        \ScanLink23[8] , \nLeftOut_53[8] , \nLeftOut_9[6] , \nLeftOut_58[3] , 
        \nLeftOut_21[8] , \nRightOut_31[7] , \nRightOut_32[4] , 
        \nLeftOut_89[6] , \nLeftOut_94[9] , \ScanLink28[3] , \nRightOut_29[5] , 
        \nRightOut_55[3] , \nRightOut_56[0] , \nRightOut_84[6] , 
        \nRightOut_87[5] , \nLeftOut_91[4] , \nRightOut_93[11] , 
        \nRightOut_0[15] , \ScanLink8[6] , \ScanLink14[14] , \nLeftOut_43[2] , 
        \ScanLink22[11] , \ScanLink30[1] , \nLeftOut_27[6] , \nRightOut_37[9] , 
        \nLeftOut_40[1] , \nLeftOut_81[13] , \nLeftOut_39[14] , 
        \nRightOut_68[10] , \nLeftOut_92[7] , \nLeftOut_59[10] , 
        \nRightOut_8[4] , \nRightOut_86[16] , \nRightOut_82[8] , 
        \nLeftOut_1[13] , \ScanLink9[14] , \ScanLink14[7] , \nRightOut_19[11] , 
        \nLeftOut_24[5] , \nLeftOut_94[14] , \nLeftOut_28[11] , 
        \nLeftOut_48[15] , \nRightOut_74[8] , \nLeftOut_85[11] , 
        \ScanLink26[13] , \nLeftOut_64[7] , \nRightOut_69[7] , 
        \nLeftOut_90[16] , \ScanLink17[4] , \nLeftOut_67[4] , \nLeftOut_79[8] , 
        \nRightOut_79[15] , \nRightOut_82[14] , \nRightOut_15[1] , 
        \nLeftOut_18[1] , \nRightOut_71[5] , \nRightOut_72[6] , 
        \ScanLink12[9] , \nRightOut_16[2] , \nLeftOut_62[9] , \nLeftOut_39[3] , 
        \nRightOut_50[7] , \nRightOut_81[2] , \nRightOut_82[1] , 
        \nRightOut_53[4] , \nRightOut_34[3] , \ScanLink6[13] , 
        \nRightOut_37[0] , \ScanLink30[8] , \nLeftOut_40[8] , 
        \nLeftOut_11[13] , \nLeftOut_21[1] , \nRightOut_56[9] , 
        \nLeftOut_47[12] , \nLeftOut_22[2] , \nLeftOut_27[16] , 
        \ScanLink29[14] , \nRightOut_35[14] , \nRightOut_48[5] , 
        \nRightOut_55[10] , \nRightOut_63[15] , \nLeftOut_52[15] , 
        \ScanLink2[11] , \nRightOut_10[5] , \ScanLink11[3] , 
        \nRightOut_16[16] , \nLeftOut_32[11] , \nLeftOut_45[5] , 
        \nLeftOut_64[10] , \nRightOut_20[13] , \nLeftOut_46[6] , 
        \nRightOut_31[16] , \nRightOut_76[12] , \nLeftOut_94[0] , 
        \nLeftOut_62[0] , \ScanLink12[0] , \nLeftOut_15[11] , 
        \nRightOut_15[8] , \nRightOut_51[12] , \nLeftOut_23[14] , 
        \nLeftOut_75[15] , \nLeftOut_43[10] , \nLeftOut_61[3] , 
        \nRightOut_12[14] , \nRightOut_24[11] , \nRightOut_72[10] , 
        \nRightOut_13[6] , \nLeftOut_18[8] , \nLeftOut_36[13] , 
        \nRightOut_44[15] , \nRightOut_89[11] , \nLeftOut_60[12] , 
        \nLeftOut_79[1] , \nLeftOut_5[11] , \nRightOut_74[1] , 
        \nRightOut_77[2] , \nRightOut_61[6] , \nRightOut_62[5] , 
        \nLeftOut_71[9] , \nLeftOut_10[0] , \ScanLink11[15] , \nLeftOut_13[3] , 
        \nLeftOut_29[12] , \nRightOut_79[4] , \nLeftOut_49[16] , 
        \ScanLink27[10] , \nRightOut_67[8] , \nLeftOut_84[12] , 
        \nLeftOut_77[7] , \nLeftOut_0[14] , \nRightOut_0[11] , 
        \nRightOut_0[5] , \nLeftOut_1[7] , \nRightOut_5[14] , 
        \nRightOut_78[16] , \nRightOut_18[12] , \nLeftOut_50[2] , 
        \nRightOut_69[13] , \nLeftOut_74[4] , \nLeftOut_82[4] , 
        \nLeftOut_91[15] , \ScanLink23[1] , \nRightOut_1[16] , \nLeftOut_2[4] , 
        \nRightOut_24[9] , \nLeftOut_80[10] , \nLeftOut_53[1] , 
        \ScanLink20[2] , \ScanLink23[12] , \ScanLink6[9] , \nRightOut_39[6] , 
        \nLeftOut_81[7] , \nRightOut_92[12] , \nLeftOut_34[6] , 
        \nRightOut_5[8] , \nLeftOut_29[9] , \nRightOut_91[8] , 
        \nLeftOut_37[5] , \nLeftOut_58[13] , \nRightOut_87[15] , 
        \nLeftOut_7[9] , \nRightOut_21[4] , \nRightOut_22[7] , 
        \nLeftOut_32[8] , \nRightOut_45[0] , \nLeftOut_48[0] , 
        \nLeftOut_87[9] , \ScanLink0[7] , \ScanLink3[4] , \nRightOut_46[3] , 
        \nRightOut_94[5] , \nRightOut_3[6] , \nRightOut_4[13] , 
        \ScanLink9[10] , \nRightOut_16[6] , \nLeftOut_18[5] , 
        \nRightOut_71[1] , \nRightOut_72[2] , \ScanLink10[12] , 
        \nRightOut_15[5] , \nLeftOut_28[15] , \nRightOut_69[3] , 
        \nLeftOut_48[11] , \nRightOut_10[8] , \ScanLink14[3] , 
        \nLeftOut_67[0] , \nLeftOut_85[15] , \nRightOut_79[11] , 
        \nRightOut_82[10] , \ScanLink14[10] , \nRightOut_19[15] , 
        \nLeftOut_40[5] , \nLeftOut_64[3] , \nRightOut_68[14] , 
        \nLeftOut_90[12] , \nLeftOut_92[3] , \ScanLink17[0] , \nLeftOut_24[1] , 
        \nRightOut_29[1] , \nLeftOut_43[6] , \ScanLink22[15] , \ScanLink30[5] , 
        \nRightOut_53[9] , \nLeftOut_91[0] , \nRightOut_93[15] , 
        \nLeftOut_94[10] , \ScanLink5[7] , \ScanLink8[2] , \nRightOut_8[0] , 
        \nLeftOut_9[2] , \nLeftOut_27[2] , \nLeftOut_59[14] , 
        \nRightOut_86[12] , \nRightOut_31[3] , \nLeftOut_39[10] , 
        \ScanLink28[7] , \nRightOut_32[0] , \nLeftOut_89[2] , \nLeftOut_45[8] , 
        \nLeftOut_58[7] , \nRightOut_40[0] , \nRightOut_48[8] , 
        \nRightOut_55[7] , \nRightOut_56[4] , \nRightOut_84[2] , 
        \nRightOut_87[1] , \nRightOut_5[5] , \nLeftOut_37[8] , \ScanLink6[4] , 
        \nRightOut_6[6] , \nLeftOut_29[4] , \nRightOut_91[5] , 
        \nRightOut_92[6] , \nRightOut_43[3] , \nRightOut_0[8] , 
        \nLeftOut_2[9] , \nRightOut_24[4] , \ScanLink3[9] , \ScanLink7[14] , 
        \nRightOut_27[7] , \nLeftOut_31[6] , \nLeftOut_82[9] , 
        \nRightOut_89[7] , \nLeftOut_10[14] , \nLeftOut_46[15] , 
        \nRightOut_94[8] , \nLeftOut_26[11] , \nLeftOut_70[10] , 
        \ScanLink28[13] , \nLeftOut_32[5] , \nRightOut_34[13] , 
        \nRightOut_58[2] , \nRightOut_62[12] , \nLeftOut_4[7] , 
        \nLeftOut_33[16] , \nLeftOut_53[12] , \nLeftOut_55[2] , 
        \nLeftOut_87[4] , \ScanLink26[1] , \nLeftOut_7[4] , \nRightOut_17[11] , 
        \nRightOut_21[9] , \nRightOut_21[14] , \nRightOut_41[10] , 
        \nLeftOut_56[1] , \ScanLink25[2] , \nRightOut_13[13] , 
        \nLeftOut_14[16] , \nRightOut_18[0] , \nRightOut_30[11] , 
        \nRightOut_66[10] , \nRightOut_77[15] , \nLeftOut_84[7] , 
        \nRightOut_50[15] , \nLeftOut_72[7] , \nLeftOut_22[13] , 
        \nLeftOut_74[12] , \nLeftOut_16[3] , \nLeftOut_71[4] , 
        \nRightOut_25[16] , \nLeftOut_15[0] , \nRightOut_45[12] , 
        \nRightOut_88[16] , \nLeftOut_37[14] , \nRightOut_62[8] , 
        \nLeftOut_57[10] , \nLeftOut_61[15] , \nRightOut_67[5] , 
        \nLeftOut_69[6] , \nLeftOut_74[9] , \ScanLink19[6] , \nLeftOut_4[16] , 
        \nRightOut_64[6] , \nRightOut_79[9] , \nRightOut_0[1] , \ScanLink0[3] , 
        \ScanLink3[0] , \nRightOut_3[2] , \nRightOut_21[0] , \nRightOut_22[3] , 
        \nLeftOut_48[4] , \ScanLink26[8] , \nLeftOut_56[8] , \nRightOut_46[7] , 
        \nRightOut_94[1] , \nLeftOut_1[3] , \nLeftOut_2[0] , \nRightOut_39[2] , 
        \nRightOut_45[4] , \nLeftOut_81[3] , \nRightOut_92[16] , 
        \nLeftOut_53[5] , \ScanLink20[6] , \ScanLink15[13] , \nLeftOut_50[6] , 
        \nLeftOut_80[14] , \ScanLink23[5] , \nRightOut_1[12] , 
        \nLeftOut_37[1] , \nLeftOut_38[13] , \nLeftOut_82[0] , 
        \nRightOut_40[9] , \nRightOut_87[11] , \nLeftOut_34[2] , 
        \nLeftOut_95[13] , \nLeftOut_10[4] , \ScanLink11[11] , 
        \nLeftOut_49[12] , \nLeftOut_84[16] , \nLeftOut_13[7] , 
        \nLeftOut_29[16] , \ScanLink27[14] , \nRightOut_79[0] , 
        \nRightOut_5[10] , \nRightOut_18[16] , \nLeftOut_74[0] , 
        \nLeftOut_91[11] , \nRightOut_78[12] , \nRightOut_83[13] , 
        \ScanLink2[15] , \nLeftOut_5[15] , \ScanLink8[13] , \nLeftOut_15[9] , 
        \nRightOut_61[2] , \nLeftOut_77[3] , \ScanLink32[13] , 
        \nRightOut_62[1] , \nRightOut_10[1] , \nRightOut_18[9] , 
        \nRightOut_13[2] , \nLeftOut_67[9] , \nLeftOut_79[5] , \ScanLink17[9] , 
        \nRightOut_74[5] , \nRightOut_77[6] , \nRightOut_8[9] , 
        \ScanLink11[7] , \ScanLink12[4] , \nLeftOut_61[7] , \nLeftOut_15[15] , 
        \nLeftOut_23[10] , \nLeftOut_43[14] , \nRightOut_31[12] , 
        \nRightOut_51[16] , \nLeftOut_75[11] , \nLeftOut_62[4] , 
        \nRightOut_12[10] , \nRightOut_44[11] , \nLeftOut_56[13] , 
        \nRightOut_67[13] , \nLeftOut_60[16] , \nRightOut_89[15] , 
        \nRightOut_71[8] , \nRightOut_16[12] , \nLeftOut_21[5] , 
        \nLeftOut_22[6] , \nRightOut_24[15] , \nRightOut_72[14] , 
        \nRightOut_35[10] , \nLeftOut_27[12] , \nRightOut_48[1] , 
        \nRightOut_55[14] , \nRightOut_63[11] , \nRightOut_87[8] , 
        \nLeftOut_47[16] , \nLeftOut_71[13] , \ScanLink29[10] , 
        \nRightOut_40[13] , \nLeftOut_46[2] , \nRightOut_76[16] , 
        \nLeftOut_94[4] , \nLeftOut_24[8] , \nLeftOut_32[15] , 
        \nRightOut_32[9] , \nLeftOut_45[1] , \nLeftOut_64[14] , 
        \nLeftOut_52[11] , \nLeftOut_39[7] , \nRightOut_53[0] , 
        \nRightOut_81[6] , \nRightOut_37[4] , \nRightOut_50[3] , 
        \nRightOut_82[5] , \nLeftOut_0[15] , \nRightOut_0[10] , 
        \nRightOut_4[12] , \ScanLink10[13] , \nRightOut_29[8] , 
        \nRightOut_34[7] , \nLeftOut_91[9] , \nLeftOut_48[10] , 
        \nRightOut_69[2] , \nLeftOut_85[14] , \nRightOut_19[14] , 
        \nLeftOut_28[14] , \ScanLink8[3] , \ScanLink9[11] , \nRightOut_10[9] , 
        \nLeftOut_64[2] , \nRightOut_79[10] , \nLeftOut_90[13] , 
        \ScanLink17[1] , \ScanLink14[2] , \nLeftOut_67[1] , \nRightOut_15[4] , 
        \nLeftOut_18[4] , \nRightOut_71[0] , \nRightOut_82[11] , 
        \nRightOut_72[3] , \nLeftOut_9[3] , \nRightOut_16[7] , 
        \nRightOut_32[1] , \nLeftOut_45[9] , \nLeftOut_58[6] , 
        \ScanLink14[11] , \nRightOut_31[2] , \nLeftOut_89[3] , \ScanLink28[6] , 
        \nLeftOut_43[7] , \nRightOut_48[9] , \nRightOut_55[6] , 
        \nRightOut_56[5] , \nRightOut_84[3] , \nRightOut_87[0] , 
        \ScanLink22[14] , \ScanLink30[4] , \nRightOut_29[0] , \nLeftOut_91[1] , 
        \nRightOut_93[14] , \nLeftOut_40[4] , \nRightOut_68[15] , 
        \nLeftOut_92[2] , \nLeftOut_81[16] , \nRightOut_8[1] , 
        \nRightOut_86[13] , \nLeftOut_24[0] , \nLeftOut_27[3] , 
        \nLeftOut_39[11] , \nLeftOut_59[15] , \nRightOut_53[8] , 
        \nLeftOut_94[11] , \nRightOut_0[9] , \nLeftOut_32[4] , 
        \nRightOut_34[12] , \nRightOut_58[3] , \ScanLink3[8] , 
        \nRightOut_54[16] , \nRightOut_62[13] , \nLeftOut_4[6] , 
        \nLeftOut_7[5] , \nLeftOut_10[15] , \nLeftOut_26[10] , 
        \nLeftOut_31[7] , \nRightOut_89[6] , \nLeftOut_70[11] , 
        \ScanLink28[12] , \nRightOut_21[15] , \nLeftOut_46[14] , 
        \nLeftOut_56[0] , \nRightOut_77[14] , \nRightOut_94[9] , 
        \ScanLink25[3] , \nRightOut_17[10] , \nRightOut_21[8] , 
        \nRightOut_41[11] , \nLeftOut_53[13] , \nLeftOut_65[16] , 
        \nLeftOut_84[6] , \nLeftOut_87[5] , \nLeftOut_55[3] , \ScanLink26[0] , 
        \ScanLink5[6] , \nRightOut_5[4] , \ScanLink6[5] , \nLeftOut_29[5] , 
        \nRightOut_91[4] , \nRightOut_6[7] , \nLeftOut_37[9] , 
        \nRightOut_43[2] , \ScanLink7[15] , \nRightOut_27[6] , 
        \nRightOut_40[1] , \nRightOut_92[7] , \nLeftOut_82[8] , 
        \nLeftOut_2[8] , \nRightOut_24[5] , \nRightOut_64[7] , 
        \nLeftOut_69[7] , \nLeftOut_74[8] , \ScanLink19[7] , \nRightOut_67[4] , 
        \nRightOut_79[8] , \nRightOut_0[0] , \nLeftOut_1[2] , 
        \nRightOut_13[12] , \nLeftOut_15[1] , \nRightOut_18[1] , 
        \nLeftOut_22[12] , \nLeftOut_42[16] , \nRightOut_30[10] , 
        \nRightOut_50[14] , \nLeftOut_71[5] , \nLeftOut_74[13] , 
        \nRightOut_66[11] , \nLeftOut_72[6] , \nRightOut_62[9] , 
        \nLeftOut_37[15] , \nLeftOut_57[11] , \nLeftOut_61[14] , 
        \nRightOut_45[13] , \nLeftOut_16[2] , \nRightOut_73[16] , 
        \nLeftOut_50[7] , \ScanLink23[4] , \nRightOut_1[13] , \nLeftOut_2[1] , 
        \ScanLink15[12] , \nRightOut_39[3] , \nRightOut_69[16] , 
        \nLeftOut_80[15] , \nLeftOut_82[1] , \nLeftOut_81[2] , 
        \nLeftOut_53[4] , \ScanLink20[7] , \nRightOut_21[1] , \nLeftOut_34[3] , 
        \nLeftOut_37[0] , \nRightOut_40[8] , \nLeftOut_95[12] , 
        \nLeftOut_58[16] , \nLeftOut_38[12] , \nRightOut_87[10] , 
        \nRightOut_22[2] , \nLeftOut_48[5] , \nLeftOut_56[9] , 
        \nRightOut_45[5] , \ScanLink26[9] , \ScanLink0[2] , \ScanLink3[1] , 
        \nRightOut_46[6] , \nRightOut_3[3] , \ScanLink8[12] , \nLeftOut_15[8] , 
        \nRightOut_94[0] , \nRightOut_61[3] , \nRightOut_62[0] , 
        \ScanLink11[10] , \nLeftOut_13[6] , \nRightOut_18[8] , 
        \nLeftOut_49[13] , \ScanLink27[15] , \nLeftOut_10[5] , 
        \nRightOut_79[1] , \ScanLink2[14] , \nRightOut_5[11] , 
        \nLeftOut_74[1] , \nLeftOut_77[2] , \nRightOut_83[12] , 
        \ScanLink32[12] , \nLeftOut_91[10] , \nRightOut_78[13] , 
        \nRightOut_10[0] , \ScanLink11[6] , \nRightOut_31[13] , 
        \nRightOut_67[12] , \nLeftOut_62[5] , \ScanLink12[5] , 
        \nLeftOut_61[6] , \nRightOut_12[11] , \nLeftOut_15[14] , 
        \nLeftOut_23[11] , \nLeftOut_75[10] , \nLeftOut_43[15] , 
        \nRightOut_24[14] , \nRightOut_71[9] , \nRightOut_72[15] , 
        \nRightOut_13[3] , \nLeftOut_36[16] , \nRightOut_44[10] , 
        \nLeftOut_56[12] , \nLeftOut_79[4] , \nRightOut_89[14] , 
        \ScanLink17[8] , \nLeftOut_67[8] , \nRightOut_77[7] , \nLeftOut_5[14] , 
        \nRightOut_8[8] , \nRightOut_74[4] , \nRightOut_82[4] , 
        \nLeftOut_24[9] , \nRightOut_50[2] , \nRightOut_53[1] , 
        \nRightOut_34[6] , \nLeftOut_39[6] , \nRightOut_81[7] , 
        \nLeftOut_1[16] , \nRightOut_29[9] , \nLeftOut_91[8] , 
        \nLeftOut_10[8] , \nLeftOut_11[16] , \nRightOut_37[5] , 
        \nRightOut_13[16] , \nLeftOut_14[13] , \nRightOut_16[13] , 
        \nLeftOut_21[4] , \nLeftOut_27[13] , \nLeftOut_71[12] , 
        \ScanLink29[11] , \nLeftOut_22[7] , \nRightOut_35[11] , 
        \nRightOut_55[15] , \nRightOut_63[10] , \nLeftOut_32[14] , 
        \nRightOut_32[8] , \nRightOut_48[0] , \nRightOut_87[9] , 
        \nLeftOut_45[0] , \nLeftOut_52[10] , \nLeftOut_64[15] , 
        \nLeftOut_94[5] , \nRightOut_18[5] , \nRightOut_20[16] , 
        \nRightOut_40[12] , \nLeftOut_46[3] , \nLeftOut_22[16] , 
        \nRightOut_30[14] , \nRightOut_66[15] , \nRightOut_50[10] , 
        \nLeftOut_72[2] , \nLeftOut_71[1] , \nLeftOut_42[12] , 
        \nLeftOut_16[6] , \nRightOut_25[13] , \nRightOut_73[12] , 
        \nLeftOut_15[5] , \nLeftOut_37[11] , \nLeftOut_57[15] , 
        \nLeftOut_61[10] , \nRightOut_88[13] , \nLeftOut_69[3] , 
        \ScanLink19[3] , \nRightOut_67[0] , \nLeftOut_0[11] , \ScanLink3[13] , 
        \nLeftOut_4[13] , \ScanLink5[2] , \nRightOut_40[5] , \nRightOut_64[3] , 
        \nRightOut_92[3] , \nRightOut_5[0] , \ScanLink6[1] , \nRightOut_6[3] , 
        \nRightOut_43[6] , \nRightOut_24[1] , \nLeftOut_29[1] , 
        \nRightOut_91[0] , \nLeftOut_53[9] , \nLeftOut_4[2] , \ScanLink7[11] , 
        \nLeftOut_10[11] , \nRightOut_27[2] , \nLeftOut_46[10] , 
        \ScanLink23[9] , \nLeftOut_26[14] , \nLeftOut_70[15] , 
        \nLeftOut_31[3] , \nRightOut_89[2] , \nLeftOut_32[0] , 
        \nRightOut_34[16] , \nRightOut_45[8] , \nRightOut_54[12] , 
        \nLeftOut_55[7] , \nRightOut_58[7] , \ScanLink26[4] , \nLeftOut_7[1] , 
        \nRightOut_17[14] , \nLeftOut_33[13] , \nLeftOut_48[8] , 
        \nLeftOut_65[12] , \nLeftOut_87[1] , \nLeftOut_84[2] , 
        \nRightOut_21[11] , \nRightOut_41[15] , \nLeftOut_56[4] , 
        \ScanLink25[7] , \ScanLink14[15] , \nRightOut_29[4] , 
        \nRightOut_37[8] , \nRightOut_77[10] , \nLeftOut_40[0] , 
        \nRightOut_68[11] , \nLeftOut_81[12] , \nLeftOut_92[6] , 
        \nLeftOut_91[5] , \nRightOut_93[10] , \nLeftOut_43[3] , 
        \nRightOut_0[14] , \ScanLink22[10] , \ScanLink30[0] , \nLeftOut_1[12] , 
        \nRightOut_4[16] , \ScanLink8[7] , \nRightOut_8[5] , \nLeftOut_24[4] , 
        \nLeftOut_27[7] , \nLeftOut_59[11] , \nLeftOut_94[15] , 
        \nLeftOut_39[15] , \nRightOut_82[9] , \ScanLink9[15] , \nLeftOut_9[7] , 
        \nRightOut_31[6] , \nLeftOut_58[2] , \nLeftOut_89[7] , 
        \nLeftOut_94[8] , \ScanLink28[2] , \ScanLink12[8] , \nLeftOut_18[0] , 
        \nLeftOut_21[9] , \nRightOut_32[5] , \nRightOut_55[2] , 
        \nRightOut_87[4] , \nRightOut_56[1] , \nRightOut_72[7] , 
        \nRightOut_84[7] , \nRightOut_71[4] , \nRightOut_16[3] , 
        \nLeftOut_62[8] , \ScanLink14[6] , \nRightOut_15[0] , 
        \nLeftOut_28[10] , \nLeftOut_48[14] , \ScanLink26[12] , 
        \nLeftOut_67[5] , \nRightOut_69[6] , \nRightOut_74[9] , 
        \nRightOut_82[15] , \nLeftOut_85[10] , \nLeftOut_64[6] , 
        \nLeftOut_79[9] , \nRightOut_79[14] , \ScanLink17[5] , \ScanLink6[12] , 
        \nLeftOut_11[12] , \nRightOut_19[10] , \nLeftOut_21[0] , 
        \nLeftOut_22[3] , \nRightOut_35[15] , \nRightOut_48[4] , 
        \nRightOut_55[11] , \nRightOut_63[14] , \nRightOut_56[8] , 
        \nLeftOut_71[16] , \ScanLink29[15] , \nRightOut_20[12] , 
        \nLeftOut_46[7] , \nLeftOut_47[13] , \nRightOut_76[13] , 
        \nLeftOut_32[10] , \nRightOut_40[16] , \nLeftOut_64[11] , 
        \nLeftOut_94[1] , \nRightOut_37[1] , \nLeftOut_39[2] , 
        \nLeftOut_45[4] , \nLeftOut_52[14] , \nLeftOut_40[9] , 
        \nRightOut_50[6] , \nRightOut_53[5] , \nRightOut_81[3] , 
        \nRightOut_82[0] , \ScanLink2[10] , \nLeftOut_5[10] , 
        \nRightOut_10[4] , \nRightOut_34[2] , \ScanLink30[9] , 
        \nRightOut_13[7] , \nRightOut_74[0] , \nLeftOut_79[0] , 
        \nLeftOut_10[1] , \ScanLink11[2] , \ScanLink12[1] , \nLeftOut_15[10] , 
        \nRightOut_77[3] , \nLeftOut_23[15] , \nLeftOut_43[11] , 
        \nLeftOut_61[2] , \nLeftOut_75[14] , \nRightOut_15[9] , 
        \nRightOut_51[13] , \nLeftOut_62[1] , \nRightOut_12[15] , 
        \nLeftOut_18[9] , \nLeftOut_56[16] , \nRightOut_67[16] , 
        \nRightOut_89[10] , \nLeftOut_36[12] , \nLeftOut_60[13] , 
        \nRightOut_44[14] , \nRightOut_24[10] , \nRightOut_72[11] , 
        \nRightOut_67[9] , \nRightOut_79[5] , \nLeftOut_84[13] , 
        \nRightOut_5[15] , \ScanLink11[14] , \nLeftOut_13[2] , 
        \nRightOut_18[13] , \nLeftOut_29[13] , \ScanLink27[11] , 
        \nLeftOut_74[5] , \nLeftOut_91[14] , \nLeftOut_77[6] , 
        \nRightOut_83[16] , \nRightOut_0[4] , \ScanLink0[6] , \ScanLink3[5] , 
        \nRightOut_3[7] , \nLeftOut_7[8] , \nRightOut_22[6] , 
        \nRightOut_61[7] , \nRightOut_62[4] , \nLeftOut_71[8] , 
        \nLeftOut_48[1] , \nLeftOut_87[8] , \nRightOut_21[5] , 
        \nRightOut_94[4] , \nRightOut_46[2] , \nLeftOut_32[9] , 
        \nLeftOut_1[6] , \nLeftOut_2[5] , \nRightOut_45[1] , \nLeftOut_53[0] , 
        \ScanLink20[3] , \nRightOut_24[8] , \ScanLink23[13] , 
        \nRightOut_39[7] , \nLeftOut_81[6] , \nRightOut_92[13] , 
        \nLeftOut_50[3] , \nRightOut_69[12] , \nLeftOut_82[5] , 
        \nLeftOut_80[11] , \ScanLink23[0] , \nRightOut_5[9] , \nLeftOut_37[4] , 
        \nLeftOut_38[16] , \nRightOut_87[14] , \ScanLink6[8] , 
        \nLeftOut_34[7] , \nLeftOut_58[12] , \nLeftOut_95[16] , 
        \nLeftOut_13[0] , \nLeftOut_29[8] , \nRightOut_91[9] , 
        \ScanLink27[13] , \nLeftOut_29[11] , \nLeftOut_49[15] , 
        \nRightOut_64[8] , \nRightOut_79[7] , \nLeftOut_10[3] , 
        \nLeftOut_84[11] , \nRightOut_83[14] , \nRightOut_0[6] , 
        \ScanLink0[4] , \nLeftOut_4[9] , \ScanLink8[14] , \nRightOut_18[11] , 
        \nLeftOut_69[8] , \nLeftOut_74[7] , \nLeftOut_77[4] , \ScanLink19[8] , 
        \ScanLink32[14] , \nLeftOut_91[16] , \nRightOut_78[15] , 
        \nRightOut_61[5] , \nRightOut_62[6] , \nRightOut_21[7] , 
        \nLeftOut_72[9] , \nRightOut_22[4] , \nLeftOut_48[3] , 
        \nLeftOut_84[9] , \nRightOut_45[3] , \nLeftOut_1[4] , \ScanLink3[7] , 
        \nRightOut_3[5] , \nRightOut_46[0] , \nRightOut_89[9] , 
        \nLeftOut_31[8] , \nRightOut_27[9] , \nRightOut_94[6] , 
        \nRightOut_1[15] , \nLeftOut_2[7] , \ScanLink15[14] , 
        \nRightOut_39[5] , \nLeftOut_50[1] , \nLeftOut_80[13] , 
        \ScanLink23[2] , \nRightOut_69[10] , \nLeftOut_82[7] , 
        \nLeftOut_81[4] , \nRightOut_92[11] , \nLeftOut_53[2] , 
        \ScanLink20[1] , \ScanLink23[11] , \ScanLink5[9] , \nRightOut_6[8] , 
        \nLeftOut_34[5] , \nLeftOut_95[14] , \nLeftOut_38[14] , 
        \nLeftOut_58[10] , \nLeftOut_11[10] , \nLeftOut_37[6] , 
        \nRightOut_87[16] , \nRightOut_92[8] , \nRightOut_16[15] , 
        \nLeftOut_21[2] , \nLeftOut_27[15] , \nLeftOut_47[11] , 
        \nLeftOut_71[14] , \nLeftOut_22[1] , \nRightOut_55[13] , 
        \nRightOut_55[9] , \nLeftOut_32[12] , \nLeftOut_45[6] , 
        \nRightOut_48[6] , \nRightOut_63[16] , \nLeftOut_52[16] , 
        \nLeftOut_58[9] , \nLeftOut_64[13] , \nRightOut_40[14] , 
        \nLeftOut_94[3] , \ScanLink28[9] , \nRightOut_20[10] , 
        \nRightOut_76[11] , \nRightOut_34[0] , \nLeftOut_39[0] , 
        \nLeftOut_46[5] , \nRightOut_50[4] , \nRightOut_82[2] , 
        \nRightOut_53[7] , \nRightOut_81[1] , \nLeftOut_43[8] , 
        \nRightOut_0[16] , \nLeftOut_1[10] , \ScanLink2[12] , \ScanLink6[10] , 
        \nRightOut_10[6] , \nRightOut_13[5] , \nRightOut_37[3] , 
        \nLeftOut_79[2] , \nRightOut_77[1] , \nLeftOut_5[12] , \ScanLink8[5] , 
        \nRightOut_8[7] , \ScanLink11[0] , \nRightOut_74[2] , \ScanLink12[3] , 
        \nRightOut_31[15] , \nLeftOut_62[3] , \nRightOut_51[11] , 
        \nRightOut_67[14] , \nLeftOut_15[12] , \nRightOut_16[8] , 
        \nLeftOut_61[0] , \nLeftOut_75[16] , \nRightOut_24[12] , 
        \nLeftOut_43[13] , \nRightOut_72[13] , \nRightOut_29[6] , 
        \nRightOut_34[9] , \nLeftOut_36[10] , \nRightOut_44[16] , 
        \nLeftOut_60[11] , \nLeftOut_43[1] , \nLeftOut_56[14] , 
        \nRightOut_89[12] , \ScanLink22[12] , \ScanLink30[2] , 
        \nLeftOut_91[7] , \nRightOut_93[12] , \nLeftOut_40[2] , 
        \nRightOut_68[13] , \nLeftOut_92[4] , \nLeftOut_81[10] , 
        \nRightOut_86[15] , \nLeftOut_24[6] , \nLeftOut_27[5] , 
        \nLeftOut_59[13] , \nLeftOut_39[9] , \nRightOut_4[14] , 
        \nLeftOut_9[5] , \nRightOut_32[7] , \nRightOut_81[8] , 
        \ScanLink10[15] , \ScanLink11[9] , \nRightOut_15[2] , \nLeftOut_18[2] , 
        \nLeftOut_22[8] , \nRightOut_31[4] , \nLeftOut_58[0] , 
        \nLeftOut_89[5] , \ScanLink28[0] , \nRightOut_56[3] , 
        \nRightOut_84[5] , \nRightOut_55[0] , \nRightOut_71[6] , 
        \nRightOut_87[6] , \nRightOut_72[5] , \nRightOut_16[1] , 
        \nLeftOut_61[9] , \nRightOut_69[4] , \nRightOut_77[8] , 
        \nLeftOut_85[12] , \nLeftOut_28[12] , \nLeftOut_48[16] , 
        \ScanLink26[10] , \ScanLink14[4] , \nRightOut_19[12] , 
        \nLeftOut_64[4] , \nRightOut_79[16] , \ScanLink17[7] , 
        \nLeftOut_90[15] , \nLeftOut_14[11] , \nLeftOut_42[10] , 
        \nLeftOut_67[7] , \nLeftOut_22[14] , \nLeftOut_74[15] , 
        \nRightOut_30[16] , \nRightOut_50[12] , \nLeftOut_71[3] , 
        \nLeftOut_72[0] , \ScanLink3[11] , \nLeftOut_4[11] , \nLeftOut_13[9] , 
        \nRightOut_13[14] , \nLeftOut_15[7] , \nRightOut_18[7] , 
        \nRightOut_88[11] , \nLeftOut_37[13] , \nLeftOut_61[12] , 
        \nLeftOut_16[4] , \nRightOut_25[11] , \nRightOut_45[15] , 
        \nRightOut_64[1] , \nLeftOut_69[1] , \nRightOut_73[10] , 
        \ScanLink19[1] , \nLeftOut_0[13] , \ScanLink5[0] , \ScanLink6[3] , 
        \nRightOut_6[1] , \nLeftOut_29[3] , \nRightOut_67[2] , 
        \nRightOut_91[2] , \nRightOut_43[4] , \nRightOut_5[2] , 
        \ScanLink7[13] , \nRightOut_27[0] , \nRightOut_40[7] , 
        \nLeftOut_50[8] , \nRightOut_92[1] , \nLeftOut_1[14] , \nLeftOut_4[0] , 
        \nLeftOut_7[3] , \nLeftOut_10[13] , \nRightOut_24[3] , \ScanLink20[8] , 
        \nLeftOut_26[16] , \nLeftOut_31[1] , \nLeftOut_32[2] , 
        \nRightOut_58[5] , \nRightOut_62[15] , \nRightOut_34[14] , 
        \nRightOut_54[10] , \nRightOut_46[9] , \nRightOut_89[0] , 
        \ScanLink28[14] , \nLeftOut_46[12] , \nRightOut_17[16] , 
        \nRightOut_21[13] , \ScanLink25[5] , \nLeftOut_56[6] , 
        \nRightOut_77[12] , \nLeftOut_33[11] , \nLeftOut_84[0] , 
        \nLeftOut_53[15] , \nLeftOut_65[10] , \nLeftOut_87[3] , 
        \nLeftOut_5[16] , \nRightOut_10[2] , \ScanLink11[4] , \ScanLink12[7] , 
        \nLeftOut_15[16] , \nLeftOut_55[5] , \ScanLink26[6] , 
        \nLeftOut_23[13] , \nLeftOut_75[12] , \nRightOut_51[15] , 
        \nLeftOut_61[4] , \nRightOut_67[10] , \nRightOut_12[13] , 
        \nRightOut_31[11] , \nLeftOut_62[7] , \nLeftOut_36[14] , 
        \nLeftOut_56[10] , \nRightOut_72[8] , \nRightOut_89[16] , 
        \nLeftOut_60[15] , \nRightOut_24[16] , \nRightOut_44[12] , 
        \nRightOut_13[1] , \ScanLink14[9] , \nLeftOut_64[9] , 
        \nRightOut_69[9] , \nRightOut_74[6] , \nLeftOut_79[6] , 
        \ScanLink6[14] , \ScanLink8[8] , \nLeftOut_27[8] , \nLeftOut_39[4] , 
        \nRightOut_77[5] , \nRightOut_53[3] , \nRightOut_81[5] , 
        \nRightOut_50[0] , \nRightOut_37[7] , \nRightOut_82[6] , 
        \nLeftOut_92[9] , \nRightOut_0[2] , \nLeftOut_1[0] , \nLeftOut_2[3] , 
        \nLeftOut_9[8] , \nLeftOut_11[14] , \nLeftOut_21[6] , \nLeftOut_22[5] , 
        \nRightOut_34[4] , \nRightOut_48[2] , \nRightOut_63[12] , 
        \nRightOut_35[13] , \nLeftOut_27[11] , \nLeftOut_71[10] , 
        \ScanLink29[13] , \nLeftOut_47[15] , \nRightOut_84[8] , 
        \nRightOut_16[11] , \nRightOut_20[14] , \nLeftOut_46[1] , 
        \nLeftOut_89[8] , \nRightOut_76[15] , \nRightOut_31[9] , 
        \nLeftOut_32[16] , \nRightOut_40[10] , \nLeftOut_94[7] , 
        \nLeftOut_45[2] , \nLeftOut_52[12] , \ScanLink15[10] , 
        \nLeftOut_53[6] , \ScanLink20[5] , \ScanLink23[15] , \nRightOut_39[1] , 
        \nLeftOut_81[0] , \nRightOut_92[15] , \nRightOut_69[14] , 
        \nLeftOut_82[3] , \nRightOut_1[11] , \nLeftOut_34[1] , 
        \nLeftOut_37[2] , \nLeftOut_50[5] , \ScanLink23[6] , 
        \nRightOut_87[12] , \nLeftOut_38[10] , \nLeftOut_58[14] , 
        \nLeftOut_95[10] , \nRightOut_43[9] , \ScanLink3[3] , 
        \nRightOut_21[3] , \nRightOut_22[0] , \nLeftOut_55[8] , 
        \nLeftOut_48[7] , \ScanLink25[8] , \nRightOut_94[2] , \nRightOut_3[1] , 
        \nRightOut_46[4] , \ScanLink0[0] , \ScanLink8[10] , \nLeftOut_16[9] , 
        \nRightOut_45[7] , \nRightOut_58[8] , \nRightOut_61[1] , 
        \nRightOut_62[2] , \nLeftOut_10[7] , \nLeftOut_84[15] , 
        \nRightOut_5[13] , \ScanLink11[12] , \nRightOut_79[3] , 
        \nLeftOut_13[4] , \nLeftOut_29[15] , \nLeftOut_49[11] , 
        \nRightOut_18[15] , \nLeftOut_74[3] , \nRightOut_78[11] , 
        \nLeftOut_77[0] , \nLeftOut_91[12] , \ScanLink32[10] , \ScanLink0[9] , 
        \nRightOut_3[8] , \nLeftOut_26[12] , \nLeftOut_46[16] , 
        \nRightOut_83[10] , \nLeftOut_70[13] , \ScanLink28[10] , 
        \nRightOut_89[4] , \nLeftOut_31[5] , \nLeftOut_32[6] , 
        \nRightOut_54[14] , \nRightOut_34[10] , \nRightOut_62[11] , 
        \nLeftOut_1[9] , \nLeftOut_4[4] , \nRightOut_22[9] , \nRightOut_58[1] , 
        \ScanLink5[4] , \nRightOut_5[6] , \nLeftOut_7[7] , \nRightOut_17[12] , 
        \nLeftOut_33[15] , \nLeftOut_53[11] , \nLeftOut_55[1] , 
        \ScanLink26[2] , \nLeftOut_65[14] , \nLeftOut_87[7] , 
        \nRightOut_41[13] , \nLeftOut_84[4] , \nRightOut_77[16] , 
        \nRightOut_40[3] , \nLeftOut_56[2] , \ScanLink25[1] , 
        \nRightOut_92[5] , \ScanLink6[7] , \nRightOut_43[0] , \nRightOut_6[5] , 
        \nRightOut_24[7] , \nLeftOut_29[7] , \nLeftOut_34[8] , 
        \nRightOut_91[6] , \nRightOut_27[4] , \nRightOut_39[8] , 
        \nLeftOut_81[9] , \nLeftOut_69[5] , \nLeftOut_77[9] , \ScanLink19[5] , 
        \nRightOut_0[12] , \ScanLink3[15] , \nRightOut_67[6] , 
        \nLeftOut_4[15] , \nRightOut_4[10] , \ScanLink10[11] , 
        \nRightOut_13[10] , \nLeftOut_14[15] , \nRightOut_18[3] , 
        \nRightOut_64[5] , \nLeftOut_22[10] , \nRightOut_30[12] , 
        \nLeftOut_72[4] , \nRightOut_50[16] , \nRightOut_66[13] , 
        \nLeftOut_71[7] , \nLeftOut_74[11] , \nLeftOut_16[0] , 
        \nRightOut_25[15] , \nLeftOut_42[14] , \nRightOut_73[14] , 
        \nRightOut_45[11] , \nLeftOut_15[3] , \nLeftOut_57[13] , 
        \nLeftOut_61[16] , \nRightOut_61[8] , \nLeftOut_28[16] , 
        \nRightOut_88[15] , \ScanLink26[14] , \nRightOut_13[8] , 
        \ScanLink14[0] , \nLeftOut_48[12] , \nRightOut_69[0] , 
        \nRightOut_82[13] , \nLeftOut_85[16] , \nLeftOut_64[0] , 
        \nLeftOut_67[3] , \ScanLink17[3] , \nLeftOut_90[11] , 
        \nRightOut_19[16] , \nRightOut_79[12] , \ScanLink9[13] , 
        \nRightOut_16[5] , \nLeftOut_18[6] , \nRightOut_72[1] , 
        \nRightOut_71[2] , \nLeftOut_9[1] , \nRightOut_15[6] , 
        \nRightOut_31[0] , \nLeftOut_46[8] , \nLeftOut_89[1] , \ScanLink28[4] , 
        \ScanLink14[13] , \nRightOut_29[2] , \nRightOut_32[3] , 
        \nLeftOut_58[4] , \nLeftOut_40[6] , \nRightOut_55[4] , 
        \nRightOut_87[2] , \nRightOut_56[7] , \nLeftOut_81[14] , 
        \nRightOut_84[1] , \nLeftOut_92[0] , \nLeftOut_91[3] , 
        \nRightOut_93[16] , \nLeftOut_43[5] , \ScanLink30[6] , 
        \nRightOut_2[14] , \nRightOut_6[16] , \ScanLink8[1] , \nLeftOut_24[2] , 
        \nLeftOut_94[13] , \nLeftOut_27[1] , \nLeftOut_39[13] , 
        \nRightOut_50[9] , \nRightOut_86[11] , \nRightOut_8[3] , 
        \nLeftOut_44[6] , \nLeftOut_47[5] , \nLeftOut_69[16] , 
        \nRightOut_80[15] , \nLeftOut_95[3] , \ScanLink29[9] , 
        \ScanLink31[15] , \nRightOut_11[6] , \nLeftOut_20[2] , 
        \nLeftOut_23[1] , \nRightOut_54[9] , \nLeftOut_59[9] , 
        \ScanLink24[12] , \nRightOut_38[12] , \nRightOut_49[6] , 
        \nRightOut_58[16] , \nRightOut_95[12] , \nLeftOut_87[10] , 
        \nRightOut_35[0] , \nRightOut_36[3] , \ScanLink32[8] , 
        \nLeftOut_38[0] , \nLeftOut_42[8] , \nRightOut_52[7] , 
        \nRightOut_80[1] , \nRightOut_51[4] , \nRightOut_83[2] , 
        \nRightOut_75[2] , \nRightOut_76[1] , \nRightOut_12[5] , 
        \nLeftOut_78[2] , \ScanLink13[3] , \nRightOut_49[13] , 
        \nLeftOut_83[12] , \nLeftOut_0[4] , \ScanLink1[13] , \ScanLink2[7] , 
        \nLeftOut_2[11] , \nRightOut_8[12] , \ScanLink10[0] , 
        \nRightOut_17[8] , \nLeftOut_60[0] , \nRightOut_91[10] , 
        \ScanLink20[10] , \ScanLink16[15] , \nLeftOut_63[3] , 
        \nLeftOut_78[13] , \nRightOut_23[11] , \nLeftOut_31[13] , 
        \nLeftOut_67[12] , \nLeftOut_75[7] , \nLeftOut_68[8] , 
        \nRightOut_75[10] , \ScanLink18[8] , \nLeftOut_76[4] , 
        \nLeftOut_11[3] , \nLeftOut_12[11] , \nRightOut_15[14] , 
        \nRightOut_43[15] , \nLeftOut_24[14] , \nLeftOut_72[15] , 
        \nLeftOut_44[10] , \nLeftOut_12[0] , \nRightOut_36[16] , 
        \nRightOut_56[12] , \nRightOut_65[8] , \nLeftOut_73[9] , 
        \nRightOut_78[7] , \nLeftOut_89[14] , \nRightOut_2[5] , 
        \ScanLink5[11] , \nRightOut_47[0] , \nRightOut_60[5] , 
        \nRightOut_63[6] , \nRightOut_88[9] , \nLeftOut_30[8] , 
        \nRightOut_95[6] , \ScanLink1[4] , \nLeftOut_6[13] , \nRightOut_44[3] , 
        \nRightOut_1[6] , \nLeftOut_3[7] , \ScanLink4[9] , \nLeftOut_5[9] , 
        \nRightOut_23[4] , \nLeftOut_49[3] , \nRightOut_11[16] , 
        \nRightOut_20[7] , \nLeftOut_85[9] , \nRightOut_71[12] , 
        \nRightOut_7[8] , \nRightOut_27[13] , \nLeftOut_35[11] , 
        \nLeftOut_36[6] , \nLeftOut_55[15] , \nRightOut_93[8] , 
        \nLeftOut_63[10] , \nLeftOut_35[5] , \nRightOut_38[5] , 
        \nRightOut_52[10] , \nLeftOut_80[4] , \nRightOut_26[9] , 
        \nRightOut_32[14] , \ScanLink21[1] , \nLeftOut_52[2] , 
        \nRightOut_64[15] , \ScanLink4[0] , \nLeftOut_9[14] , \nLeftOut_14[7] , 
        \nLeftOut_16[13] , \nLeftOut_51[1] , \ScanLink22[2] , \nLeftOut_17[4] , 
        \nLeftOut_20[16] , \nLeftOut_40[12] , \ScanLink18[11] , 
        \nLeftOut_83[7] , \nRightOut_85[14] , \nLeftOut_19[14] , 
        \nRightOut_28[14] , \nRightOut_48[10] , \nRightOut_19[7] , 
        \nLeftOut_73[0] , \nLeftOut_79[10] , \ScanLink21[13] , 
        \nRightOut_66[2] , \nLeftOut_70[3] , \nLeftOut_82[11] , 
        \nRightOut_90[13] , \nLeftOut_12[9] , \nRightOut_65[1] , 
        \nRightOut_25[3] , \nLeftOut_68[1] , \ScanLink18[1] , \ScanLink21[8] , 
        \nRightOut_26[0] , \nLeftOut_51[8] , \nRightOut_4[2] , \nLeftOut_5[0] , 
        \ScanLink7[3] , \nRightOut_7[1] , \nLeftOut_28[3] , \nRightOut_41[7] , 
        \nRightOut_93[1] , \nRightOut_90[2] , \nRightOut_7[15] , 
        \nRightOut_42[4] , \nLeftOut_86[3] , \nLeftOut_6[3] , \nLeftOut_54[5] , 
        \nLeftOut_93[14] , \ScanLink27[6] , \nLeftOut_7[10] , \ScanLink9[5] , 
        \nRightOut_9[7] , \ScanLink13[14] , \nLeftOut_30[1] , \nLeftOut_57[6] , 
        \nLeftOut_68[15] , \ScanLink24[5] , \nRightOut_81[16] , 
        \nLeftOut_85[0] , \nLeftOut_86[13] , \nLeftOut_33[2] , 
        \nRightOut_39[11] , \nRightOut_47[9] , \nRightOut_88[0] , 
        \nRightOut_59[15] , \nRightOut_59[5] , \nRightOut_94[11] , 
        \ScanLink25[11] , \nLeftOut_25[6] , \nLeftOut_34[12] , 
        \nLeftOut_38[9] , \nLeftOut_62[13] , \nLeftOut_54[16] , 
        \nRightOut_80[8] , \nRightOut_10[15] , \nLeftOut_26[5] , 
        \nRightOut_26[10] , \nRightOut_70[11] , \nLeftOut_17[10] , 
        \nLeftOut_21[15] , \nRightOut_46[14] , \nLeftOut_77[14] , 
        \nLeftOut_93[4] , \nLeftOut_41[11] , \ScanLink19[12] , 
        \nLeftOut_23[8] , \nRightOut_28[6] , \nRightOut_35[9] , 
        \nLeftOut_41[2] , \ScanLink32[1] , \nLeftOut_42[1] , 
        \nRightOut_65[16] , \ScanLink31[2] , \nRightOut_53[13] , 
        \nLeftOut_90[7] , \nRightOut_54[0] , \ScanLink0[10] , 
        \nRightOut_86[6] , \nRightOut_57[3] , \nRightOut_85[5] , 
        \nLeftOut_0[0] , \nLeftOut_3[12] , \ScanLink4[12] , \nLeftOut_8[5] , 
        \nRightOut_30[4] , \nLeftOut_88[5] , \ScanLink29[0] , 
        \nRightOut_33[7] , \nRightOut_17[1] , \nLeftOut_59[0] , 
        \nLeftOut_60[9] , \nRightOut_9[11] , \ScanLink10[9] , 
        \nRightOut_14[2] , \nLeftOut_19[2] , \nRightOut_70[6] , 
        \nRightOut_73[5] , \nRightOut_11[12] , \nLeftOut_13[12] , 
        \ScanLink15[4] , \nRightOut_22[12] , \nRightOut_42[16] , 
        \ScanLink16[7] , \nLeftOut_30[10] , \nLeftOut_50[14] , 
        \nLeftOut_66[7] , \nRightOut_74[13] , \nLeftOut_66[11] , 
        \nRightOut_37[15] , \nRightOut_57[11] , \nLeftOut_65[4] , 
        \nRightOut_68[4] , \nRightOut_61[14] , \nLeftOut_45[13] , 
        \nRightOut_76[8] , \nLeftOut_35[15] , \nLeftOut_35[1] , 
        \nLeftOut_73[16] , \nRightOut_42[9] , \nLeftOut_36[2] , 
        \nLeftOut_55[11] , \nLeftOut_63[14] , \nRightOut_71[16] , 
        \nLeftOut_20[12] , \nRightOut_47[13] , \nLeftOut_76[13] , 
        \nLeftOut_83[3] , \nLeftOut_40[16] , \ScanLink18[15] , \ScanLink1[0] , 
        \nRightOut_1[2] , \nLeftOut_3[3] , \nLeftOut_51[5] , \ScanLink22[6] , 
        \nRightOut_64[11] , \nRightOut_32[10] , \ScanLink21[5] , 
        \nRightOut_38[1] , \nLeftOut_52[6] , \nRightOut_52[14] , 
        \nLeftOut_80[0] , \ScanLink2[3] , \nRightOut_44[7] , \nRightOut_59[8] , 
        \nRightOut_95[2] , \nLeftOut_2[15] , \nRightOut_2[1] , \ScanLink5[15] , 
        \nRightOut_20[3] , \nRightOut_47[4] , \ScanLink24[8] , 
        \nRightOut_23[0] , \nLeftOut_54[8] , \nLeftOut_49[7] , 
        \nRightOut_2[10] , \nRightOut_8[16] , \nRightOut_15[10] , 
        \nLeftOut_17[9] , \nRightOut_60[1] , \nRightOut_63[2] , 
        \nLeftOut_11[7] , \nLeftOut_12[4] , \nRightOut_23[15] , 
        \nRightOut_43[11] , \nRightOut_36[12] , \nLeftOut_51[13] , 
        \nRightOut_75[14] , \nLeftOut_76[0] , \nRightOut_56[16] , 
        \nLeftOut_67[16] , \nLeftOut_75[3] , \nRightOut_78[3] , 
        \nLeftOut_89[10] , \nRightOut_60[13] , \nLeftOut_12[15] , 
        \nLeftOut_44[14] , \nLeftOut_24[10] , \nLeftOut_72[11] , 
        \nRightOut_73[8] , \nRightOut_84[13] , \ScanLink10[4] , 
        \ScanLink16[11] , \nLeftOut_18[13] , \nRightOut_29[13] , 
        \ScanLink20[14] , \ScanLink13[7] , \nLeftOut_63[7] , 
        \nRightOut_91[14] , \nRightOut_6[12] , \nLeftOut_8[13] , 
        \nLeftOut_60[4] , \nLeftOut_83[16] , \nRightOut_76[5] , 
        \nLeftOut_8[8] , \ScanLink9[8] , \nRightOut_11[2] , \nRightOut_12[1] , 
        \nRightOut_68[9] , \nRightOut_75[6] , \nLeftOut_65[9] , 
        \nLeftOut_78[6] , \ScanLink15[9] , \nLeftOut_26[8] , \nRightOut_35[4] , 
        \nRightOut_36[7] , \nLeftOut_93[9] , \nRightOut_51[0] , 
        \nLeftOut_38[4] , \nRightOut_83[6] , \nRightOut_52[3] , 
        \nRightOut_80[5] , \nLeftOut_20[6] , \nRightOut_30[9] , 
        \nLeftOut_44[2] , \nLeftOut_92[13] , \nLeftOut_47[1] , 
        \nLeftOut_69[12] , \nLeftOut_88[8] , \ScanLink31[11] , 
        \nRightOut_80[11] , \nLeftOut_95[7] , \nLeftOut_87[14] , 
        \nRightOut_38[16] , \nRightOut_58[12] , \nRightOut_85[8] , 
        \nRightOut_95[16] , \nRightOut_49[2] , \ScanLink0[14] , 
        \nLeftOut_3[16] , \nRightOut_9[15] , \ScanLink12[13] , 
        \nLeftOut_23[5] , \nRightOut_12[8] , \ScanLink16[3] , \nLeftOut_65[0] , 
        \ScanLink15[0] , \nLeftOut_30[14] , \nLeftOut_66[15] , 
        \nLeftOut_50[10] , \nRightOut_22[16] , \nLeftOut_66[3] , 
        \nLeftOut_13[16] , \nRightOut_14[13] , \nRightOut_42[12] , 
        \nLeftOut_25[13] , \nLeftOut_73[12] , \nRightOut_14[6] , 
        \nRightOut_37[11] , \nRightOut_57[15] , \nRightOut_61[10] , 
        \nRightOut_68[0] , \nLeftOut_88[13] , \nRightOut_17[5] , 
        \nLeftOut_19[6] , \nRightOut_70[2] , \nRightOut_73[1] , 
        \nRightOut_57[7] , \nRightOut_85[1] , \nLeftOut_7[14] , 
        \nRightOut_86[2] , \nLeftOut_8[1] , \nRightOut_54[4] , 
        \nRightOut_30[0] , \nRightOut_33[3] , \nLeftOut_59[4] , 
        \nLeftOut_47[8] , \nLeftOut_88[1] , \ScanLink29[4] , \nLeftOut_0[9] , 
        \ScanLink1[9] , \nLeftOut_5[4] , \nLeftOut_6[7] , \ScanLink9[1] , 
        \nRightOut_10[11] , \nRightOut_46[10] , \nLeftOut_26[1] , 
        \nRightOut_26[14] , \nRightOut_51[9] , \nRightOut_70[15] , 
        \nRightOut_9[3] , \nLeftOut_17[14] , \nLeftOut_25[2] , 
        \nLeftOut_34[16] , \nLeftOut_54[12] , \nRightOut_28[2] , 
        \nRightOut_33[13] , \nLeftOut_90[3] , \ScanLink31[6] , 
        \nLeftOut_41[6] , \nLeftOut_42[5] , \nRightOut_65[12] , 
        \ScanLink32[5] , \nLeftOut_21[11] , \nLeftOut_41[15] , 
        \nLeftOut_77[10] , \nRightOut_81[12] , \nLeftOut_93[0] , 
        \nLeftOut_85[4] , \nRightOut_23[9] , \nLeftOut_57[2] , 
        \nLeftOut_68[11] , \ScanLink24[1] , \ScanLink30[12] , 
        \nRightOut_7[11] , \nLeftOut_54[1] , \nLeftOut_93[10] , 
        \ScanLink27[2] , \ScanLink13[10] , \nLeftOut_86[7] , \nLeftOut_33[6] , 
        \ScanLink25[15] , \nRightOut_2[8] , \nRightOut_39[15] , 
        \nRightOut_59[11] , \nRightOut_59[1] , \nRightOut_94[15] , 
        \nRightOut_88[4] , \nRightOut_26[4] , \nLeftOut_30[5] , \ScanLink4[4] , 
        \nRightOut_4[6] , \ScanLink7[7] , \nRightOut_25[7] , \nRightOut_38[8] , 
        \nRightOut_42[0] , \nLeftOut_80[9] , \nRightOut_7[5] , 
        \nLeftOut_28[7] , \nLeftOut_35[8] , \nRightOut_90[6] , 
        \nRightOut_41[3] , \nRightOut_93[5] , \nRightOut_1[9] , \ScanLink2[8] , 
        \nRightOut_3[13] , \nLeftOut_9[10] , \nRightOut_65[5] , 
        \nRightOut_28[10] , \nRightOut_66[6] , \nLeftOut_68[5] , 
        \nLeftOut_76[9] , \ScanLink18[5] , \nLeftOut_5[6] , \nRightOut_7[13] , 
        \nLeftOut_14[3] , \nRightOut_48[14] , \nLeftOut_17[0] , 
        \nLeftOut_19[10] , \nRightOut_19[3] , \nRightOut_60[8] , 
        \nLeftOut_70[7] , \nLeftOut_82[15] , \nRightOut_85[10] , 
        \nLeftOut_73[4] , \nLeftOut_79[14] , \ScanLink17[12] , 
        \nLeftOut_86[5] , \nLeftOut_54[3] , \nLeftOut_93[12] , \ScanLink27[0] , 
        \nLeftOut_6[5] , \nLeftOut_57[0] , \ScanLink30[10] , \ScanLink24[3] , 
        \nRightOut_20[8] , \nLeftOut_68[13] , \nRightOut_81[10] , 
        \nLeftOut_85[6] , \nLeftOut_30[7] , \nLeftOut_33[4] , 
        \nRightOut_59[13] , \nLeftOut_86[15] , \nRightOut_88[6] , 
        \nRightOut_59[3] , \nRightOut_95[9] , \nLeftOut_3[8] , 
        \ScanLink13[12] , \ScanLink4[6] , \nRightOut_4[4] , \nRightOut_25[5] , 
        \nRightOut_26[6] , \nLeftOut_36[9] , \nLeftOut_83[8] , 
        \nLeftOut_3[14] , \nRightOut_3[11] , \ScanLink7[5] , \nLeftOut_28[5] , 
        \nRightOut_41[1] , \nRightOut_93[7] , \nRightOut_90[4] , 
        \nRightOut_7[7] , \nLeftOut_9[12] , \nRightOut_42[2] , 
        \nRightOut_66[4] , \nLeftOut_14[1] , \nLeftOut_17[2] , 
        \nRightOut_65[7] , \nLeftOut_68[7] , \nLeftOut_75[8] , 
        \nRightOut_78[8] , \nRightOut_85[12] , \ScanLink18[7] , 
        \nRightOut_63[9] , \ScanLink4[14] , \nRightOut_11[9] , 
        \nLeftOut_19[12] , \nRightOut_28[12] , \nRightOut_48[16] , 
        \ScanLink17[10] , \nRightOut_19[1] , \nLeftOut_73[6] , 
        \nLeftOut_79[16] , \ScanLink21[15] , \nRightOut_42[10] , 
        \nLeftOut_70[5] , \nRightOut_90[15] , \nLeftOut_13[14] , 
        \nRightOut_14[11] , \ScanLink15[2] , \nRightOut_22[14] , 
        \nLeftOut_66[1] , \nRightOut_74[15] , \ScanLink16[1] , 
        \nLeftOut_30[16] , \nLeftOut_50[12] , \nLeftOut_65[2] , 
        \nRightOut_37[13] , \nRightOut_68[2] , \nLeftOut_88[11] , 
        \nRightOut_61[12] , \nRightOut_17[7] , \nLeftOut_25[11] , 
        \nLeftOut_45[15] , \nLeftOut_73[10] , \nLeftOut_7[16] , 
        \nRightOut_14[4] , \nLeftOut_19[4] , \nRightOut_54[6] , 
        \nRightOut_70[0] , \nRightOut_73[3] , \nRightOut_49[9] , 
        \nRightOut_57[5] , \nRightOut_85[3] , \nRightOut_86[0] , 
        \ScanLink29[6] , \nRightOut_2[12] , \nLeftOut_8[3] , \nRightOut_30[2] , 
        \nLeftOut_88[3] , \nRightOut_33[1] , \nLeftOut_44[9] , 
        \nLeftOut_59[6] , \ScanLink9[3] , \nLeftOut_25[0] , \nLeftOut_34[14] , 
        \nRightOut_52[8] , \nLeftOut_62[15] , \nLeftOut_54[10] , 
        \nRightOut_9[1] , \nRightOut_10[13] , \nLeftOut_26[3] , 
        \nRightOut_26[16] , \nRightOut_46[12] , \nLeftOut_17[16] , 
        \nLeftOut_21[13] , \nLeftOut_77[12] , \nLeftOut_93[2] , 
        \nRightOut_28[0] , \nRightOut_33[11] , \nLeftOut_41[4] , 
        \ScanLink19[14] , \nLeftOut_42[7] , \ScanLink32[7] , 
        \nRightOut_53[15] , \nRightOut_65[10] , \ScanLink31[4] , 
        \nLeftOut_90[1] , \nRightOut_29[11] , \nLeftOut_8[11] , 
        \ScanLink10[6] , \ScanLink13[5] , \nRightOut_49[15] , \nLeftOut_60[6] , 
        \nRightOut_70[9] , \nRightOut_84[11] , \nLeftOut_83[14] , 
        \nLeftOut_63[5] , \nLeftOut_78[15] , \nRightOut_91[16] , 
        \ScanLink16[13] , \nLeftOut_18[11] , \nRightOut_75[4] , 
        \nRightOut_9[8] , \nRightOut_11[0] , \nLeftOut_66[8] , 
        \nRightOut_76[7] , \nRightOut_12[3] , \ScanLink16[8] , 
        \nLeftOut_78[4] , \nLeftOut_25[9] , \nRightOut_28[9] , 
        \nRightOut_35[6] , \nRightOut_36[5] , \nRightOut_52[1] , 
        \nLeftOut_90[8] , \nLeftOut_38[6] , \nRightOut_80[7] , 
        \nRightOut_83[4] , \nRightOut_51[2] , \nRightOut_80[13] , 
        \nLeftOut_95[5] , \nRightOut_6[10] , \nRightOut_33[8] , 
        \nLeftOut_47[3] , \nLeftOut_69[10] , \ScanLink31[13] , 
        \nLeftOut_44[0] , \nLeftOut_92[11] , \nRightOut_11[10] , 
        \ScanLink12[11] , \nLeftOut_20[4] , \nLeftOut_23[7] , 
        \nRightOut_38[14] , \nRightOut_49[0] , \ScanLink24[14] , 
        \nRightOut_58[10] , \nRightOut_86[9] , \nRightOut_95[14] , 
        \nRightOut_41[8] , \nLeftOut_87[16] , \nRightOut_27[15] , 
        \nLeftOut_36[0] , \nRightOut_47[11] , \nRightOut_71[14] , \nEnable[0] , 
        \nLeftOut_0[2] , \nLeftOut_3[1] , \nRightOut_32[12] , \nLeftOut_35[3] , 
        \nLeftOut_55[13] , \nLeftOut_63[16] , \nRightOut_38[3] , 
        \nLeftOut_52[4] , \nRightOut_52[16] , \nLeftOut_80[2] , 
        \nRightOut_64[13] , \ScanLink21[7] , \nLeftOut_51[7] , \ScanLink22[4] , 
        \ScanLink1[15] , \ScanLink2[1] , \nLeftOut_16[15] , \nLeftOut_40[14] , 
        \nLeftOut_20[10] , \nLeftOut_76[11] , \nLeftOut_83[1] , 
        \nRightOut_47[6] , \nRightOut_2[3] , \nRightOut_95[0] , \ScanLink1[2] , 
        \nRightOut_1[0] , \nLeftOut_6[15] , \nRightOut_44[5] , 
        \nRightOut_20[1] , \nRightOut_23[2] , \nLeftOut_49[5] , 
        \ScanLink27[9] , \nLeftOut_57[9] , \ScanLink0[12] , \nRightOut_8[14] , 
        \nLeftOut_14[8] , \nRightOut_19[8] , \nRightOut_60[3] , 
        \nRightOut_15[12] , \nLeftOut_31[15] , \nRightOut_63[0] , 
        \nLeftOut_75[1] , \nLeftOut_51[11] , \nLeftOut_67[14] , 
        \nRightOut_75[16] , \nLeftOut_76[2] , \ScanLink9[7] , \nRightOut_9[5] , 
        \nLeftOut_11[5] , \nLeftOut_24[12] , \nRightOut_43[13] , 
        \nLeftOut_72[13] , \nLeftOut_44[16] , \nLeftOut_12[6] , 
        \nRightOut_60[11] , \nLeftOut_26[7] , \nRightOut_36[10] , 
        \nRightOut_46[16] , \nRightOut_56[14] , \nRightOut_78[1] , 
        \nLeftOut_89[12] , \nRightOut_26[12] , \nRightOut_70[13] , 
        \nRightOut_83[9] , \nLeftOut_17[12] , \nLeftOut_25[4] , 
        \nLeftOut_34[10] , \nLeftOut_54[14] , \nLeftOut_62[11] , 
        \nRightOut_28[4] , \nRightOut_33[15] , \nLeftOut_42[3] , 
        \nRightOut_53[11] , \nLeftOut_90[5] , \nRightOut_65[14] , 
        \nRightOut_36[8] , \ScanLink31[0] , \nLeftOut_41[13] , 
        \nLeftOut_41[0] , \ScanLink32[3] , \ScanLink19[10] , \nLeftOut_20[9] , 
        \nRightOut_57[1] , \nLeftOut_77[16] , \nLeftOut_93[6] , 
        \nRightOut_85[7] , \nLeftOut_7[12] , \nRightOut_86[4] , 
        \nLeftOut_8[7] , \nRightOut_54[2] , \nLeftOut_59[2] , 
        \nRightOut_30[6] , \nRightOut_33[5] , \nLeftOut_88[7] , 
        \nLeftOut_3[10] , \nRightOut_14[0] , \nLeftOut_63[8] , 
        \nLeftOut_95[8] , \ScanLink29[2] , \nRightOut_3[15] , \ScanLink4[10] , 
        \nRightOut_9[13] , \ScanLink13[8] , \nRightOut_14[15] , 
        \ScanLink15[6] , \ScanLink16[5] , \nRightOut_17[3] , \nLeftOut_19[0] , 
        \nRightOut_70[4] , \nRightOut_73[7] , \nLeftOut_65[6] , 
        \nLeftOut_30[12] , \nLeftOut_50[16] , \nLeftOut_66[13] , 
        \nLeftOut_78[9] , \nLeftOut_66[5] , \nRightOut_22[10] , 
        \nRightOut_74[11] , \nLeftOut_13[10] , \nLeftOut_25[15] , 
        \nRightOut_42[14] , \nLeftOut_73[14] , \nLeftOut_45[11] , 
        \nRightOut_28[16] , \nRightOut_57[13] , \nRightOut_61[16] , 
        \nRightOut_68[6] , \nRightOut_75[9] , \nLeftOut_88[15] , 
        \ScanLink4[2] , \ScanLink7[1] , \nRightOut_7[3] , \nLeftOut_9[16] , 
        \nLeftOut_14[5] , \nRightOut_48[12] , \nLeftOut_17[6] , 
        \nLeftOut_19[16] , \nRightOut_19[5] , \nLeftOut_70[1] , 
        \nRightOut_85[16] , \nLeftOut_82[13] , \nRightOut_90[11] , 
        \nLeftOut_73[2] , \nLeftOut_79[12] , \ScanLink21[11] , 
        \nRightOut_65[3] , \ScanLink17[14] , \nLeftOut_11[8] , 
        \nRightOut_25[1] , \nRightOut_26[2] , \nRightOut_66[0] , 
        \nLeftOut_68[3] , \ScanLink18[3] , \ScanLink22[9] , \nRightOut_42[6] , 
        \nLeftOut_52[9] , \nLeftOut_28[1] , \nRightOut_90[0] , 
        \nRightOut_41[5] , \nRightOut_93[3] , \nLeftOut_0[6] , \ScanLink1[11] , 
        \ScanLink1[6] , \nLeftOut_2[13] , \nRightOut_4[0] , \ScanLink5[13] , 
        \nLeftOut_5[2] , \nLeftOut_6[1] , \nLeftOut_57[4] , \nRightOut_81[14] , 
        \nLeftOut_85[2] , \ScanLink24[7] , \ScanLink30[14] , \nLeftOut_54[7] , 
        \nLeftOut_93[16] , \ScanLink27[4] , \nRightOut_8[10] , 
        \nLeftOut_30[3] , \nLeftOut_33[0] , \nRightOut_44[8] , 
        \nLeftOut_49[8] , \nLeftOut_86[1] , \nRightOut_39[13] , 
        \nRightOut_59[7] , \ScanLink25[13] , \nRightOut_94[13] , 
        \nRightOut_88[2] , \nLeftOut_86[11] , \nLeftOut_11[1] , 
        \nLeftOut_12[2] , \nRightOut_15[16] , \nRightOut_23[13] , 
        \nRightOut_75[12] , \nLeftOut_76[6] , \nLeftOut_31[11] , 
        \nLeftOut_51[15] , \nLeftOut_67[10] , \nRightOut_56[10] , 
        \nLeftOut_75[5] , \nRightOut_78[5] , \nLeftOut_89[16] , 
        \nRightOut_36[14] , \nRightOut_60[15] , \nRightOut_66[9] , 
        \nLeftOut_12[13] , \nLeftOut_24[16] , \nLeftOut_44[12] , 
        \nLeftOut_70[8] , \nRightOut_60[7] , \nRightOut_63[4] , 
        \nRightOut_1[4] , \nLeftOut_33[9] , \nLeftOut_6[11] , 
        \nRightOut_44[1] , \ScanLink2[5] , \nRightOut_2[7] , \nRightOut_95[4] , 
        \nRightOut_4[9] , \nLeftOut_6[8] , \nRightOut_47[2] , \ScanLink7[8] , 
        \nRightOut_20[5] , \nRightOut_23[6] , \nLeftOut_35[7] , 
        \nLeftOut_49[1] , \nLeftOut_86[8] , \nRightOut_27[11] , 
        \nLeftOut_28[8] , \nLeftOut_35[13] , \nLeftOut_63[12] , 
        \nLeftOut_36[4] , \nRightOut_71[10] , \nRightOut_90[9] , 
        \nRightOut_11[14] , \nRightOut_47[15] , \nLeftOut_16[11] , 
        \nLeftOut_20[14] , \nLeftOut_76[15] , \nLeftOut_83[5] , 
        \nLeftOut_40[10] , \nLeftOut_51[3] , \ScanLink18[13] , \ScanLink22[0] , 
        \nRightOut_2[16] , \nLeftOut_3[5] , \nRightOut_32[16] , 
        \nLeftOut_52[0] , \ScanLink21[3] , \nRightOut_6[14] , 
        \nRightOut_25[8] , \nRightOut_38[7] , \nRightOut_52[12] , 
        \nLeftOut_80[6] , \nLeftOut_8[15] , \ScanLink12[15] , \nLeftOut_20[0] , 
        \nLeftOut_44[4] , \nLeftOut_47[7] , \nLeftOut_92[15] , 
        \nLeftOut_69[14] , \nLeftOut_95[1] , \nLeftOut_23[3] , 
        \nRightOut_38[10] , \nRightOut_57[8] , \nLeftOut_87[12] , 
        \nRightOut_49[4] , \nRightOut_58[14] , \nRightOut_95[10] , 
        \ScanLink24[10] , \nRightOut_35[2] , \ScanLink31[9] , 
        \nRightOut_36[1] , \nLeftOut_41[9] , \nLeftOut_38[2] , 
        \nRightOut_51[6] , \nRightOut_83[0] , \nRightOut_52[5] , 
        \nRightOut_80[3] , \nRightOut_76[3] , \nRightOut_11[4] , 
        \nRightOut_12[7] , \nRightOut_75[0] , \nLeftOut_78[0] , 
        \nRightOut_84[15] , \ScanLink10[2] , \nRightOut_14[9] , 
        \nLeftOut_19[9] , \nRightOut_49[11] , \nRightOut_29[15] , 
        \nLeftOut_18[15] , \nLeftOut_63[1] , \nLeftOut_78[11] , 
        \ScanLink20[12] , \nLeftOut_60[2] , \nRightOut_91[12] , 
        \ScanLink13[1] , \nLeftOut_83[10] ;
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink4[15] , \ScanLink4[14] , \ScanLink4[13] , 
        \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , \ScanLink4[9] , 
        \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , \ScanLink4[5] , 
        \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , \ScanLink4[1] , 
        \ScanLink4[0] }), .ScanOut({\ScanLink5[15] , \ScanLink5[14] , 
        \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , 
        \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_4[16] , \nLeftOut_4[15] , \nLeftOut_4[14] , \nLeftOut_4[13] , 
        \nLeftOut_4[12] , \nLeftOut_4[11] , \nLeftOut_4[10] , \nLeftOut_4[9] , 
        \nLeftOut_4[8] , \nLeftOut_4[7] , \nLeftOut_4[6] , \nLeftOut_4[5] , 
        \nLeftOut_4[4] , \nLeftOut_4[3] , \nLeftOut_4[2] , \nLeftOut_4[1] , 
        \nLeftOut_4[0] }), .inright({\nRightOut_4[16] , \nRightOut_4[15] , 
        \nRightOut_4[14] , \nRightOut_4[13] , \nRightOut_4[12] , 
        \nRightOut_4[11] , \nRightOut_4[10] , \nRightOut_4[9] , 
        \nRightOut_4[8] , \nRightOut_4[7] , \nRightOut_4[6] , \nRightOut_4[5] , 
        \nRightOut_4[4] , \nRightOut_4[3] , \nRightOut_4[2] , \nRightOut_4[1] , 
        \nRightOut_4[0] }), .outleft({\nLeftOut_4[16] , \nLeftOut_4[15] , 
        \nLeftOut_4[14] , \nLeftOut_4[13] , \nLeftOut_4[12] , \nLeftOut_4[11] , 
        \nLeftOut_4[10] , \nLeftOut_4[9] , \nLeftOut_4[8] , \nLeftOut_4[7] , 
        \nLeftOut_4[6] , \nLeftOut_4[5] , \nLeftOut_4[4] , \nLeftOut_4[3] , 
        \nLeftOut_4[2] , \nLeftOut_4[1] , \nLeftOut_4[0] }), .outright({
        \nRightOut_4[16] , \nRightOut_4[15] , \nRightOut_4[14] , 
        \nRightOut_4[13] , \nRightOut_4[12] , \nRightOut_4[11] , 
        \nRightOut_4[10] , \nRightOut_4[9] , \nRightOut_4[8] , 
        \nRightOut_4[7] , \nRightOut_4[6] , \nRightOut_4[5] , \nRightOut_4[4] , 
        \nRightOut_4[3] , \nRightOut_4[2] , \nRightOut_4[1] , \nRightOut_4[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_10 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink10[15] , \ScanLink10[14] , \ScanLink10[13] , 
        \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , \ScanLink10[9] , 
        \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , \ScanLink10[5] , 
        \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , \ScanLink10[1] , 
        \ScanLink10[0] }), .ScanOut({\ScanLink11[15] , \ScanLink11[14] , 
        \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , 
        \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , 
        \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , 
        \ScanLink11[1] , \ScanLink11[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_10[16] , \nLeftOut_10[15] , \nLeftOut_10[14] , 
        \nLeftOut_10[13] , \nLeftOut_10[12] , \nLeftOut_10[11] , 
        \nLeftOut_10[10] , \nLeftOut_10[9] , \nLeftOut_10[8] , 
        \nLeftOut_10[7] , \nLeftOut_10[6] , \nLeftOut_10[5] , \nLeftOut_10[4] , 
        \nLeftOut_10[3] , \nLeftOut_10[2] , \nLeftOut_10[1] , \nLeftOut_10[0] 
        }), .inright({\nRightOut_10[16] , \nRightOut_10[15] , 
        \nRightOut_10[14] , \nRightOut_10[13] , \nRightOut_10[12] , 
        \nRightOut_10[11] , \nRightOut_10[10] , \nRightOut_10[9] , 
        \nRightOut_10[8] , \nRightOut_10[7] , \nRightOut_10[6] , 
        \nRightOut_10[5] , \nRightOut_10[4] , \nRightOut_10[3] , 
        \nRightOut_10[2] , \nRightOut_10[1] , \nRightOut_10[0] }), .outleft({
        \nLeftOut_10[16] , \nLeftOut_10[15] , \nLeftOut_10[14] , 
        \nLeftOut_10[13] , \nLeftOut_10[12] , \nLeftOut_10[11] , 
        \nLeftOut_10[10] , \nLeftOut_10[9] , \nLeftOut_10[8] , 
        \nLeftOut_10[7] , \nLeftOut_10[6] , \nLeftOut_10[5] , \nLeftOut_10[4] , 
        \nLeftOut_10[3] , \nLeftOut_10[2] , \nLeftOut_10[1] , \nLeftOut_10[0] 
        }), .outright({\nRightOut_10[16] , \nRightOut_10[15] , 
        \nRightOut_10[14] , \nRightOut_10[13] , \nRightOut_10[12] , 
        \nRightOut_10[11] , \nRightOut_10[10] , \nRightOut_10[9] , 
        \nRightOut_10[8] , \nRightOut_10[7] , \nRightOut_10[6] , 
        \nRightOut_10[5] , \nRightOut_10[4] , \nRightOut_10[3] , 
        \nRightOut_10[2] , \nRightOut_10[1] , \nRightOut_10[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_37 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_20[16] , \nRightOut_20[15] , \nRightOut_20[14] , 
        \nRightOut_20[13] , \nRightOut_20[12] , \nRightOut_20[11] , 
        \nRightOut_20[10] , \nRightOut_20[9] , \nRightOut_20[8] , 
        \nRightOut_20[7] , \nRightOut_20[6] , \nRightOut_20[5] , 
        \nRightOut_20[4] , \nRightOut_20[3] , \nRightOut_20[2] , 
        \nRightOut_20[1] , \nRightOut_20[0] }), .inright({\nRightOut_21[16] , 
        \nRightOut_21[15] , \nRightOut_21[14] , \nRightOut_21[13] , 
        \nRightOut_21[12] , \nRightOut_21[11] , \nRightOut_21[10] , 
        \nRightOut_21[9] , \nRightOut_21[8] , \nRightOut_21[7] , 
        \nRightOut_21[6] , \nRightOut_21[5] , \nRightOut_21[4] , 
        \nRightOut_21[3] , \nRightOut_21[2] , \nRightOut_21[1] , 
        \nRightOut_21[0] }), .outleft({\nLeftOut_37[16] , \nLeftOut_37[15] , 
        \nLeftOut_37[14] , \nLeftOut_37[13] , \nLeftOut_37[12] , 
        \nLeftOut_37[11] , \nLeftOut_37[10] , \nLeftOut_37[9] , 
        \nLeftOut_37[8] , \nLeftOut_37[7] , \nLeftOut_37[6] , \nLeftOut_37[5] , 
        \nLeftOut_37[4] , \nLeftOut_37[3] , \nLeftOut_37[2] , \nLeftOut_37[1] , 
        \nLeftOut_37[0] }), .outright({\nRightOut_37[16] , \nRightOut_37[15] , 
        \nRightOut_37[14] , \nRightOut_37[13] , \nRightOut_37[12] , 
        \nRightOut_37[11] , \nRightOut_37[10] , \nRightOut_37[9] , 
        \nRightOut_37[8] , \nRightOut_37[7] , \nRightOut_37[6] , 
        \nRightOut_37[5] , \nRightOut_37[4] , \nRightOut_37[3] , 
        \nRightOut_37[2] , \nRightOut_37[1] , \nRightOut_37[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_42 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_26[16] , \nLeftOut_26[15] , \nLeftOut_26[14] , 
        \nLeftOut_26[13] , \nLeftOut_26[12] , \nLeftOut_26[11] , 
        \nLeftOut_26[10] , \nLeftOut_26[9] , \nLeftOut_26[8] , 
        \nLeftOut_26[7] , \nLeftOut_26[6] , \nLeftOut_26[5] , \nLeftOut_26[4] , 
        \nLeftOut_26[3] , \nLeftOut_26[2] , \nLeftOut_26[1] , \nLeftOut_26[0] 
        }), .inright({\nLeftOut_27[16] , \nLeftOut_27[15] , \nLeftOut_27[14] , 
        \nLeftOut_27[13] , \nLeftOut_27[12] , \nLeftOut_27[11] , 
        \nLeftOut_27[10] , \nLeftOut_27[9] , \nLeftOut_27[8] , 
        \nLeftOut_27[7] , \nLeftOut_27[6] , \nLeftOut_27[5] , \nLeftOut_27[4] , 
        \nLeftOut_27[3] , \nLeftOut_27[2] , \nLeftOut_27[1] , \nLeftOut_27[0] 
        }), .outleft({\nLeftOut_42[16] , \nLeftOut_42[15] , \nLeftOut_42[14] , 
        \nLeftOut_42[13] , \nLeftOut_42[12] , \nLeftOut_42[11] , 
        \nLeftOut_42[10] , \nLeftOut_42[9] , \nLeftOut_42[8] , 
        \nLeftOut_42[7] , \nLeftOut_42[6] , \nLeftOut_42[5] , \nLeftOut_42[4] , 
        \nLeftOut_42[3] , \nLeftOut_42[2] , \nLeftOut_42[1] , \nLeftOut_42[0] 
        }), .outright({\nRightOut_42[16] , \nRightOut_42[15] , 
        \nRightOut_42[14] , \nRightOut_42[13] , \nRightOut_42[12] , 
        \nRightOut_42[11] , \nRightOut_42[10] , \nRightOut_42[9] , 
        \nRightOut_42[8] , \nRightOut_42[7] , \nRightOut_42[6] , 
        \nRightOut_42[5] , \nRightOut_42[4] , \nRightOut_42[3] , 
        \nRightOut_42[2] , \nRightOut_42[1] , \nRightOut_42[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s2_SCAN1 node_65 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_49[16] , \nLeftOut_49[15] , \nLeftOut_49[14] , 
        \nLeftOut_49[13] , \nLeftOut_49[12] , \nLeftOut_49[11] , 
        \nLeftOut_49[10] , \nLeftOut_49[9] , \nLeftOut_49[8] , 
        \nLeftOut_49[7] , \nLeftOut_49[6] , \nLeftOut_49[5] , \nLeftOut_49[4] , 
        \nLeftOut_49[3] , \nLeftOut_49[2] , \nLeftOut_49[1] , \nLeftOut_49[0] 
        }), .inright({\nLeftOut_53[16] , \nLeftOut_53[15] , \nLeftOut_53[14] , 
        \nLeftOut_53[13] , \nLeftOut_53[12] , \nLeftOut_53[11] , 
        \nLeftOut_53[10] , \nLeftOut_53[9] , \nLeftOut_53[8] , 
        \nLeftOut_53[7] , \nLeftOut_53[6] , \nLeftOut_53[5] , \nLeftOut_53[4] , 
        \nLeftOut_53[3] , \nLeftOut_53[2] , \nLeftOut_53[1] , \nLeftOut_53[0] 
        }), .outleft({\nLeftOut_65[16] , \nLeftOut_65[15] , \nLeftOut_65[14] , 
        \nLeftOut_65[13] , \nLeftOut_65[12] , \nLeftOut_65[11] , 
        \nLeftOut_65[10] , \nLeftOut_65[9] , \nLeftOut_65[8] , 
        \nLeftOut_65[7] , \nLeftOut_65[6] , \nLeftOut_65[5] , \nLeftOut_65[4] , 
        \nLeftOut_65[3] , \nLeftOut_65[2] , \nLeftOut_65[1] , \nLeftOut_65[0] 
        }), .outright({\nRightOut_65[16] , \nRightOut_65[15] , 
        \nRightOut_65[14] , \nRightOut_65[13] , \nRightOut_65[12] , 
        \nRightOut_65[11] , \nRightOut_65[10] , \nRightOut_65[9] , 
        \nRightOut_65[8] , \nRightOut_65[7] , \nRightOut_65[6] , 
        \nRightOut_65[5] , \nRightOut_65[4] , \nRightOut_65[3] , 
        \nRightOut_65[2] , \nRightOut_65[1] , \nRightOut_65[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_80 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_64[16] , \nLeftOut_64[15] , \nLeftOut_64[14] , 
        \nLeftOut_64[13] , \nLeftOut_64[12] , \nLeftOut_64[11] , 
        \nLeftOut_64[10] , \nLeftOut_64[9] , \nLeftOut_64[8] , 
        \nLeftOut_64[7] , \nLeftOut_64[6] , \nLeftOut_64[5] , \nLeftOut_64[4] , 
        \nLeftOut_64[3] , \nLeftOut_64[2] , \nLeftOut_64[1] , \nLeftOut_64[0] 
        }), .inright({\nLeftOut_72[16] , \nLeftOut_72[15] , \nLeftOut_72[14] , 
        \nLeftOut_72[13] , \nLeftOut_72[12] , \nLeftOut_72[11] , 
        \nLeftOut_72[10] , \nLeftOut_72[9] , \nLeftOut_72[8] , 
        \nLeftOut_72[7] , \nLeftOut_72[6] , \nLeftOut_72[5] , \nLeftOut_72[4] , 
        \nLeftOut_72[3] , \nLeftOut_72[2] , \nLeftOut_72[1] , \nLeftOut_72[0] 
        }), .outleft({\nLeftOut_80[16] , \nLeftOut_80[15] , \nLeftOut_80[14] , 
        \nLeftOut_80[13] , \nLeftOut_80[12] , \nLeftOut_80[11] , 
        \nLeftOut_80[10] , \nLeftOut_80[9] , \nLeftOut_80[8] , 
        \nLeftOut_80[7] , \nLeftOut_80[6] , \nLeftOut_80[5] , \nLeftOut_80[4] , 
        \nLeftOut_80[3] , \nLeftOut_80[2] , \nLeftOut_80[1] , \nLeftOut_80[0] 
        }), .outright({\nRightOut_80[16] , \nRightOut_80[15] , 
        \nRightOut_80[14] , \nRightOut_80[13] , \nRightOut_80[12] , 
        \nRightOut_80[11] , \nRightOut_80[10] , \nRightOut_80[9] , 
        \nRightOut_80[8] , \nRightOut_80[7] , \nRightOut_80[6] , 
        \nRightOut_80[5] , \nRightOut_80[4] , \nRightOut_80[3] , 
        \nRightOut_80[2] , \nRightOut_80[1] , \nRightOut_80[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_100 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink20[15] , \ScanLink20[14] , \ScanLink20[13] , 
        \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , \ScanLink20[9] , 
        \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , \ScanLink20[5] , 
        \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , \ScanLink20[1] , 
        \ScanLink20[0] }), .ScanOut({\ScanLink21[15] , \ScanLink21[14] , 
        \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , 
        \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , 
        \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , 
        \ScanLink21[1] , \ScanLink21[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_88[16] , \nLeftOut_88[15] , \nLeftOut_88[14] , 
        \nLeftOut_88[13] , \nLeftOut_88[12] , \nLeftOut_88[11] , 
        \nLeftOut_88[10] , \nLeftOut_88[9] , \nLeftOut_88[8] , 
        \nLeftOut_88[7] , \nLeftOut_88[6] , \nLeftOut_88[5] , \nLeftOut_88[4] , 
        \nLeftOut_88[3] , \nLeftOut_88[2] , \nLeftOut_88[1] , \nLeftOut_88[0] 
        }), .inright({\nLeftOut_89[16] , \nLeftOut_89[15] , \nLeftOut_89[14] , 
        \nLeftOut_89[13] , \nLeftOut_89[12] , \nLeftOut_89[11] , 
        \nLeftOut_89[10] , \nLeftOut_89[9] , \nLeftOut_89[8] , 
        \nLeftOut_89[7] , \nLeftOut_89[6] , \nLeftOut_89[5] , \nLeftOut_89[4] , 
        \nLeftOut_89[3] , \nLeftOut_89[2] , \nLeftOut_89[1] , \nLeftOut_89[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s12_SCAN1 node_59 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_41[16] , \nRightOut_41[15] , \nRightOut_41[14] , 
        \nRightOut_41[13] , \nRightOut_41[12] , \nRightOut_41[11] , 
        \nRightOut_41[10] , \nRightOut_41[9] , \nRightOut_41[8] , 
        \nRightOut_41[7] , \nRightOut_41[6] , \nRightOut_41[5] , 
        \nRightOut_41[4] , \nRightOut_41[3] , \nRightOut_41[2] , 
        \nRightOut_41[1] , \nRightOut_41[0] }), .inright({\nRightOut_43[16] , 
        \nRightOut_43[15] , \nRightOut_43[14] , \nRightOut_43[13] , 
        \nRightOut_43[12] , \nRightOut_43[11] , \nRightOut_43[10] , 
        \nRightOut_43[9] , \nRightOut_43[8] , \nRightOut_43[7] , 
        \nRightOut_43[6] , \nRightOut_43[5] , \nRightOut_43[4] , 
        \nRightOut_43[3] , \nRightOut_43[2] , \nRightOut_43[1] , 
        \nRightOut_43[0] }), .outleft({\nLeftOut_59[16] , \nLeftOut_59[15] , 
        \nLeftOut_59[14] , \nLeftOut_59[13] , \nLeftOut_59[12] , 
        \nLeftOut_59[11] , \nLeftOut_59[10] , \nLeftOut_59[9] , 
        \nLeftOut_59[8] , \nLeftOut_59[7] , \nLeftOut_59[6] , \nLeftOut_59[5] , 
        \nLeftOut_59[4] , \nLeftOut_59[3] , \nLeftOut_59[2] , \nLeftOut_59[1] , 
        \nLeftOut_59[0] }), .outright({\nRightOut_59[16] , \nRightOut_59[15] , 
        \nRightOut_59[14] , \nRightOut_59[13] , \nRightOut_59[12] , 
        \nRightOut_59[11] , \nRightOut_59[10] , \nRightOut_59[9] , 
        \nRightOut_59[8] , \nRightOut_59[7] , \nRightOut_59[6] , 
        \nRightOut_59[5] , \nRightOut_59[4] , \nRightOut_59[3] , 
        \nRightOut_59[2] , \nRightOut_59[1] , \nRightOut_59[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink0[15] , \ScanLink0[14] , \ScanLink0[13] , 
        \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , \ScanLink0[9] , 
        \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , \ScanLink0[5] , 
        \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , \ScanLink0[1] , 
        \ScanLink0[0] }), .ScanOut({\ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_0[16] , \nLeftOut_0[15] , \nLeftOut_0[14] , \nLeftOut_0[13] , 
        \nLeftOut_0[12] , \nLeftOut_0[11] , \nLeftOut_0[10] , \nLeftOut_0[9] , 
        \nLeftOut_0[8] , \nLeftOut_0[7] , \nLeftOut_0[6] , \nLeftOut_0[5] , 
        \nLeftOut_0[4] , \nLeftOut_0[3] , \nLeftOut_0[2] , \nLeftOut_0[1] , 
        \nLeftOut_0[0] }), .inright({\nRightOut_0[16] , \nRightOut_0[15] , 
        \nRightOut_0[14] , \nRightOut_0[13] , \nRightOut_0[12] , 
        \nRightOut_0[11] , \nRightOut_0[10] , \nRightOut_0[9] , 
        \nRightOut_0[8] , \nRightOut_0[7] , \nRightOut_0[6] , \nRightOut_0[5] , 
        \nRightOut_0[4] , \nRightOut_0[3] , \nRightOut_0[2] , \nRightOut_0[1] , 
        \nRightOut_0[0] }), .outleft({\nLeftOut_0[16] , \nLeftOut_0[15] , 
        \nLeftOut_0[14] , \nLeftOut_0[13] , \nLeftOut_0[12] , \nLeftOut_0[11] , 
        \nLeftOut_0[10] , \nLeftOut_0[9] , \nLeftOut_0[8] , \nLeftOut_0[7] , 
        \nLeftOut_0[6] , \nLeftOut_0[5] , \nLeftOut_0[4] , \nLeftOut_0[3] , 
        \nLeftOut_0[2] , \nLeftOut_0[1] , \nLeftOut_0[0] }), .outright({
        \nRightOut_0[16] , \nRightOut_0[15] , \nRightOut_0[14] , 
        \nRightOut_0[13] , \nRightOut_0[12] , \nRightOut_0[11] , 
        \nRightOut_0[10] , \nRightOut_0[9] , \nRightOut_0[8] , 
        \nRightOut_0[7] , \nRightOut_0[6] , \nRightOut_0[5] , \nRightOut_0[4] , 
        \nRightOut_0[3] , \nRightOut_0[2] , \nRightOut_0[1] , \nRightOut_0[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink2[15] , \ScanLink2[14] , \ScanLink2[13] , 
        \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , \ScanLink2[9] , 
        \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , \ScanLink2[5] , 
        \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , \ScanLink2[1] , 
        \ScanLink2[0] }), .ScanOut({\ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_2[16] , \nLeftOut_2[15] , \nLeftOut_2[14] , \nLeftOut_2[13] , 
        \nLeftOut_2[12] , \nLeftOut_2[11] , \nLeftOut_2[10] , \nLeftOut_2[9] , 
        \nLeftOut_2[8] , \nLeftOut_2[7] , \nLeftOut_2[6] , \nLeftOut_2[5] , 
        \nLeftOut_2[4] , \nLeftOut_2[3] , \nLeftOut_2[2] , \nLeftOut_2[1] , 
        \nLeftOut_2[0] }), .inright({\nRightOut_2[16] , \nRightOut_2[15] , 
        \nRightOut_2[14] , \nRightOut_2[13] , \nRightOut_2[12] , 
        \nRightOut_2[11] , \nRightOut_2[10] , \nRightOut_2[9] , 
        \nRightOut_2[8] , \nRightOut_2[7] , \nRightOut_2[6] , \nRightOut_2[5] , 
        \nRightOut_2[4] , \nRightOut_2[3] , \nRightOut_2[2] , \nRightOut_2[1] , 
        \nRightOut_2[0] }), .outleft({\nLeftOut_2[16] , \nLeftOut_2[15] , 
        \nLeftOut_2[14] , \nLeftOut_2[13] , \nLeftOut_2[12] , \nLeftOut_2[11] , 
        \nLeftOut_2[10] , \nLeftOut_2[9] , \nLeftOut_2[8] , \nLeftOut_2[7] , 
        \nLeftOut_2[6] , \nLeftOut_2[5] , \nLeftOut_2[4] , \nLeftOut_2[3] , 
        \nLeftOut_2[2] , \nLeftOut_2[1] , \nLeftOut_2[0] }), .outright({
        \nRightOut_2[16] , \nRightOut_2[15] , \nRightOut_2[14] , 
        \nRightOut_2[13] , \nRightOut_2[12] , \nRightOut_2[11] , 
        \nRightOut_2[10] , \nRightOut_2[9] , \nRightOut_2[8] , 
        \nRightOut_2[7] , \nRightOut_2[6] , \nRightOut_2[5] , \nRightOut_2[4] , 
        \nRightOut_2[3] , \nRightOut_2[2] , \nRightOut_2[1] , \nRightOut_2[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink3[15] , \ScanLink3[14] , \ScanLink3[13] , 
        \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , \ScanLink3[9] , 
        \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , \ScanLink3[5] , 
        \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , \ScanLink3[1] , 
        \ScanLink3[0] }), .ScanOut({\ScanLink4[15] , \ScanLink4[14] , 
        \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , 
        \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_3[16] , \nLeftOut_3[15] , \nLeftOut_3[14] , \nLeftOut_3[13] , 
        \nLeftOut_3[12] , \nLeftOut_3[11] , \nLeftOut_3[10] , \nLeftOut_3[9] , 
        \nLeftOut_3[8] , \nLeftOut_3[7] , \nLeftOut_3[6] , \nLeftOut_3[5] , 
        \nLeftOut_3[4] , \nLeftOut_3[3] , \nLeftOut_3[2] , \nLeftOut_3[1] , 
        \nLeftOut_3[0] }), .inright({\nRightOut_3[16] , \nRightOut_3[15] , 
        \nRightOut_3[14] , \nRightOut_3[13] , \nRightOut_3[12] , 
        \nRightOut_3[11] , \nRightOut_3[10] , \nRightOut_3[9] , 
        \nRightOut_3[8] , \nRightOut_3[7] , \nRightOut_3[6] , \nRightOut_3[5] , 
        \nRightOut_3[4] , \nRightOut_3[3] , \nRightOut_3[2] , \nRightOut_3[1] , 
        \nRightOut_3[0] }), .outleft({\nLeftOut_3[16] , \nLeftOut_3[15] , 
        \nLeftOut_3[14] , \nLeftOut_3[13] , \nLeftOut_3[12] , \nLeftOut_3[11] , 
        \nLeftOut_3[10] , \nLeftOut_3[9] , \nLeftOut_3[8] , \nLeftOut_3[7] , 
        \nLeftOut_3[6] , \nLeftOut_3[5] , \nLeftOut_3[4] , \nLeftOut_3[3] , 
        \nLeftOut_3[2] , \nLeftOut_3[1] , \nLeftOut_3[0] }), .outright({
        \nRightOut_3[16] , \nRightOut_3[15] , \nRightOut_3[14] , 
        \nRightOut_3[13] , \nRightOut_3[12] , \nRightOut_3[11] , 
        \nRightOut_3[10] , \nRightOut_3[9] , \nRightOut_3[8] , 
        \nRightOut_3[7] , \nRightOut_3[6] , \nRightOut_3[5] , \nRightOut_3[4] , 
        \nRightOut_3[3] , \nRightOut_3[2] , \nRightOut_3[1] , \nRightOut_3[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_19 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_3[16] , \nLeftOut_3[15] , \nLeftOut_3[14] , \nLeftOut_3[13] , 
        \nLeftOut_3[12] , \nLeftOut_3[11] , \nLeftOut_3[10] , \nLeftOut_3[9] , 
        \nLeftOut_3[8] , \nLeftOut_3[7] , \nLeftOut_3[6] , \nLeftOut_3[5] , 
        \nLeftOut_3[4] , \nLeftOut_3[3] , \nLeftOut_3[2] , \nLeftOut_3[1] , 
        \nLeftOut_3[0] }), .inright({\nRightOut_3[16] , \nRightOut_3[15] , 
        \nRightOut_3[14] , \nRightOut_3[13] , \nRightOut_3[12] , 
        \nRightOut_3[11] , \nRightOut_3[10] , \nRightOut_3[9] , 
        \nRightOut_3[8] , \nRightOut_3[7] , \nRightOut_3[6] , \nRightOut_3[5] , 
        \nRightOut_3[4] , \nRightOut_3[3] , \nRightOut_3[2] , \nRightOut_3[1] , 
        \nRightOut_3[0] }), .outleft({\nLeftOut_19[16] , \nLeftOut_19[15] , 
        \nLeftOut_19[14] , \nLeftOut_19[13] , \nLeftOut_19[12] , 
        \nLeftOut_19[11] , \nLeftOut_19[10] , \nLeftOut_19[9] , 
        \nLeftOut_19[8] , \nLeftOut_19[7] , \nLeftOut_19[6] , \nLeftOut_19[5] , 
        \nLeftOut_19[4] , \nLeftOut_19[3] , \nLeftOut_19[2] , \nLeftOut_19[1] , 
        \nLeftOut_19[0] }), .outright({\nRightOut_19[16] , \nRightOut_19[15] , 
        \nRightOut_19[14] , \nRightOut_19[13] , \nRightOut_19[12] , 
        \nRightOut_19[11] , \nRightOut_19[10] , \nRightOut_19[9] , 
        \nRightOut_19[8] , \nRightOut_19[7] , \nRightOut_19[6] , 
        \nRightOut_19[5] , \nRightOut_19[4] , \nRightOut_19[3] , 
        \nRightOut_19[2] , \nRightOut_19[1] , \nRightOut_19[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_25 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_9[16] , \nLeftOut_9[15] , \nLeftOut_9[14] , \nLeftOut_9[13] , 
        \nLeftOut_9[12] , \nLeftOut_9[11] , \nLeftOut_9[10] , \nLeftOut_9[9] , 
        \nLeftOut_9[8] , \nLeftOut_9[7] , \nLeftOut_9[6] , \nLeftOut_9[5] , 
        \nLeftOut_9[4] , \nLeftOut_9[3] , \nLeftOut_9[2] , \nLeftOut_9[1] , 
        \nLeftOut_9[0] }), .inright({\nRightOut_9[16] , \nRightOut_9[15] , 
        \nRightOut_9[14] , \nRightOut_9[13] , \nRightOut_9[12] , 
        \nRightOut_9[11] , \nRightOut_9[10] , \nRightOut_9[9] , 
        \nRightOut_9[8] , \nRightOut_9[7] , \nRightOut_9[6] , \nRightOut_9[5] , 
        \nRightOut_9[4] , \nRightOut_9[3] , \nRightOut_9[2] , \nRightOut_9[1] , 
        \nRightOut_9[0] }), .outleft({\nLeftOut_25[16] , \nLeftOut_25[15] , 
        \nLeftOut_25[14] , \nLeftOut_25[13] , \nLeftOut_25[12] , 
        \nLeftOut_25[11] , \nLeftOut_25[10] , \nLeftOut_25[9] , 
        \nLeftOut_25[8] , \nLeftOut_25[7] , \nLeftOut_25[6] , \nLeftOut_25[5] , 
        \nLeftOut_25[4] , \nLeftOut_25[3] , \nLeftOut_25[2] , \nLeftOut_25[1] , 
        \nLeftOut_25[0] }), .outright({\nRightOut_25[16] , \nRightOut_25[15] , 
        \nRightOut_25[14] , \nRightOut_25[13] , \nRightOut_25[12] , 
        \nRightOut_25[11] , \nRightOut_25[10] , \nRightOut_25[9] , 
        \nRightOut_25[8] , \nRightOut_25[7] , \nRightOut_25[6] , 
        \nRightOut_25[5] , \nRightOut_25[4] , \nRightOut_25[3] , 
        \nRightOut_25[2] , \nRightOut_25[1] , \nRightOut_25[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s9_SCAN1 node_89 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_65[16] , \nRightOut_65[15] , \nRightOut_65[14] , 
        \nRightOut_65[13] , \nRightOut_65[12] , \nRightOut_65[11] , 
        \nRightOut_65[10] , \nRightOut_65[9] , \nRightOut_65[8] , 
        \nRightOut_65[7] , \nRightOut_65[6] , \nRightOut_65[5] , 
        \nRightOut_65[4] , \nRightOut_65[3] , \nRightOut_65[2] , 
        \nRightOut_65[1] , \nRightOut_65[0] }), .inright({\nRightOut_73[16] , 
        \nRightOut_73[15] , \nRightOut_73[14] , \nRightOut_73[13] , 
        \nRightOut_73[12] , \nRightOut_73[11] , \nRightOut_73[10] , 
        \nRightOut_73[9] , \nRightOut_73[8] , \nRightOut_73[7] , 
        \nRightOut_73[6] , \nRightOut_73[5] , \nRightOut_73[4] , 
        \nRightOut_73[3] , \nRightOut_73[2] , \nRightOut_73[1] , 
        \nRightOut_73[0] }), .outleft({\nLeftOut_89[16] , \nLeftOut_89[15] , 
        \nLeftOut_89[14] , \nLeftOut_89[13] , \nLeftOut_89[12] , 
        \nLeftOut_89[11] , \nLeftOut_89[10] , \nLeftOut_89[9] , 
        \nLeftOut_89[8] , \nLeftOut_89[7] , \nLeftOut_89[6] , \nLeftOut_89[5] , 
        \nLeftOut_89[4] , \nLeftOut_89[3] , \nLeftOut_89[2] , \nLeftOut_89[1] , 
        \nLeftOut_89[0] }), .outright({\nRightOut_89[16] , \nRightOut_89[15] , 
        \nRightOut_89[14] , \nRightOut_89[13] , \nRightOut_89[12] , 
        \nRightOut_89[11] , \nRightOut_89[10] , \nRightOut_89[9] , 
        \nRightOut_89[8] , \nRightOut_89[7] , \nRightOut_89[6] , 
        \nRightOut_89[5] , \nRightOut_89[4] , \nRightOut_89[3] , 
        \nRightOut_89[2] , \nRightOut_89[1] , \nRightOut_89[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_109 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink29[15] , \ScanLink29[14] , \ScanLink29[13] , 
        \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , \ScanLink29[9] , 
        \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , \ScanLink29[5] , 
        \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , \ScanLink29[1] , 
        \ScanLink29[0] }), .ScanOut({\ScanLink30[15] , \ScanLink30[14] , 
        \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , 
        \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , 
        \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , 
        \ScanLink30[1] , \ScanLink30[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_90[16] , \nRightOut_90[15] , \nRightOut_90[14] , 
        \nRightOut_90[13] , \nRightOut_90[12] , \nRightOut_90[11] , 
        \nRightOut_90[10] , \nRightOut_90[9] , \nRightOut_90[8] , 
        \nRightOut_90[7] , \nRightOut_90[6] , \nRightOut_90[5] , 
        \nRightOut_90[4] , \nRightOut_90[3] , \nRightOut_90[2] , 
        \nRightOut_90[1] , \nRightOut_90[0] }), .inright({\nRightOut_91[16] , 
        \nRightOut_91[15] , \nRightOut_91[14] , \nRightOut_91[13] , 
        \nRightOut_91[12] , \nRightOut_91[11] , \nRightOut_91[10] , 
        \nRightOut_91[9] , \nRightOut_91[8] , \nRightOut_91[7] , 
        \nRightOut_91[6] , \nRightOut_91[5] , \nRightOut_91[4] , 
        \nRightOut_91[3] , \nRightOut_91[2] , \nRightOut_91[1] , 
        \nRightOut_91[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_22 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_6[16] , \nLeftOut_6[15] , \nLeftOut_6[14] , \nLeftOut_6[13] , 
        \nLeftOut_6[12] , \nLeftOut_6[11] , \nLeftOut_6[10] , \nLeftOut_6[9] , 
        \nLeftOut_6[8] , \nLeftOut_6[7] , \nLeftOut_6[6] , \nLeftOut_6[5] , 
        \nLeftOut_6[4] , \nLeftOut_6[3] , \nLeftOut_6[2] , \nLeftOut_6[1] , 
        \nLeftOut_6[0] }), .inright({\nRightOut_6[16] , \nRightOut_6[15] , 
        \nRightOut_6[14] , \nRightOut_6[13] , \nRightOut_6[12] , 
        \nRightOut_6[11] , \nRightOut_6[10] , \nRightOut_6[9] , 
        \nRightOut_6[8] , \nRightOut_6[7] , \nRightOut_6[6] , \nRightOut_6[5] , 
        \nRightOut_6[4] , \nRightOut_6[3] , \nRightOut_6[2] , \nRightOut_6[1] , 
        \nRightOut_6[0] }), .outleft({\nLeftOut_22[16] , \nLeftOut_22[15] , 
        \nLeftOut_22[14] , \nLeftOut_22[13] , \nLeftOut_22[12] , 
        \nLeftOut_22[11] , \nLeftOut_22[10] , \nLeftOut_22[9] , 
        \nLeftOut_22[8] , \nLeftOut_22[7] , \nLeftOut_22[6] , \nLeftOut_22[5] , 
        \nLeftOut_22[4] , \nLeftOut_22[3] , \nLeftOut_22[2] , \nLeftOut_22[1] , 
        \nLeftOut_22[0] }), .outright({\nRightOut_22[16] , \nRightOut_22[15] , 
        \nRightOut_22[14] , \nRightOut_22[13] , \nRightOut_22[12] , 
        \nRightOut_22[11] , \nRightOut_22[10] , \nRightOut_22[9] , 
        \nRightOut_22[8] , \nRightOut_22[7] , \nRightOut_22[6] , 
        \nRightOut_22[5] , \nRightOut_22[4] , \nRightOut_22[3] , 
        \nRightOut_22[2] , \nRightOut_22[1] , \nRightOut_22[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_39 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_22[16] , \nRightOut_22[15] , \nRightOut_22[14] , 
        \nRightOut_22[13] , \nRightOut_22[12] , \nRightOut_22[11] , 
        \nRightOut_22[10] , \nRightOut_22[9] , \nRightOut_22[8] , 
        \nRightOut_22[7] , \nRightOut_22[6] , \nRightOut_22[5] , 
        \nRightOut_22[4] , \nRightOut_22[3] , \nRightOut_22[2] , 
        \nRightOut_22[1] , \nRightOut_22[0] }), .inright({\nRightOut_23[16] , 
        \nRightOut_23[15] , \nRightOut_23[14] , \nRightOut_23[13] , 
        \nRightOut_23[12] , \nRightOut_23[11] , \nRightOut_23[10] , 
        \nRightOut_23[9] , \nRightOut_23[8] , \nRightOut_23[7] , 
        \nRightOut_23[6] , \nRightOut_23[5] , \nRightOut_23[4] , 
        \nRightOut_23[3] , \nRightOut_23[2] , \nRightOut_23[1] , 
        \nRightOut_23[0] }), .outleft({\nLeftOut_39[16] , \nLeftOut_39[15] , 
        \nLeftOut_39[14] , \nLeftOut_39[13] , \nLeftOut_39[12] , 
        \nLeftOut_39[11] , \nLeftOut_39[10] , \nLeftOut_39[9] , 
        \nLeftOut_39[8] , \nLeftOut_39[7] , \nLeftOut_39[6] , \nLeftOut_39[5] , 
        \nLeftOut_39[4] , \nLeftOut_39[3] , \nLeftOut_39[2] , \nLeftOut_39[1] , 
        \nLeftOut_39[0] }), .outright({\nRightOut_39[16] , \nRightOut_39[15] , 
        \nRightOut_39[14] , \nRightOut_39[13] , \nRightOut_39[12] , 
        \nRightOut_39[11] , \nRightOut_39[10] , \nRightOut_39[9] , 
        \nRightOut_39[8] , \nRightOut_39[7] , \nRightOut_39[6] , 
        \nRightOut_39[5] , \nRightOut_39[4] , \nRightOut_39[3] , 
        \nRightOut_39[2] , \nRightOut_39[1] , \nRightOut_39[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_50 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_32[16] , \nRightOut_32[15] , \nRightOut_32[14] , 
        \nRightOut_32[13] , \nRightOut_32[12] , \nRightOut_32[11] , 
        \nRightOut_32[10] , \nRightOut_32[9] , \nRightOut_32[8] , 
        \nRightOut_32[7] , \nRightOut_32[6] , \nRightOut_32[5] , 
        \nRightOut_32[4] , \nRightOut_32[3] , \nRightOut_32[2] , 
        \nRightOut_32[1] , \nRightOut_32[0] }), .inright({\nRightOut_34[16] , 
        \nRightOut_34[15] , \nRightOut_34[14] , \nRightOut_34[13] , 
        \nRightOut_34[12] , \nRightOut_34[11] , \nRightOut_34[10] , 
        \nRightOut_34[9] , \nRightOut_34[8] , \nRightOut_34[7] , 
        \nRightOut_34[6] , \nRightOut_34[5] , \nRightOut_34[4] , 
        \nRightOut_34[3] , \nRightOut_34[2] , \nRightOut_34[1] , 
        \nRightOut_34[0] }), .outleft({\nLeftOut_50[16] , \nLeftOut_50[15] , 
        \nLeftOut_50[14] , \nLeftOut_50[13] , \nLeftOut_50[12] , 
        \nLeftOut_50[11] , \nLeftOut_50[10] , \nLeftOut_50[9] , 
        \nLeftOut_50[8] , \nLeftOut_50[7] , \nLeftOut_50[6] , \nLeftOut_50[5] , 
        \nLeftOut_50[4] , \nLeftOut_50[3] , \nLeftOut_50[2] , \nLeftOut_50[1] , 
        \nLeftOut_50[0] }), .outright({\nRightOut_50[16] , \nRightOut_50[15] , 
        \nRightOut_50[14] , \nRightOut_50[13] , \nRightOut_50[12] , 
        \nRightOut_50[11] , \nRightOut_50[10] , \nRightOut_50[9] , 
        \nRightOut_50[8] , \nRightOut_50[7] , \nRightOut_50[6] , 
        \nRightOut_50[5] , \nRightOut_50[4] , \nRightOut_50[3] , 
        \nRightOut_50[2] , \nRightOut_50[1] , \nRightOut_50[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s12_SCAN1 node_92 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_68[16] , \nRightOut_68[15] , \nRightOut_68[14] , 
        \nRightOut_68[13] , \nRightOut_68[12] , \nRightOut_68[11] , 
        \nRightOut_68[10] , \nRightOut_68[9] , \nRightOut_68[8] , 
        \nRightOut_68[7] , \nRightOut_68[6] , \nRightOut_68[5] , 
        \nRightOut_68[4] , \nRightOut_68[3] , \nRightOut_68[2] , 
        \nRightOut_68[1] , \nRightOut_68[0] }), .inright({\nRightOut_76[16] , 
        \nRightOut_76[15] , \nRightOut_76[14] , \nRightOut_76[13] , 
        \nRightOut_76[12] , \nRightOut_76[11] , \nRightOut_76[10] , 
        \nRightOut_76[9] , \nRightOut_76[8] , \nRightOut_76[7] , 
        \nRightOut_76[6] , \nRightOut_76[5] , \nRightOut_76[4] , 
        \nRightOut_76[3] , \nRightOut_76[2] , \nRightOut_76[1] , 
        \nRightOut_76[0] }), .outleft({\nLeftOut_92[16] , \nLeftOut_92[15] , 
        \nLeftOut_92[14] , \nLeftOut_92[13] , \nLeftOut_92[12] , 
        \nLeftOut_92[11] , \nLeftOut_92[10] , \nLeftOut_92[9] , 
        \nLeftOut_92[8] , \nLeftOut_92[7] , \nLeftOut_92[6] , \nLeftOut_92[5] , 
        \nLeftOut_92[4] , \nLeftOut_92[3] , \nLeftOut_92[2] , \nLeftOut_92[1] , 
        \nLeftOut_92[0] }), .outright({\nRightOut_92[16] , \nRightOut_92[15] , 
        \nRightOut_92[14] , \nRightOut_92[13] , \nRightOut_92[12] , 
        \nRightOut_92[11] , \nRightOut_92[10] , \nRightOut_92[9] , 
        \nRightOut_92[8] , \nRightOut_92[7] , \nRightOut_92[6] , 
        \nRightOut_92[5] , \nRightOut_92[4] , \nRightOut_92[3] , 
        \nRightOut_92[2] , \nRightOut_92[1] , \nRightOut_92[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s4_SCAN1 node_57 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_41[16] , \nLeftOut_41[15] , \nLeftOut_41[14] , 
        \nLeftOut_41[13] , \nLeftOut_41[12] , \nLeftOut_41[11] , 
        \nLeftOut_41[10] , \nLeftOut_41[9] , \nLeftOut_41[8] , 
        \nLeftOut_41[7] , \nLeftOut_41[6] , \nLeftOut_41[5] , \nLeftOut_41[4] , 
        \nLeftOut_41[3] , \nLeftOut_41[2] , \nLeftOut_41[1] , \nLeftOut_41[0] 
        }), .inright({\nLeftOut_43[16] , \nLeftOut_43[15] , \nLeftOut_43[14] , 
        \nLeftOut_43[13] , \nLeftOut_43[12] , \nLeftOut_43[11] , 
        \nLeftOut_43[10] , \nLeftOut_43[9] , \nLeftOut_43[8] , 
        \nLeftOut_43[7] , \nLeftOut_43[6] , \nLeftOut_43[5] , \nLeftOut_43[4] , 
        \nLeftOut_43[3] , \nLeftOut_43[2] , \nLeftOut_43[1] , \nLeftOut_43[0] 
        }), .outleft({\nLeftOut_57[16] , \nLeftOut_57[15] , \nLeftOut_57[14] , 
        \nLeftOut_57[13] , \nLeftOut_57[12] , \nLeftOut_57[11] , 
        \nLeftOut_57[10] , \nLeftOut_57[9] , \nLeftOut_57[8] , 
        \nLeftOut_57[7] , \nLeftOut_57[6] , \nLeftOut_57[5] , \nLeftOut_57[4] , 
        \nLeftOut_57[3] , \nLeftOut_57[2] , \nLeftOut_57[1] , \nLeftOut_57[0] 
        }), .outright({\nRightOut_57[16] , \nRightOut_57[15] , 
        \nRightOut_57[14] , \nRightOut_57[13] , \nRightOut_57[12] , 
        \nRightOut_57[11] , \nRightOut_57[10] , \nRightOut_57[9] , 
        \nRightOut_57[8] , \nRightOut_57[7] , \nRightOut_57[6] , 
        \nRightOut_57[5] , \nRightOut_57[4] , \nRightOut_57[3] , 
        \nRightOut_57[2] , \nRightOut_57[1] , \nRightOut_57[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s12_SCAN1 node_70 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_50[16] , \nRightOut_50[15] , \nRightOut_50[14] , 
        \nRightOut_50[13] , \nRightOut_50[12] , \nRightOut_50[11] , 
        \nRightOut_50[10] , \nRightOut_50[9] , \nRightOut_50[8] , 
        \nRightOut_50[7] , \nRightOut_50[6] , \nRightOut_50[5] , 
        \nRightOut_50[4] , \nRightOut_50[3] , \nRightOut_50[2] , 
        \nRightOut_50[1] , \nRightOut_50[0] }), .inright({\nRightOut_54[16] , 
        \nRightOut_54[15] , \nRightOut_54[14] , \nRightOut_54[13] , 
        \nRightOut_54[12] , \nRightOut_54[11] , \nRightOut_54[10] , 
        \nRightOut_54[9] , \nRightOut_54[8] , \nRightOut_54[7] , 
        \nRightOut_54[6] , \nRightOut_54[5] , \nRightOut_54[4] , 
        \nRightOut_54[3] , \nRightOut_54[2] , \nRightOut_54[1] , 
        \nRightOut_54[0] }), .outleft({\nLeftOut_70[16] , \nLeftOut_70[15] , 
        \nLeftOut_70[14] , \nLeftOut_70[13] , \nLeftOut_70[12] , 
        \nLeftOut_70[11] , \nLeftOut_70[10] , \nLeftOut_70[9] , 
        \nLeftOut_70[8] , \nLeftOut_70[7] , \nLeftOut_70[6] , \nLeftOut_70[5] , 
        \nLeftOut_70[4] , \nLeftOut_70[3] , \nLeftOut_70[2] , \nLeftOut_70[1] , 
        \nLeftOut_70[0] }), .outright({\nRightOut_70[16] , \nRightOut_70[15] , 
        \nRightOut_70[14] , \nRightOut_70[13] , \nRightOut_70[12] , 
        \nRightOut_70[11] , \nRightOut_70[10] , \nRightOut_70[9] , 
        \nRightOut_70[8] , \nRightOut_70[7] , \nRightOut_70[6] , 
        \nRightOut_70[5] , \nRightOut_70[4] , \nRightOut_70[3] , 
        \nRightOut_70[2] , \nRightOut_70[1] , \nRightOut_70[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s10_SCAN1 node_77 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_57[16] , \nRightOut_57[15] , \nRightOut_57[14] , 
        \nRightOut_57[13] , \nRightOut_57[12] , \nRightOut_57[11] , 
        \nRightOut_57[10] , \nRightOut_57[9] , \nRightOut_57[8] , 
        \nRightOut_57[7] , \nRightOut_57[6] , \nRightOut_57[5] , 
        \nRightOut_57[4] , \nRightOut_57[3] , \nRightOut_57[2] , 
        \nRightOut_57[1] , \nRightOut_57[0] }), .inright({\nRightOut_61[16] , 
        \nRightOut_61[15] , \nRightOut_61[14] , \nRightOut_61[13] , 
        \nRightOut_61[12] , \nRightOut_61[11] , \nRightOut_61[10] , 
        \nRightOut_61[9] , \nRightOut_61[8] , \nRightOut_61[7] , 
        \nRightOut_61[6] , \nRightOut_61[5] , \nRightOut_61[4] , 
        \nRightOut_61[3] , \nRightOut_61[2] , \nRightOut_61[1] , 
        \nRightOut_61[0] }), .outleft({\nLeftOut_77[16] , \nLeftOut_77[15] , 
        \nLeftOut_77[14] , \nLeftOut_77[13] , \nLeftOut_77[12] , 
        \nLeftOut_77[11] , \nLeftOut_77[10] , \nLeftOut_77[9] , 
        \nLeftOut_77[8] , \nLeftOut_77[7] , \nLeftOut_77[6] , \nLeftOut_77[5] , 
        \nLeftOut_77[4] , \nLeftOut_77[3] , \nLeftOut_77[2] , \nLeftOut_77[1] , 
        \nLeftOut_77[0] }), .outright({\nRightOut_77[16] , \nRightOut_77[15] , 
        \nRightOut_77[14] , \nRightOut_77[13] , \nRightOut_77[12] , 
        \nRightOut_77[11] , \nRightOut_77[10] , \nRightOut_77[9] , 
        \nRightOut_77[8] , \nRightOut_77[7] , \nRightOut_77[6] , 
        \nRightOut_77[5] , \nRightOut_77[4] , \nRightOut_77[3] , 
        \nRightOut_77[2] , \nRightOut_77[1] , \nRightOut_77[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s15_SCAN1 node_95 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_71[16] , \nRightOut_71[15] , \nRightOut_71[14] , 
        \nRightOut_71[13] , \nRightOut_71[12] , \nRightOut_71[11] , 
        \nRightOut_71[10] , \nRightOut_71[9] , \nRightOut_71[8] , 
        \nRightOut_71[7] , \nRightOut_71[6] , \nRightOut_71[5] , 
        \nRightOut_71[4] , \nRightOut_71[3] , \nRightOut_71[2] , 
        \nRightOut_71[1] , \nRightOut_71[0] }), .inright({\nRightOut_79[16] , 
        \nRightOut_79[15] , \nRightOut_79[14] , \nRightOut_79[13] , 
        \nRightOut_79[12] , \nRightOut_79[11] , \nRightOut_79[10] , 
        \nRightOut_79[9] , \nRightOut_79[8] , \nRightOut_79[7] , 
        \nRightOut_79[6] , \nRightOut_79[5] , \nRightOut_79[4] , 
        \nRightOut_79[3] , \nRightOut_79[2] , \nRightOut_79[1] , 
        \nRightOut_79[0] }), .outleft({\nLeftOut_95[16] , \nLeftOut_95[15] , 
        \nLeftOut_95[14] , \nLeftOut_95[13] , \nLeftOut_95[12] , 
        \nLeftOut_95[11] , \nLeftOut_95[10] , \nLeftOut_95[9] , 
        \nLeftOut_95[8] , \nLeftOut_95[7] , \nLeftOut_95[6] , \nLeftOut_95[5] , 
        \nLeftOut_95[4] , \nLeftOut_95[3] , \nLeftOut_95[2] , \nLeftOut_95[1] , 
        \nLeftOut_95[0] }), .outright({\nRightOut_95[16] , \nRightOut_95[15] , 
        \nRightOut_95[14] , \nRightOut_95[13] , \nRightOut_95[12] , 
        \nRightOut_95[11] , \nRightOut_95[10] , \nRightOut_95[9] , 
        \nRightOut_95[8] , \nRightOut_95[7] , \nRightOut_95[6] , 
        \nRightOut_95[5] , \nRightOut_95[4] , \nRightOut_95[3] , 
        \nRightOut_95[2] , \nRightOut_95[1] , \nRightOut_95[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_16 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_0[16] , \nLeftOut_0[15] , \nLeftOut_0[14] , \nLeftOut_0[13] , 
        \nLeftOut_0[12] , \nLeftOut_0[11] , \nLeftOut_0[10] , \nLeftOut_0[9] , 
        \nLeftOut_0[8] , \nLeftOut_0[7] , \nLeftOut_0[6] , \nLeftOut_0[5] , 
        \nLeftOut_0[4] , \nLeftOut_0[3] , \nLeftOut_0[2] , \nLeftOut_0[1] , 
        \nLeftOut_0[0] }), .inright({\nRightOut_0[16] , \nRightOut_0[15] , 
        \nRightOut_0[14] , \nRightOut_0[13] , \nRightOut_0[12] , 
        \nRightOut_0[11] , \nRightOut_0[10] , \nRightOut_0[9] , 
        \nRightOut_0[8] , \nRightOut_0[7] , \nRightOut_0[6] , \nRightOut_0[5] , 
        \nRightOut_0[4] , \nRightOut_0[3] , \nRightOut_0[2] , \nRightOut_0[1] , 
        \nRightOut_0[0] }), .outleft({\nLeftOut_16[16] , \nLeftOut_16[15] , 
        \nLeftOut_16[14] , \nLeftOut_16[13] , \nLeftOut_16[12] , 
        \nLeftOut_16[11] , \nLeftOut_16[10] , \nLeftOut_16[9] , 
        \nLeftOut_16[8] , \nLeftOut_16[7] , \nLeftOut_16[6] , \nLeftOut_16[5] , 
        \nLeftOut_16[4] , \nLeftOut_16[3] , \nLeftOut_16[2] , \nLeftOut_16[1] , 
        \nLeftOut_16[0] }), .outright({\nRightOut_16[16] , \nRightOut_16[15] , 
        \nRightOut_16[14] , \nRightOut_16[13] , \nRightOut_16[12] , 
        \nRightOut_16[11] , \nRightOut_16[10] , \nRightOut_16[9] , 
        \nRightOut_16[8] , \nRightOut_16[7] , \nRightOut_16[6] , 
        \nRightOut_16[5] , \nRightOut_16[4] , \nRightOut_16[3] , 
        \nRightOut_16[2] , \nRightOut_16[1] , \nRightOut_16[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_17 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_1[16] , \nLeftOut_1[15] , \nLeftOut_1[14] , \nLeftOut_1[13] , 
        \nLeftOut_1[12] , \nLeftOut_1[11] , \nLeftOut_1[10] , \nLeftOut_1[9] , 
        \nLeftOut_1[8] , \nLeftOut_1[7] , \nLeftOut_1[6] , \nLeftOut_1[5] , 
        \nLeftOut_1[4] , \nLeftOut_1[3] , \nLeftOut_1[2] , \nLeftOut_1[1] , 
        \nLeftOut_1[0] }), .inright({\nRightOut_1[16] , \nRightOut_1[15] , 
        \nRightOut_1[14] , \nRightOut_1[13] , \nRightOut_1[12] , 
        \nRightOut_1[11] , \nRightOut_1[10] , \nRightOut_1[9] , 
        \nRightOut_1[8] , \nRightOut_1[7] , \nRightOut_1[6] , \nRightOut_1[5] , 
        \nRightOut_1[4] , \nRightOut_1[3] , \nRightOut_1[2] , \nRightOut_1[1] , 
        \nRightOut_1[0] }), .outleft({\nLeftOut_17[16] , \nLeftOut_17[15] , 
        \nLeftOut_17[14] , \nLeftOut_17[13] , \nLeftOut_17[12] , 
        \nLeftOut_17[11] , \nLeftOut_17[10] , \nLeftOut_17[9] , 
        \nLeftOut_17[8] , \nLeftOut_17[7] , \nLeftOut_17[6] , \nLeftOut_17[5] , 
        \nLeftOut_17[4] , \nLeftOut_17[3] , \nLeftOut_17[2] , \nLeftOut_17[1] , 
        \nLeftOut_17[0] }), .outright({\nRightOut_17[16] , \nRightOut_17[15] , 
        \nRightOut_17[14] , \nRightOut_17[13] , \nRightOut_17[12] , 
        \nRightOut_17[11] , \nRightOut_17[10] , \nRightOut_17[9] , 
        \nRightOut_17[8] , \nRightOut_17[7] , \nRightOut_17[6] , 
        \nRightOut_17[5] , \nRightOut_17[4] , \nRightOut_17[3] , 
        \nRightOut_17[2] , \nRightOut_17[1] , \nRightOut_17[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s14_SCAN1 node_79 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_59[16] , \nRightOut_59[15] , \nRightOut_59[14] , 
        \nRightOut_59[13] , \nRightOut_59[12] , \nRightOut_59[11] , 
        \nRightOut_59[10] , \nRightOut_59[9] , \nRightOut_59[8] , 
        \nRightOut_59[7] , \nRightOut_59[6] , \nRightOut_59[5] , 
        \nRightOut_59[4] , \nRightOut_59[3] , \nRightOut_59[2] , 
        \nRightOut_59[1] , \nRightOut_59[0] }), .inright({\nRightOut_63[16] , 
        \nRightOut_63[15] , \nRightOut_63[14] , \nRightOut_63[13] , 
        \nRightOut_63[12] , \nRightOut_63[11] , \nRightOut_63[10] , 
        \nRightOut_63[9] , \nRightOut_63[8] , \nRightOut_63[7] , 
        \nRightOut_63[6] , \nRightOut_63[5] , \nRightOut_63[4] , 
        \nRightOut_63[3] , \nRightOut_63[2] , \nRightOut_63[1] , 
        \nRightOut_63[0] }), .outleft({\nLeftOut_79[16] , \nLeftOut_79[15] , 
        \nLeftOut_79[14] , \nLeftOut_79[13] , \nLeftOut_79[12] , 
        \nLeftOut_79[11] , \nLeftOut_79[10] , \nLeftOut_79[9] , 
        \nLeftOut_79[8] , \nLeftOut_79[7] , \nLeftOut_79[6] , \nLeftOut_79[5] , 
        \nLeftOut_79[4] , \nLeftOut_79[3] , \nLeftOut_79[2] , \nLeftOut_79[1] , 
        \nLeftOut_79[0] }), .outright({\nRightOut_79[16] , \nRightOut_79[15] , 
        \nRightOut_79[14] , \nRightOut_79[13] , \nRightOut_79[12] , 
        \nRightOut_79[11] , \nRightOut_79[10] , \nRightOut_79[9] , 
        \nRightOut_79[8] , \nRightOut_79[7] , \nRightOut_79[6] , 
        \nRightOut_79[5] , \nRightOut_79[4] , \nRightOut_79[3] , 
        \nRightOut_79[2] , \nRightOut_79[1] , \nRightOut_79[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_23 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_7[16] , \nLeftOut_7[15] , \nLeftOut_7[14] , \nLeftOut_7[13] , 
        \nLeftOut_7[12] , \nLeftOut_7[11] , \nLeftOut_7[10] , \nLeftOut_7[9] , 
        \nLeftOut_7[8] , \nLeftOut_7[7] , \nLeftOut_7[6] , \nLeftOut_7[5] , 
        \nLeftOut_7[4] , \nLeftOut_7[3] , \nLeftOut_7[2] , \nLeftOut_7[1] , 
        \nLeftOut_7[0] }), .inright({\nRightOut_7[16] , \nRightOut_7[15] , 
        \nRightOut_7[14] , \nRightOut_7[13] , \nRightOut_7[12] , 
        \nRightOut_7[11] , \nRightOut_7[10] , \nRightOut_7[9] , 
        \nRightOut_7[8] , \nRightOut_7[7] , \nRightOut_7[6] , \nRightOut_7[5] , 
        \nRightOut_7[4] , \nRightOut_7[3] , \nRightOut_7[2] , \nRightOut_7[1] , 
        \nRightOut_7[0] }), .outleft({\nLeftOut_23[16] , \nLeftOut_23[15] , 
        \nLeftOut_23[14] , \nLeftOut_23[13] , \nLeftOut_23[12] , 
        \nLeftOut_23[11] , \nLeftOut_23[10] , \nLeftOut_23[9] , 
        \nLeftOut_23[8] , \nLeftOut_23[7] , \nLeftOut_23[6] , \nLeftOut_23[5] , 
        \nLeftOut_23[4] , \nLeftOut_23[3] , \nLeftOut_23[2] , \nLeftOut_23[1] , 
        \nLeftOut_23[0] }), .outright({\nRightOut_23[16] , \nRightOut_23[15] , 
        \nRightOut_23[14] , \nRightOut_23[13] , \nRightOut_23[12] , 
        \nRightOut_23[11] , \nRightOut_23[10] , \nRightOut_23[9] , 
        \nRightOut_23[8] , \nRightOut_23[7] , \nRightOut_23[6] , 
        \nRightOut_23[5] , \nRightOut_23[4] , \nRightOut_23[3] , 
        \nRightOut_23[2] , \nRightOut_23[1] , \nRightOut_23[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_30 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_14[16] , \nLeftOut_14[15] , \nLeftOut_14[14] , 
        \nLeftOut_14[13] , \nLeftOut_14[12] , \nLeftOut_14[11] , 
        \nLeftOut_14[10] , \nLeftOut_14[9] , \nLeftOut_14[8] , 
        \nLeftOut_14[7] , \nLeftOut_14[6] , \nLeftOut_14[5] , \nLeftOut_14[4] , 
        \nLeftOut_14[3] , \nLeftOut_14[2] , \nLeftOut_14[1] , \nLeftOut_14[0] 
        }), .inright({\nRightOut_14[16] , \nRightOut_14[15] , 
        \nRightOut_14[14] , \nRightOut_14[13] , \nRightOut_14[12] , 
        \nRightOut_14[11] , \nRightOut_14[10] , \nRightOut_14[9] , 
        \nRightOut_14[8] , \nRightOut_14[7] , \nRightOut_14[6] , 
        \nRightOut_14[5] , \nRightOut_14[4] , \nRightOut_14[3] , 
        \nRightOut_14[2] , \nRightOut_14[1] , \nRightOut_14[0] }), .outleft({
        \nLeftOut_30[16] , \nLeftOut_30[15] , \nLeftOut_30[14] , 
        \nLeftOut_30[13] , \nLeftOut_30[12] , \nLeftOut_30[11] , 
        \nLeftOut_30[10] , \nLeftOut_30[9] , \nLeftOut_30[8] , 
        \nLeftOut_30[7] , \nLeftOut_30[6] , \nLeftOut_30[5] , \nLeftOut_30[4] , 
        \nLeftOut_30[3] , \nLeftOut_30[2] , \nLeftOut_30[1] , \nLeftOut_30[0] 
        }), .outright({\nRightOut_30[16] , \nRightOut_30[15] , 
        \nRightOut_30[14] , \nRightOut_30[13] , \nRightOut_30[12] , 
        \nRightOut_30[11] , \nRightOut_30[10] , \nRightOut_30[9] , 
        \nRightOut_30[8] , \nRightOut_30[7] , \nRightOut_30[6] , 
        \nRightOut_30[5] , \nRightOut_30[4] , \nRightOut_30[3] , 
        \nRightOut_30[2] , \nRightOut_30[1] , \nRightOut_30[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_45 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_28[16] , \nRightOut_28[15] , \nRightOut_28[14] , 
        \nRightOut_28[13] , \nRightOut_28[12] , \nRightOut_28[11] , 
        \nRightOut_28[10] , \nRightOut_28[9] , \nRightOut_28[8] , 
        \nRightOut_28[7] , \nRightOut_28[6] , \nRightOut_28[5] , 
        \nRightOut_28[4] , \nRightOut_28[3] , \nRightOut_28[2] , 
        \nRightOut_28[1] , \nRightOut_28[0] }), .inright({\nRightOut_29[16] , 
        \nRightOut_29[15] , \nRightOut_29[14] , \nRightOut_29[13] , 
        \nRightOut_29[12] , \nRightOut_29[11] , \nRightOut_29[10] , 
        \nRightOut_29[9] , \nRightOut_29[8] , \nRightOut_29[7] , 
        \nRightOut_29[6] , \nRightOut_29[5] , \nRightOut_29[4] , 
        \nRightOut_29[3] , \nRightOut_29[2] , \nRightOut_29[1] , 
        \nRightOut_29[0] }), .outleft({\nLeftOut_45[16] , \nLeftOut_45[15] , 
        \nLeftOut_45[14] , \nLeftOut_45[13] , \nLeftOut_45[12] , 
        \nLeftOut_45[11] , \nLeftOut_45[10] , \nLeftOut_45[9] , 
        \nLeftOut_45[8] , \nLeftOut_45[7] , \nLeftOut_45[6] , \nLeftOut_45[5] , 
        \nLeftOut_45[4] , \nLeftOut_45[3] , \nLeftOut_45[2] , \nLeftOut_45[1] , 
        \nLeftOut_45[0] }), .outright({\nRightOut_45[16] , \nRightOut_45[15] , 
        \nRightOut_45[14] , \nRightOut_45[13] , \nRightOut_45[12] , 
        \nRightOut_45[11] , \nRightOut_45[10] , \nRightOut_45[9] , 
        \nRightOut_45[8] , \nRightOut_45[7] , \nRightOut_45[6] , 
        \nRightOut_45[5] , \nRightOut_45[4] , \nRightOut_45[3] , 
        \nRightOut_45[2] , \nRightOut_45[1] , \nRightOut_45[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_62 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_44[16] , \nRightOut_44[15] , \nRightOut_44[14] , 
        \nRightOut_44[13] , \nRightOut_44[12] , \nRightOut_44[11] , 
        \nRightOut_44[10] , \nRightOut_44[9] , \nRightOut_44[8] , 
        \nRightOut_44[7] , \nRightOut_44[6] , \nRightOut_44[5] , 
        \nRightOut_44[4] , \nRightOut_44[3] , \nRightOut_44[2] , 
        \nRightOut_44[1] , \nRightOut_44[0] }), .inright({\nRightOut_46[16] , 
        \nRightOut_46[15] , \nRightOut_46[14] , \nRightOut_46[13] , 
        \nRightOut_46[12] , \nRightOut_46[11] , \nRightOut_46[10] , 
        \nRightOut_46[9] , \nRightOut_46[8] , \nRightOut_46[7] , 
        \nRightOut_46[6] , \nRightOut_46[5] , \nRightOut_46[4] , 
        \nRightOut_46[3] , \nRightOut_46[2] , \nRightOut_46[1] , 
        \nRightOut_46[0] }), .outleft({\nLeftOut_62[16] , \nLeftOut_62[15] , 
        \nLeftOut_62[14] , \nLeftOut_62[13] , \nLeftOut_62[12] , 
        \nLeftOut_62[11] , \nLeftOut_62[10] , \nLeftOut_62[9] , 
        \nLeftOut_62[8] , \nLeftOut_62[7] , \nLeftOut_62[6] , \nLeftOut_62[5] , 
        \nLeftOut_62[4] , \nLeftOut_62[3] , \nLeftOut_62[2] , \nLeftOut_62[1] , 
        \nLeftOut_62[0] }), .outright({\nRightOut_62[16] , \nRightOut_62[15] , 
        \nRightOut_62[14] , \nRightOut_62[13] , \nRightOut_62[12] , 
        \nRightOut_62[11] , \nRightOut_62[10] , \nRightOut_62[9] , 
        \nRightOut_62[8] , \nRightOut_62[7] , \nRightOut_62[6] , 
        \nRightOut_62[5] , \nRightOut_62[4] , \nRightOut_62[3] , 
        \nRightOut_62[2] , \nRightOut_62[1] , \nRightOut_62[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s7_SCAN1 node_87 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_71[16] , \nLeftOut_71[15] , \nLeftOut_71[14] , 
        \nLeftOut_71[13] , \nLeftOut_71[12] , \nLeftOut_71[11] , 
        \nLeftOut_71[10] , \nLeftOut_71[9] , \nLeftOut_71[8] , 
        \nLeftOut_71[7] , \nLeftOut_71[6] , \nLeftOut_71[5] , \nLeftOut_71[4] , 
        \nLeftOut_71[3] , \nLeftOut_71[2] , \nLeftOut_71[1] , \nLeftOut_71[0] 
        }), .inright({\nLeftOut_79[16] , \nLeftOut_79[15] , \nLeftOut_79[14] , 
        \nLeftOut_79[13] , \nLeftOut_79[12] , \nLeftOut_79[11] , 
        \nLeftOut_79[10] , \nLeftOut_79[9] , \nLeftOut_79[8] , 
        \nLeftOut_79[7] , \nLeftOut_79[6] , \nLeftOut_79[5] , \nLeftOut_79[4] , 
        \nLeftOut_79[3] , \nLeftOut_79[2] , \nLeftOut_79[1] , \nLeftOut_79[0] 
        }), .outleft({\nLeftOut_87[16] , \nLeftOut_87[15] , \nLeftOut_87[14] , 
        \nLeftOut_87[13] , \nLeftOut_87[12] , \nLeftOut_87[11] , 
        \nLeftOut_87[10] , \nLeftOut_87[9] , \nLeftOut_87[8] , 
        \nLeftOut_87[7] , \nLeftOut_87[6] , \nLeftOut_87[5] , \nLeftOut_87[4] , 
        \nLeftOut_87[3] , \nLeftOut_87[2] , \nLeftOut_87[1] , \nLeftOut_87[0] 
        }), .outright({\nRightOut_87[16] , \nRightOut_87[15] , 
        \nRightOut_87[14] , \nRightOut_87[13] , \nRightOut_87[12] , 
        \nRightOut_87[11] , \nRightOut_87[10] , \nRightOut_87[9] , 
        \nRightOut_87[8] , \nRightOut_87[7] , \nRightOut_87[6] , 
        \nRightOut_87[5] , \nRightOut_87[4] , \nRightOut_87[3] , 
        \nRightOut_87[2] , \nRightOut_87[1] , \nRightOut_87[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_107 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink27[15] , \ScanLink27[14] , \ScanLink27[13] , 
        \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , \ScanLink27[9] , 
        \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , \ScanLink27[5] , 
        \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , \ScanLink27[1] , 
        \ScanLink27[0] }), .ScanOut({\ScanLink28[15] , \ScanLink28[14] , 
        \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , 
        \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , 
        \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , 
        \ScanLink28[1] , \ScanLink28[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_86[16] , \nRightOut_86[15] , \nRightOut_86[14] , 
        \nRightOut_86[13] , \nRightOut_86[12] , \nRightOut_86[11] , 
        \nRightOut_86[10] , \nRightOut_86[9] , \nRightOut_86[8] , 
        \nRightOut_86[7] , \nRightOut_86[6] , \nRightOut_86[5] , 
        \nRightOut_86[4] , \nRightOut_86[3] , \nRightOut_86[2] , 
        \nRightOut_86[1] , \nRightOut_86[0] }), .inright({\nRightOut_87[16] , 
        \nRightOut_87[15] , \nRightOut_87[14] , \nRightOut_87[13] , 
        \nRightOut_87[12] , \nRightOut_87[11] , \nRightOut_87[10] , 
        \nRightOut_87[9] , \nRightOut_87[8] , \nRightOut_87[7] , 
        \nRightOut_87[6] , \nRightOut_87[5] , \nRightOut_87[4] , 
        \nRightOut_87[3] , \nRightOut_87[2] , \nRightOut_87[1] , 
        \nRightOut_87[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_38 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_22[16] , \nLeftOut_22[15] , \nLeftOut_22[14] , 
        \nLeftOut_22[13] , \nLeftOut_22[12] , \nLeftOut_22[11] , 
        \nLeftOut_22[10] , \nLeftOut_22[9] , \nLeftOut_22[8] , 
        \nLeftOut_22[7] , \nLeftOut_22[6] , \nLeftOut_22[5] , \nLeftOut_22[4] , 
        \nLeftOut_22[3] , \nLeftOut_22[2] , \nLeftOut_22[1] , \nLeftOut_22[0] 
        }), .inright({\nLeftOut_23[16] , \nLeftOut_23[15] , \nLeftOut_23[14] , 
        \nLeftOut_23[13] , \nLeftOut_23[12] , \nLeftOut_23[11] , 
        \nLeftOut_23[10] , \nLeftOut_23[9] , \nLeftOut_23[8] , 
        \nLeftOut_23[7] , \nLeftOut_23[6] , \nLeftOut_23[5] , \nLeftOut_23[4] , 
        \nLeftOut_23[3] , \nLeftOut_23[2] , \nLeftOut_23[1] , \nLeftOut_23[0] 
        }), .outleft({\nLeftOut_38[16] , \nLeftOut_38[15] , \nLeftOut_38[14] , 
        \nLeftOut_38[13] , \nLeftOut_38[12] , \nLeftOut_38[11] , 
        \nLeftOut_38[10] , \nLeftOut_38[9] , \nLeftOut_38[8] , 
        \nLeftOut_38[7] , \nLeftOut_38[6] , \nLeftOut_38[5] , \nLeftOut_38[4] , 
        \nLeftOut_38[3] , \nLeftOut_38[2] , \nLeftOut_38[1] , \nLeftOut_38[0] 
        }), .outright({\nRightOut_38[16] , \nRightOut_38[15] , 
        \nRightOut_38[14] , \nRightOut_38[13] , \nRightOut_38[12] , 
        \nRightOut_38[11] , \nRightOut_38[10] , \nRightOut_38[9] , 
        \nRightOut_38[8] , \nRightOut_38[7] , \nRightOut_38[6] , 
        \nRightOut_38[5] , \nRightOut_38[4] , \nRightOut_38[3] , 
        \nRightOut_38[2] , \nRightOut_38[1] , \nRightOut_38[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_44 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_28[16] , \nLeftOut_28[15] , \nLeftOut_28[14] , 
        \nLeftOut_28[13] , \nLeftOut_28[12] , \nLeftOut_28[11] , 
        \nLeftOut_28[10] , \nLeftOut_28[9] , \nLeftOut_28[8] , 
        \nLeftOut_28[7] , \nLeftOut_28[6] , \nLeftOut_28[5] , \nLeftOut_28[4] , 
        \nLeftOut_28[3] , \nLeftOut_28[2] , \nLeftOut_28[1] , \nLeftOut_28[0] 
        }), .inright({\nLeftOut_29[16] , \nLeftOut_29[15] , \nLeftOut_29[14] , 
        \nLeftOut_29[13] , \nLeftOut_29[12] , \nLeftOut_29[11] , 
        \nLeftOut_29[10] , \nLeftOut_29[9] , \nLeftOut_29[8] , 
        \nLeftOut_29[7] , \nLeftOut_29[6] , \nLeftOut_29[5] , \nLeftOut_29[4] , 
        \nLeftOut_29[3] , \nLeftOut_29[2] , \nLeftOut_29[1] , \nLeftOut_29[0] 
        }), .outleft({\nLeftOut_44[16] , \nLeftOut_44[15] , \nLeftOut_44[14] , 
        \nLeftOut_44[13] , \nLeftOut_44[12] , \nLeftOut_44[11] , 
        \nLeftOut_44[10] , \nLeftOut_44[9] , \nLeftOut_44[8] , 
        \nLeftOut_44[7] , \nLeftOut_44[6] , \nLeftOut_44[5] , \nLeftOut_44[4] , 
        \nLeftOut_44[3] , \nLeftOut_44[2] , \nLeftOut_44[1] , \nLeftOut_44[0] 
        }), .outright({\nRightOut_44[16] , \nRightOut_44[15] , 
        \nRightOut_44[14] , \nRightOut_44[13] , \nRightOut_44[12] , 
        \nRightOut_44[11] , \nRightOut_44[10] , \nRightOut_44[9] , 
        \nRightOut_44[8] , \nRightOut_44[7] , \nRightOut_44[6] , 
        \nRightOut_44[5] , \nRightOut_44[4] , \nRightOut_44[3] , 
        \nRightOut_44[2] , \nRightOut_44[1] , \nRightOut_44[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_56 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_40[16] , \nLeftOut_40[15] , \nLeftOut_40[14] , 
        \nLeftOut_40[13] , \nLeftOut_40[12] , \nLeftOut_40[11] , 
        \nLeftOut_40[10] , \nLeftOut_40[9] , \nLeftOut_40[8] , 
        \nLeftOut_40[7] , \nLeftOut_40[6] , \nLeftOut_40[5] , \nLeftOut_40[4] , 
        \nLeftOut_40[3] , \nLeftOut_40[2] , \nLeftOut_40[1] , \nLeftOut_40[0] 
        }), .inright({\nLeftOut_42[16] , \nLeftOut_42[15] , \nLeftOut_42[14] , 
        \nLeftOut_42[13] , \nLeftOut_42[12] , \nLeftOut_42[11] , 
        \nLeftOut_42[10] , \nLeftOut_42[9] , \nLeftOut_42[8] , 
        \nLeftOut_42[7] , \nLeftOut_42[6] , \nLeftOut_42[5] , \nLeftOut_42[4] , 
        \nLeftOut_42[3] , \nLeftOut_42[2] , \nLeftOut_42[1] , \nLeftOut_42[0] 
        }), .outleft({\nLeftOut_56[16] , \nLeftOut_56[15] , \nLeftOut_56[14] , 
        \nLeftOut_56[13] , \nLeftOut_56[12] , \nLeftOut_56[11] , 
        \nLeftOut_56[10] , \nLeftOut_56[9] , \nLeftOut_56[8] , 
        \nLeftOut_56[7] , \nLeftOut_56[6] , \nLeftOut_56[5] , \nLeftOut_56[4] , 
        \nLeftOut_56[3] , \nLeftOut_56[2] , \nLeftOut_56[1] , \nLeftOut_56[0] 
        }), .outright({\nRightOut_56[16] , \nRightOut_56[15] , 
        \nRightOut_56[14] , \nRightOut_56[13] , \nRightOut_56[12] , 
        \nRightOut_56[11] , \nRightOut_56[10] , \nRightOut_56[9] , 
        \nRightOut_56[8] , \nRightOut_56[7] , \nRightOut_56[6] , 
        \nRightOut_56[5] , \nRightOut_56[4] , \nRightOut_56[3] , 
        \nRightOut_56[2] , \nRightOut_56[1] , \nRightOut_56[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s14_SCAN1 node_71 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_51[16] , \nRightOut_51[15] , \nRightOut_51[14] , 
        \nRightOut_51[13] , \nRightOut_51[12] , \nRightOut_51[11] , 
        \nRightOut_51[10] , \nRightOut_51[9] , \nRightOut_51[8] , 
        \nRightOut_51[7] , \nRightOut_51[6] , \nRightOut_51[5] , 
        \nRightOut_51[4] , \nRightOut_51[3] , \nRightOut_51[2] , 
        \nRightOut_51[1] , \nRightOut_51[0] }), .inright({\nRightOut_55[16] , 
        \nRightOut_55[15] , \nRightOut_55[14] , \nRightOut_55[13] , 
        \nRightOut_55[12] , \nRightOut_55[11] , \nRightOut_55[10] , 
        \nRightOut_55[9] , \nRightOut_55[8] , \nRightOut_55[7] , 
        \nRightOut_55[6] , \nRightOut_55[5] , \nRightOut_55[4] , 
        \nRightOut_55[3] , \nRightOut_55[2] , \nRightOut_55[1] , 
        \nRightOut_55[0] }), .outleft({\nLeftOut_71[16] , \nLeftOut_71[15] , 
        \nLeftOut_71[14] , \nLeftOut_71[13] , \nLeftOut_71[12] , 
        \nLeftOut_71[11] , \nLeftOut_71[10] , \nLeftOut_71[9] , 
        \nLeftOut_71[8] , \nLeftOut_71[7] , \nLeftOut_71[6] , \nLeftOut_71[5] , 
        \nLeftOut_71[4] , \nLeftOut_71[3] , \nLeftOut_71[2] , \nLeftOut_71[1] , 
        \nLeftOut_71[0] }), .outright({\nRightOut_71[16] , \nRightOut_71[15] , 
        \nRightOut_71[14] , \nRightOut_71[13] , \nRightOut_71[12] , 
        \nRightOut_71[11] , \nRightOut_71[10] , \nRightOut_71[9] , 
        \nRightOut_71[8] , \nRightOut_71[7] , \nRightOut_71[6] , 
        \nRightOut_71[5] , \nRightOut_71[4] , \nRightOut_71[3] , 
        \nRightOut_71[2] , \nRightOut_71[1] , \nRightOut_71[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s14_SCAN1 node_94 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_70[16] , \nRightOut_70[15] , \nRightOut_70[14] , 
        \nRightOut_70[13] , \nRightOut_70[12] , \nRightOut_70[11] , 
        \nRightOut_70[10] , \nRightOut_70[9] , \nRightOut_70[8] , 
        \nRightOut_70[7] , \nRightOut_70[6] , \nRightOut_70[5] , 
        \nRightOut_70[4] , \nRightOut_70[3] , \nRightOut_70[2] , 
        \nRightOut_70[1] , \nRightOut_70[0] }), .inright({\nRightOut_78[16] , 
        \nRightOut_78[15] , \nRightOut_78[14] , \nRightOut_78[13] , 
        \nRightOut_78[12] , \nRightOut_78[11] , \nRightOut_78[10] , 
        \nRightOut_78[9] , \nRightOut_78[8] , \nRightOut_78[7] , 
        \nRightOut_78[6] , \nRightOut_78[5] , \nRightOut_78[4] , 
        \nRightOut_78[3] , \nRightOut_78[2] , \nRightOut_78[1] , 
        \nRightOut_78[0] }), .outleft({\nLeftOut_94[16] , \nLeftOut_94[15] , 
        \nLeftOut_94[14] , \nLeftOut_94[13] , \nLeftOut_94[12] , 
        \nLeftOut_94[11] , \nLeftOut_94[10] , \nLeftOut_94[9] , 
        \nLeftOut_94[8] , \nLeftOut_94[7] , \nLeftOut_94[6] , \nLeftOut_94[5] , 
        \nLeftOut_94[4] , \nLeftOut_94[3] , \nLeftOut_94[2] , \nLeftOut_94[1] , 
        \nLeftOut_94[0] }), .outright({\nRightOut_94[16] , \nRightOut_94[15] , 
        \nRightOut_94[14] , \nRightOut_94[13] , \nRightOut_94[12] , 
        \nRightOut_94[11] , \nRightOut_94[10] , \nRightOut_94[9] , 
        \nRightOut_94[8] , \nRightOut_94[7] , \nRightOut_94[6] , 
        \nRightOut_94[5] , \nRightOut_94[4] , \nRightOut_94[3] , 
        \nRightOut_94[2] , \nRightOut_94[1] , \nRightOut_94[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s12_SCAN1 node_63 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_45[16] , \nRightOut_45[15] , \nRightOut_45[14] , 
        \nRightOut_45[13] , \nRightOut_45[12] , \nRightOut_45[11] , 
        \nRightOut_45[10] , \nRightOut_45[9] , \nRightOut_45[8] , 
        \nRightOut_45[7] , \nRightOut_45[6] , \nRightOut_45[5] , 
        \nRightOut_45[4] , \nRightOut_45[3] , \nRightOut_45[2] , 
        \nRightOut_45[1] , \nRightOut_45[0] }), .inright({\nRightOut_47[16] , 
        \nRightOut_47[15] , \nRightOut_47[14] , \nRightOut_47[13] , 
        \nRightOut_47[12] , \nRightOut_47[11] , \nRightOut_47[10] , 
        \nRightOut_47[9] , \nRightOut_47[8] , \nRightOut_47[7] , 
        \nRightOut_47[6] , \nRightOut_47[5] , \nRightOut_47[4] , 
        \nRightOut_47[3] , \nRightOut_47[2] , \nRightOut_47[1] , 
        \nRightOut_47[0] }), .outleft({\nLeftOut_63[16] , \nLeftOut_63[15] , 
        \nLeftOut_63[14] , \nLeftOut_63[13] , \nLeftOut_63[12] , 
        \nLeftOut_63[11] , \nLeftOut_63[10] , \nLeftOut_63[9] , 
        \nLeftOut_63[8] , \nLeftOut_63[7] , \nLeftOut_63[6] , \nLeftOut_63[5] , 
        \nLeftOut_63[4] , \nLeftOut_63[3] , \nLeftOut_63[2] , \nLeftOut_63[1] , 
        \nLeftOut_63[0] }), .outright({\nRightOut_63[16] , \nRightOut_63[15] , 
        \nRightOut_63[14] , \nRightOut_63[13] , \nRightOut_63[12] , 
        \nRightOut_63[11] , \nRightOut_63[10] , \nRightOut_63[9] , 
        \nRightOut_63[8] , \nRightOut_63[7] , \nRightOut_63[6] , 
        \nRightOut_63[5] , \nRightOut_63[4] , \nRightOut_63[3] , 
        \nRightOut_63[2] , \nRightOut_63[1] , \nRightOut_63[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s6_SCAN1 node_86 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_70[16] , \nLeftOut_70[15] , \nLeftOut_70[14] , 
        \nLeftOut_70[13] , \nLeftOut_70[12] , \nLeftOut_70[11] , 
        \nLeftOut_70[10] , \nLeftOut_70[9] , \nLeftOut_70[8] , 
        \nLeftOut_70[7] , \nLeftOut_70[6] , \nLeftOut_70[5] , \nLeftOut_70[4] , 
        \nLeftOut_70[3] , \nLeftOut_70[2] , \nLeftOut_70[1] , \nLeftOut_70[0] 
        }), .inright({\nLeftOut_78[16] , \nLeftOut_78[15] , \nLeftOut_78[14] , 
        \nLeftOut_78[13] , \nLeftOut_78[12] , \nLeftOut_78[11] , 
        \nLeftOut_78[10] , \nLeftOut_78[9] , \nLeftOut_78[8] , 
        \nLeftOut_78[7] , \nLeftOut_78[6] , \nLeftOut_78[5] , \nLeftOut_78[4] , 
        \nLeftOut_78[3] , \nLeftOut_78[2] , \nLeftOut_78[1] , \nLeftOut_78[0] 
        }), .outleft({\nLeftOut_86[16] , \nLeftOut_86[15] , \nLeftOut_86[14] , 
        \nLeftOut_86[13] , \nLeftOut_86[12] , \nLeftOut_86[11] , 
        \nLeftOut_86[10] , \nLeftOut_86[9] , \nLeftOut_86[8] , 
        \nLeftOut_86[7] , \nLeftOut_86[6] , \nLeftOut_86[5] , \nLeftOut_86[4] , 
        \nLeftOut_86[3] , \nLeftOut_86[2] , \nLeftOut_86[1] , \nLeftOut_86[0] 
        }), .outright({\nRightOut_86[16] , \nRightOut_86[15] , 
        \nRightOut_86[14] , \nRightOut_86[13] , \nRightOut_86[12] , 
        \nRightOut_86[11] , \nRightOut_86[10] , \nRightOut_86[9] , 
        \nRightOut_86[8] , \nRightOut_86[7] , \nRightOut_86[6] , 
        \nRightOut_86[5] , \nRightOut_86[4] , \nRightOut_86[3] , 
        \nRightOut_86[2] , \nRightOut_86[1] , \nRightOut_86[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_106 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink26[15] , \ScanLink26[14] , \ScanLink26[13] , 
        \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , \ScanLink26[9] , 
        \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , \ScanLink26[5] , 
        \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , \ScanLink26[1] , 
        \ScanLink26[0] }), .ScanOut({\ScanLink27[15] , \ScanLink27[14] , 
        \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , 
        \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , 
        \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , 
        \ScanLink27[1] , \ScanLink27[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_84[16] , \nRightOut_84[15] , \nRightOut_84[14] , 
        \nRightOut_84[13] , \nRightOut_84[12] , \nRightOut_84[11] , 
        \nRightOut_84[10] , \nRightOut_84[9] , \nRightOut_84[8] , 
        \nRightOut_84[7] , \nRightOut_84[6] , \nRightOut_84[5] , 
        \nRightOut_84[4] , \nRightOut_84[3] , \nRightOut_84[2] , 
        \nRightOut_84[1] , \nRightOut_84[0] }), .inright({\nRightOut_85[16] , 
        \nRightOut_85[15] , \nRightOut_85[14] , \nRightOut_85[13] , 
        \nRightOut_85[12] , \nRightOut_85[11] , \nRightOut_85[10] , 
        \nRightOut_85[9] , \nRightOut_85[8] , \nRightOut_85[7] , 
        \nRightOut_85[6] , \nRightOut_85[5] , \nRightOut_85[4] , 
        \nRightOut_85[3] , \nRightOut_85[2] , \nRightOut_85[1] , 
        \nRightOut_85[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_31 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_15[16] , \nLeftOut_15[15] , \nLeftOut_15[14] , 
        \nLeftOut_15[13] , \nLeftOut_15[12] , \nLeftOut_15[11] , 
        \nLeftOut_15[10] , \nLeftOut_15[9] , \nLeftOut_15[8] , 
        \nLeftOut_15[7] , \nLeftOut_15[6] , \nLeftOut_15[5] , \nLeftOut_15[4] , 
        \nLeftOut_15[3] , \nLeftOut_15[2] , \nLeftOut_15[1] , \nLeftOut_15[0] 
        }), .inright({\nRightOut_15[16] , \nRightOut_15[15] , 
        \nRightOut_15[14] , \nRightOut_15[13] , \nRightOut_15[12] , 
        \nRightOut_15[11] , \nRightOut_15[10] , \nRightOut_15[9] , 
        \nRightOut_15[8] , \nRightOut_15[7] , \nRightOut_15[6] , 
        \nRightOut_15[5] , \nRightOut_15[4] , \nRightOut_15[3] , 
        \nRightOut_15[2] , \nRightOut_15[1] , \nRightOut_15[0] }), .outleft({
        \nLeftOut_31[16] , \nLeftOut_31[15] , \nLeftOut_31[14] , 
        \nLeftOut_31[13] , \nLeftOut_31[12] , \nLeftOut_31[11] , 
        \nLeftOut_31[10] , \nLeftOut_31[9] , \nLeftOut_31[8] , 
        \nLeftOut_31[7] , \nLeftOut_31[6] , \nLeftOut_31[5] , \nLeftOut_31[4] , 
        \nLeftOut_31[3] , \nLeftOut_31[2] , \nLeftOut_31[1] , \nLeftOut_31[0] 
        }), .outright({\nRightOut_31[16] , \nRightOut_31[15] , 
        \nRightOut_31[14] , \nRightOut_31[13] , \nRightOut_31[12] , 
        \nRightOut_31[11] , \nRightOut_31[10] , \nRightOut_31[9] , 
        \nRightOut_31[8] , \nRightOut_31[7] , \nRightOut_31[6] , 
        \nRightOut_31[5] , \nRightOut_31[4] , \nRightOut_31[3] , 
        \nRightOut_31[2] , \nRightOut_31[1] , \nRightOut_31[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s12_SCAN1 node_78 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_58[16] , \nRightOut_58[15] , \nRightOut_58[14] , 
        \nRightOut_58[13] , \nRightOut_58[12] , \nRightOut_58[11] , 
        \nRightOut_58[10] , \nRightOut_58[9] , \nRightOut_58[8] , 
        \nRightOut_58[7] , \nRightOut_58[6] , \nRightOut_58[5] , 
        \nRightOut_58[4] , \nRightOut_58[3] , \nRightOut_58[2] , 
        \nRightOut_58[1] , \nRightOut_58[0] }), .inright({\nRightOut_62[16] , 
        \nRightOut_62[15] , \nRightOut_62[14] , \nRightOut_62[13] , 
        \nRightOut_62[12] , \nRightOut_62[11] , \nRightOut_62[10] , 
        \nRightOut_62[9] , \nRightOut_62[8] , \nRightOut_62[7] , 
        \nRightOut_62[6] , \nRightOut_62[5] , \nRightOut_62[4] , 
        \nRightOut_62[3] , \nRightOut_62[2] , \nRightOut_62[1] , 
        \nRightOut_62[0] }), .outleft({\nLeftOut_78[16] , \nLeftOut_78[15] , 
        \nLeftOut_78[14] , \nLeftOut_78[13] , \nLeftOut_78[12] , 
        \nLeftOut_78[11] , \nLeftOut_78[10] , \nLeftOut_78[9] , 
        \nLeftOut_78[8] , \nLeftOut_78[7] , \nLeftOut_78[6] , \nLeftOut_78[5] , 
        \nLeftOut_78[4] , \nLeftOut_78[3] , \nLeftOut_78[2] , \nLeftOut_78[1] , 
        \nLeftOut_78[0] }), .outright({\nRightOut_78[16] , \nRightOut_78[15] , 
        \nRightOut_78[14] , \nRightOut_78[13] , \nRightOut_78[12] , 
        \nRightOut_78[11] , \nRightOut_78[10] , \nRightOut_78[9] , 
        \nRightOut_78[8] , \nRightOut_78[7] , \nRightOut_78[6] , 
        \nRightOut_78[5] , \nRightOut_78[4] , \nRightOut_78[3] , 
        \nRightOut_78[2] , \nRightOut_78[1] , \nRightOut_78[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink5[15] , \ScanLink5[14] , \ScanLink5[13] , 
        \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , \ScanLink5[9] , 
        \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , \ScanLink5[5] , 
        \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , \ScanLink5[1] , 
        \ScanLink5[0] }), .ScanOut({\ScanLink6[15] , \ScanLink6[14] , 
        \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , 
        \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_5[16] , \nLeftOut_5[15] , \nLeftOut_5[14] , \nLeftOut_5[13] , 
        \nLeftOut_5[12] , \nLeftOut_5[11] , \nLeftOut_5[10] , \nLeftOut_5[9] , 
        \nLeftOut_5[8] , \nLeftOut_5[7] , \nLeftOut_5[6] , \nLeftOut_5[5] , 
        \nLeftOut_5[4] , \nLeftOut_5[3] , \nLeftOut_5[2] , \nLeftOut_5[1] , 
        \nLeftOut_5[0] }), .inright({\nRightOut_5[16] , \nRightOut_5[15] , 
        \nRightOut_5[14] , \nRightOut_5[13] , \nRightOut_5[12] , 
        \nRightOut_5[11] , \nRightOut_5[10] , \nRightOut_5[9] , 
        \nRightOut_5[8] , \nRightOut_5[7] , \nRightOut_5[6] , \nRightOut_5[5] , 
        \nRightOut_5[4] , \nRightOut_5[3] , \nRightOut_5[2] , \nRightOut_5[1] , 
        \nRightOut_5[0] }), .outleft({\nLeftOut_5[16] , \nLeftOut_5[15] , 
        \nLeftOut_5[14] , \nLeftOut_5[13] , \nLeftOut_5[12] , \nLeftOut_5[11] , 
        \nLeftOut_5[10] , \nLeftOut_5[9] , \nLeftOut_5[8] , \nLeftOut_5[7] , 
        \nLeftOut_5[6] , \nLeftOut_5[5] , \nLeftOut_5[4] , \nLeftOut_5[3] , 
        \nLeftOut_5[2] , \nLeftOut_5[1] , \nLeftOut_5[0] }), .outright({
        \nRightOut_5[16] , \nRightOut_5[15] , \nRightOut_5[14] , 
        \nRightOut_5[13] , \nRightOut_5[12] , \nRightOut_5[11] , 
        \nRightOut_5[10] , \nRightOut_5[9] , \nRightOut_5[8] , 
        \nRightOut_5[7] , \nRightOut_5[6] , \nRightOut_5[5] , \nRightOut_5[4] , 
        \nRightOut_5[3] , \nRightOut_5[2] , \nRightOut_5[1] , \nRightOut_5[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink7[15] , \ScanLink7[14] , \ScanLink7[13] , 
        \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , \ScanLink7[9] , 
        \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , \ScanLink7[5] , 
        \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , \ScanLink7[1] , 
        \ScanLink7[0] }), .ScanOut({\ScanLink8[15] , \ScanLink8[14] , 
        \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , 
        \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_7[16] , \nLeftOut_7[15] , \nLeftOut_7[14] , \nLeftOut_7[13] , 
        \nLeftOut_7[12] , \nLeftOut_7[11] , \nLeftOut_7[10] , \nLeftOut_7[9] , 
        \nLeftOut_7[8] , \nLeftOut_7[7] , \nLeftOut_7[6] , \nLeftOut_7[5] , 
        \nLeftOut_7[4] , \nLeftOut_7[3] , \nLeftOut_7[2] , \nLeftOut_7[1] , 
        \nLeftOut_7[0] }), .inright({\nRightOut_7[16] , \nRightOut_7[15] , 
        \nRightOut_7[14] , \nRightOut_7[13] , \nRightOut_7[12] , 
        \nRightOut_7[11] , \nRightOut_7[10] , \nRightOut_7[9] , 
        \nRightOut_7[8] , \nRightOut_7[7] , \nRightOut_7[6] , \nRightOut_7[5] , 
        \nRightOut_7[4] , \nRightOut_7[3] , \nRightOut_7[2] , \nRightOut_7[1] , 
        \nRightOut_7[0] }), .outleft({\nLeftOut_7[16] , \nLeftOut_7[15] , 
        \nLeftOut_7[14] , \nLeftOut_7[13] , \nLeftOut_7[12] , \nLeftOut_7[11] , 
        \nLeftOut_7[10] , \nLeftOut_7[9] , \nLeftOut_7[8] , \nLeftOut_7[7] , 
        \nLeftOut_7[6] , \nLeftOut_7[5] , \nLeftOut_7[4] , \nLeftOut_7[3] , 
        \nLeftOut_7[2] , \nLeftOut_7[1] , \nLeftOut_7[0] }), .outright({
        \nRightOut_7[16] , \nRightOut_7[15] , \nRightOut_7[14] , 
        \nRightOut_7[13] , \nRightOut_7[12] , \nRightOut_7[11] , 
        \nRightOut_7[10] , \nRightOut_7[9] , \nRightOut_7[8] , 
        \nRightOut_7[7] , \nRightOut_7[6] , \nRightOut_7[5] , \nRightOut_7[4] , 
        \nRightOut_7[3] , \nRightOut_7[2] , \nRightOut_7[1] , \nRightOut_7[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_11 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink11[15] , \ScanLink11[14] , \ScanLink11[13] , 
        \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , \ScanLink11[9] , 
        \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , \ScanLink11[5] , 
        \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , \ScanLink11[1] , 
        \ScanLink11[0] }), .ScanOut({\ScanLink12[15] , \ScanLink12[14] , 
        \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , 
        \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , 
        \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , 
        \ScanLink12[1] , \ScanLink12[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_11[16] , \nLeftOut_11[15] , \nLeftOut_11[14] , 
        \nLeftOut_11[13] , \nLeftOut_11[12] , \nLeftOut_11[11] , 
        \nLeftOut_11[10] , \nLeftOut_11[9] , \nLeftOut_11[8] , 
        \nLeftOut_11[7] , \nLeftOut_11[6] , \nLeftOut_11[5] , \nLeftOut_11[4] , 
        \nLeftOut_11[3] , \nLeftOut_11[2] , \nLeftOut_11[1] , \nLeftOut_11[0] 
        }), .inright({\nRightOut_11[16] , \nRightOut_11[15] , 
        \nRightOut_11[14] , \nRightOut_11[13] , \nRightOut_11[12] , 
        \nRightOut_11[11] , \nRightOut_11[10] , \nRightOut_11[9] , 
        \nRightOut_11[8] , \nRightOut_11[7] , \nRightOut_11[6] , 
        \nRightOut_11[5] , \nRightOut_11[4] , \nRightOut_11[3] , 
        \nRightOut_11[2] , \nRightOut_11[1] , \nRightOut_11[0] }), .outleft({
        \nLeftOut_11[16] , \nLeftOut_11[15] , \nLeftOut_11[14] , 
        \nLeftOut_11[13] , \nLeftOut_11[12] , \nLeftOut_11[11] , 
        \nLeftOut_11[10] , \nLeftOut_11[9] , \nLeftOut_11[8] , 
        \nLeftOut_11[7] , \nLeftOut_11[6] , \nLeftOut_11[5] , \nLeftOut_11[4] , 
        \nLeftOut_11[3] , \nLeftOut_11[2] , \nLeftOut_11[1] , \nLeftOut_11[0] 
        }), .outright({\nRightOut_11[16] , \nRightOut_11[15] , 
        \nRightOut_11[14] , \nRightOut_11[13] , \nRightOut_11[12] , 
        \nRightOut_11[11] , \nRightOut_11[10] , \nRightOut_11[9] , 
        \nRightOut_11[8] , \nRightOut_11[7] , \nRightOut_11[6] , 
        \nRightOut_11[5] , \nRightOut_11[4] , \nRightOut_11[3] , 
        \nRightOut_11[2] , \nRightOut_11[1] , \nRightOut_11[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_36 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_20[16] , \nLeftOut_20[15] , \nLeftOut_20[14] , 
        \nLeftOut_20[13] , \nLeftOut_20[12] , \nLeftOut_20[11] , 
        \nLeftOut_20[10] , \nLeftOut_20[9] , \nLeftOut_20[8] , 
        \nLeftOut_20[7] , \nLeftOut_20[6] , \nLeftOut_20[5] , \nLeftOut_20[4] , 
        \nLeftOut_20[3] , \nLeftOut_20[2] , \nLeftOut_20[1] , \nLeftOut_20[0] 
        }), .inright({\nLeftOut_21[16] , \nLeftOut_21[15] , \nLeftOut_21[14] , 
        \nLeftOut_21[13] , \nLeftOut_21[12] , \nLeftOut_21[11] , 
        \nLeftOut_21[10] , \nLeftOut_21[9] , \nLeftOut_21[8] , 
        \nLeftOut_21[7] , \nLeftOut_21[6] , \nLeftOut_21[5] , \nLeftOut_21[4] , 
        \nLeftOut_21[3] , \nLeftOut_21[2] , \nLeftOut_21[1] , \nLeftOut_21[0] 
        }), .outleft({\nLeftOut_36[16] , \nLeftOut_36[15] , \nLeftOut_36[14] , 
        \nLeftOut_36[13] , \nLeftOut_36[12] , \nLeftOut_36[11] , 
        \nLeftOut_36[10] , \nLeftOut_36[9] , \nLeftOut_36[8] , 
        \nLeftOut_36[7] , \nLeftOut_36[6] , \nLeftOut_36[5] , \nLeftOut_36[4] , 
        \nLeftOut_36[3] , \nLeftOut_36[2] , \nLeftOut_36[1] , \nLeftOut_36[0] 
        }), .outright({\nRightOut_36[16] , \nRightOut_36[15] , 
        \nRightOut_36[14] , \nRightOut_36[13] , \nRightOut_36[12] , 
        \nRightOut_36[11] , \nRightOut_36[10] , \nRightOut_36[9] , 
        \nRightOut_36[8] , \nRightOut_36[7] , \nRightOut_36[6] , 
        \nRightOut_36[5] , \nRightOut_36[4] , \nRightOut_36[3] , 
        \nRightOut_36[2] , \nRightOut_36[1] , \nRightOut_36[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_58 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_40[16] , \nRightOut_40[15] , \nRightOut_40[14] , 
        \nRightOut_40[13] , \nRightOut_40[12] , \nRightOut_40[11] , 
        \nRightOut_40[10] , \nRightOut_40[9] , \nRightOut_40[8] , 
        \nRightOut_40[7] , \nRightOut_40[6] , \nRightOut_40[5] , 
        \nRightOut_40[4] , \nRightOut_40[3] , \nRightOut_40[2] , 
        \nRightOut_40[1] , \nRightOut_40[0] }), .inright({\nRightOut_42[16] , 
        \nRightOut_42[15] , \nRightOut_42[14] , \nRightOut_42[13] , 
        \nRightOut_42[12] , \nRightOut_42[11] , \nRightOut_42[10] , 
        \nRightOut_42[9] , \nRightOut_42[8] , \nRightOut_42[7] , 
        \nRightOut_42[6] , \nRightOut_42[5] , \nRightOut_42[4] , 
        \nRightOut_42[3] , \nRightOut_42[2] , \nRightOut_42[1] , 
        \nRightOut_42[0] }), .outleft({\nLeftOut_58[16] , \nLeftOut_58[15] , 
        \nLeftOut_58[14] , \nLeftOut_58[13] , \nLeftOut_58[12] , 
        \nLeftOut_58[11] , \nLeftOut_58[10] , \nLeftOut_58[9] , 
        \nLeftOut_58[8] , \nLeftOut_58[7] , \nLeftOut_58[6] , \nLeftOut_58[5] , 
        \nLeftOut_58[4] , \nLeftOut_58[3] , \nLeftOut_58[2] , \nLeftOut_58[1] , 
        \nLeftOut_58[0] }), .outright({\nRightOut_58[16] , \nRightOut_58[15] , 
        \nRightOut_58[14] , \nRightOut_58[13] , \nRightOut_58[12] , 
        \nRightOut_58[11] , \nRightOut_58[10] , \nRightOut_58[9] , 
        \nRightOut_58[8] , \nRightOut_58[7] , \nRightOut_58[6] , 
        \nRightOut_58[5] , \nRightOut_58[4] , \nRightOut_58[3] , 
        \nRightOut_58[2] , \nRightOut_58[1] , \nRightOut_58[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_13 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink13[15] , \ScanLink13[14] , \ScanLink13[13] , 
        \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , \ScanLink13[9] , 
        \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , \ScanLink13[5] , 
        \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , \ScanLink13[1] , 
        \ScanLink13[0] }), .ScanOut({\ScanLink14[15] , \ScanLink14[14] , 
        \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , 
        \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , 
        \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , 
        \ScanLink14[1] , \ScanLink14[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_13[16] , \nLeftOut_13[15] , \nLeftOut_13[14] , 
        \nLeftOut_13[13] , \nLeftOut_13[12] , \nLeftOut_13[11] , 
        \nLeftOut_13[10] , \nLeftOut_13[9] , \nLeftOut_13[8] , 
        \nLeftOut_13[7] , \nLeftOut_13[6] , \nLeftOut_13[5] , \nLeftOut_13[4] , 
        \nLeftOut_13[3] , \nLeftOut_13[2] , \nLeftOut_13[1] , \nLeftOut_13[0] 
        }), .inright({\nRightOut_13[16] , \nRightOut_13[15] , 
        \nRightOut_13[14] , \nRightOut_13[13] , \nRightOut_13[12] , 
        \nRightOut_13[11] , \nRightOut_13[10] , \nRightOut_13[9] , 
        \nRightOut_13[8] , \nRightOut_13[7] , \nRightOut_13[6] , 
        \nRightOut_13[5] , \nRightOut_13[4] , \nRightOut_13[3] , 
        \nRightOut_13[2] , \nRightOut_13[1] , \nRightOut_13[0] }), .outleft({
        \nLeftOut_13[16] , \nLeftOut_13[15] , \nLeftOut_13[14] , 
        \nLeftOut_13[13] , \nLeftOut_13[12] , \nLeftOut_13[11] , 
        \nLeftOut_13[10] , \nLeftOut_13[9] , \nLeftOut_13[8] , 
        \nLeftOut_13[7] , \nLeftOut_13[6] , \nLeftOut_13[5] , \nLeftOut_13[4] , 
        \nLeftOut_13[3] , \nLeftOut_13[2] , \nLeftOut_13[1] , \nLeftOut_13[0] 
        }), .outright({\nRightOut_13[16] , \nRightOut_13[15] , 
        \nRightOut_13[14] , \nRightOut_13[13] , \nRightOut_13[12] , 
        \nRightOut_13[11] , \nRightOut_13[10] , \nRightOut_13[9] , 
        \nRightOut_13[8] , \nRightOut_13[7] , \nRightOut_13[6] , 
        \nRightOut_13[5] , \nRightOut_13[4] , \nRightOut_13[3] , 
        \nRightOut_13[2] , \nRightOut_13[1] , \nRightOut_13[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_18 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_2[16] , \nLeftOut_2[15] , \nLeftOut_2[14] , \nLeftOut_2[13] , 
        \nLeftOut_2[12] , \nLeftOut_2[11] , \nLeftOut_2[10] , \nLeftOut_2[9] , 
        \nLeftOut_2[8] , \nLeftOut_2[7] , \nLeftOut_2[6] , \nLeftOut_2[5] , 
        \nLeftOut_2[4] , \nLeftOut_2[3] , \nLeftOut_2[2] , \nLeftOut_2[1] , 
        \nLeftOut_2[0] }), .inright({\nRightOut_2[16] , \nRightOut_2[15] , 
        \nRightOut_2[14] , \nRightOut_2[13] , \nRightOut_2[12] , 
        \nRightOut_2[11] , \nRightOut_2[10] , \nRightOut_2[9] , 
        \nRightOut_2[8] , \nRightOut_2[7] , \nRightOut_2[6] , \nRightOut_2[5] , 
        \nRightOut_2[4] , \nRightOut_2[3] , \nRightOut_2[2] , \nRightOut_2[1] , 
        \nRightOut_2[0] }), .outleft({\nLeftOut_18[16] , \nLeftOut_18[15] , 
        \nLeftOut_18[14] , \nLeftOut_18[13] , \nLeftOut_18[12] , 
        \nLeftOut_18[11] , \nLeftOut_18[10] , \nLeftOut_18[9] , 
        \nLeftOut_18[8] , \nLeftOut_18[7] , \nLeftOut_18[6] , \nLeftOut_18[5] , 
        \nLeftOut_18[4] , \nLeftOut_18[3] , \nLeftOut_18[2] , \nLeftOut_18[1] , 
        \nLeftOut_18[0] }), .outright({\nRightOut_18[16] , \nRightOut_18[15] , 
        \nRightOut_18[14] , \nRightOut_18[13] , \nRightOut_18[12] , 
        \nRightOut_18[11] , \nRightOut_18[10] , \nRightOut_18[9] , 
        \nRightOut_18[8] , \nRightOut_18[7] , \nRightOut_18[6] , 
        \nRightOut_18[5] , \nRightOut_18[4] , \nRightOut_18[3] , 
        \nRightOut_18[2] , \nRightOut_18[1] , \nRightOut_18[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_43 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_26[16] , \nRightOut_26[15] , \nRightOut_26[14] , 
        \nRightOut_26[13] , \nRightOut_26[12] , \nRightOut_26[11] , 
        \nRightOut_26[10] , \nRightOut_26[9] , \nRightOut_26[8] , 
        \nRightOut_26[7] , \nRightOut_26[6] , \nRightOut_26[5] , 
        \nRightOut_26[4] , \nRightOut_26[3] , \nRightOut_26[2] , 
        \nRightOut_26[1] , \nRightOut_26[0] }), .inright({\nRightOut_27[16] , 
        \nRightOut_27[15] , \nRightOut_27[14] , \nRightOut_27[13] , 
        \nRightOut_27[12] , \nRightOut_27[11] , \nRightOut_27[10] , 
        \nRightOut_27[9] , \nRightOut_27[8] , \nRightOut_27[7] , 
        \nRightOut_27[6] , \nRightOut_27[5] , \nRightOut_27[4] , 
        \nRightOut_27[3] , \nRightOut_27[2] , \nRightOut_27[1] , 
        \nRightOut_27[0] }), .outleft({\nLeftOut_43[16] , \nLeftOut_43[15] , 
        \nLeftOut_43[14] , \nLeftOut_43[13] , \nLeftOut_43[12] , 
        \nLeftOut_43[11] , \nLeftOut_43[10] , \nLeftOut_43[9] , 
        \nLeftOut_43[8] , \nLeftOut_43[7] , \nLeftOut_43[6] , \nLeftOut_43[5] , 
        \nLeftOut_43[4] , \nLeftOut_43[3] , \nLeftOut_43[2] , \nLeftOut_43[1] , 
        \nLeftOut_43[0] }), .outright({\nRightOut_43[16] , \nRightOut_43[15] , 
        \nRightOut_43[14] , \nRightOut_43[13] , \nRightOut_43[12] , 
        \nRightOut_43[11] , \nRightOut_43[10] , \nRightOut_43[9] , 
        \nRightOut_43[8] , \nRightOut_43[7] , \nRightOut_43[6] , 
        \nRightOut_43[5] , \nRightOut_43[4] , \nRightOut_43[3] , 
        \nRightOut_43[2] , \nRightOut_43[1] , \nRightOut_43[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s1_SCAN1 node_81 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_65[16] , \nLeftOut_65[15] , \nLeftOut_65[14] , 
        \nLeftOut_65[13] , \nLeftOut_65[12] , \nLeftOut_65[11] , 
        \nLeftOut_65[10] , \nLeftOut_65[9] , \nLeftOut_65[8] , 
        \nLeftOut_65[7] , \nLeftOut_65[6] , \nLeftOut_65[5] , \nLeftOut_65[4] , 
        \nLeftOut_65[3] , \nLeftOut_65[2] , \nLeftOut_65[1] , \nLeftOut_65[0] 
        }), .inright({\nLeftOut_73[16] , \nLeftOut_73[15] , \nLeftOut_73[14] , 
        \nLeftOut_73[13] , \nLeftOut_73[12] , \nLeftOut_73[11] , 
        \nLeftOut_73[10] , \nLeftOut_73[9] , \nLeftOut_73[8] , 
        \nLeftOut_73[7] , \nLeftOut_73[6] , \nLeftOut_73[5] , \nLeftOut_73[4] , 
        \nLeftOut_73[3] , \nLeftOut_73[2] , \nLeftOut_73[1] , \nLeftOut_73[0] 
        }), .outleft({\nLeftOut_81[16] , \nLeftOut_81[15] , \nLeftOut_81[14] , 
        \nLeftOut_81[13] , \nLeftOut_81[12] , \nLeftOut_81[11] , 
        \nLeftOut_81[10] , \nLeftOut_81[9] , \nLeftOut_81[8] , 
        \nLeftOut_81[7] , \nLeftOut_81[6] , \nLeftOut_81[5] , \nLeftOut_81[4] , 
        \nLeftOut_81[3] , \nLeftOut_81[2] , \nLeftOut_81[1] , \nLeftOut_81[0] 
        }), .outright({\nRightOut_81[16] , \nRightOut_81[15] , 
        \nRightOut_81[14] , \nRightOut_81[13] , \nRightOut_81[12] , 
        \nRightOut_81[11] , \nRightOut_81[10] , \nRightOut_81[9] , 
        \nRightOut_81[8] , \nRightOut_81[7] , \nRightOut_81[6] , 
        \nRightOut_81[5] , \nRightOut_81[4] , \nRightOut_81[3] , 
        \nRightOut_81[2] , \nRightOut_81[1] , \nRightOut_81[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_101 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink21[15] , \ScanLink21[14] , \ScanLink21[13] , 
        \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , \ScanLink21[9] , 
        \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , \ScanLink21[5] , 
        \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , \ScanLink21[1] , 
        \ScanLink21[0] }), .ScanOut({\ScanLink22[15] , \ScanLink22[14] , 
        \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , 
        \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , 
        \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , 
        \ScanLink22[1] , \ScanLink22[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_90[16] , \nLeftOut_90[15] , \nLeftOut_90[14] , 
        \nLeftOut_90[13] , \nLeftOut_90[12] , \nLeftOut_90[11] , 
        \nLeftOut_90[10] , \nLeftOut_90[9] , \nLeftOut_90[8] , 
        \nLeftOut_90[7] , \nLeftOut_90[6] , \nLeftOut_90[5] , \nLeftOut_90[4] , 
        \nLeftOut_90[3] , \nLeftOut_90[2] , \nLeftOut_90[1] , \nLeftOut_90[0] 
        }), .inright({\nLeftOut_91[16] , \nLeftOut_91[15] , \nLeftOut_91[14] , 
        \nLeftOut_91[13] , \nLeftOut_91[12] , \nLeftOut_91[11] , 
        \nLeftOut_91[10] , \nLeftOut_91[9] , \nLeftOut_91[8] , 
        \nLeftOut_91[7] , \nLeftOut_91[6] , \nLeftOut_91[5] , \nLeftOut_91[4] , 
        \nLeftOut_91[3] , \nLeftOut_91[2] , \nLeftOut_91[1] , \nLeftOut_91[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s12_SCAN1 node_51 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_33[16] , \nRightOut_33[15] , \nRightOut_33[14] , 
        \nRightOut_33[13] , \nRightOut_33[12] , \nRightOut_33[11] , 
        \nRightOut_33[10] , \nRightOut_33[9] , \nRightOut_33[8] , 
        \nRightOut_33[7] , \nRightOut_33[6] , \nRightOut_33[5] , 
        \nRightOut_33[4] , \nRightOut_33[3] , \nRightOut_33[2] , 
        \nRightOut_33[1] , \nRightOut_33[0] }), .inright({\nRightOut_35[16] , 
        \nRightOut_35[15] , \nRightOut_35[14] , \nRightOut_35[13] , 
        \nRightOut_35[12] , \nRightOut_35[11] , \nRightOut_35[10] , 
        \nRightOut_35[9] , \nRightOut_35[8] , \nRightOut_35[7] , 
        \nRightOut_35[6] , \nRightOut_35[5] , \nRightOut_35[4] , 
        \nRightOut_35[3] , \nRightOut_35[2] , \nRightOut_35[1] , 
        \nRightOut_35[0] }), .outleft({\nLeftOut_51[16] , \nLeftOut_51[15] , 
        \nLeftOut_51[14] , \nLeftOut_51[13] , \nLeftOut_51[12] , 
        \nLeftOut_51[11] , \nLeftOut_51[10] , \nLeftOut_51[9] , 
        \nLeftOut_51[8] , \nLeftOut_51[7] , \nLeftOut_51[6] , \nLeftOut_51[5] , 
        \nLeftOut_51[4] , \nLeftOut_51[3] , \nLeftOut_51[2] , \nLeftOut_51[1] , 
        \nLeftOut_51[0] }), .outright({\nRightOut_51[16] , \nRightOut_51[15] , 
        \nRightOut_51[14] , \nRightOut_51[13] , \nRightOut_51[12] , 
        \nRightOut_51[11] , \nRightOut_51[10] , \nRightOut_51[9] , 
        \nRightOut_51[8] , \nRightOut_51[7] , \nRightOut_51[6] , 
        \nRightOut_51[5] , \nRightOut_51[4] , \nRightOut_51[3] , 
        \nRightOut_51[2] , \nRightOut_51[1] , \nRightOut_51[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_64 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_48[16] , \nLeftOut_48[15] , \nLeftOut_48[14] , 
        \nLeftOut_48[13] , \nLeftOut_48[12] , \nLeftOut_48[11] , 
        \nLeftOut_48[10] , \nLeftOut_48[9] , \nLeftOut_48[8] , 
        \nLeftOut_48[7] , \nLeftOut_48[6] , \nLeftOut_48[5] , \nLeftOut_48[4] , 
        \nLeftOut_48[3] , \nLeftOut_48[2] , \nLeftOut_48[1] , \nLeftOut_48[0] 
        }), .inright({\nLeftOut_52[16] , \nLeftOut_52[15] , \nLeftOut_52[14] , 
        \nLeftOut_52[13] , \nLeftOut_52[12] , \nLeftOut_52[11] , 
        \nLeftOut_52[10] , \nLeftOut_52[9] , \nLeftOut_52[8] , 
        \nLeftOut_52[7] , \nLeftOut_52[6] , \nLeftOut_52[5] , \nLeftOut_52[4] , 
        \nLeftOut_52[3] , \nLeftOut_52[2] , \nLeftOut_52[1] , \nLeftOut_52[0] 
        }), .outleft({\nLeftOut_64[16] , \nLeftOut_64[15] , \nLeftOut_64[14] , 
        \nLeftOut_64[13] , \nLeftOut_64[12] , \nLeftOut_64[11] , 
        \nLeftOut_64[10] , \nLeftOut_64[9] , \nLeftOut_64[8] , 
        \nLeftOut_64[7] , \nLeftOut_64[6] , \nLeftOut_64[5] , \nLeftOut_64[4] , 
        \nLeftOut_64[3] , \nLeftOut_64[2] , \nLeftOut_64[1] , \nLeftOut_64[0] 
        }), .outright({\nRightOut_64[16] , \nRightOut_64[15] , 
        \nRightOut_64[14] , \nRightOut_64[13] , \nRightOut_64[12] , 
        \nRightOut_64[11] , \nRightOut_64[10] , \nRightOut_64[9] , 
        \nRightOut_64[8] , \nRightOut_64[7] , \nRightOut_64[6] , 
        \nRightOut_64[5] , \nRightOut_64[4] , \nRightOut_64[3] , 
        \nRightOut_64[2] , \nRightOut_64[1] , \nRightOut_64[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_76 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_56[16] , \nRightOut_56[15] , \nRightOut_56[14] , 
        \nRightOut_56[13] , \nRightOut_56[12] , \nRightOut_56[11] , 
        \nRightOut_56[10] , \nRightOut_56[9] , \nRightOut_56[8] , 
        \nRightOut_56[7] , \nRightOut_56[6] , \nRightOut_56[5] , 
        \nRightOut_56[4] , \nRightOut_56[3] , \nRightOut_56[2] , 
        \nRightOut_56[1] , \nRightOut_56[0] }), .inright({\nRightOut_60[16] , 
        \nRightOut_60[15] , \nRightOut_60[14] , \nRightOut_60[13] , 
        \nRightOut_60[12] , \nRightOut_60[11] , \nRightOut_60[10] , 
        \nRightOut_60[9] , \nRightOut_60[8] , \nRightOut_60[7] , 
        \nRightOut_60[6] , \nRightOut_60[5] , \nRightOut_60[4] , 
        \nRightOut_60[3] , \nRightOut_60[2] , \nRightOut_60[1] , 
        \nRightOut_60[0] }), .outleft({\nLeftOut_76[16] , \nLeftOut_76[15] , 
        \nLeftOut_76[14] , \nLeftOut_76[13] , \nLeftOut_76[12] , 
        \nLeftOut_76[11] , \nLeftOut_76[10] , \nLeftOut_76[9] , 
        \nLeftOut_76[8] , \nLeftOut_76[7] , \nLeftOut_76[6] , \nLeftOut_76[5] , 
        \nLeftOut_76[4] , \nLeftOut_76[3] , \nLeftOut_76[2] , \nLeftOut_76[1] , 
        \nLeftOut_76[0] }), .outright({\nRightOut_76[16] , \nRightOut_76[15] , 
        \nRightOut_76[14] , \nRightOut_76[13] , \nRightOut_76[12] , 
        \nRightOut_76[11] , \nRightOut_76[10] , \nRightOut_76[9] , 
        \nRightOut_76[8] , \nRightOut_76[7] , \nRightOut_76[6] , 
        \nRightOut_76[5] , \nRightOut_76[4] , \nRightOut_76[3] , 
        \nRightOut_76[2] , \nRightOut_76[1] , \nRightOut_76[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_24 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_8[16] , \nLeftOut_8[15] , \nLeftOut_8[14] , \nLeftOut_8[13] , 
        \nLeftOut_8[12] , \nLeftOut_8[11] , \nLeftOut_8[10] , \nLeftOut_8[9] , 
        \nLeftOut_8[8] , \nLeftOut_8[7] , \nLeftOut_8[6] , \nLeftOut_8[5] , 
        \nLeftOut_8[4] , \nLeftOut_8[3] , \nLeftOut_8[2] , \nLeftOut_8[1] , 
        \nLeftOut_8[0] }), .inright({\nRightOut_8[16] , \nRightOut_8[15] , 
        \nRightOut_8[14] , \nRightOut_8[13] , \nRightOut_8[12] , 
        \nRightOut_8[11] , \nRightOut_8[10] , \nRightOut_8[9] , 
        \nRightOut_8[8] , \nRightOut_8[7] , \nRightOut_8[6] , \nRightOut_8[5] , 
        \nRightOut_8[4] , \nRightOut_8[3] , \nRightOut_8[2] , \nRightOut_8[1] , 
        \nRightOut_8[0] }), .outleft({\nLeftOut_24[16] , \nLeftOut_24[15] , 
        \nLeftOut_24[14] , \nLeftOut_24[13] , \nLeftOut_24[12] , 
        \nLeftOut_24[11] , \nLeftOut_24[10] , \nLeftOut_24[9] , 
        \nLeftOut_24[8] , \nLeftOut_24[7] , \nLeftOut_24[6] , \nLeftOut_24[5] , 
        \nLeftOut_24[4] , \nLeftOut_24[3] , \nLeftOut_24[2] , \nLeftOut_24[1] , 
        \nLeftOut_24[0] }), .outright({\nRightOut_24[16] , \nRightOut_24[15] , 
        \nRightOut_24[14] , \nRightOut_24[13] , \nRightOut_24[12] , 
        \nRightOut_24[11] , \nRightOut_24[10] , \nRightOut_24[9] , 
        \nRightOut_24[8] , \nRightOut_24[7] , \nRightOut_24[6] , 
        \nRightOut_24[5] , \nRightOut_24[4] , \nRightOut_24[3] , 
        \nRightOut_24[2] , \nRightOut_24[1] , \nRightOut_24[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_88 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_64[16] , \nRightOut_64[15] , \nRightOut_64[14] , 
        \nRightOut_64[13] , \nRightOut_64[12] , \nRightOut_64[11] , 
        \nRightOut_64[10] , \nRightOut_64[9] , \nRightOut_64[8] , 
        \nRightOut_64[7] , \nRightOut_64[6] , \nRightOut_64[5] , 
        \nRightOut_64[4] , \nRightOut_64[3] , \nRightOut_64[2] , 
        \nRightOut_64[1] , \nRightOut_64[0] }), .inright({\nRightOut_72[16] , 
        \nRightOut_72[15] , \nRightOut_72[14] , \nRightOut_72[13] , 
        \nRightOut_72[12] , \nRightOut_72[11] , \nRightOut_72[10] , 
        \nRightOut_72[9] , \nRightOut_72[8] , \nRightOut_72[7] , 
        \nRightOut_72[6] , \nRightOut_72[5] , \nRightOut_72[4] , 
        \nRightOut_72[3] , \nRightOut_72[2] , \nRightOut_72[1] , 
        \nRightOut_72[0] }), .outleft({\nLeftOut_88[16] , \nLeftOut_88[15] , 
        \nLeftOut_88[14] , \nLeftOut_88[13] , \nLeftOut_88[12] , 
        \nLeftOut_88[11] , \nLeftOut_88[10] , \nLeftOut_88[9] , 
        \nLeftOut_88[8] , \nLeftOut_88[7] , \nLeftOut_88[6] , \nLeftOut_88[5] , 
        \nLeftOut_88[4] , \nLeftOut_88[3] , \nLeftOut_88[2] , \nLeftOut_88[1] , 
        \nLeftOut_88[0] }), .outright({\nRightOut_88[16] , \nRightOut_88[15] , 
        \nRightOut_88[14] , \nRightOut_88[13] , \nRightOut_88[12] , 
        \nRightOut_88[11] , \nRightOut_88[10] , \nRightOut_88[9] , 
        \nRightOut_88[8] , \nRightOut_88[7] , \nRightOut_88[6] , 
        \nRightOut_88[5] , \nRightOut_88[4] , \nRightOut_88[3] , 
        \nRightOut_88[2] , \nRightOut_88[1] , \nRightOut_88[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s13_SCAN1 node_93 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_69[16] , \nRightOut_69[15] , \nRightOut_69[14] , 
        \nRightOut_69[13] , \nRightOut_69[12] , \nRightOut_69[11] , 
        \nRightOut_69[10] , \nRightOut_69[9] , \nRightOut_69[8] , 
        \nRightOut_69[7] , \nRightOut_69[6] , \nRightOut_69[5] , 
        \nRightOut_69[4] , \nRightOut_69[3] , \nRightOut_69[2] , 
        \nRightOut_69[1] , \nRightOut_69[0] }), .inright({\nRightOut_77[16] , 
        \nRightOut_77[15] , \nRightOut_77[14] , \nRightOut_77[13] , 
        \nRightOut_77[12] , \nRightOut_77[11] , \nRightOut_77[10] , 
        \nRightOut_77[9] , \nRightOut_77[8] , \nRightOut_77[7] , 
        \nRightOut_77[6] , \nRightOut_77[5] , \nRightOut_77[4] , 
        \nRightOut_77[3] , \nRightOut_77[2] , \nRightOut_77[1] , 
        \nRightOut_77[0] }), .outleft({\nLeftOut_93[16] , \nLeftOut_93[15] , 
        \nLeftOut_93[14] , \nLeftOut_93[13] , \nLeftOut_93[12] , 
        \nLeftOut_93[11] , \nLeftOut_93[10] , \nLeftOut_93[9] , 
        \nLeftOut_93[8] , \nLeftOut_93[7] , \nLeftOut_93[6] , \nLeftOut_93[5] , 
        \nLeftOut_93[4] , \nLeftOut_93[3] , \nLeftOut_93[2] , \nLeftOut_93[1] , 
        \nLeftOut_93[0] }), .outright({\nRightOut_93[16] , \nRightOut_93[15] , 
        \nRightOut_93[14] , \nRightOut_93[13] , \nRightOut_93[12] , 
        \nRightOut_93[11] , \nRightOut_93[10] , \nRightOut_93[9] , 
        \nRightOut_93[8] , \nRightOut_93[7] , \nRightOut_93[6] , 
        \nRightOut_93[5] , \nRightOut_93[4] , \nRightOut_93[3] , 
        \nRightOut_93[2] , \nRightOut_93[1] , \nRightOut_93[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_108 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink28[15] , \ScanLink28[14] , \ScanLink28[13] , 
        \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , \ScanLink28[9] , 
        \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , \ScanLink28[5] , 
        \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , \ScanLink28[1] , 
        \ScanLink28[0] }), .ScanOut({\ScanLink29[15] , \ScanLink29[14] , 
        \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , 
        \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , 
        \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , 
        \ScanLink29[1] , \ScanLink29[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_88[16] , \nRightOut_88[15] , \nRightOut_88[14] , 
        \nRightOut_88[13] , \nRightOut_88[12] , \nRightOut_88[11] , 
        \nRightOut_88[10] , \nRightOut_88[9] , \nRightOut_88[8] , 
        \nRightOut_88[7] , \nRightOut_88[6] , \nRightOut_88[5] , 
        \nRightOut_88[4] , \nRightOut_88[3] , \nRightOut_88[2] , 
        \nRightOut_88[1] , \nRightOut_88[0] }), .inright({\nRightOut_89[16] , 
        \nRightOut_89[15] , \nRightOut_89[14] , \nRightOut_89[13] , 
        \nRightOut_89[12] , \nRightOut_89[11] , \nRightOut_89[10] , 
        \nRightOut_89[9] , \nRightOut_89[8] , \nRightOut_89[7] , 
        \nRightOut_89[6] , \nRightOut_89[5] , \nRightOut_89[4] , 
        \nRightOut_89[3] , \nRightOut_89[2] , \nRightOut_89[1] , 
        \nRightOut_89[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_41 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_24[16] , \nRightOut_24[15] , \nRightOut_24[14] , 
        \nRightOut_24[13] , \nRightOut_24[12] , \nRightOut_24[11] , 
        \nRightOut_24[10] , \nRightOut_24[9] , \nRightOut_24[8] , 
        \nRightOut_24[7] , \nRightOut_24[6] , \nRightOut_24[5] , 
        \nRightOut_24[4] , \nRightOut_24[3] , \nRightOut_24[2] , 
        \nRightOut_24[1] , \nRightOut_24[0] }), .inright({\nRightOut_25[16] , 
        \nRightOut_25[15] , \nRightOut_25[14] , \nRightOut_25[13] , 
        \nRightOut_25[12] , \nRightOut_25[11] , \nRightOut_25[10] , 
        \nRightOut_25[9] , \nRightOut_25[8] , \nRightOut_25[7] , 
        \nRightOut_25[6] , \nRightOut_25[5] , \nRightOut_25[4] , 
        \nRightOut_25[3] , \nRightOut_25[2] , \nRightOut_25[1] , 
        \nRightOut_25[0] }), .outleft({\nLeftOut_41[16] , \nLeftOut_41[15] , 
        \nLeftOut_41[14] , \nLeftOut_41[13] , \nLeftOut_41[12] , 
        \nLeftOut_41[11] , \nLeftOut_41[10] , \nLeftOut_41[9] , 
        \nLeftOut_41[8] , \nLeftOut_41[7] , \nLeftOut_41[6] , \nLeftOut_41[5] , 
        \nLeftOut_41[4] , \nLeftOut_41[3] , \nLeftOut_41[2] , \nLeftOut_41[1] , 
        \nLeftOut_41[0] }), .outright({\nRightOut_41[16] , \nRightOut_41[15] , 
        \nRightOut_41[14] , \nRightOut_41[13] , \nRightOut_41[12] , 
        \nRightOut_41[11] , \nRightOut_41[10] , \nRightOut_41[9] , 
        \nRightOut_41[8] , \nRightOut_41[7] , \nRightOut_41[6] , 
        \nRightOut_41[5] , \nRightOut_41[4] , \nRightOut_41[3] , 
        \nRightOut_41[2] , \nRightOut_41[1] , \nRightOut_41[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s4_SCAN1 node_66 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_50[16] , \nLeftOut_50[15] , \nLeftOut_50[14] , 
        \nLeftOut_50[13] , \nLeftOut_50[12] , \nLeftOut_50[11] , 
        \nLeftOut_50[10] , \nLeftOut_50[9] , \nLeftOut_50[8] , 
        \nLeftOut_50[7] , \nLeftOut_50[6] , \nLeftOut_50[5] , \nLeftOut_50[4] , 
        \nLeftOut_50[3] , \nLeftOut_50[2] , \nLeftOut_50[1] , \nLeftOut_50[0] 
        }), .inright({\nLeftOut_54[16] , \nLeftOut_54[15] , \nLeftOut_54[14] , 
        \nLeftOut_54[13] , \nLeftOut_54[12] , \nLeftOut_54[11] , 
        \nLeftOut_54[10] , \nLeftOut_54[9] , \nLeftOut_54[8] , 
        \nLeftOut_54[7] , \nLeftOut_54[6] , \nLeftOut_54[5] , \nLeftOut_54[4] , 
        \nLeftOut_54[3] , \nLeftOut_54[2] , \nLeftOut_54[1] , \nLeftOut_54[0] 
        }), .outleft({\nLeftOut_66[16] , \nLeftOut_66[15] , \nLeftOut_66[14] , 
        \nLeftOut_66[13] , \nLeftOut_66[12] , \nLeftOut_66[11] , 
        \nLeftOut_66[10] , \nLeftOut_66[9] , \nLeftOut_66[8] , 
        \nLeftOut_66[7] , \nLeftOut_66[6] , \nLeftOut_66[5] , \nLeftOut_66[4] , 
        \nLeftOut_66[3] , \nLeftOut_66[2] , \nLeftOut_66[1] , \nLeftOut_66[0] 
        }), .outright({\nRightOut_66[16] , \nRightOut_66[15] , 
        \nRightOut_66[14] , \nRightOut_66[13] , \nRightOut_66[12] , 
        \nRightOut_66[11] , \nRightOut_66[10] , \nRightOut_66[9] , 
        \nRightOut_66[8] , \nRightOut_66[7] , \nRightOut_66[6] , 
        \nRightOut_66[5] , \nRightOut_66[4] , \nRightOut_66[3] , 
        \nRightOut_66[2] , \nRightOut_66[1] , \nRightOut_66[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s3_SCAN1 node_83 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_67[16] , \nLeftOut_67[15] , \nLeftOut_67[14] , 
        \nLeftOut_67[13] , \nLeftOut_67[12] , \nLeftOut_67[11] , 
        \nLeftOut_67[10] , \nLeftOut_67[9] , \nLeftOut_67[8] , 
        \nLeftOut_67[7] , \nLeftOut_67[6] , \nLeftOut_67[5] , \nLeftOut_67[4] , 
        \nLeftOut_67[3] , \nLeftOut_67[2] , \nLeftOut_67[1] , \nLeftOut_67[0] 
        }), .inright({\nLeftOut_75[16] , \nLeftOut_75[15] , \nLeftOut_75[14] , 
        \nLeftOut_75[13] , \nLeftOut_75[12] , \nLeftOut_75[11] , 
        \nLeftOut_75[10] , \nLeftOut_75[9] , \nLeftOut_75[8] , 
        \nLeftOut_75[7] , \nLeftOut_75[6] , \nLeftOut_75[5] , \nLeftOut_75[4] , 
        \nLeftOut_75[3] , \nLeftOut_75[2] , \nLeftOut_75[1] , \nLeftOut_75[0] 
        }), .outleft({\nLeftOut_83[16] , \nLeftOut_83[15] , \nLeftOut_83[14] , 
        \nLeftOut_83[13] , \nLeftOut_83[12] , \nLeftOut_83[11] , 
        \nLeftOut_83[10] , \nLeftOut_83[9] , \nLeftOut_83[8] , 
        \nLeftOut_83[7] , \nLeftOut_83[6] , \nLeftOut_83[5] , \nLeftOut_83[4] , 
        \nLeftOut_83[3] , \nLeftOut_83[2] , \nLeftOut_83[1] , \nLeftOut_83[0] 
        }), .outright({\nRightOut_83[16] , \nRightOut_83[15] , 
        \nRightOut_83[14] , \nRightOut_83[13] , \nRightOut_83[12] , 
        \nRightOut_83[11] , \nRightOut_83[10] , \nRightOut_83[9] , 
        \nRightOut_83[8] , \nRightOut_83[7] , \nRightOut_83[6] , 
        \nRightOut_83[5] , \nRightOut_83[4] , \nRightOut_83[3] , 
        \nRightOut_83[2] , \nRightOut_83[1] , \nRightOut_83[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_103 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink23[15] , \ScanLink23[14] , \ScanLink23[13] , 
        \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , \ScanLink23[9] , 
        \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , \ScanLink23[5] , 
        \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , \ScanLink23[1] , 
        \ScanLink23[0] }), .ScanOut({\ScanLink24[15] , \ScanLink24[14] , 
        \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , 
        \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , 
        \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , 
        \ScanLink24[1] , \ScanLink24[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_94[16] , \nLeftOut_94[15] , \nLeftOut_94[14] , 
        \nLeftOut_94[13] , \nLeftOut_94[12] , \nLeftOut_94[11] , 
        \nLeftOut_94[10] , \nLeftOut_94[9] , \nLeftOut_94[8] , 
        \nLeftOut_94[7] , \nLeftOut_94[6] , \nLeftOut_94[5] , \nLeftOut_94[4] , 
        \nLeftOut_94[3] , \nLeftOut_94[2] , \nLeftOut_94[1] , \nLeftOut_94[0] 
        }), .inright({\nLeftOut_95[16] , \nLeftOut_95[15] , \nLeftOut_95[14] , 
        \nLeftOut_95[13] , \nLeftOut_95[12] , \nLeftOut_95[11] , 
        \nLeftOut_95[10] , \nLeftOut_95[9] , \nLeftOut_95[8] , 
        \nLeftOut_95[7] , \nLeftOut_95[6] , \nLeftOut_95[5] , \nLeftOut_95[4] , 
        \nLeftOut_95[3] , \nLeftOut_95[2] , \nLeftOut_95[1] , \nLeftOut_95[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_98 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink18[15] , \ScanLink18[14] , \ScanLink18[13] , 
        \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , \ScanLink18[9] , 
        \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , \ScanLink18[5] , 
        \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , \ScanLink18[1] , 
        \ScanLink18[0] }), .ScanOut({\ScanLink19[15] , \ScanLink19[14] , 
        \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , 
        \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , 
        \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , 
        \ScanLink19[1] , \ScanLink19[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_84[16] , \nLeftOut_84[15] , \nLeftOut_84[14] , 
        \nLeftOut_84[13] , \nLeftOut_84[12] , \nLeftOut_84[11] , 
        \nLeftOut_84[10] , \nLeftOut_84[9] , \nLeftOut_84[8] , 
        \nLeftOut_84[7] , \nLeftOut_84[6] , \nLeftOut_84[5] , \nLeftOut_84[4] , 
        \nLeftOut_84[3] , \nLeftOut_84[2] , \nLeftOut_84[1] , \nLeftOut_84[0] 
        }), .inright({\nLeftOut_85[16] , \nLeftOut_85[15] , \nLeftOut_85[14] , 
        \nLeftOut_85[13] , \nLeftOut_85[12] , \nLeftOut_85[11] , 
        \nLeftOut_85[10] , \nLeftOut_85[9] , \nLeftOut_85[8] , 
        \nLeftOut_85[7] , \nLeftOut_85[6] , \nLeftOut_85[5] , \nLeftOut_85[4] , 
        \nLeftOut_85[3] , \nLeftOut_85[2] , \nLeftOut_85[1] , \nLeftOut_85[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_34 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_18[16] , \nLeftOut_18[15] , \nLeftOut_18[14] , 
        \nLeftOut_18[13] , \nLeftOut_18[12] , \nLeftOut_18[11] , 
        \nLeftOut_18[10] , \nLeftOut_18[9] , \nLeftOut_18[8] , 
        \nLeftOut_18[7] , \nLeftOut_18[6] , \nLeftOut_18[5] , \nLeftOut_18[4] , 
        \nLeftOut_18[3] , \nLeftOut_18[2] , \nLeftOut_18[1] , \nLeftOut_18[0] 
        }), .inright({\nLeftOut_19[16] , \nLeftOut_19[15] , \nLeftOut_19[14] , 
        \nLeftOut_19[13] , \nLeftOut_19[12] , \nLeftOut_19[11] , 
        \nLeftOut_19[10] , \nLeftOut_19[9] , \nLeftOut_19[8] , 
        \nLeftOut_19[7] , \nLeftOut_19[6] , \nLeftOut_19[5] , \nLeftOut_19[4] , 
        \nLeftOut_19[3] , \nLeftOut_19[2] , \nLeftOut_19[1] , \nLeftOut_19[0] 
        }), .outleft({\nLeftOut_34[16] , \nLeftOut_34[15] , \nLeftOut_34[14] , 
        \nLeftOut_34[13] , \nLeftOut_34[12] , \nLeftOut_34[11] , 
        \nLeftOut_34[10] , \nLeftOut_34[9] , \nLeftOut_34[8] , 
        \nLeftOut_34[7] , \nLeftOut_34[6] , \nLeftOut_34[5] , \nLeftOut_34[4] , 
        \nLeftOut_34[3] , \nLeftOut_34[2] , \nLeftOut_34[1] , \nLeftOut_34[0] 
        }), .outright({\nRightOut_34[16] , \nRightOut_34[15] , 
        \nRightOut_34[14] , \nRightOut_34[13] , \nRightOut_34[12] , 
        \nRightOut_34[11] , \nRightOut_34[10] , \nRightOut_34[9] , 
        \nRightOut_34[8] , \nRightOut_34[7] , \nRightOut_34[6] , 
        \nRightOut_34[5] , \nRightOut_34[4] , \nRightOut_34[3] , 
        \nRightOut_34[2] , \nRightOut_34[1] , \nRightOut_34[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink9[15] , \ScanLink9[14] , \ScanLink9[13] , 
        \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , \ScanLink9[9] , 
        \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , \ScanLink9[5] , 
        \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , \ScanLink9[1] , 
        \ScanLink9[0] }), .ScanOut({\ScanLink10[15] , \ScanLink10[14] , 
        \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , 
        \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , 
        \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , 
        \ScanLink10[1] , \ScanLink10[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_9[16] , \nLeftOut_9[15] , \nLeftOut_9[14] , \nLeftOut_9[13] , 
        \nLeftOut_9[12] , \nLeftOut_9[11] , \nLeftOut_9[10] , \nLeftOut_9[9] , 
        \nLeftOut_9[8] , \nLeftOut_9[7] , \nLeftOut_9[6] , \nLeftOut_9[5] , 
        \nLeftOut_9[4] , \nLeftOut_9[3] , \nLeftOut_9[2] , \nLeftOut_9[1] , 
        \nLeftOut_9[0] }), .inright({\nRightOut_9[16] , \nRightOut_9[15] , 
        \nRightOut_9[14] , \nRightOut_9[13] , \nRightOut_9[12] , 
        \nRightOut_9[11] , \nRightOut_9[10] , \nRightOut_9[9] , 
        \nRightOut_9[8] , \nRightOut_9[7] , \nRightOut_9[6] , \nRightOut_9[5] , 
        \nRightOut_9[4] , \nRightOut_9[3] , \nRightOut_9[2] , \nRightOut_9[1] , 
        \nRightOut_9[0] }), .outleft({\nLeftOut_9[16] , \nLeftOut_9[15] , 
        \nLeftOut_9[14] , \nLeftOut_9[13] , \nLeftOut_9[12] , \nLeftOut_9[11] , 
        \nLeftOut_9[10] , \nLeftOut_9[9] , \nLeftOut_9[8] , \nLeftOut_9[7] , 
        \nLeftOut_9[6] , \nLeftOut_9[5] , \nLeftOut_9[4] , \nLeftOut_9[3] , 
        \nLeftOut_9[2] , \nLeftOut_9[1] , \nLeftOut_9[0] }), .outright({
        \nRightOut_9[16] , \nRightOut_9[15] , \nRightOut_9[14] , 
        \nRightOut_9[13] , \nRightOut_9[12] , \nRightOut_9[11] , 
        \nRightOut_9[10] , \nRightOut_9[9] , \nRightOut_9[8] , 
        \nRightOut_9[7] , \nRightOut_9[6] , \nRightOut_9[5] , \nRightOut_9[4] , 
        \nRightOut_9[3] , \nRightOut_9[2] , \nRightOut_9[1] , \nRightOut_9[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_26 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_10[16] , \nLeftOut_10[15] , \nLeftOut_10[14] , 
        \nLeftOut_10[13] , \nLeftOut_10[12] , \nLeftOut_10[11] , 
        \nLeftOut_10[10] , \nLeftOut_10[9] , \nLeftOut_10[8] , 
        \nLeftOut_10[7] , \nLeftOut_10[6] , \nLeftOut_10[5] , \nLeftOut_10[4] , 
        \nLeftOut_10[3] , \nLeftOut_10[2] , \nLeftOut_10[1] , \nLeftOut_10[0] 
        }), .inright({\nRightOut_10[16] , \nRightOut_10[15] , 
        \nRightOut_10[14] , \nRightOut_10[13] , \nRightOut_10[12] , 
        \nRightOut_10[11] , \nRightOut_10[10] , \nRightOut_10[9] , 
        \nRightOut_10[8] , \nRightOut_10[7] , \nRightOut_10[6] , 
        \nRightOut_10[5] , \nRightOut_10[4] , \nRightOut_10[3] , 
        \nRightOut_10[2] , \nRightOut_10[1] , \nRightOut_10[0] }), .outleft({
        \nLeftOut_26[16] , \nLeftOut_26[15] , \nLeftOut_26[14] , 
        \nLeftOut_26[13] , \nLeftOut_26[12] , \nLeftOut_26[11] , 
        \nLeftOut_26[10] , \nLeftOut_26[9] , \nLeftOut_26[8] , 
        \nLeftOut_26[7] , \nLeftOut_26[6] , \nLeftOut_26[5] , \nLeftOut_26[4] , 
        \nLeftOut_26[3] , \nLeftOut_26[2] , \nLeftOut_26[1] , \nLeftOut_26[0] 
        }), .outright({\nRightOut_26[16] , \nRightOut_26[15] , 
        \nRightOut_26[14] , \nRightOut_26[13] , \nRightOut_26[12] , 
        \nRightOut_26[11] , \nRightOut_26[10] , \nRightOut_26[9] , 
        \nRightOut_26[8] , \nRightOut_26[7] , \nRightOut_26[6] , 
        \nRightOut_26[5] , \nRightOut_26[4] , \nRightOut_26[3] , 
        \nRightOut_26[2] , \nRightOut_26[1] , \nRightOut_26[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_48 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_32[16] , \nLeftOut_32[15] , \nLeftOut_32[14] , 
        \nLeftOut_32[13] , \nLeftOut_32[12] , \nLeftOut_32[11] , 
        \nLeftOut_32[10] , \nLeftOut_32[9] , \nLeftOut_32[8] , 
        \nLeftOut_32[7] , \nLeftOut_32[6] , \nLeftOut_32[5] , \nLeftOut_32[4] , 
        \nLeftOut_32[3] , \nLeftOut_32[2] , \nLeftOut_32[1] , \nLeftOut_32[0] 
        }), .inright({\nLeftOut_34[16] , \nLeftOut_34[15] , \nLeftOut_34[14] , 
        \nLeftOut_34[13] , \nLeftOut_34[12] , \nLeftOut_34[11] , 
        \nLeftOut_34[10] , \nLeftOut_34[9] , \nLeftOut_34[8] , 
        \nLeftOut_34[7] , \nLeftOut_34[6] , \nLeftOut_34[5] , \nLeftOut_34[4] , 
        \nLeftOut_34[3] , \nLeftOut_34[2] , \nLeftOut_34[1] , \nLeftOut_34[0] 
        }), .outleft({\nLeftOut_48[16] , \nLeftOut_48[15] , \nLeftOut_48[14] , 
        \nLeftOut_48[13] , \nLeftOut_48[12] , \nLeftOut_48[11] , 
        \nLeftOut_48[10] , \nLeftOut_48[9] , \nLeftOut_48[8] , 
        \nLeftOut_48[7] , \nLeftOut_48[6] , \nLeftOut_48[5] , \nLeftOut_48[4] , 
        \nLeftOut_48[3] , \nLeftOut_48[2] , \nLeftOut_48[1] , \nLeftOut_48[0] 
        }), .outright({\nRightOut_48[16] , \nRightOut_48[15] , 
        \nRightOut_48[14] , \nRightOut_48[13] , \nRightOut_48[12] , 
        \nRightOut_48[11] , \nRightOut_48[10] , \nRightOut_48[9] , 
        \nRightOut_48[8] , \nRightOut_48[7] , \nRightOut_48[6] , 
        \nRightOut_48[5] , \nRightOut_48[4] , \nRightOut_48[3] , 
        \nRightOut_48[2] , \nRightOut_48[1] , \nRightOut_48[0] }) );
    FFT_Control_SIZE16_IDWIDTH1_SCAN1 node_Control ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink32[15] , \ScanLink32[14] , \ScanLink32[13] , 
        \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , \ScanLink32[9] , 
        \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , \ScanLink32[5] , 
        \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , \ScanLink32[1] , 
        \ScanLink32[0] }), .ScanOut({\ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), 
        .ScanId(1'b1), .Id(1'b0), .Enable(\nEnable[0] ) );
    FFT_Node_SIZE16_IDWIDTH1_s4_SCAN1 node_53 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_37[16] , \nLeftOut_37[15] , \nLeftOut_37[14] , 
        \nLeftOut_37[13] , \nLeftOut_37[12] , \nLeftOut_37[11] , 
        \nLeftOut_37[10] , \nLeftOut_37[9] , \nLeftOut_37[8] , 
        \nLeftOut_37[7] , \nLeftOut_37[6] , \nLeftOut_37[5] , \nLeftOut_37[4] , 
        \nLeftOut_37[3] , \nLeftOut_37[2] , \nLeftOut_37[1] , \nLeftOut_37[0] 
        }), .inright({\nLeftOut_39[16] , \nLeftOut_39[15] , \nLeftOut_39[14] , 
        \nLeftOut_39[13] , \nLeftOut_39[12] , \nLeftOut_39[11] , 
        \nLeftOut_39[10] , \nLeftOut_39[9] , \nLeftOut_39[8] , 
        \nLeftOut_39[7] , \nLeftOut_39[6] , \nLeftOut_39[5] , \nLeftOut_39[4] , 
        \nLeftOut_39[3] , \nLeftOut_39[2] , \nLeftOut_39[1] , \nLeftOut_39[0] 
        }), .outleft({\nLeftOut_53[16] , \nLeftOut_53[15] , \nLeftOut_53[14] , 
        \nLeftOut_53[13] , \nLeftOut_53[12] , \nLeftOut_53[11] , 
        \nLeftOut_53[10] , \nLeftOut_53[9] , \nLeftOut_53[8] , 
        \nLeftOut_53[7] , \nLeftOut_53[6] , \nLeftOut_53[5] , \nLeftOut_53[4] , 
        \nLeftOut_53[3] , \nLeftOut_53[2] , \nLeftOut_53[1] , \nLeftOut_53[0] 
        }), .outright({\nRightOut_53[16] , \nRightOut_53[15] , 
        \nRightOut_53[14] , \nRightOut_53[13] , \nRightOut_53[12] , 
        \nRightOut_53[11] , \nRightOut_53[10] , \nRightOut_53[9] , 
        \nRightOut_53[8] , \nRightOut_53[7] , \nRightOut_53[6] , 
        \nRightOut_53[5] , \nRightOut_53[4] , \nRightOut_53[3] , 
        \nRightOut_53[2] , \nRightOut_53[1] , \nRightOut_53[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s4_SCAN1 node_74 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_58[16] , \nLeftOut_58[15] , \nLeftOut_58[14] , 
        \nLeftOut_58[13] , \nLeftOut_58[12] , \nLeftOut_58[11] , 
        \nLeftOut_58[10] , \nLeftOut_58[9] , \nLeftOut_58[8] , 
        \nLeftOut_58[7] , \nLeftOut_58[6] , \nLeftOut_58[5] , \nLeftOut_58[4] , 
        \nLeftOut_58[3] , \nLeftOut_58[2] , \nLeftOut_58[1] , \nLeftOut_58[0] 
        }), .inright({\nLeftOut_62[16] , \nLeftOut_62[15] , \nLeftOut_62[14] , 
        \nLeftOut_62[13] , \nLeftOut_62[12] , \nLeftOut_62[11] , 
        \nLeftOut_62[10] , \nLeftOut_62[9] , \nLeftOut_62[8] , 
        \nLeftOut_62[7] , \nLeftOut_62[6] , \nLeftOut_62[5] , \nLeftOut_62[4] , 
        \nLeftOut_62[3] , \nLeftOut_62[2] , \nLeftOut_62[1] , \nLeftOut_62[0] 
        }), .outleft({\nLeftOut_74[16] , \nLeftOut_74[15] , \nLeftOut_74[14] , 
        \nLeftOut_74[13] , \nLeftOut_74[12] , \nLeftOut_74[11] , 
        \nLeftOut_74[10] , \nLeftOut_74[9] , \nLeftOut_74[8] , 
        \nLeftOut_74[7] , \nLeftOut_74[6] , \nLeftOut_74[5] , \nLeftOut_74[4] , 
        \nLeftOut_74[3] , \nLeftOut_74[2] , \nLeftOut_74[1] , \nLeftOut_74[0] 
        }), .outright({\nRightOut_74[16] , \nRightOut_74[15] , 
        \nRightOut_74[14] , \nRightOut_74[13] , \nRightOut_74[12] , 
        \nRightOut_74[11] , \nRightOut_74[10] , \nRightOut_74[9] , 
        \nRightOut_74[8] , \nRightOut_74[7] , \nRightOut_74[6] , 
        \nRightOut_74[5] , \nRightOut_74[4] , \nRightOut_74[3] , 
        \nRightOut_74[2] , \nRightOut_74[1] , \nRightOut_74[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s11_SCAN1 node_91 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_67[16] , \nRightOut_67[15] , \nRightOut_67[14] , 
        \nRightOut_67[13] , \nRightOut_67[12] , \nRightOut_67[11] , 
        \nRightOut_67[10] , \nRightOut_67[9] , \nRightOut_67[8] , 
        \nRightOut_67[7] , \nRightOut_67[6] , \nRightOut_67[5] , 
        \nRightOut_67[4] , \nRightOut_67[3] , \nRightOut_67[2] , 
        \nRightOut_67[1] , \nRightOut_67[0] }), .inright({\nRightOut_75[16] , 
        \nRightOut_75[15] , \nRightOut_75[14] , \nRightOut_75[13] , 
        \nRightOut_75[12] , \nRightOut_75[11] , \nRightOut_75[10] , 
        \nRightOut_75[9] , \nRightOut_75[8] , \nRightOut_75[7] , 
        \nRightOut_75[6] , \nRightOut_75[5] , \nRightOut_75[4] , 
        \nRightOut_75[3] , \nRightOut_75[2] , \nRightOut_75[1] , 
        \nRightOut_75[0] }), .outleft({\nLeftOut_91[16] , \nLeftOut_91[15] , 
        \nLeftOut_91[14] , \nLeftOut_91[13] , \nLeftOut_91[12] , 
        \nLeftOut_91[11] , \nLeftOut_91[10] , \nLeftOut_91[9] , 
        \nLeftOut_91[8] , \nLeftOut_91[7] , \nLeftOut_91[6] , \nLeftOut_91[5] , 
        \nLeftOut_91[4] , \nLeftOut_91[3] , \nLeftOut_91[2] , \nLeftOut_91[1] , 
        \nLeftOut_91[0] }), .outright({\nRightOut_91[16] , \nRightOut_91[15] , 
        \nRightOut_91[14] , \nRightOut_91[13] , \nRightOut_91[12] , 
        \nRightOut_91[11] , \nRightOut_91[10] , \nRightOut_91[9] , 
        \nRightOut_91[8] , \nRightOut_91[7] , \nRightOut_91[6] , 
        \nRightOut_91[5] , \nRightOut_91[4] , \nRightOut_91[3] , 
        \nRightOut_91[2] , \nRightOut_91[1] , \nRightOut_91[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_111 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink31[15] , \ScanLink31[14] , \ScanLink31[13] , 
        \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , \ScanLink31[9] , 
        \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , \ScanLink31[5] , 
        \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , \ScanLink31[1] , 
        \ScanLink31[0] }), .ScanOut({\ScanLink32[15] , \ScanLink32[14] , 
        \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , 
        \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , 
        \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , 
        \ScanLink32[1] , \ScanLink32[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_94[16] , \nRightOut_94[15] , \nRightOut_94[14] , 
        \nRightOut_94[13] , \nRightOut_94[12] , \nRightOut_94[11] , 
        \nRightOut_94[10] , \nRightOut_94[9] , \nRightOut_94[8] , 
        \nRightOut_94[7] , \nRightOut_94[6] , \nRightOut_94[5] , 
        \nRightOut_94[4] , \nRightOut_94[3] , \nRightOut_94[2] , 
        \nRightOut_94[1] , \nRightOut_94[0] }), .inright({\nRightOut_95[16] , 
        \nRightOut_95[15] , \nRightOut_95[14] , \nRightOut_95[13] , 
        \nRightOut_95[12] , \nRightOut_95[11] , \nRightOut_95[10] , 
        \nRightOut_95[9] , \nRightOut_95[8] , \nRightOut_95[7] , 
        \nRightOut_95[6] , \nRightOut_95[5] , \nRightOut_95[4] , 
        \nRightOut_95[3] , \nRightOut_95[2] , \nRightOut_95[1] , 
        \nRightOut_95[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_54 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_36[16] , \nRightOut_36[15] , \nRightOut_36[14] , 
        \nRightOut_36[13] , \nRightOut_36[12] , \nRightOut_36[11] , 
        \nRightOut_36[10] , \nRightOut_36[9] , \nRightOut_36[8] , 
        \nRightOut_36[7] , \nRightOut_36[6] , \nRightOut_36[5] , 
        \nRightOut_36[4] , \nRightOut_36[3] , \nRightOut_36[2] , 
        \nRightOut_36[1] , \nRightOut_36[0] }), .inright({\nRightOut_38[16] , 
        \nRightOut_38[15] , \nRightOut_38[14] , \nRightOut_38[13] , 
        \nRightOut_38[12] , \nRightOut_38[11] , \nRightOut_38[10] , 
        \nRightOut_38[9] , \nRightOut_38[8] , \nRightOut_38[7] , 
        \nRightOut_38[6] , \nRightOut_38[5] , \nRightOut_38[4] , 
        \nRightOut_38[3] , \nRightOut_38[2] , \nRightOut_38[1] , 
        \nRightOut_38[0] }), .outleft({\nLeftOut_54[16] , \nLeftOut_54[15] , 
        \nLeftOut_54[14] , \nLeftOut_54[13] , \nLeftOut_54[12] , 
        \nLeftOut_54[11] , \nLeftOut_54[10] , \nLeftOut_54[9] , 
        \nLeftOut_54[8] , \nLeftOut_54[7] , \nLeftOut_54[6] , \nLeftOut_54[5] , 
        \nLeftOut_54[4] , \nLeftOut_54[3] , \nLeftOut_54[2] , \nLeftOut_54[1] , 
        \nLeftOut_54[0] }), .outright({\nRightOut_54[16] , \nRightOut_54[15] , 
        \nRightOut_54[14] , \nRightOut_54[13] , \nRightOut_54[12] , 
        \nRightOut_54[11] , \nRightOut_54[10] , \nRightOut_54[9] , 
        \nRightOut_54[8] , \nRightOut_54[7] , \nRightOut_54[6] , 
        \nRightOut_54[5] , \nRightOut_54[4] , \nRightOut_54[3] , 
        \nRightOut_54[2] , \nRightOut_54[1] , \nRightOut_54[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s2_SCAN1 node_73 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_57[16] , \nLeftOut_57[15] , \nLeftOut_57[14] , 
        \nLeftOut_57[13] , \nLeftOut_57[12] , \nLeftOut_57[11] , 
        \nLeftOut_57[10] , \nLeftOut_57[9] , \nLeftOut_57[8] , 
        \nLeftOut_57[7] , \nLeftOut_57[6] , \nLeftOut_57[5] , \nLeftOut_57[4] , 
        \nLeftOut_57[3] , \nLeftOut_57[2] , \nLeftOut_57[1] , \nLeftOut_57[0] 
        }), .inright({\nLeftOut_61[16] , \nLeftOut_61[15] , \nLeftOut_61[14] , 
        \nLeftOut_61[13] , \nLeftOut_61[12] , \nLeftOut_61[11] , 
        \nLeftOut_61[10] , \nLeftOut_61[9] , \nLeftOut_61[8] , 
        \nLeftOut_61[7] , \nLeftOut_61[6] , \nLeftOut_61[5] , \nLeftOut_61[4] , 
        \nLeftOut_61[3] , \nLeftOut_61[2] , \nLeftOut_61[1] , \nLeftOut_61[0] 
        }), .outleft({\nLeftOut_73[16] , \nLeftOut_73[15] , \nLeftOut_73[14] , 
        \nLeftOut_73[13] , \nLeftOut_73[12] , \nLeftOut_73[11] , 
        \nLeftOut_73[10] , \nLeftOut_73[9] , \nLeftOut_73[8] , 
        \nLeftOut_73[7] , \nLeftOut_73[6] , \nLeftOut_73[5] , \nLeftOut_73[4] , 
        \nLeftOut_73[3] , \nLeftOut_73[2] , \nLeftOut_73[1] , \nLeftOut_73[0] 
        }), .outright({\nRightOut_73[16] , \nRightOut_73[15] , 
        \nRightOut_73[14] , \nRightOut_73[13] , \nRightOut_73[12] , 
        \nRightOut_73[11] , \nRightOut_73[10] , \nRightOut_73[9] , 
        \nRightOut_73[8] , \nRightOut_73[7] , \nRightOut_73[6] , 
        \nRightOut_73[5] , \nRightOut_73[4] , \nRightOut_73[3] , 
        \nRightOut_73[2] , \nRightOut_73[1] , \nRightOut_73[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_21 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_5[16] , \nLeftOut_5[15] , \nLeftOut_5[14] , \nLeftOut_5[13] , 
        \nLeftOut_5[12] , \nLeftOut_5[11] , \nLeftOut_5[10] , \nLeftOut_5[9] , 
        \nLeftOut_5[8] , \nLeftOut_5[7] , \nLeftOut_5[6] , \nLeftOut_5[5] , 
        \nLeftOut_5[4] , \nLeftOut_5[3] , \nLeftOut_5[2] , \nLeftOut_5[1] , 
        \nLeftOut_5[0] }), .inright({\nRightOut_5[16] , \nRightOut_5[15] , 
        \nRightOut_5[14] , \nRightOut_5[13] , \nRightOut_5[12] , 
        \nRightOut_5[11] , \nRightOut_5[10] , \nRightOut_5[9] , 
        \nRightOut_5[8] , \nRightOut_5[7] , \nRightOut_5[6] , \nRightOut_5[5] , 
        \nRightOut_5[4] , \nRightOut_5[3] , \nRightOut_5[2] , \nRightOut_5[1] , 
        \nRightOut_5[0] }), .outleft({\nLeftOut_21[16] , \nLeftOut_21[15] , 
        \nLeftOut_21[14] , \nLeftOut_21[13] , \nLeftOut_21[12] , 
        \nLeftOut_21[11] , \nLeftOut_21[10] , \nLeftOut_21[9] , 
        \nLeftOut_21[8] , \nLeftOut_21[7] , \nLeftOut_21[6] , \nLeftOut_21[5] , 
        \nLeftOut_21[4] , \nLeftOut_21[3] , \nLeftOut_21[2] , \nLeftOut_21[1] , 
        \nLeftOut_21[0] }), .outright({\nRightOut_21[16] , \nRightOut_21[15] , 
        \nRightOut_21[14] , \nRightOut_21[13] , \nRightOut_21[12] , 
        \nRightOut_21[11] , \nRightOut_21[10] , \nRightOut_21[9] , 
        \nRightOut_21[8] , \nRightOut_21[7] , \nRightOut_21[6] , 
        \nRightOut_21[5] , \nRightOut_21[4] , \nRightOut_21[3] , 
        \nRightOut_21[2] , \nRightOut_21[1] , \nRightOut_21[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_96 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink16[15] , \ScanLink16[14] , \ScanLink16[13] , 
        \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , \ScanLink16[9] , 
        \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , \ScanLink16[5] , 
        \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , \ScanLink16[1] , 
        \ScanLink16[0] }), .ScanOut({\ScanLink17[15] , \ScanLink17[14] , 
        \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , 
        \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , 
        \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , 
        \ScanLink17[1] , \ScanLink17[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_80[16] , \nLeftOut_80[15] , \nLeftOut_80[14] , 
        \nLeftOut_80[13] , \nLeftOut_80[12] , \nLeftOut_80[11] , 
        \nLeftOut_80[10] , \nLeftOut_80[9] , \nLeftOut_80[8] , 
        \nLeftOut_80[7] , \nLeftOut_80[6] , \nLeftOut_80[5] , \nLeftOut_80[4] , 
        \nLeftOut_80[3] , \nLeftOut_80[2] , \nLeftOut_80[1] , \nLeftOut_80[0] 
        }), .inright({\nLeftOut_81[16] , \nLeftOut_81[15] , \nLeftOut_81[14] , 
        \nLeftOut_81[13] , \nLeftOut_81[12] , \nLeftOut_81[11] , 
        \nLeftOut_81[10] , \nLeftOut_81[9] , \nLeftOut_81[8] , 
        \nLeftOut_81[7] , \nLeftOut_81[6] , \nLeftOut_81[5] , \nLeftOut_81[4] , 
        \nLeftOut_81[3] , \nLeftOut_81[2] , \nLeftOut_81[1] , \nLeftOut_81[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_68 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_48[16] , \nRightOut_48[15] , \nRightOut_48[14] , 
        \nRightOut_48[13] , \nRightOut_48[12] , \nRightOut_48[11] , 
        \nRightOut_48[10] , \nRightOut_48[9] , \nRightOut_48[8] , 
        \nRightOut_48[7] , \nRightOut_48[6] , \nRightOut_48[5] , 
        \nRightOut_48[4] , \nRightOut_48[3] , \nRightOut_48[2] , 
        \nRightOut_48[1] , \nRightOut_48[0] }), .inright({\nRightOut_52[16] , 
        \nRightOut_52[15] , \nRightOut_52[14] , \nRightOut_52[13] , 
        \nRightOut_52[12] , \nRightOut_52[11] , \nRightOut_52[10] , 
        \nRightOut_52[9] , \nRightOut_52[8] , \nRightOut_52[7] , 
        \nRightOut_52[6] , \nRightOut_52[5] , \nRightOut_52[4] , 
        \nRightOut_52[3] , \nRightOut_52[2] , \nRightOut_52[1] , 
        \nRightOut_52[0] }), .outleft({\nLeftOut_68[16] , \nLeftOut_68[15] , 
        \nLeftOut_68[14] , \nLeftOut_68[13] , \nLeftOut_68[12] , 
        \nLeftOut_68[11] , \nLeftOut_68[10] , \nLeftOut_68[9] , 
        \nLeftOut_68[8] , \nLeftOut_68[7] , \nLeftOut_68[6] , \nLeftOut_68[5] , 
        \nLeftOut_68[4] , \nLeftOut_68[3] , \nLeftOut_68[2] , \nLeftOut_68[1] , 
        \nLeftOut_68[0] }), .outright({\nRightOut_68[16] , \nRightOut_68[15] , 
        \nRightOut_68[14] , \nRightOut_68[13] , \nRightOut_68[12] , 
        \nRightOut_68[11] , \nRightOut_68[10] , \nRightOut_68[9] , 
        \nRightOut_68[8] , \nRightOut_68[7] , \nRightOut_68[6] , 
        \nRightOut_68[5] , \nRightOut_68[4] , \nRightOut_68[3] , 
        \nRightOut_68[2] , \nRightOut_68[1] , \nRightOut_68[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink1[15] , \ScanLink1[14] , \ScanLink1[13] , 
        \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , \ScanLink1[9] , 
        \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , \ScanLink1[5] , 
        \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , \ScanLink1[1] , 
        \ScanLink1[0] }), .ScanOut({\ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_1[16] , \nLeftOut_1[15] , \nLeftOut_1[14] , \nLeftOut_1[13] , 
        \nLeftOut_1[12] , \nLeftOut_1[11] , \nLeftOut_1[10] , \nLeftOut_1[9] , 
        \nLeftOut_1[8] , \nLeftOut_1[7] , \nLeftOut_1[6] , \nLeftOut_1[5] , 
        \nLeftOut_1[4] , \nLeftOut_1[3] , \nLeftOut_1[2] , \nLeftOut_1[1] , 
        \nLeftOut_1[0] }), .inright({\nRightOut_1[16] , \nRightOut_1[15] , 
        \nRightOut_1[14] , \nRightOut_1[13] , \nRightOut_1[12] , 
        \nRightOut_1[11] , \nRightOut_1[10] , \nRightOut_1[9] , 
        \nRightOut_1[8] , \nRightOut_1[7] , \nRightOut_1[6] , \nRightOut_1[5] , 
        \nRightOut_1[4] , \nRightOut_1[3] , \nRightOut_1[2] , \nRightOut_1[1] , 
        \nRightOut_1[0] }), .outleft({\nLeftOut_1[16] , \nLeftOut_1[15] , 
        \nLeftOut_1[14] , \nLeftOut_1[13] , \nLeftOut_1[12] , \nLeftOut_1[11] , 
        \nLeftOut_1[10] , \nLeftOut_1[9] , \nLeftOut_1[8] , \nLeftOut_1[7] , 
        \nLeftOut_1[6] , \nLeftOut_1[5] , \nLeftOut_1[4] , \nLeftOut_1[3] , 
        \nLeftOut_1[2] , \nLeftOut_1[1] , \nLeftOut_1[0] }), .outright({
        \nRightOut_1[16] , \nRightOut_1[15] , \nRightOut_1[14] , 
        \nRightOut_1[13] , \nRightOut_1[12] , \nRightOut_1[11] , 
        \nRightOut_1[10] , \nRightOut_1[9] , \nRightOut_1[8] , 
        \nRightOut_1[7] , \nRightOut_1[6] , \nRightOut_1[5] , \nRightOut_1[4] , 
        \nRightOut_1[3] , \nRightOut_1[2] , \nRightOut_1[1] , \nRightOut_1[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink8[15] , \ScanLink8[14] , \ScanLink8[13] , 
        \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , \ScanLink8[9] , 
        \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , \ScanLink8[5] , 
        \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , \ScanLink8[1] , 
        \ScanLink8[0] }), .ScanOut({\ScanLink9[15] , \ScanLink9[14] , 
        \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , 
        \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , 
        \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , 
        \ScanLink9[1] , \ScanLink9[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_8[16] , \nLeftOut_8[15] , \nLeftOut_8[14] , \nLeftOut_8[13] , 
        \nLeftOut_8[12] , \nLeftOut_8[11] , \nLeftOut_8[10] , \nLeftOut_8[9] , 
        \nLeftOut_8[8] , \nLeftOut_8[7] , \nLeftOut_8[6] , \nLeftOut_8[5] , 
        \nLeftOut_8[4] , \nLeftOut_8[3] , \nLeftOut_8[2] , \nLeftOut_8[1] , 
        \nLeftOut_8[0] }), .inright({\nRightOut_8[16] , \nRightOut_8[15] , 
        \nRightOut_8[14] , \nRightOut_8[13] , \nRightOut_8[12] , 
        \nRightOut_8[11] , \nRightOut_8[10] , \nRightOut_8[9] , 
        \nRightOut_8[8] , \nRightOut_8[7] , \nRightOut_8[6] , \nRightOut_8[5] , 
        \nRightOut_8[4] , \nRightOut_8[3] , \nRightOut_8[2] , \nRightOut_8[1] , 
        \nRightOut_8[0] }), .outleft({\nLeftOut_8[16] , \nLeftOut_8[15] , 
        \nLeftOut_8[14] , \nLeftOut_8[13] , \nLeftOut_8[12] , \nLeftOut_8[11] , 
        \nLeftOut_8[10] , \nLeftOut_8[9] , \nLeftOut_8[8] , \nLeftOut_8[7] , 
        \nLeftOut_8[6] , \nLeftOut_8[5] , \nLeftOut_8[4] , \nLeftOut_8[3] , 
        \nLeftOut_8[2] , \nLeftOut_8[1] , \nLeftOut_8[0] }), .outright({
        \nRightOut_8[16] , \nRightOut_8[15] , \nRightOut_8[14] , 
        \nRightOut_8[13] , \nRightOut_8[12] , \nRightOut_8[11] , 
        \nRightOut_8[10] , \nRightOut_8[9] , \nRightOut_8[8] , 
        \nRightOut_8[7] , \nRightOut_8[6] , \nRightOut_8[5] , \nRightOut_8[4] , 
        \nRightOut_8[3] , \nRightOut_8[2] , \nRightOut_8[1] , \nRightOut_8[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_14 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink14[15] , \ScanLink14[14] , \ScanLink14[13] , 
        \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , \ScanLink14[9] , 
        \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , \ScanLink14[5] , 
        \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , \ScanLink14[1] , 
        \ScanLink14[0] }), .ScanOut({\ScanLink15[15] , \ScanLink15[14] , 
        \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , 
        \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , 
        \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , 
        \ScanLink15[1] , \ScanLink15[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_14[16] , \nLeftOut_14[15] , \nLeftOut_14[14] , 
        \nLeftOut_14[13] , \nLeftOut_14[12] , \nLeftOut_14[11] , 
        \nLeftOut_14[10] , \nLeftOut_14[9] , \nLeftOut_14[8] , 
        \nLeftOut_14[7] , \nLeftOut_14[6] , \nLeftOut_14[5] , \nLeftOut_14[4] , 
        \nLeftOut_14[3] , \nLeftOut_14[2] , \nLeftOut_14[1] , \nLeftOut_14[0] 
        }), .inright({\nRightOut_14[16] , \nRightOut_14[15] , 
        \nRightOut_14[14] , \nRightOut_14[13] , \nRightOut_14[12] , 
        \nRightOut_14[11] , \nRightOut_14[10] , \nRightOut_14[9] , 
        \nRightOut_14[8] , \nRightOut_14[7] , \nRightOut_14[6] , 
        \nRightOut_14[5] , \nRightOut_14[4] , \nRightOut_14[3] , 
        \nRightOut_14[2] , \nRightOut_14[1] , \nRightOut_14[0] }), .outleft({
        \nLeftOut_14[16] , \nLeftOut_14[15] , \nLeftOut_14[14] , 
        \nLeftOut_14[13] , \nLeftOut_14[12] , \nLeftOut_14[11] , 
        \nLeftOut_14[10] , \nLeftOut_14[9] , \nLeftOut_14[8] , 
        \nLeftOut_14[7] , \nLeftOut_14[6] , \nLeftOut_14[5] , \nLeftOut_14[4] , 
        \nLeftOut_14[3] , \nLeftOut_14[2] , \nLeftOut_14[1] , \nLeftOut_14[0] 
        }), .outright({\nRightOut_14[16] , \nRightOut_14[15] , 
        \nRightOut_14[14] , \nRightOut_14[13] , \nRightOut_14[12] , 
        \nRightOut_14[11] , \nRightOut_14[10] , \nRightOut_14[9] , 
        \nRightOut_14[8] , \nRightOut_14[7] , \nRightOut_14[6] , 
        \nRightOut_14[5] , \nRightOut_14[4] , \nRightOut_14[3] , 
        \nRightOut_14[2] , \nRightOut_14[1] , \nRightOut_14[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_33 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_16[16] , \nRightOut_16[15] , \nRightOut_16[14] , 
        \nRightOut_16[13] , \nRightOut_16[12] , \nRightOut_16[11] , 
        \nRightOut_16[10] , \nRightOut_16[9] , \nRightOut_16[8] , 
        \nRightOut_16[7] , \nRightOut_16[6] , \nRightOut_16[5] , 
        \nRightOut_16[4] , \nRightOut_16[3] , \nRightOut_16[2] , 
        \nRightOut_16[1] , \nRightOut_16[0] }), .inright({\nRightOut_17[16] , 
        \nRightOut_17[15] , \nRightOut_17[14] , \nRightOut_17[13] , 
        \nRightOut_17[12] , \nRightOut_17[11] , \nRightOut_17[10] , 
        \nRightOut_17[9] , \nRightOut_17[8] , \nRightOut_17[7] , 
        \nRightOut_17[6] , \nRightOut_17[5] , \nRightOut_17[4] , 
        \nRightOut_17[3] , \nRightOut_17[2] , \nRightOut_17[1] , 
        \nRightOut_17[0] }), .outleft({\nLeftOut_33[16] , \nLeftOut_33[15] , 
        \nLeftOut_33[14] , \nLeftOut_33[13] , \nLeftOut_33[12] , 
        \nLeftOut_33[11] , \nLeftOut_33[10] , \nLeftOut_33[9] , 
        \nLeftOut_33[8] , \nLeftOut_33[7] , \nLeftOut_33[6] , \nLeftOut_33[5] , 
        \nLeftOut_33[4] , \nLeftOut_33[3] , \nLeftOut_33[2] , \nLeftOut_33[1] , 
        \nLeftOut_33[0] }), .outright({\nRightOut_33[16] , \nRightOut_33[15] , 
        \nRightOut_33[14] , \nRightOut_33[13] , \nRightOut_33[12] , 
        \nRightOut_33[11] , \nRightOut_33[10] , \nRightOut_33[9] , 
        \nRightOut_33[8] , \nRightOut_33[7] , \nRightOut_33[6] , 
        \nRightOut_33[5] , \nRightOut_33[4] , \nRightOut_33[3] , 
        \nRightOut_33[2] , \nRightOut_33[1] , \nRightOut_33[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_20 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_4[16] , \nLeftOut_4[15] , \nLeftOut_4[14] , \nLeftOut_4[13] , 
        \nLeftOut_4[12] , \nLeftOut_4[11] , \nLeftOut_4[10] , \nLeftOut_4[9] , 
        \nLeftOut_4[8] , \nLeftOut_4[7] , \nLeftOut_4[6] , \nLeftOut_4[5] , 
        \nLeftOut_4[4] , \nLeftOut_4[3] , \nLeftOut_4[2] , \nLeftOut_4[1] , 
        \nLeftOut_4[0] }), .inright({\nRightOut_4[16] , \nRightOut_4[15] , 
        \nRightOut_4[14] , \nRightOut_4[13] , \nRightOut_4[12] , 
        \nRightOut_4[11] , \nRightOut_4[10] , \nRightOut_4[9] , 
        \nRightOut_4[8] , \nRightOut_4[7] , \nRightOut_4[6] , \nRightOut_4[5] , 
        \nRightOut_4[4] , \nRightOut_4[3] , \nRightOut_4[2] , \nRightOut_4[1] , 
        \nRightOut_4[0] }), .outleft({\nLeftOut_20[16] , \nLeftOut_20[15] , 
        \nLeftOut_20[14] , \nLeftOut_20[13] , \nLeftOut_20[12] , 
        \nLeftOut_20[11] , \nLeftOut_20[10] , \nLeftOut_20[9] , 
        \nLeftOut_20[8] , \nLeftOut_20[7] , \nLeftOut_20[6] , \nLeftOut_20[5] , 
        \nLeftOut_20[4] , \nLeftOut_20[3] , \nLeftOut_20[2] , \nLeftOut_20[1] , 
        \nLeftOut_20[0] }), .outright({\nRightOut_20[16] , \nRightOut_20[15] , 
        \nRightOut_20[14] , \nRightOut_20[13] , \nRightOut_20[12] , 
        \nRightOut_20[11] , \nRightOut_20[10] , \nRightOut_20[9] , 
        \nRightOut_20[8] , \nRightOut_20[7] , \nRightOut_20[6] , 
        \nRightOut_20[5] , \nRightOut_20[4] , \nRightOut_20[3] , 
        \nRightOut_20[2] , \nRightOut_20[1] , \nRightOut_20[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_28 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_12[16] , \nLeftOut_12[15] , \nLeftOut_12[14] , 
        \nLeftOut_12[13] , \nLeftOut_12[12] , \nLeftOut_12[11] , 
        \nLeftOut_12[10] , \nLeftOut_12[9] , \nLeftOut_12[8] , 
        \nLeftOut_12[7] , \nLeftOut_12[6] , \nLeftOut_12[5] , \nLeftOut_12[4] , 
        \nLeftOut_12[3] , \nLeftOut_12[2] , \nLeftOut_12[1] , \nLeftOut_12[0] 
        }), .inright({\nRightOut_12[16] , \nRightOut_12[15] , 
        \nRightOut_12[14] , \nRightOut_12[13] , \nRightOut_12[12] , 
        \nRightOut_12[11] , \nRightOut_12[10] , \nRightOut_12[9] , 
        \nRightOut_12[8] , \nRightOut_12[7] , \nRightOut_12[6] , 
        \nRightOut_12[5] , \nRightOut_12[4] , \nRightOut_12[3] , 
        \nRightOut_12[2] , \nRightOut_12[1] , \nRightOut_12[0] }), .outleft({
        \nLeftOut_28[16] , \nLeftOut_28[15] , \nLeftOut_28[14] , 
        \nLeftOut_28[13] , \nLeftOut_28[12] , \nLeftOut_28[11] , 
        \nLeftOut_28[10] , \nLeftOut_28[9] , \nLeftOut_28[8] , 
        \nLeftOut_28[7] , \nLeftOut_28[6] , \nLeftOut_28[5] , \nLeftOut_28[4] , 
        \nLeftOut_28[3] , \nLeftOut_28[2] , \nLeftOut_28[1] , \nLeftOut_28[0] 
        }), .outright({\nRightOut_28[16] , \nRightOut_28[15] , 
        \nRightOut_28[14] , \nRightOut_28[13] , \nRightOut_28[12] , 
        \nRightOut_28[11] , \nRightOut_28[10] , \nRightOut_28[9] , 
        \nRightOut_28[8] , \nRightOut_28[7] , \nRightOut_28[6] , 
        \nRightOut_28[5] , \nRightOut_28[4] , \nRightOut_28[3] , 
        \nRightOut_28[2] , \nRightOut_28[1] , \nRightOut_28[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_104 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink24[15] , \ScanLink24[14] , \ScanLink24[13] , 
        \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , \ScanLink24[9] , 
        \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , \ScanLink24[5] , 
        \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , \ScanLink24[1] , 
        \ScanLink24[0] }), .ScanOut({\ScanLink25[15] , \ScanLink25[14] , 
        \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , 
        \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , 
        \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , 
        \ScanLink25[1] , \ScanLink25[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_80[16] , \nRightOut_80[15] , \nRightOut_80[14] , 
        \nRightOut_80[13] , \nRightOut_80[12] , \nRightOut_80[11] , 
        \nRightOut_80[10] , \nRightOut_80[9] , \nRightOut_80[8] , 
        \nRightOut_80[7] , \nRightOut_80[6] , \nRightOut_80[5] , 
        \nRightOut_80[4] , \nRightOut_80[3] , \nRightOut_80[2] , 
        \nRightOut_80[1] , \nRightOut_80[0] }), .inright({\nRightOut_81[16] , 
        \nRightOut_81[15] , \nRightOut_81[14] , \nRightOut_81[13] , 
        \nRightOut_81[12] , \nRightOut_81[11] , \nRightOut_81[10] , 
        \nRightOut_81[9] , \nRightOut_81[8] , \nRightOut_81[7] , 
        \nRightOut_81[6] , \nRightOut_81[5] , \nRightOut_81[4] , 
        \nRightOut_81[3] , \nRightOut_81[2] , \nRightOut_81[1] , 
        \nRightOut_81[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_46 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_30[16] , \nLeftOut_30[15] , \nLeftOut_30[14] , 
        \nLeftOut_30[13] , \nLeftOut_30[12] , \nLeftOut_30[11] , 
        \nLeftOut_30[10] , \nLeftOut_30[9] , \nLeftOut_30[8] , 
        \nLeftOut_30[7] , \nLeftOut_30[6] , \nLeftOut_30[5] , \nLeftOut_30[4] , 
        \nLeftOut_30[3] , \nLeftOut_30[2] , \nLeftOut_30[1] , \nLeftOut_30[0] 
        }), .inright({\nLeftOut_31[16] , \nLeftOut_31[15] , \nLeftOut_31[14] , 
        \nLeftOut_31[13] , \nLeftOut_31[12] , \nLeftOut_31[11] , 
        \nLeftOut_31[10] , \nLeftOut_31[9] , \nLeftOut_31[8] , 
        \nLeftOut_31[7] , \nLeftOut_31[6] , \nLeftOut_31[5] , \nLeftOut_31[4] , 
        \nLeftOut_31[3] , \nLeftOut_31[2] , \nLeftOut_31[1] , \nLeftOut_31[0] 
        }), .outleft({\nLeftOut_46[16] , \nLeftOut_46[15] , \nLeftOut_46[14] , 
        \nLeftOut_46[13] , \nLeftOut_46[12] , \nLeftOut_46[11] , 
        \nLeftOut_46[10] , \nLeftOut_46[9] , \nLeftOut_46[8] , 
        \nLeftOut_46[7] , \nLeftOut_46[6] , \nLeftOut_46[5] , \nLeftOut_46[4] , 
        \nLeftOut_46[3] , \nLeftOut_46[2] , \nLeftOut_46[1] , \nLeftOut_46[0] 
        }), .outright({\nRightOut_46[16] , \nRightOut_46[15] , 
        \nRightOut_46[14] , \nRightOut_46[13] , \nRightOut_46[12] , 
        \nRightOut_46[11] , \nRightOut_46[10] , \nRightOut_46[9] , 
        \nRightOut_46[8] , \nRightOut_46[7] , \nRightOut_46[6] , 
        \nRightOut_46[5] , \nRightOut_46[4] , \nRightOut_46[3] , 
        \nRightOut_46[2] , \nRightOut_46[1] , \nRightOut_46[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s4_SCAN1 node_84 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_68[16] , \nLeftOut_68[15] , \nLeftOut_68[14] , 
        \nLeftOut_68[13] , \nLeftOut_68[12] , \nLeftOut_68[11] , 
        \nLeftOut_68[10] , \nLeftOut_68[9] , \nLeftOut_68[8] , 
        \nLeftOut_68[7] , \nLeftOut_68[6] , \nLeftOut_68[5] , \nLeftOut_68[4] , 
        \nLeftOut_68[3] , \nLeftOut_68[2] , \nLeftOut_68[1] , \nLeftOut_68[0] 
        }), .inright({\nLeftOut_76[16] , \nLeftOut_76[15] , \nLeftOut_76[14] , 
        \nLeftOut_76[13] , \nLeftOut_76[12] , \nLeftOut_76[11] , 
        \nLeftOut_76[10] , \nLeftOut_76[9] , \nLeftOut_76[8] , 
        \nLeftOut_76[7] , \nLeftOut_76[6] , \nLeftOut_76[5] , \nLeftOut_76[4] , 
        \nLeftOut_76[3] , \nLeftOut_76[2] , \nLeftOut_76[1] , \nLeftOut_76[0] 
        }), .outleft({\nLeftOut_84[16] , \nLeftOut_84[15] , \nLeftOut_84[14] , 
        \nLeftOut_84[13] , \nLeftOut_84[12] , \nLeftOut_84[11] , 
        \nLeftOut_84[10] , \nLeftOut_84[9] , \nLeftOut_84[8] , 
        \nLeftOut_84[7] , \nLeftOut_84[6] , \nLeftOut_84[5] , \nLeftOut_84[4] , 
        \nLeftOut_84[3] , \nLeftOut_84[2] , \nLeftOut_84[1] , \nLeftOut_84[0] 
        }), .outright({\nRightOut_84[16] , \nRightOut_84[15] , 
        \nRightOut_84[14] , \nRightOut_84[13] , \nRightOut_84[12] , 
        \nRightOut_84[11] , \nRightOut_84[10] , \nRightOut_84[9] , 
        \nRightOut_84[8] , \nRightOut_84[7] , \nRightOut_84[6] , 
        \nRightOut_84[5] , \nRightOut_84[4] , \nRightOut_84[3] , 
        \nRightOut_84[2] , \nRightOut_84[1] , \nRightOut_84[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s4_SCAN1 node_61 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_45[16] , \nLeftOut_45[15] , \nLeftOut_45[14] , 
        \nLeftOut_45[13] , \nLeftOut_45[12] , \nLeftOut_45[11] , 
        \nLeftOut_45[10] , \nLeftOut_45[9] , \nLeftOut_45[8] , 
        \nLeftOut_45[7] , \nLeftOut_45[6] , \nLeftOut_45[5] , \nLeftOut_45[4] , 
        \nLeftOut_45[3] , \nLeftOut_45[2] , \nLeftOut_45[1] , \nLeftOut_45[0] 
        }), .inright({\nLeftOut_47[16] , \nLeftOut_47[15] , \nLeftOut_47[14] , 
        \nLeftOut_47[13] , \nLeftOut_47[12] , \nLeftOut_47[11] , 
        \nLeftOut_47[10] , \nLeftOut_47[9] , \nLeftOut_47[8] , 
        \nLeftOut_47[7] , \nLeftOut_47[6] , \nLeftOut_47[5] , \nLeftOut_47[4] , 
        \nLeftOut_47[3] , \nLeftOut_47[2] , \nLeftOut_47[1] , \nLeftOut_47[0] 
        }), .outleft({\nLeftOut_61[16] , \nLeftOut_61[15] , \nLeftOut_61[14] , 
        \nLeftOut_61[13] , \nLeftOut_61[12] , \nLeftOut_61[11] , 
        \nLeftOut_61[10] , \nLeftOut_61[9] , \nLeftOut_61[8] , 
        \nLeftOut_61[7] , \nLeftOut_61[6] , \nLeftOut_61[5] , \nLeftOut_61[4] , 
        \nLeftOut_61[3] , \nLeftOut_61[2] , \nLeftOut_61[1] , \nLeftOut_61[0] 
        }), .outright({\nRightOut_61[16] , \nRightOut_61[15] , 
        \nRightOut_61[14] , \nRightOut_61[13] , \nRightOut_61[12] , 
        \nRightOut_61[11] , \nRightOut_61[10] , \nRightOut_61[9] , 
        \nRightOut_61[8] , \nRightOut_61[7] , \nRightOut_61[6] , 
        \nRightOut_61[5] , \nRightOut_61[4] , \nRightOut_61[3] , 
        \nRightOut_61[2] , \nRightOut_61[1] , \nRightOut_61[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s10_SCAN1 node_69 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_49[16] , \nRightOut_49[15] , \nRightOut_49[14] , 
        \nRightOut_49[13] , \nRightOut_49[12] , \nRightOut_49[11] , 
        \nRightOut_49[10] , \nRightOut_49[9] , \nRightOut_49[8] , 
        \nRightOut_49[7] , \nRightOut_49[6] , \nRightOut_49[5] , 
        \nRightOut_49[4] , \nRightOut_49[3] , \nRightOut_49[2] , 
        \nRightOut_49[1] , \nRightOut_49[0] }), .inright({\nRightOut_53[16] , 
        \nRightOut_53[15] , \nRightOut_53[14] , \nRightOut_53[13] , 
        \nRightOut_53[12] , \nRightOut_53[11] , \nRightOut_53[10] , 
        \nRightOut_53[9] , \nRightOut_53[8] , \nRightOut_53[7] , 
        \nRightOut_53[6] , \nRightOut_53[5] , \nRightOut_53[4] , 
        \nRightOut_53[3] , \nRightOut_53[2] , \nRightOut_53[1] , 
        \nRightOut_53[0] }), .outleft({\nLeftOut_69[16] , \nLeftOut_69[15] , 
        \nLeftOut_69[14] , \nLeftOut_69[13] , \nLeftOut_69[12] , 
        \nLeftOut_69[11] , \nLeftOut_69[10] , \nLeftOut_69[9] , 
        \nLeftOut_69[8] , \nLeftOut_69[7] , \nLeftOut_69[6] , \nLeftOut_69[5] , 
        \nLeftOut_69[4] , \nLeftOut_69[3] , \nLeftOut_69[2] , \nLeftOut_69[1] , 
        \nLeftOut_69[0] }), .outright({\nRightOut_69[16] , \nRightOut_69[15] , 
        \nRightOut_69[14] , \nRightOut_69[13] , \nRightOut_69[12] , 
        \nRightOut_69[11] , \nRightOut_69[10] , \nRightOut_69[9] , 
        \nRightOut_69[8] , \nRightOut_69[7] , \nRightOut_69[6] , 
        \nRightOut_69[5] , \nRightOut_69[4] , \nRightOut_69[3] , 
        \nRightOut_69[2] , \nRightOut_69[1] , \nRightOut_69[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s12_SCAN1 node_55 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_37[16] , \nRightOut_37[15] , \nRightOut_37[14] , 
        \nRightOut_37[13] , \nRightOut_37[12] , \nRightOut_37[11] , 
        \nRightOut_37[10] , \nRightOut_37[9] , \nRightOut_37[8] , 
        \nRightOut_37[7] , \nRightOut_37[6] , \nRightOut_37[5] , 
        \nRightOut_37[4] , \nRightOut_37[3] , \nRightOut_37[2] , 
        \nRightOut_37[1] , \nRightOut_37[0] }), .inright({\nRightOut_39[16] , 
        \nRightOut_39[15] , \nRightOut_39[14] , \nRightOut_39[13] , 
        \nRightOut_39[12] , \nRightOut_39[11] , \nRightOut_39[10] , 
        \nRightOut_39[9] , \nRightOut_39[8] , \nRightOut_39[7] , 
        \nRightOut_39[6] , \nRightOut_39[5] , \nRightOut_39[4] , 
        \nRightOut_39[3] , \nRightOut_39[2] , \nRightOut_39[1] , 
        \nRightOut_39[0] }), .outleft({\nLeftOut_55[16] , \nLeftOut_55[15] , 
        \nLeftOut_55[14] , \nLeftOut_55[13] , \nLeftOut_55[12] , 
        \nLeftOut_55[11] , \nLeftOut_55[10] , \nLeftOut_55[9] , 
        \nLeftOut_55[8] , \nLeftOut_55[7] , \nLeftOut_55[6] , \nLeftOut_55[5] , 
        \nLeftOut_55[4] , \nLeftOut_55[3] , \nLeftOut_55[2] , \nLeftOut_55[1] , 
        \nLeftOut_55[0] }), .outright({\nRightOut_55[16] , \nRightOut_55[15] , 
        \nRightOut_55[14] , \nRightOut_55[13] , \nRightOut_55[12] , 
        \nRightOut_55[11] , \nRightOut_55[10] , \nRightOut_55[9] , 
        \nRightOut_55[8] , \nRightOut_55[7] , \nRightOut_55[6] , 
        \nRightOut_55[5] , \nRightOut_55[4] , \nRightOut_55[3] , 
        \nRightOut_55[2] , \nRightOut_55[1] , \nRightOut_55[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_97 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink17[15] , \ScanLink17[14] , \ScanLink17[13] , 
        \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , \ScanLink17[9] , 
        \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , \ScanLink17[5] , 
        \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , \ScanLink17[1] , 
        \ScanLink17[0] }), .ScanOut({\ScanLink18[15] , \ScanLink18[14] , 
        \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , 
        \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , 
        \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , 
        \ScanLink18[1] , \ScanLink18[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_82[16] , \nLeftOut_82[15] , \nLeftOut_82[14] , 
        \nLeftOut_82[13] , \nLeftOut_82[12] , \nLeftOut_82[11] , 
        \nLeftOut_82[10] , \nLeftOut_82[9] , \nLeftOut_82[8] , 
        \nLeftOut_82[7] , \nLeftOut_82[6] , \nLeftOut_82[5] , \nLeftOut_82[4] , 
        \nLeftOut_82[3] , \nLeftOut_82[2] , \nLeftOut_82[1] , \nLeftOut_82[0] 
        }), .inright({\nLeftOut_83[16] , \nLeftOut_83[15] , \nLeftOut_83[14] , 
        \nLeftOut_83[13] , \nLeftOut_83[12] , \nLeftOut_83[11] , 
        \nLeftOut_83[10] , \nLeftOut_83[9] , \nLeftOut_83[8] , 
        \nLeftOut_83[7] , \nLeftOut_83[6] , \nLeftOut_83[5] , \nLeftOut_83[4] , 
        \nLeftOut_83[3] , \nLeftOut_83[2] , \nLeftOut_83[1] , \nLeftOut_83[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_15 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink15[15] , \ScanLink15[14] , \ScanLink15[13] , 
        \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , \ScanLink15[9] , 
        \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , \ScanLink15[5] , 
        \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , \ScanLink15[1] , 
        \ScanLink15[0] }), .ScanOut({\ScanLink16[15] , \ScanLink16[14] , 
        \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , 
        \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , 
        \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , 
        \ScanLink16[1] , \ScanLink16[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_15[16] , \nLeftOut_15[15] , \nLeftOut_15[14] , 
        \nLeftOut_15[13] , \nLeftOut_15[12] , \nLeftOut_15[11] , 
        \nLeftOut_15[10] , \nLeftOut_15[9] , \nLeftOut_15[8] , 
        \nLeftOut_15[7] , \nLeftOut_15[6] , \nLeftOut_15[5] , \nLeftOut_15[4] , 
        \nLeftOut_15[3] , \nLeftOut_15[2] , \nLeftOut_15[1] , \nLeftOut_15[0] 
        }), .inright({\nRightOut_15[16] , \nRightOut_15[15] , 
        \nRightOut_15[14] , \nRightOut_15[13] , \nRightOut_15[12] , 
        \nRightOut_15[11] , \nRightOut_15[10] , \nRightOut_15[9] , 
        \nRightOut_15[8] , \nRightOut_15[7] , \nRightOut_15[6] , 
        \nRightOut_15[5] , \nRightOut_15[4] , \nRightOut_15[3] , 
        \nRightOut_15[2] , \nRightOut_15[1] , \nRightOut_15[0] }), .outleft({
        \nLeftOut_15[16] , \nLeftOut_15[15] , \nLeftOut_15[14] , 
        \nLeftOut_15[13] , \nLeftOut_15[12] , \nLeftOut_15[11] , 
        \nLeftOut_15[10] , \nLeftOut_15[9] , \nLeftOut_15[8] , 
        \nLeftOut_15[7] , \nLeftOut_15[6] , \nLeftOut_15[5] , \nLeftOut_15[4] , 
        \nLeftOut_15[3] , \nLeftOut_15[2] , \nLeftOut_15[1] , \nLeftOut_15[0] 
        }), .outright({\nRightOut_15[16] , \nRightOut_15[15] , 
        \nRightOut_15[14] , \nRightOut_15[13] , \nRightOut_15[12] , 
        \nRightOut_15[11] , \nRightOut_15[10] , \nRightOut_15[9] , 
        \nRightOut_15[8] , \nRightOut_15[7] , \nRightOut_15[6] , 
        \nRightOut_15[5] , \nRightOut_15[4] , \nRightOut_15[3] , 
        \nRightOut_15[2] , \nRightOut_15[1] , \nRightOut_15[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_29 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_13[16] , \nLeftOut_13[15] , \nLeftOut_13[14] , 
        \nLeftOut_13[13] , \nLeftOut_13[12] , \nLeftOut_13[11] , 
        \nLeftOut_13[10] , \nLeftOut_13[9] , \nLeftOut_13[8] , 
        \nLeftOut_13[7] , \nLeftOut_13[6] , \nLeftOut_13[5] , \nLeftOut_13[4] , 
        \nLeftOut_13[3] , \nLeftOut_13[2] , \nLeftOut_13[1] , \nLeftOut_13[0] 
        }), .inright({\nRightOut_13[16] , \nRightOut_13[15] , 
        \nRightOut_13[14] , \nRightOut_13[13] , \nRightOut_13[12] , 
        \nRightOut_13[11] , \nRightOut_13[10] , \nRightOut_13[9] , 
        \nRightOut_13[8] , \nRightOut_13[7] , \nRightOut_13[6] , 
        \nRightOut_13[5] , \nRightOut_13[4] , \nRightOut_13[3] , 
        \nRightOut_13[2] , \nRightOut_13[1] , \nRightOut_13[0] }), .outleft({
        \nLeftOut_29[16] , \nLeftOut_29[15] , \nLeftOut_29[14] , 
        \nLeftOut_29[13] , \nLeftOut_29[12] , \nLeftOut_29[11] , 
        \nLeftOut_29[10] , \nLeftOut_29[9] , \nLeftOut_29[8] , 
        \nLeftOut_29[7] , \nLeftOut_29[6] , \nLeftOut_29[5] , \nLeftOut_29[4] , 
        \nLeftOut_29[3] , \nLeftOut_29[2] , \nLeftOut_29[1] , \nLeftOut_29[0] 
        }), .outright({\nRightOut_29[16] , \nRightOut_29[15] , 
        \nRightOut_29[14] , \nRightOut_29[13] , \nRightOut_29[12] , 
        \nRightOut_29[11] , \nRightOut_29[10] , \nRightOut_29[9] , 
        \nRightOut_29[8] , \nRightOut_29[7] , \nRightOut_29[6] , 
        \nRightOut_29[5] , \nRightOut_29[4] , \nRightOut_29[3] , 
        \nRightOut_29[2] , \nRightOut_29[1] , \nRightOut_29[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_47 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_30[16] , \nRightOut_30[15] , \nRightOut_30[14] , 
        \nRightOut_30[13] , \nRightOut_30[12] , \nRightOut_30[11] , 
        \nRightOut_30[10] , \nRightOut_30[9] , \nRightOut_30[8] , 
        \nRightOut_30[7] , \nRightOut_30[6] , \nRightOut_30[5] , 
        \nRightOut_30[4] , \nRightOut_30[3] , \nRightOut_30[2] , 
        \nRightOut_30[1] , \nRightOut_30[0] }), .inright({\nRightOut_31[16] , 
        \nRightOut_31[15] , \nRightOut_31[14] , \nRightOut_31[13] , 
        \nRightOut_31[12] , \nRightOut_31[11] , \nRightOut_31[10] , 
        \nRightOut_31[9] , \nRightOut_31[8] , \nRightOut_31[7] , 
        \nRightOut_31[6] , \nRightOut_31[5] , \nRightOut_31[4] , 
        \nRightOut_31[3] , \nRightOut_31[2] , \nRightOut_31[1] , 
        \nRightOut_31[0] }), .outleft({\nLeftOut_47[16] , \nLeftOut_47[15] , 
        \nLeftOut_47[14] , \nLeftOut_47[13] , \nLeftOut_47[12] , 
        \nLeftOut_47[11] , \nLeftOut_47[10] , \nLeftOut_47[9] , 
        \nLeftOut_47[8] , \nLeftOut_47[7] , \nLeftOut_47[6] , \nLeftOut_47[5] , 
        \nLeftOut_47[4] , \nLeftOut_47[3] , \nLeftOut_47[2] , \nLeftOut_47[1] , 
        \nLeftOut_47[0] }), .outright({\nRightOut_47[16] , \nRightOut_47[15] , 
        \nRightOut_47[14] , \nRightOut_47[13] , \nRightOut_47[12] , 
        \nRightOut_47[11] , \nRightOut_47[10] , \nRightOut_47[9] , 
        \nRightOut_47[8] , \nRightOut_47[7] , \nRightOut_47[6] , 
        \nRightOut_47[5] , \nRightOut_47[4] , \nRightOut_47[3] , 
        \nRightOut_47[2] , \nRightOut_47[1] , \nRightOut_47[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_72 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_56[16] , \nLeftOut_56[15] , \nLeftOut_56[14] , 
        \nLeftOut_56[13] , \nLeftOut_56[12] , \nLeftOut_56[11] , 
        \nLeftOut_56[10] , \nLeftOut_56[9] , \nLeftOut_56[8] , 
        \nLeftOut_56[7] , \nLeftOut_56[6] , \nLeftOut_56[5] , \nLeftOut_56[4] , 
        \nLeftOut_56[3] , \nLeftOut_56[2] , \nLeftOut_56[1] , \nLeftOut_56[0] 
        }), .inright({\nLeftOut_60[16] , \nLeftOut_60[15] , \nLeftOut_60[14] , 
        \nLeftOut_60[13] , \nLeftOut_60[12] , \nLeftOut_60[11] , 
        \nLeftOut_60[10] , \nLeftOut_60[9] , \nLeftOut_60[8] , 
        \nLeftOut_60[7] , \nLeftOut_60[6] , \nLeftOut_60[5] , \nLeftOut_60[4] , 
        \nLeftOut_60[3] , \nLeftOut_60[2] , \nLeftOut_60[1] , \nLeftOut_60[0] 
        }), .outleft({\nLeftOut_72[16] , \nLeftOut_72[15] , \nLeftOut_72[14] , 
        \nLeftOut_72[13] , \nLeftOut_72[12] , \nLeftOut_72[11] , 
        \nLeftOut_72[10] , \nLeftOut_72[9] , \nLeftOut_72[8] , 
        \nLeftOut_72[7] , \nLeftOut_72[6] , \nLeftOut_72[5] , \nLeftOut_72[4] , 
        \nLeftOut_72[3] , \nLeftOut_72[2] , \nLeftOut_72[1] , \nLeftOut_72[0] 
        }), .outright({\nRightOut_72[16] , \nRightOut_72[15] , 
        \nRightOut_72[14] , \nRightOut_72[13] , \nRightOut_72[12] , 
        \nRightOut_72[11] , \nRightOut_72[10] , \nRightOut_72[9] , 
        \nRightOut_72[8] , \nRightOut_72[7] , \nRightOut_72[6] , 
        \nRightOut_72[5] , \nRightOut_72[4] , \nRightOut_72[3] , 
        \nRightOut_72[2] , \nRightOut_72[1] , \nRightOut_72[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_60 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_44[16] , \nLeftOut_44[15] , \nLeftOut_44[14] , 
        \nLeftOut_44[13] , \nLeftOut_44[12] , \nLeftOut_44[11] , 
        \nLeftOut_44[10] , \nLeftOut_44[9] , \nLeftOut_44[8] , 
        \nLeftOut_44[7] , \nLeftOut_44[6] , \nLeftOut_44[5] , \nLeftOut_44[4] , 
        \nLeftOut_44[3] , \nLeftOut_44[2] , \nLeftOut_44[1] , \nLeftOut_44[0] 
        }), .inright({\nLeftOut_46[16] , \nLeftOut_46[15] , \nLeftOut_46[14] , 
        \nLeftOut_46[13] , \nLeftOut_46[12] , \nLeftOut_46[11] , 
        \nLeftOut_46[10] , \nLeftOut_46[9] , \nLeftOut_46[8] , 
        \nLeftOut_46[7] , \nLeftOut_46[6] , \nLeftOut_46[5] , \nLeftOut_46[4] , 
        \nLeftOut_46[3] , \nLeftOut_46[2] , \nLeftOut_46[1] , \nLeftOut_46[0] 
        }), .outleft({\nLeftOut_60[16] , \nLeftOut_60[15] , \nLeftOut_60[14] , 
        \nLeftOut_60[13] , \nLeftOut_60[12] , \nLeftOut_60[11] , 
        \nLeftOut_60[10] , \nLeftOut_60[9] , \nLeftOut_60[8] , 
        \nLeftOut_60[7] , \nLeftOut_60[6] , \nLeftOut_60[5] , \nLeftOut_60[4] , 
        \nLeftOut_60[3] , \nLeftOut_60[2] , \nLeftOut_60[1] , \nLeftOut_60[0] 
        }), .outright({\nRightOut_60[16] , \nRightOut_60[15] , 
        \nRightOut_60[14] , \nRightOut_60[13] , \nRightOut_60[12] , 
        \nRightOut_60[11] , \nRightOut_60[10] , \nRightOut_60[9] , 
        \nRightOut_60[8] , \nRightOut_60[7] , \nRightOut_60[6] , 
        \nRightOut_60[5] , \nRightOut_60[4] , \nRightOut_60[3] , 
        \nRightOut_60[2] , \nRightOut_60[1] , \nRightOut_60[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_105 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink25[15] , \ScanLink25[14] , \ScanLink25[13] , 
        \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , \ScanLink25[9] , 
        \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , \ScanLink25[5] , 
        \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , \ScanLink25[1] , 
        \ScanLink25[0] }), .ScanOut({\ScanLink26[15] , \ScanLink26[14] , 
        \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , 
        \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , 
        \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , 
        \ScanLink26[1] , \ScanLink26[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_82[16] , \nRightOut_82[15] , \nRightOut_82[14] , 
        \nRightOut_82[13] , \nRightOut_82[12] , \nRightOut_82[11] , 
        \nRightOut_82[10] , \nRightOut_82[9] , \nRightOut_82[8] , 
        \nRightOut_82[7] , \nRightOut_82[6] , \nRightOut_82[5] , 
        \nRightOut_82[4] , \nRightOut_82[3] , \nRightOut_82[2] , 
        \nRightOut_82[1] , \nRightOut_82[0] }), .inright({\nRightOut_83[16] , 
        \nRightOut_83[15] , \nRightOut_83[14] , \nRightOut_83[13] , 
        \nRightOut_83[12] , \nRightOut_83[11] , \nRightOut_83[10] , 
        \nRightOut_83[9] , \nRightOut_83[8] , \nRightOut_83[7] , 
        \nRightOut_83[6] , \nRightOut_83[5] , \nRightOut_83[4] , 
        \nRightOut_83[3] , \nRightOut_83[2] , \nRightOut_83[1] , 
        \nRightOut_83[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_32 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_16[16] , \nLeftOut_16[15] , \nLeftOut_16[14] , 
        \nLeftOut_16[13] , \nLeftOut_16[12] , \nLeftOut_16[11] , 
        \nLeftOut_16[10] , \nLeftOut_16[9] , \nLeftOut_16[8] , 
        \nLeftOut_16[7] , \nLeftOut_16[6] , \nLeftOut_16[5] , \nLeftOut_16[4] , 
        \nLeftOut_16[3] , \nLeftOut_16[2] , \nLeftOut_16[1] , \nLeftOut_16[0] 
        }), .inright({\nLeftOut_17[16] , \nLeftOut_17[15] , \nLeftOut_17[14] , 
        \nLeftOut_17[13] , \nLeftOut_17[12] , \nLeftOut_17[11] , 
        \nLeftOut_17[10] , \nLeftOut_17[9] , \nLeftOut_17[8] , 
        \nLeftOut_17[7] , \nLeftOut_17[6] , \nLeftOut_17[5] , \nLeftOut_17[4] , 
        \nLeftOut_17[3] , \nLeftOut_17[2] , \nLeftOut_17[1] , \nLeftOut_17[0] 
        }), .outleft({\nLeftOut_32[16] , \nLeftOut_32[15] , \nLeftOut_32[14] , 
        \nLeftOut_32[13] , \nLeftOut_32[12] , \nLeftOut_32[11] , 
        \nLeftOut_32[10] , \nLeftOut_32[9] , \nLeftOut_32[8] , 
        \nLeftOut_32[7] , \nLeftOut_32[6] , \nLeftOut_32[5] , \nLeftOut_32[4] , 
        \nLeftOut_32[3] , \nLeftOut_32[2] , \nLeftOut_32[1] , \nLeftOut_32[0] 
        }), .outright({\nRightOut_32[16] , \nRightOut_32[15] , 
        \nRightOut_32[14] , \nRightOut_32[13] , \nRightOut_32[12] , 
        \nRightOut_32[11] , \nRightOut_32[10] , \nRightOut_32[9] , 
        \nRightOut_32[8] , \nRightOut_32[7] , \nRightOut_32[6] , 
        \nRightOut_32[5] , \nRightOut_32[4] , \nRightOut_32[3] , 
        \nRightOut_32[2] , \nRightOut_32[1] , \nRightOut_32[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s5_SCAN1 node_85 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_69[16] , \nLeftOut_69[15] , \nLeftOut_69[14] , 
        \nLeftOut_69[13] , \nLeftOut_69[12] , \nLeftOut_69[11] , 
        \nLeftOut_69[10] , \nLeftOut_69[9] , \nLeftOut_69[8] , 
        \nLeftOut_69[7] , \nLeftOut_69[6] , \nLeftOut_69[5] , \nLeftOut_69[4] , 
        \nLeftOut_69[3] , \nLeftOut_69[2] , \nLeftOut_69[1] , \nLeftOut_69[0] 
        }), .inright({\nLeftOut_77[16] , \nLeftOut_77[15] , \nLeftOut_77[14] , 
        \nLeftOut_77[13] , \nLeftOut_77[12] , \nLeftOut_77[11] , 
        \nLeftOut_77[10] , \nLeftOut_77[9] , \nLeftOut_77[8] , 
        \nLeftOut_77[7] , \nLeftOut_77[6] , \nLeftOut_77[5] , \nLeftOut_77[4] , 
        \nLeftOut_77[3] , \nLeftOut_77[2] , \nLeftOut_77[1] , \nLeftOut_77[0] 
        }), .outleft({\nLeftOut_85[16] , \nLeftOut_85[15] , \nLeftOut_85[14] , 
        \nLeftOut_85[13] , \nLeftOut_85[12] , \nLeftOut_85[11] , 
        \nLeftOut_85[10] , \nLeftOut_85[9] , \nLeftOut_85[8] , 
        \nLeftOut_85[7] , \nLeftOut_85[6] , \nLeftOut_85[5] , \nLeftOut_85[4] , 
        \nLeftOut_85[3] , \nLeftOut_85[2] , \nLeftOut_85[1] , \nLeftOut_85[0] 
        }), .outright({\nRightOut_85[16] , \nRightOut_85[15] , 
        \nRightOut_85[14] , \nRightOut_85[13] , \nRightOut_85[12] , 
        \nRightOut_85[11] , \nRightOut_85[10] , \nRightOut_85[9] , 
        \nRightOut_85[8] , \nRightOut_85[7] , \nRightOut_85[6] , 
        \nRightOut_85[5] , \nRightOut_85[4] , \nRightOut_85[3] , 
        \nRightOut_85[2] , \nRightOut_85[1] , \nRightOut_85[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink6[15] , \ScanLink6[14] , \ScanLink6[13] , 
        \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , \ScanLink6[9] , 
        \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , \ScanLink6[5] , 
        \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , \ScanLink6[1] , 
        \ScanLink6[0] }), .ScanOut({\ScanLink7[15] , \ScanLink7[14] , 
        \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , 
        \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_6[16] , \nLeftOut_6[15] , \nLeftOut_6[14] , \nLeftOut_6[13] , 
        \nLeftOut_6[12] , \nLeftOut_6[11] , \nLeftOut_6[10] , \nLeftOut_6[9] , 
        \nLeftOut_6[8] , \nLeftOut_6[7] , \nLeftOut_6[6] , \nLeftOut_6[5] , 
        \nLeftOut_6[4] , \nLeftOut_6[3] , \nLeftOut_6[2] , \nLeftOut_6[1] , 
        \nLeftOut_6[0] }), .inright({\nRightOut_6[16] , \nRightOut_6[15] , 
        \nRightOut_6[14] , \nRightOut_6[13] , \nRightOut_6[12] , 
        \nRightOut_6[11] , \nRightOut_6[10] , \nRightOut_6[9] , 
        \nRightOut_6[8] , \nRightOut_6[7] , \nRightOut_6[6] , \nRightOut_6[5] , 
        \nRightOut_6[4] , \nRightOut_6[3] , \nRightOut_6[2] , \nRightOut_6[1] , 
        \nRightOut_6[0] }), .outleft({\nLeftOut_6[16] , \nLeftOut_6[15] , 
        \nLeftOut_6[14] , \nLeftOut_6[13] , \nLeftOut_6[12] , \nLeftOut_6[11] , 
        \nLeftOut_6[10] , \nLeftOut_6[9] , \nLeftOut_6[8] , \nLeftOut_6[7] , 
        \nLeftOut_6[6] , \nLeftOut_6[5] , \nLeftOut_6[4] , \nLeftOut_6[3] , 
        \nLeftOut_6[2] , \nLeftOut_6[1] , \nLeftOut_6[0] }), .outright({
        \nRightOut_6[16] , \nRightOut_6[15] , \nRightOut_6[14] , 
        \nRightOut_6[13] , \nRightOut_6[12] , \nRightOut_6[11] , 
        \nRightOut_6[10] , \nRightOut_6[9] , \nRightOut_6[8] , 
        \nRightOut_6[7] , \nRightOut_6[6] , \nRightOut_6[5] , \nRightOut_6[4] , 
        \nRightOut_6[3] , \nRightOut_6[2] , \nRightOut_6[1] , \nRightOut_6[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_12 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink12[15] , \ScanLink12[14] , \ScanLink12[13] , 
        \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , \ScanLink12[9] , 
        \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , \ScanLink12[5] , 
        \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , \ScanLink12[1] , 
        \ScanLink12[0] }), .ScanOut({\ScanLink13[15] , \ScanLink13[14] , 
        \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , 
        \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , 
        \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , 
        \ScanLink13[1] , \ScanLink13[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_12[16] , \nLeftOut_12[15] , \nLeftOut_12[14] , 
        \nLeftOut_12[13] , \nLeftOut_12[12] , \nLeftOut_12[11] , 
        \nLeftOut_12[10] , \nLeftOut_12[9] , \nLeftOut_12[8] , 
        \nLeftOut_12[7] , \nLeftOut_12[6] , \nLeftOut_12[5] , \nLeftOut_12[4] , 
        \nLeftOut_12[3] , \nLeftOut_12[2] , \nLeftOut_12[1] , \nLeftOut_12[0] 
        }), .inright({\nRightOut_12[16] , \nRightOut_12[15] , 
        \nRightOut_12[14] , \nRightOut_12[13] , \nRightOut_12[12] , 
        \nRightOut_12[11] , \nRightOut_12[10] , \nRightOut_12[9] , 
        \nRightOut_12[8] , \nRightOut_12[7] , \nRightOut_12[6] , 
        \nRightOut_12[5] , \nRightOut_12[4] , \nRightOut_12[3] , 
        \nRightOut_12[2] , \nRightOut_12[1] , \nRightOut_12[0] }), .outleft({
        \nLeftOut_12[16] , \nLeftOut_12[15] , \nLeftOut_12[14] , 
        \nLeftOut_12[13] , \nLeftOut_12[12] , \nLeftOut_12[11] , 
        \nLeftOut_12[10] , \nLeftOut_12[9] , \nLeftOut_12[8] , 
        \nLeftOut_12[7] , \nLeftOut_12[6] , \nLeftOut_12[5] , \nLeftOut_12[4] , 
        \nLeftOut_12[3] , \nLeftOut_12[2] , \nLeftOut_12[1] , \nLeftOut_12[0] 
        }), .outright({\nRightOut_12[16] , \nRightOut_12[15] , 
        \nRightOut_12[14] , \nRightOut_12[13] , \nRightOut_12[12] , 
        \nRightOut_12[11] , \nRightOut_12[10] , \nRightOut_12[9] , 
        \nRightOut_12[8] , \nRightOut_12[7] , \nRightOut_12[6] , 
        \nRightOut_12[5] , \nRightOut_12[4] , \nRightOut_12[3] , 
        \nRightOut_12[2] , \nRightOut_12[1] , \nRightOut_12[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_99 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink19[15] , \ScanLink19[14] , \ScanLink19[13] , 
        \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , \ScanLink19[9] , 
        \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , \ScanLink19[5] , 
        \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , \ScanLink19[1] , 
        \ScanLink19[0] }), .ScanOut({\ScanLink20[15] , \ScanLink20[14] , 
        \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , 
        \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , 
        \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , 
        \ScanLink20[1] , \ScanLink20[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_86[16] , \nLeftOut_86[15] , \nLeftOut_86[14] , 
        \nLeftOut_86[13] , \nLeftOut_86[12] , \nLeftOut_86[11] , 
        \nLeftOut_86[10] , \nLeftOut_86[9] , \nLeftOut_86[8] , 
        \nLeftOut_86[7] , \nLeftOut_86[6] , \nLeftOut_86[5] , \nLeftOut_86[4] , 
        \nLeftOut_86[3] , \nLeftOut_86[2] , \nLeftOut_86[1] , \nLeftOut_86[0] 
        }), .inright({\nLeftOut_87[16] , \nLeftOut_87[15] , \nLeftOut_87[14] , 
        \nLeftOut_87[13] , \nLeftOut_87[12] , \nLeftOut_87[11] , 
        \nLeftOut_87[10] , \nLeftOut_87[9] , \nLeftOut_87[8] , 
        \nLeftOut_87[7] , \nLeftOut_87[6] , \nLeftOut_87[5] , \nLeftOut_87[4] , 
        \nLeftOut_87[3] , \nLeftOut_87[2] , \nLeftOut_87[1] , \nLeftOut_87[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_27 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_11[16] , \nLeftOut_11[15] , \nLeftOut_11[14] , 
        \nLeftOut_11[13] , \nLeftOut_11[12] , \nLeftOut_11[11] , 
        \nLeftOut_11[10] , \nLeftOut_11[9] , \nLeftOut_11[8] , 
        \nLeftOut_11[7] , \nLeftOut_11[6] , \nLeftOut_11[5] , \nLeftOut_11[4] , 
        \nLeftOut_11[3] , \nLeftOut_11[2] , \nLeftOut_11[1] , \nLeftOut_11[0] 
        }), .inright({\nRightOut_11[16] , \nRightOut_11[15] , 
        \nRightOut_11[14] , \nRightOut_11[13] , \nRightOut_11[12] , 
        \nRightOut_11[11] , \nRightOut_11[10] , \nRightOut_11[9] , 
        \nRightOut_11[8] , \nRightOut_11[7] , \nRightOut_11[6] , 
        \nRightOut_11[5] , \nRightOut_11[4] , \nRightOut_11[3] , 
        \nRightOut_11[2] , \nRightOut_11[1] , \nRightOut_11[0] }), .outleft({
        \nLeftOut_27[16] , \nLeftOut_27[15] , \nLeftOut_27[14] , 
        \nLeftOut_27[13] , \nLeftOut_27[12] , \nLeftOut_27[11] , 
        \nLeftOut_27[10] , \nLeftOut_27[9] , \nLeftOut_27[8] , 
        \nLeftOut_27[7] , \nLeftOut_27[6] , \nLeftOut_27[5] , \nLeftOut_27[4] , 
        \nLeftOut_27[3] , \nLeftOut_27[2] , \nLeftOut_27[1] , \nLeftOut_27[0] 
        }), .outright({\nRightOut_27[16] , \nRightOut_27[15] , 
        \nRightOut_27[14] , \nRightOut_27[13] , \nRightOut_27[12] , 
        \nRightOut_27[11] , \nRightOut_27[10] , \nRightOut_27[9] , 
        \nRightOut_27[8] , \nRightOut_27[7] , \nRightOut_27[6] , 
        \nRightOut_27[5] , \nRightOut_27[4] , \nRightOut_27[3] , 
        \nRightOut_27[2] , \nRightOut_27[1] , \nRightOut_27[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s8_SCAN1 node_35 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_18[16] , \nRightOut_18[15] , \nRightOut_18[14] , 
        \nRightOut_18[13] , \nRightOut_18[12] , \nRightOut_18[11] , 
        \nRightOut_18[10] , \nRightOut_18[9] , \nRightOut_18[8] , 
        \nRightOut_18[7] , \nRightOut_18[6] , \nRightOut_18[5] , 
        \nRightOut_18[4] , \nRightOut_18[3] , \nRightOut_18[2] , 
        \nRightOut_18[1] , \nRightOut_18[0] }), .inright({\nRightOut_19[16] , 
        \nRightOut_19[15] , \nRightOut_19[14] , \nRightOut_19[13] , 
        \nRightOut_19[12] , \nRightOut_19[11] , \nRightOut_19[10] , 
        \nRightOut_19[9] , \nRightOut_19[8] , \nRightOut_19[7] , 
        \nRightOut_19[6] , \nRightOut_19[5] , \nRightOut_19[4] , 
        \nRightOut_19[3] , \nRightOut_19[2] , \nRightOut_19[1] , 
        \nRightOut_19[0] }), .outleft({\nLeftOut_35[16] , \nLeftOut_35[15] , 
        \nLeftOut_35[14] , \nLeftOut_35[13] , \nLeftOut_35[12] , 
        \nLeftOut_35[11] , \nLeftOut_35[10] , \nLeftOut_35[9] , 
        \nLeftOut_35[8] , \nLeftOut_35[7] , \nLeftOut_35[6] , \nLeftOut_35[5] , 
        \nLeftOut_35[4] , \nLeftOut_35[3] , \nLeftOut_35[2] , \nLeftOut_35[1] , 
        \nLeftOut_35[0] }), .outright({\nRightOut_35[16] , \nRightOut_35[15] , 
        \nRightOut_35[14] , \nRightOut_35[13] , \nRightOut_35[12] , 
        \nRightOut_35[11] , \nRightOut_35[10] , \nRightOut_35[9] , 
        \nRightOut_35[8] , \nRightOut_35[7] , \nRightOut_35[6] , 
        \nRightOut_35[5] , \nRightOut_35[4] , \nRightOut_35[3] , 
        \nRightOut_35[2] , \nRightOut_35[1] , \nRightOut_35[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_40 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_24[16] , \nLeftOut_24[15] , \nLeftOut_24[14] , 
        \nLeftOut_24[13] , \nLeftOut_24[12] , \nLeftOut_24[11] , 
        \nLeftOut_24[10] , \nLeftOut_24[9] , \nLeftOut_24[8] , 
        \nLeftOut_24[7] , \nLeftOut_24[6] , \nLeftOut_24[5] , \nLeftOut_24[4] , 
        \nLeftOut_24[3] , \nLeftOut_24[2] , \nLeftOut_24[1] , \nLeftOut_24[0] 
        }), .inright({\nLeftOut_25[16] , \nLeftOut_25[15] , \nLeftOut_25[14] , 
        \nLeftOut_25[13] , \nLeftOut_25[12] , \nLeftOut_25[11] , 
        \nLeftOut_25[10] , \nLeftOut_25[9] , \nLeftOut_25[8] , 
        \nLeftOut_25[7] , \nLeftOut_25[6] , \nLeftOut_25[5] , \nLeftOut_25[4] , 
        \nLeftOut_25[3] , \nLeftOut_25[2] , \nLeftOut_25[1] , \nLeftOut_25[0] 
        }), .outleft({\nLeftOut_40[16] , \nLeftOut_40[15] , \nLeftOut_40[14] , 
        \nLeftOut_40[13] , \nLeftOut_40[12] , \nLeftOut_40[11] , 
        \nLeftOut_40[10] , \nLeftOut_40[9] , \nLeftOut_40[8] , 
        \nLeftOut_40[7] , \nLeftOut_40[6] , \nLeftOut_40[5] , \nLeftOut_40[4] , 
        \nLeftOut_40[3] , \nLeftOut_40[2] , \nLeftOut_40[1] , \nLeftOut_40[0] 
        }), .outright({\nRightOut_40[16] , \nRightOut_40[15] , 
        \nRightOut_40[14] , \nRightOut_40[13] , \nRightOut_40[12] , 
        \nRightOut_40[11] , \nRightOut_40[10] , \nRightOut_40[9] , 
        \nRightOut_40[8] , \nRightOut_40[7] , \nRightOut_40[6] , 
        \nRightOut_40[5] , \nRightOut_40[4] , \nRightOut_40[3] , 
        \nRightOut_40[2] , \nRightOut_40[1] , \nRightOut_40[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s6_SCAN1 node_67 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_51[16] , \nLeftOut_51[15] , \nLeftOut_51[14] , 
        \nLeftOut_51[13] , \nLeftOut_51[12] , \nLeftOut_51[11] , 
        \nLeftOut_51[10] , \nLeftOut_51[9] , \nLeftOut_51[8] , 
        \nLeftOut_51[7] , \nLeftOut_51[6] , \nLeftOut_51[5] , \nLeftOut_51[4] , 
        \nLeftOut_51[3] , \nLeftOut_51[2] , \nLeftOut_51[1] , \nLeftOut_51[0] 
        }), .inright({\nLeftOut_55[16] , \nLeftOut_55[15] , \nLeftOut_55[14] , 
        \nLeftOut_55[13] , \nLeftOut_55[12] , \nLeftOut_55[11] , 
        \nLeftOut_55[10] , \nLeftOut_55[9] , \nLeftOut_55[8] , 
        \nLeftOut_55[7] , \nLeftOut_55[6] , \nLeftOut_55[5] , \nLeftOut_55[4] , 
        \nLeftOut_55[3] , \nLeftOut_55[2] , \nLeftOut_55[1] , \nLeftOut_55[0] 
        }), .outleft({\nLeftOut_67[16] , \nLeftOut_67[15] , \nLeftOut_67[14] , 
        \nLeftOut_67[13] , \nLeftOut_67[12] , \nLeftOut_67[11] , 
        \nLeftOut_67[10] , \nLeftOut_67[9] , \nLeftOut_67[8] , 
        \nLeftOut_67[7] , \nLeftOut_67[6] , \nLeftOut_67[5] , \nLeftOut_67[4] , 
        \nLeftOut_67[3] , \nLeftOut_67[2] , \nLeftOut_67[1] , \nLeftOut_67[0] 
        }), .outright({\nRightOut_67[16] , \nRightOut_67[15] , 
        \nRightOut_67[14] , \nRightOut_67[13] , \nRightOut_67[12] , 
        \nRightOut_67[11] , \nRightOut_67[10] , \nRightOut_67[9] , 
        \nRightOut_67[8] , \nRightOut_67[7] , \nRightOut_67[6] , 
        \nRightOut_67[5] , \nRightOut_67[4] , \nRightOut_67[3] , 
        \nRightOut_67[2] , \nRightOut_67[1] , \nRightOut_67[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s2_SCAN1 node_82 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_66[16] , \nLeftOut_66[15] , \nLeftOut_66[14] , 
        \nLeftOut_66[13] , \nLeftOut_66[12] , \nLeftOut_66[11] , 
        \nLeftOut_66[10] , \nLeftOut_66[9] , \nLeftOut_66[8] , 
        \nLeftOut_66[7] , \nLeftOut_66[6] , \nLeftOut_66[5] , \nLeftOut_66[4] , 
        \nLeftOut_66[3] , \nLeftOut_66[2] , \nLeftOut_66[1] , \nLeftOut_66[0] 
        }), .inright({\nLeftOut_74[16] , \nLeftOut_74[15] , \nLeftOut_74[14] , 
        \nLeftOut_74[13] , \nLeftOut_74[12] , \nLeftOut_74[11] , 
        \nLeftOut_74[10] , \nLeftOut_74[9] , \nLeftOut_74[8] , 
        \nLeftOut_74[7] , \nLeftOut_74[6] , \nLeftOut_74[5] , \nLeftOut_74[4] , 
        \nLeftOut_74[3] , \nLeftOut_74[2] , \nLeftOut_74[1] , \nLeftOut_74[0] 
        }), .outleft({\nLeftOut_82[16] , \nLeftOut_82[15] , \nLeftOut_82[14] , 
        \nLeftOut_82[13] , \nLeftOut_82[12] , \nLeftOut_82[11] , 
        \nLeftOut_82[10] , \nLeftOut_82[9] , \nLeftOut_82[8] , 
        \nLeftOut_82[7] , \nLeftOut_82[6] , \nLeftOut_82[5] , \nLeftOut_82[4] , 
        \nLeftOut_82[3] , \nLeftOut_82[2] , \nLeftOut_82[1] , \nLeftOut_82[0] 
        }), .outright({\nRightOut_82[16] , \nRightOut_82[15] , 
        \nRightOut_82[14] , \nRightOut_82[13] , \nRightOut_82[12] , 
        \nRightOut_82[11] , \nRightOut_82[10] , \nRightOut_82[9] , 
        \nRightOut_82[8] , \nRightOut_82[7] , \nRightOut_82[6] , 
        \nRightOut_82[5] , \nRightOut_82[4] , \nRightOut_82[3] , 
        \nRightOut_82[2] , \nRightOut_82[1] , \nRightOut_82[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_102 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink22[15] , \ScanLink22[14] , \ScanLink22[13] , 
        \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , \ScanLink22[9] , 
        \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , \ScanLink22[5] , 
        \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , \ScanLink22[1] , 
        \ScanLink22[0] }), .ScanOut({\ScanLink23[15] , \ScanLink23[14] , 
        \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , 
        \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , 
        \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , 
        \ScanLink23[1] , \ScanLink23[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_92[16] , \nLeftOut_92[15] , \nLeftOut_92[14] , 
        \nLeftOut_92[13] , \nLeftOut_92[12] , \nLeftOut_92[11] , 
        \nLeftOut_92[10] , \nLeftOut_92[9] , \nLeftOut_92[8] , 
        \nLeftOut_92[7] , \nLeftOut_92[6] , \nLeftOut_92[5] , \nLeftOut_92[4] , 
        \nLeftOut_92[3] , \nLeftOut_92[2] , \nLeftOut_92[1] , \nLeftOut_92[0] 
        }), .inright({\nLeftOut_93[16] , \nLeftOut_93[15] , \nLeftOut_93[14] , 
        \nLeftOut_93[13] , \nLeftOut_93[12] , \nLeftOut_93[11] , 
        \nLeftOut_93[10] , \nLeftOut_93[9] , \nLeftOut_93[8] , 
        \nLeftOut_93[7] , \nLeftOut_93[6] , \nLeftOut_93[5] , \nLeftOut_93[4] , 
        \nLeftOut_93[3] , \nLeftOut_93[2] , \nLeftOut_93[1] , \nLeftOut_93[0] 
        }) );
    FFT_Node_SIZE16_IDWIDTH1_s0_SCAN1 node_52 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_36[16] , \nLeftOut_36[15] , \nLeftOut_36[14] , 
        \nLeftOut_36[13] , \nLeftOut_36[12] , \nLeftOut_36[11] , 
        \nLeftOut_36[10] , \nLeftOut_36[9] , \nLeftOut_36[8] , 
        \nLeftOut_36[7] , \nLeftOut_36[6] , \nLeftOut_36[5] , \nLeftOut_36[4] , 
        \nLeftOut_36[3] , \nLeftOut_36[2] , \nLeftOut_36[1] , \nLeftOut_36[0] 
        }), .inright({\nLeftOut_38[16] , \nLeftOut_38[15] , \nLeftOut_38[14] , 
        \nLeftOut_38[13] , \nLeftOut_38[12] , \nLeftOut_38[11] , 
        \nLeftOut_38[10] , \nLeftOut_38[9] , \nLeftOut_38[8] , 
        \nLeftOut_38[7] , \nLeftOut_38[6] , \nLeftOut_38[5] , \nLeftOut_38[4] , 
        \nLeftOut_38[3] , \nLeftOut_38[2] , \nLeftOut_38[1] , \nLeftOut_38[0] 
        }), .outleft({\nLeftOut_52[16] , \nLeftOut_52[15] , \nLeftOut_52[14] , 
        \nLeftOut_52[13] , \nLeftOut_52[12] , \nLeftOut_52[11] , 
        \nLeftOut_52[10] , \nLeftOut_52[9] , \nLeftOut_52[8] , 
        \nLeftOut_52[7] , \nLeftOut_52[6] , \nLeftOut_52[5] , \nLeftOut_52[4] , 
        \nLeftOut_52[3] , \nLeftOut_52[2] , \nLeftOut_52[1] , \nLeftOut_52[0] 
        }), .outright({\nRightOut_52[16] , \nRightOut_52[15] , 
        \nRightOut_52[14] , \nRightOut_52[13] , \nRightOut_52[12] , 
        \nRightOut_52[11] , \nRightOut_52[10] , \nRightOut_52[9] , 
        \nRightOut_52[8] , \nRightOut_52[7] , \nRightOut_52[6] , 
        \nRightOut_52[5] , \nRightOut_52[4] , \nRightOut_52[3] , 
        \nRightOut_52[2] , \nRightOut_52[1] , \nRightOut_52[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s6_SCAN1 node_75 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_59[16] , \nLeftOut_59[15] , \nLeftOut_59[14] , 
        \nLeftOut_59[13] , \nLeftOut_59[12] , \nLeftOut_59[11] , 
        \nLeftOut_59[10] , \nLeftOut_59[9] , \nLeftOut_59[8] , 
        \nLeftOut_59[7] , \nLeftOut_59[6] , \nLeftOut_59[5] , \nLeftOut_59[4] , 
        \nLeftOut_59[3] , \nLeftOut_59[2] , \nLeftOut_59[1] , \nLeftOut_59[0] 
        }), .inright({\nLeftOut_63[16] , \nLeftOut_63[15] , \nLeftOut_63[14] , 
        \nLeftOut_63[13] , \nLeftOut_63[12] , \nLeftOut_63[11] , 
        \nLeftOut_63[10] , \nLeftOut_63[9] , \nLeftOut_63[8] , 
        \nLeftOut_63[7] , \nLeftOut_63[6] , \nLeftOut_63[5] , \nLeftOut_63[4] , 
        \nLeftOut_63[3] , \nLeftOut_63[2] , \nLeftOut_63[1] , \nLeftOut_63[0] 
        }), .outleft({\nLeftOut_75[16] , \nLeftOut_75[15] , \nLeftOut_75[14] , 
        \nLeftOut_75[13] , \nLeftOut_75[12] , \nLeftOut_75[11] , 
        \nLeftOut_75[10] , \nLeftOut_75[9] , \nLeftOut_75[8] , 
        \nLeftOut_75[7] , \nLeftOut_75[6] , \nLeftOut_75[5] , \nLeftOut_75[4] , 
        \nLeftOut_75[3] , \nLeftOut_75[2] , \nLeftOut_75[1] , \nLeftOut_75[0] 
        }), .outright({\nRightOut_75[16] , \nRightOut_75[15] , 
        \nRightOut_75[14] , \nRightOut_75[13] , \nRightOut_75[12] , 
        \nRightOut_75[11] , \nRightOut_75[10] , \nRightOut_75[9] , 
        \nRightOut_75[8] , \nRightOut_75[7] , \nRightOut_75[6] , 
        \nRightOut_75[5] , \nRightOut_75[4] , \nRightOut_75[3] , 
        \nRightOut_75[2] , \nRightOut_75[1] , \nRightOut_75[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s10_SCAN1 node_90 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_66[16] , \nRightOut_66[15] , \nRightOut_66[14] , 
        \nRightOut_66[13] , \nRightOut_66[12] , \nRightOut_66[11] , 
        \nRightOut_66[10] , \nRightOut_66[9] , \nRightOut_66[8] , 
        \nRightOut_66[7] , \nRightOut_66[6] , \nRightOut_66[5] , 
        \nRightOut_66[4] , \nRightOut_66[3] , \nRightOut_66[2] , 
        \nRightOut_66[1] , \nRightOut_66[0] }), .inright({\nRightOut_74[16] , 
        \nRightOut_74[15] , \nRightOut_74[14] , \nRightOut_74[13] , 
        \nRightOut_74[12] , \nRightOut_74[11] , \nRightOut_74[10] , 
        \nRightOut_74[9] , \nRightOut_74[8] , \nRightOut_74[7] , 
        \nRightOut_74[6] , \nRightOut_74[5] , \nRightOut_74[4] , 
        \nRightOut_74[3] , \nRightOut_74[2] , \nRightOut_74[1] , 
        \nRightOut_74[0] }), .outleft({\nLeftOut_90[16] , \nLeftOut_90[15] , 
        \nLeftOut_90[14] , \nLeftOut_90[13] , \nLeftOut_90[12] , 
        \nLeftOut_90[11] , \nLeftOut_90[10] , \nLeftOut_90[9] , 
        \nLeftOut_90[8] , \nLeftOut_90[7] , \nLeftOut_90[6] , \nLeftOut_90[5] , 
        \nLeftOut_90[4] , \nLeftOut_90[3] , \nLeftOut_90[2] , \nLeftOut_90[1] , 
        \nLeftOut_90[0] }), .outright({\nRightOut_90[16] , \nRightOut_90[15] , 
        \nRightOut_90[14] , \nRightOut_90[13] , \nRightOut_90[12] , 
        \nRightOut_90[11] , \nRightOut_90[10] , \nRightOut_90[9] , 
        \nRightOut_90[8] , \nRightOut_90[7] , \nRightOut_90[6] , 
        \nRightOut_90[5] , \nRightOut_90[4] , \nRightOut_90[3] , 
        \nRightOut_90[2] , \nRightOut_90[1] , \nRightOut_90[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s33_SCAN1 node_110 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink30[15] , \ScanLink30[14] , \ScanLink30[13] , 
        \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , \ScanLink30[9] , 
        \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , \ScanLink30[5] , 
        \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , \ScanLink30[1] , 
        \ScanLink30[0] }), .ScanOut({\ScanLink31[15] , \ScanLink31[14] , 
        \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , 
        \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , 
        \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , 
        \ScanLink31[1] , \ScanLink31[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_92[16] , \nRightOut_92[15] , \nRightOut_92[14] , 
        \nRightOut_92[13] , \nRightOut_92[12] , \nRightOut_92[11] , 
        \nRightOut_92[10] , \nRightOut_92[9] , \nRightOut_92[8] , 
        \nRightOut_92[7] , \nRightOut_92[6] , \nRightOut_92[5] , 
        \nRightOut_92[4] , \nRightOut_92[3] , \nRightOut_92[2] , 
        \nRightOut_92[1] , \nRightOut_92[0] }), .inright({\nRightOut_93[16] , 
        \nRightOut_93[15] , \nRightOut_93[14] , \nRightOut_93[13] , 
        \nRightOut_93[12] , \nRightOut_93[11] , \nRightOut_93[10] , 
        \nRightOut_93[9] , \nRightOut_93[8] , \nRightOut_93[7] , 
        \nRightOut_93[6] , \nRightOut_93[5] , \nRightOut_93[4] , 
        \nRightOut_93[3] , \nRightOut_93[2] , \nRightOut_93[1] , 
        \nRightOut_93[0] }) );
    FFT_Node_SIZE16_IDWIDTH1_s4_SCAN1 node_49 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), .Idl(1'b0), 
        .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_33[16] , \nLeftOut_33[15] , \nLeftOut_33[14] , 
        \nLeftOut_33[13] , \nLeftOut_33[12] , \nLeftOut_33[11] , 
        \nLeftOut_33[10] , \nLeftOut_33[9] , \nLeftOut_33[8] , 
        \nLeftOut_33[7] , \nLeftOut_33[6] , \nLeftOut_33[5] , \nLeftOut_33[4] , 
        \nLeftOut_33[3] , \nLeftOut_33[2] , \nLeftOut_33[1] , \nLeftOut_33[0] 
        }), .inright({\nLeftOut_35[16] , \nLeftOut_35[15] , \nLeftOut_35[14] , 
        \nLeftOut_35[13] , \nLeftOut_35[12] , \nLeftOut_35[11] , 
        \nLeftOut_35[10] , \nLeftOut_35[9] , \nLeftOut_35[8] , 
        \nLeftOut_35[7] , \nLeftOut_35[6] , \nLeftOut_35[5] , \nLeftOut_35[4] , 
        \nLeftOut_35[3] , \nLeftOut_35[2] , \nLeftOut_35[1] , \nLeftOut_35[0] 
        }), .outleft({\nLeftOut_49[16] , \nLeftOut_49[15] , \nLeftOut_49[14] , 
        \nLeftOut_49[13] , \nLeftOut_49[12] , \nLeftOut_49[11] , 
        \nLeftOut_49[10] , \nLeftOut_49[9] , \nLeftOut_49[8] , 
        \nLeftOut_49[7] , \nLeftOut_49[6] , \nLeftOut_49[5] , \nLeftOut_49[4] , 
        \nLeftOut_49[3] , \nLeftOut_49[2] , \nLeftOut_49[1] , \nLeftOut_49[0] 
        }), .outright({\nRightOut_49[16] , \nRightOut_49[15] , 
        \nRightOut_49[14] , \nRightOut_49[13] , \nRightOut_49[12] , 
        \nRightOut_49[11] , \nRightOut_49[10] , \nRightOut_49[9] , 
        \nRightOut_49[8] , \nRightOut_49[7] , \nRightOut_49[6] , 
        \nRightOut_49[5] , \nRightOut_49[4] , \nRightOut_49[3] , 
        \nRightOut_49[2] , \nRightOut_49[1] , \nRightOut_49[0] }) );
endmodule

