
module IntMatMul_Control_pVectorSize8_pWordSize8_pScan1_DW01_cmp2_15_0 ( A, B, 
    LEQ, TC, LT_LE, GE_GT );
input  [14:0] A;
input  [14:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17;
    VMW_NOR5 U3 ( .A(n15), .B(n16), .C(A[3]), .D(A[5]), .E(A[4]), .Z(LT_LE) );
    VMW_OR4 U5 ( .A(A[11]), .B(A[10]), .C(A[9]), .D(n17), .Z(n15) );
    VMW_OR3 U6 ( .A(A[8]), .B(A[7]), .C(A[6]), .Z(n16) );
    VMW_OR3 U4 ( .A(A[14]), .B(A[13]), .C(A[12]), .Z(n17) );
endmodule


module IntMatMul_Control_pVectorSize8_pWordSize8_pScan1 ( Clk, Reset, RD, WR, 
    Addr, DataIn, DataOut, vectorInput, matrixInput, cOutput );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
output [63:0] vectorInput;
input  [63:0] cOutput;
output [511:0] matrixInput;
input  Clk, Reset, RD, WR;
    wire n9673, n9768, n9886, n9916, n10150, n10260, n10247, n10177, n9931, 
        n10229, n10089, n10119, n9978, n9696, n9706, n10332, n9844, n10192, 
        n10002, n10025, n9863, n10315, n9721, n10285, n9754, n10347, n10329, 
        n9878, n10189, n10019, n10215, n9963, n10125, n9944, n10102, n9796, 
        n10092, n10232, n9773, n9831, n10077, n9761, n9816, n9986, \holder[0] , 
        n10050, n9823, n10065, n9746, n9994, n10269, n9804, n10042, n9938, 
        n10159, n10207, n9971, n10137, n9956, n10080, n10110, n10220, n9784, 
        n9728, Logic11, n9684, n10320, n10297, n9714, n10180, n9856, n10010, 
        n9871, \holder[4] , n10037, n10307, n9733, n10349, n9894, n9904, 
        n10142, n10272, n10255, n9923, n10165, n10059, n9838, n9924, n10162, 
        n10252, n10275, n10145, n9893, n9903, n10079, n9683, n10290, n10300, 
        n9818, n9988, n9734, n9876, n10030, \holder[6] , n10187, n9851, n10017, 
        n9713, n10327, n9698, n10227, n9783, n9798, n9951, n10087, n10117, 
        n9976, n10130, n10200, n9708, n9741, n9803, n9993, n10045, n9766, 
        n9824, n10062, n9888, n9918, n10249, n10179, n9753, n9811, n9981, 
        n10057, n9691, n10299, n10340, n9774, n9836, \holder[2] , n9858, 
        n10070, n10039, n10309, n10235, n9791, n9943, n10095, n10105, n10282, 
        n9964, n10122, n10212, n10209, n10139, n9958, n10312, n9864, n9726, 
        n10022, n10195, n10005, n9843, n10335, n9701, n9748, n9674, n9936, 
        n10170, n10240, n10267, n9881, n9911, n10157, n9992, n10044, n9802, 
        n9740, n9767, n9825, n9889, n9919, n10063, n10248, n9699, n10178, 
        n10226, n9782, n9950, n10086, n10116, n9977, n10131, n10201, n9709, 
        n9682, n10291, n9735, n10301, n10186, n9850, n9877, n10016, n10031, 
        n10326, n9712, n9799, n9749, n10348, n9925, n10163, n10253, n10274, 
        n9902, n9892, n10144, n10078, n9819, n9989, n9675, n9937, n10171, 
        n10241, n10208, n9880, n10266, n9910, n10156, n10138, n9959, n10283, 
        n10313, n9865, n10023, n9727, n9842, n10194, n10004, n9690, n9700, 
        n10334, n9859, n10298, n10308, n10038, n10234, n9790, n10104, n9942, 
        n9965, n10094, n10123, n10213, n9752, n9810, n9980, n10056, n10341, 
        n9775, n9837, n10071, n9830, n10076, n9755, n10346, n9772, n9697, 
        n9817, n9987, n10051, n9879, n10328, n10188, n10018, n10214, n10124, 
        n9962, n9945, n10093, n10103, n9797, n10233, n10228, n9979, n10088, 
        n10118, n10333, n9707, n10003, n10193, n9845, n9862, n10024, n10284, 
        n9720, n10314, n9769, n9887, n9917, n10151, n10261, n9672, n9685, 
        n9895, n9930, n10246, n10176, n10143, n9905, n10273, n10254, n10321, 
        n9839, n9922, n10058, n10164, n9715, n10296, n10306, n10181, n9857, 
        n10011, n9870, n10036, n9732, n10206, n9957, n9970, n10081, n10111, 
        n10136, n10221, n9785, n9760, n9729, n9822, n10064, n9747, n9695, 
        n9805, n10268, n9939, n9995, n10043, n10158, n10244, n9932, n10174, 
        n10331, n10286, n9885, n9915, n10153, n10263, n9829, n9860, n10048, 
        n10026, n10316, n9722, n9705, n10191, n10001, n9847, n9947, n10091, 
        n10101, n10216, n9795, n10231, n9960, n10126, n9739, n9757, n10344, 
        n9985, n10053, n9815, n9832, n10074, n10278, n9770, n9929, n10148, 
        n9745, n9679, n9762, n9807, n9997, n10041, n9820, n10066, n10198, 
        n10008, n10338, n9869, n10113, n10083, n9955, n10223, n9787, n10204, 
        n9972, n10134, n9969, n9759, n9687, n10238, n10098, n10108, n10034, 
        n9872, n10294, n10304, n9730, n9717, n164, n10323, n10183, n9855, 
        n10013, n9779, n9897, n9920, n10256, n10141, n10166, n9907, n10271, 
        n10276, n9680, n9890, n9900, n10146, n9927, n10161, n10218, n9949, 
        n10251, n10128, n10014, n10324, n10184, n9852, n10288, n10293, n9710, 
        n10303, n9737, n9875, n10028, n10033, n10318, n9849, n10133, n10203, 
        n9975, n10224, n9780, n9952, n10084, n10114, n9765, n9827, n10061, 
        n9742, n9800, n9990, n10046, n9750, n10343, n9777, n10073, n9835, 
        n9812, n9982, n10054, n9689, n10258, n10168, n9899, n9909, n9967, 
        n10121, n10211, n9792, n10236, n9940, n10106, n10096, n9719, n9692, 
        n9702, n10196, n9840, n10006, n10281, n10336, n10311, n9725, n9867, 
        n10021, n9743, n9764, n9677, n9789, n10264, n9882, n10154, n9912, 
        n9935, n10173, n9809, n10243, n9999, n10068, n9826, n10060, 
        \holder[3] , n9801, n9991, n10047, n10289, n10319, n10029, n9848, 
        n9974, n10132, n10202, n10225, n9781, n9948, n9953, n10085, n10115, 
        n9758, n9681, n10219, n10129, n10185, n9853, n10015, n10325, n9711, 
        n10292, n10302, n10032, n9736, n9874, n9676, n10277, n9891, n10147, 
        n9901, n9926, n10160, n10250, n10265, n9913, n9883, n10155, n10172, 
        n9934, n9693, n10242, n9808, n9998, n10197, n10007, n10069, n9841, 
        n9703, n10280, n10337, n9724, n10310, n9866, \holder[7] , n10020, 
        n9788, n9966, n10120, n10210, n9793, n10237, n9941, n10097, n10107, 
        n9751, n9688, n10342, n9776, n9718, n9834, n10072, n10055, n9813, 
        n9983, n9756, n10259, n9898, n9908, n10169, n10345, n9814, n9984, 
        n10052, n9833, n10075, n10279, n9771, n10149, n9928, n9946, n10100, 
        n10090, n9794, n10230, n10217, n9961, n10127, Logic01, n9694, n9704, 
        n10287, n10317, n9861, n10027, n9738, n10330, n9723, n10190, n9846, 
        n10000, \holder[5] , n9671, n10245, n9933, n10175, n9884, n10152, 
        n9914, n10262, n9828, n10049, n9778, n9686, n10257, n9921, n10167, 
        n9896, n9906, n10140, n10270, n10239, n9968, n9873, n10099, n10109, 
        n10295, n10035, n9731, n10305, n10339, n10322, n9716, n10012, n10182, 
        n9854, n10199, n10009, n9868, n9954, n10082, n10112, n10222, n9786, 
        n10205, n10135, n9973, n9744, n9678, n9806, n9996, n10040, \holder[1] , 
        n9821, n10067, n9763;
    tri \DataOut[31] , \DataOut[27]1 , \DataOut[14]1 , \DataOut[26]1 , 
        \DataOut[15]1 , \DataOut[18]1 , \DataOut[0]1 , \DataOut[19]1 , 
        \DataOut[1]1 , \DataOut[23]1 , \DataOut[22]1 , \DataOut[11]1 , 
        \DataOut[10]1 , \DataOut[9]1 , \DataOut[8]1 , \DataOut[5]1 , 
        \DataOut[4]1 , \DataOut[21]1 , \DataOut[20]1 , \DataOut[13]1 , 
        \DataOut[12]1 , \DataOut[7]1 , \DataOut[6]1 , \DataOut[25]1 , 
        \DataOut[16]1 , \DataOut[24]1 , \DataOut[17]1 , \DataOut[29]1 , 
        \DataOut[30]1 , \DataOut[2]1 , \DataOut[28]1 , \DataOut[3]1 ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 ;
    assign DataOut[31] = \DataOut[31] ;
    assign DataOut[30] = \DataOut[30]1 ;
    assign DataOut[29] = \DataOut[29]1 ;
    assign DataOut[28] = \DataOut[28]1 ;
    assign DataOut[27] = \DataOut[27]1 ;
    assign DataOut[26] = \DataOut[26]1 ;
    assign DataOut[25] = \DataOut[25]1 ;
    assign DataOut[24] = \DataOut[24]1 ;
    assign DataOut[23] = \DataOut[23]1 ;
    assign DataOut[22] = \DataOut[22]1 ;
    assign DataOut[21] = \DataOut[21]1 ;
    assign DataOut[20] = \DataOut[20]1 ;
    assign DataOut[19] = \DataOut[19]1 ;
    assign DataOut[18] = \DataOut[18]1 ;
    assign DataOut[17] = \DataOut[17]1 ;
    assign DataOut[16] = \DataOut[16]1 ;
    assign DataOut[15] = \DataOut[15]1 ;
    assign DataOut[14] = \DataOut[14]1 ;
    assign DataOut[13] = \DataOut[13]1 ;
    assign DataOut[12] = \DataOut[12]1 ;
    assign DataOut[11] = \DataOut[11]1 ;
    assign DataOut[10] = \DataOut[10]1 ;
    assign DataOut[9] = \DataOut[9]1 ;
    assign DataOut[8] = \DataOut[8]1 ;
    assign DataOut[7] = \DataOut[7]1 ;
    assign DataOut[6] = \DataOut[6]1 ;
    assign DataOut[5] = \DataOut[5]1 ;
    assign DataOut[4] = \DataOut[4]1 ;
    assign DataOut[3] = \DataOut[3]1 ;
    assign DataOut[2] = \DataOut[2]1 ;
    assign DataOut[1] = \DataOut[1]1 ;
    assign DataOut[0] = \DataOut[0]1 ;
    VMW_PULLDOWN U256 ( .Z(n9754) );
    VMW_AO22 U338 ( .A(vectorInput[27]), .B(n9706), .C(vectorInput[19]), .D(
        n9696), .Z(n10321) );
    VMW_AO22 U394 ( .A(matrixInput[67]), .B(n9707), .C(matrixInput[59]), .D(
        n9697), .Z(n10217) );
    VMW_AO22 U415 ( .A(matrixInput[508]), .B(n9707), .C(matrixInput[500]), .D(
        n9697), .Z(n9776) );
    VMW_AO22 U432 ( .A(matrixInput[494]), .B(n9707), .C(matrixInput[486]), .D(
        n9697), .Z(n9790) );
    VMW_FD \matrixInput_reg[3]  ( .D(n10273), .CP(Clk), .Q(matrixInput[3]) );
    VMW_AO22 U692 ( .A(matrixInput[259]), .B(n9707), .C(matrixInput[251]), .D(
        n9697), .Z(n10025) );
    VMW_AO22 U840 ( .A(matrixInput[126]), .B(n9707), .C(matrixInput[118]), .D(
        n9697), .Z(n10158) );
    VMW_AO22 U702 ( .A(matrixInput[250]), .B(n9707), .C(matrixInput[242]), .D(
        n9697), .Z(n10034) );
    VMW_AO22 U725 ( .A(matrixInput[229]), .B(n9707), .C(matrixInput[221]), .D(
        n9697), .Z(n10055) );
    VMW_FD \vectorInput_reg[59]  ( .D(n10281), .CP(Clk), .Q(vectorInput[59])
         );
    VMW_FD \vectorInput_reg[40]  ( .D(n10300), .CP(Clk), .Q(vectorInput[40])
         );
    VMW_AO22 U529 ( .A(matrixInput[407]), .B(n9707), .C(matrixInput[399]), .D(
        n9697), .Z(n9877) );
    VMW_AO22 U585 ( .A(matrixInput[356]), .B(n9707), .C(matrixInput[348]), .D(
        n9697), .Z(n9928) );
    VMW_AO22 U867 ( .A(cOutput[46]), .B(n9699), .C(cOutput[14]), .D(n9698), 
        .Z(n9714) );
    VMW_AO22 U356 ( .A(matrixInput[101]), .B(n9707), .C(matrixInput[93]), .D(
        n9697), .Z(n10183) );
    VMW_AO22 U371 ( .A(matrixInput[15]), .B(n9707), .C(matrixInput[7]), .D(
        n9697), .Z(n10269) );
    VMW_AO22 U560 ( .A(matrixInput[378]), .B(n9707), .C(matrixInput[370]), .D(
        n9697), .Z(n9906) );
    VMW_AO22 U619 ( .A(matrixInput[325]), .B(n9707), .C(matrixInput[317]), .D(
        n9697), .Z(n9959) );
    VMW_AO22 U650 ( .A(matrixInput[36]), .B(n9707), .C(matrixInput[28]), .D(
        n9697), .Z(n10248) );
    VMW_AO22 U789 ( .A(matrixInput[172]), .B(n9707), .C(matrixInput[164]), .D(
        n9697), .Z(n10112) );
    VMW_FD \matrixInput_reg[370]  ( .D(n9906), .CP(Clk), .Q(matrixInput[370])
         );
    VMW_FD \matrixInput_reg[369]  ( .D(n9907), .CP(Clk), .Q(matrixInput[369])
         );
    VMW_FD \matrixInput_reg[343]  ( .D(n9933), .CP(Clk), .Q(matrixInput[343])
         );
    VMW_FD \matrixInput_reg[11]  ( .D(n10265), .CP(Clk), .Q(matrixInput[11])
         );
    VMW_AO22 U882 ( .A(cOutput[50]), .B(n9702), .C(cOutput[18]), .D(n9701), 
        .Z(n9729) );
    VMW_INV U912 ( .A(n9697), .Z(n9707) );
    VMW_FD \matrixInput_reg[22]  ( .D(n10254), .CP(Clk), .Q(matrixInput[22])
         );
    VMW_AO22 U447 ( .A(matrixInput[480]), .B(n9707), .C(matrixInput[472]), .D(
        n9697), .Z(n9804) );
    VMW_AO22 U547 ( .A(matrixInput[390]), .B(n9707), .C(matrixInput[382]), .D(
        n9697), .Z(n9894) );
    VMW_AO22 U677 ( .A(matrixInput[273]), .B(n9707), .C(matrixInput[265]), .D(
        n9697), .Z(n10011) );
    VMW_BUFIZ U935 ( .A(n9750), .E(RD), .Z(\DataOut[21]1 ) );
    VMW_AO22 U777 ( .A(matrixInput[183]), .B(n9707), .C(matrixInput[175]), .D(
        n9697), .Z(n10101) );
    VMW_AO22 U809 ( .A(matrixInput[154]), .B(n9707), .C(matrixInput[146]), .D(
        n9697), .Z(n10130) );
    VMW_FD \matrixInput_reg[232]  ( .D(n10044), .CP(Clk), .Q(matrixInput[232])
         );
    VMW_FD \matrixInput_reg[218]  ( .D(n10058), .CP(Clk), .Q(matrixInput[218])
         );
    VMW_FD \matrixInput_reg[201]  ( .D(n10075), .CP(Clk), .Q(matrixInput[201])
         );
    VMW_FD \matrixInput_reg[102]  ( .D(n10174), .CP(Clk), .Q(matrixInput[102])
         );
    VMW_FD \matrixInput_reg[425]  ( .D(n9851), .CP(Clk), .Q(matrixInput[425])
         );
    VMW_FD \matrixInput_reg[416]  ( .D(n9860), .CP(Clk), .Q(matrixInput[416])
         );
    VMW_FD \matrixInput_reg[131]  ( .D(n10145), .CP(Clk), .Q(matrixInput[131])
         );
    VMW_FD \matrixInput_reg[128]  ( .D(n10148), .CP(Clk), .Q(matrixInput[128])
         );
    VMW_FD \matrixInput_reg[391]  ( .D(n9885), .CP(Clk), .Q(matrixInput[391])
         );
    VMW_FD \matrixInput_reg[388]  ( .D(n9888), .CP(Clk), .Q(matrixInput[388])
         );
    VMW_FD \vectorInput_reg[5]  ( .D(n10335), .CP(Clk), .Q(vectorInput[5]) );
    VMW_OAI211 U271 ( .A(n9671), .B(n9675), .C(n9676), .D(n9677), .Z(n10347)
         );
    VMW_AO22 U835 ( .A(matrixInput[130]), .B(n9707), .C(matrixInput[122]), .D(
        n9697), .Z(n10154) );
    VMW_AO22 U294 ( .A(DataIn[3]), .B(n9706), .C(vectorInput[59]), .D(n9696), 
        .Z(n10281) );
    VMW_AO22 U304 ( .A(vectorInput[12]), .B(n9706), .C(vectorInput[4]), .D(
        n9696), .Z(n10336) );
    VMW_AO22 U460 ( .A(matrixInput[468]), .B(n9707), .C(matrixInput[460]), .D(
        n9697), .Z(n9816) );
    VMW_AO22 U485 ( .A(matrixInput[446]), .B(n9707), .C(matrixInput[438]), .D(
        n9697), .Z(n9838) );
    VMW_AO22 U750 ( .A(matrixInput[27]), .B(n9707), .C(matrixInput[19]), .D(
        n9697), .Z(n10257) );
    VMW_AO22 U812 ( .A(matrixInput[151]), .B(n9707), .C(matrixInput[143]), .D(
        n9697), .Z(n10133) );
    VMW_FD \matrixInput_reg[32]  ( .D(n10244), .CP(Clk), .Q(matrixInput[32])
         );
    VMW_FD \matrixInput_reg[18]  ( .D(n10258), .CP(Clk), .Q(matrixInput[18])
         );
    VMW_OAI21 U899 ( .A(n9716), .B(n9717), .C(n9703), .Z(n9689) );
    VMW_OAI21 U909 ( .A(n9736), .B(n9737), .C(n9703), .Z(n9674) );
    VMW_FD \matrixInput_reg[435]  ( .D(n9841), .CP(Clk), .Q(matrixInput[435])
         );
    VMW_FD \matrixInput_reg[406]  ( .D(n9870), .CP(Clk), .Q(matrixInput[406])
         );
    VMW_FD \matrixInput_reg[398]  ( .D(n9878), .CP(Clk), .Q(matrixInput[398])
         );
    VMW_FD \matrixInput_reg[381]  ( .D(n9895), .CP(Clk), .Q(matrixInput[381])
         );
    VMW_FD \matrixInput_reg[222]  ( .D(n10054), .CP(Clk), .Q(matrixInput[222])
         );
    VMW_FD \matrixInput_reg[211]  ( .D(n10065), .CP(Clk), .Q(matrixInput[211])
         );
    VMW_FD \matrixInput_reg[208]  ( .D(n10068), .CP(Clk), .Q(matrixInput[208])
         );
    VMW_FD \matrixInput_reg[138]  ( .D(n10138), .CP(Clk), .Q(matrixInput[138])
         );
    VMW_FD \matrixInput_reg[121]  ( .D(n10155), .CP(Clk), .Q(matrixInput[121])
         );
    VMW_FD \matrixInput_reg[112]  ( .D(n10164), .CP(Clk), .Q(matrixInput[112])
         );
    VMW_FD \vectorInput_reg[63]  ( .D(n10277), .CP(Clk), .Q(vectorInput[63])
         );
    VMW_AO22 U515 ( .A(matrixInput[418]), .B(n9707), .C(matrixInput[410]), .D(
        n9697), .Z(n9866) );
    VMW_AO22 U323 ( .A(vectorInput[40]), .B(n9706), .C(vectorInput[32]), .D(
        n9696), .Z(n10308) );
    VMW_AO22 U532 ( .A(matrixInput[404]), .B(n9707), .C(matrixInput[396]), .D(
        n9697), .Z(n9880) );
    VMW_AO22 U602 ( .A(matrixInput[340]), .B(n9707), .C(matrixInput[332]), .D(
        n9697), .Z(n9944) );
    VMW_AO22 U625 ( .A(matrixInput[319]), .B(n9707), .C(matrixInput[311]), .D(
        n9697), .Z(n9965) );
    VMW_FD \vectorInput_reg[50]  ( .D(n10290), .CP(Clk), .Q(vectorInput[50])
         );
    VMW_FD \vectorInput_reg[49]  ( .D(n10291), .CP(Clk), .Q(vectorInput[49])
         );
    VMW_AO22 U792 ( .A(matrixInput[169]), .B(n9707), .C(matrixInput[161]), .D(
        n9697), .Z(n10115) );
    VMW_AO22 U429 ( .A(matrixInput[497]), .B(n9707), .C(matrixInput[489]), .D(
        n9697), .Z(n9787) );
    VMW_AO22 U689 ( .A(matrixInput[262]), .B(n9707), .C(matrixInput[254]), .D(
        n9697), .Z(n10022) );
    VMW_BUFIZ U940 ( .A(n9753), .E(RD), .Z(\DataOut[13]1 ) );
    VMW_FD \matrixInput_reg[379]  ( .D(n9897), .CP(Clk), .Q(matrixInput[379])
         );
    VMW_FD \matrixInput_reg[360]  ( .D(n9916), .CP(Clk), .Q(matrixInput[360])
         );
    VMW_FD \matrixInput_reg[353]  ( .D(n9923), .CP(Clk), .Q(matrixInput[353])
         );
    VMW_AO22 U719 ( .A(matrixInput[235]), .B(n9707), .C(matrixInput[227]), .D(
        n9697), .Z(n10049) );
    VMW_FD \matrixInput_reg[438]  ( .D(n9838), .CP(Clk), .Q(matrixInput[438])
         );
    VMW_FD \matrixInput_reg[412]  ( .D(n9864), .CP(Clk), .Q(matrixInput[412])
         );
    VMW_FD \matrixInput_reg[395]  ( .D(n9881), .CP(Clk), .Q(matrixInput[395])
         );
    VMW_FD \vectorInput_reg[1]  ( .D(n10339), .CP(Clk), .Q(vectorInput[1]) );
    VMW_FD \matrixInput_reg[421]  ( .D(n9855), .CP(Clk), .Q(matrixInput[421])
         );
    VMW_PULLDOWN U243 ( .Z(n9741) );
    VMW_PULLDOWN U244 ( .Z(n9742) );
    VMW_AO22 U286 ( .A(vectorInput[16]), .B(n9706), .C(vectorInput[8]), .D(
        n9696), .Z(n10332) );
    VMW_AO22 U507 ( .A(matrixInput[426]), .B(n9707), .C(matrixInput[418]), .D(
        n9697), .Z(n9858) );
    VMW_AO22 U849 ( .A(matrixInput[18]), .B(n9707), .C(matrixInput[10]), .D(
        n9697), .Z(n10266) );
    VMW_FD \matrixInput_reg[205]  ( .D(n10071), .CP(Clk), .Q(matrixInput[205])
         );
    VMW_FD \matrixInput_reg[106]  ( .D(n10170), .CP(Clk), .Q(matrixInput[106])
         );
    VMW_FD \matrixInput_reg[135]  ( .D(n10141), .CP(Clk), .Q(matrixInput[135])
         );
    VMW_FD \matrixInput_reg[236]  ( .D(n10040), .CP(Clk), .Q(matrixInput[236])
         );
    VMW_AO22 U316 ( .A(vectorInput[47]), .B(n9706), .C(vectorInput[39]), .D(
        n9696), .Z(n10301) );
    VMW_AO22 U497 ( .A(matrixInput[435]), .B(n9707), .C(matrixInput[427]), .D(
        n9697), .Z(n9849) );
    VMW_AO22 U331 ( .A(vectorInput[33]), .B(n9706), .C(vectorInput[25]), .D(
        n9696), .Z(n10315) );
    VMW_AO22 U610 ( .A(matrixInput[333]), .B(n9707), .C(matrixInput[325]), .D(
        n9697), .Z(n9951) );
    VMW_AO22 U637 ( .A(matrixInput[308]), .B(n9707), .C(matrixInput[300]), .D(
        n9697), .Z(n9976) );
    VMW_AO22 U780 ( .A(matrixInput[180]), .B(n9707), .C(matrixInput[172]), .D(
        n9697), .Z(n10104) );
    VMW_BUFIZ U952 ( .A(n9762), .E(RD), .Z(\DataOut[18]1 ) );
    VMW_FD \matrixInput_reg[26]  ( .D(n10250), .CP(Clk), .Q(matrixInput[26])
         );
    VMW_FD \matrixInput_reg[15]  ( .D(n10261), .CP(Clk), .Q(matrixInput[15])
         );
    VMW_AO22 U378 ( .A(matrixInput[81]), .B(n9707), .C(matrixInput[73]), .D(
        n9697), .Z(n10203) );
    VMW_AO22 U520 ( .A(matrixInput[414]), .B(n9707), .C(matrixInput[406]), .D(
        n9697), .Z(n9870) );
    VMW_FD \matrixInput_reg[374]  ( .D(n9902), .CP(Clk), .Q(matrixInput[374])
         );
    VMW_FD \matrixInput_reg[347]  ( .D(n9929), .CP(Clk), .Q(matrixInput[347])
         );
    VMW_AO22 U569 ( .A(matrixInput[370]), .B(n9707), .C(matrixInput[362]), .D(
        n9697), .Z(n9914) );
    VMW_AO22 U659 ( .A(matrixInput[289]), .B(n9707), .C(matrixInput[281]), .D(
        n9697), .Z(n9995) );
    VMW_AO22 U765 ( .A(matrixInput[194]), .B(n9707), .C(matrixInput[186]), .D(
        n9697), .Z(n10090) );
    VMW_AO22 U827 ( .A(matrixInput[20]), .B(n9707), .C(matrixInput[12]), .D(
        n9697), .Z(n10264) );
    VMW_FD \vectorInput_reg[44]  ( .D(n10296), .CP(Clk), .Q(vectorInput[44])
         );
    VMW_PULLDOWN U258 ( .Z(n9756) );
    VMW_PULLDOWN U263 ( .Z(n9761) );
    VMW_AO22 U455 ( .A(matrixInput[473]), .B(n9707), .C(matrixInput[465]), .D(
        n9697), .Z(n9811) );
    VMW_AO22 U472 ( .A(matrixInput[52]), .B(n9707), .C(matrixInput[44]), .D(
        n9697), .Z(n10232) );
    VMW_AO22 U800 ( .A(matrixInput[162]), .B(n9707), .C(matrixInput[154]), .D(
        n9697), .Z(n10122) );
    VMW_AND4 U278 ( .A(RD), .B(n164), .C(n9696), .D(n9697), .Z(n9671) );
    VMW_AO22 U469 ( .A(matrixInput[460]), .B(n9707), .C(matrixInput[452]), .D(
        n9697), .Z(n9824) );
    VMW_AO22 U742 ( .A(matrixInput[214]), .B(n9707), .C(matrixInput[206]), .D(
        n9697), .Z(n10070) );
    VMW_FD \matrixInput_reg[7]  ( .D(n10269), .CP(Clk), .Q(matrixInput[7]) );
    VMW_AO22 U759 ( .A(matrixInput[199]), .B(n9707), .C(matrixInput[191]), .D(
        n9697), .Z(n10085) );
    VMW_AO22 U344 ( .A(vectorInput[21]), .B(n9706), .C(vectorInput[13]), .D(
        n9696), .Z(n10327) );
    VMW_AO22 U363 ( .A(matrixInput[95]), .B(n9707), .C(matrixInput[87]), .D(
        n9697), .Z(n10189) );
    VMW_AO22 U642 ( .A(matrixInput[305]), .B(n9707), .C(matrixInput[297]), .D(
        n9697), .Z(n9979) );
    VMW_FD \matrixInput_reg[364]  ( .D(n9912), .CP(Clk), .Q(matrixInput[364])
         );
    VMW_FD \matrixInput_reg[357]  ( .D(n9919), .CP(Clk), .Q(matrixInput[357])
         );
    VMW_AO22 U890 ( .A(cOutput[48]), .B(n9702), .C(cOutput[16]), .D(n9701), 
        .Z(n9737) );
    VMW_OAI21 U900 ( .A(n9718), .B(n9719), .C(n9705), .Z(n9688) );
    VMW_AO22 U555 ( .A(matrixInput[383]), .B(n9707), .C(matrixInput[375]), .D(
        n9697), .Z(n9901) );
    VMW_AO22 U572 ( .A(matrixInput[43]), .B(n9707), .C(matrixInput[35]), .D(
        n9697), .Z(n10241) );
    VMW_BUFIZ U927 ( .A(n9744), .E(RD), .Z(\DataOut[10]1 ) );
    VMW_AO22 U381 ( .A(matrixInput[78]), .B(n9707), .C(matrixInput[70]), .D(
        n9697), .Z(n10206) );
    VMW_AO22 U386 ( .A(matrixInput[74]), .B(n9707), .C(matrixInput[66]), .D(
        n9697), .Z(n10210) );
    VMW_AO22 U407 ( .A(DataIn[4]), .B(n9707), .C(matrixInput[508]), .D(n9697), 
        .Z(n9768) );
    VMW_AO22 U420 ( .A(matrixInput[505]), .B(n9707), .C(matrixInput[497]), .D(
        n9697), .Z(n9779) );
    VMW_AO22 U665 ( .A(matrixInput[284]), .B(n9707), .C(matrixInput[276]), .D(
        n9697), .Z(n10000) );
    VMW_AO22 U852 ( .A(matrixInput[115]), .B(n9707), .C(matrixInput[107]), .D(
        n9697), .Z(n10169) );
    VMW_BUFIZ U949 ( .A(\holder[7] ), .E(RD), .Z(\DataOut[7]1 ) );
    VMW_FD \matrixInput_reg[125]  ( .D(n10151), .CP(Clk), .Q(matrixInput[125])
         );
    VMW_FD \vectorInput_reg[54]  ( .D(n10286), .CP(Clk), .Q(vectorInput[54])
         );
    VMW_FD \matrixInput_reg[431]  ( .D(n9845), .CP(Clk), .Q(matrixInput[431])
         );
    VMW_FD \matrixInput_reg[226]  ( .D(n10050), .CP(Clk), .Q(matrixInput[226])
         );
    VMW_FD \matrixInput_reg[215]  ( .D(n10061), .CP(Clk), .Q(matrixInput[215])
         );
    VMW_FD \matrixInput_reg[116]  ( .D(n10160), .CP(Clk), .Q(matrixInput[116])
         );
    VMW_FD \vectorInput_reg[8]  ( .D(n10332), .CP(Clk), .Q(vectorInput[8]) );
    VMW_FD \matrixInput_reg[428]  ( .D(n9848), .CP(Clk), .Q(matrixInput[428])
         );
    VMW_FD \matrixInput_reg[402]  ( .D(n9874), .CP(Clk), .Q(matrixInput[402])
         );
    VMW_FD \matrixInput_reg[385]  ( .D(n9891), .CP(Clk), .Q(matrixInput[385])
         );
    VMW_FD \matrixInput_reg[36]  ( .D(n10240), .CP(Clk), .Q(matrixInput[36])
         );
    VMW_AO22 U597 ( .A(matrixInput[345]), .B(n9707), .C(matrixInput[337]), .D(
        n9697), .Z(n9939) );
    VMW_AO22 U680 ( .A(matrixInput[270]), .B(n9707), .C(matrixInput[262]), .D(
        n9697), .Z(n10014) );
    VMW_AO22 U710 ( .A(matrixInput[243]), .B(n9707), .C(matrixInput[235]), .D(
        n9697), .Z(n10041) );
    VMW_AO22 U737 ( .A(matrixInput[218]), .B(n9707), .C(matrixInput[210]), .D(
        n9697), .Z(n10066) );
    VMW_AO22 U875 ( .A(cOutput[44]), .B(n9699), .C(cOutput[12]), .D(n9698), 
        .Z(n9722) );
    VMW_FD \matrixInput_reg[433]  ( .D(n9843), .CP(Clk), .Q(matrixInput[433])
         );
    VMW_FD \matrixInput_reg[224]  ( .D(n10052), .CP(Clk), .Q(matrixInput[224])
         );
    VMW_FD \matrixInput_reg[217]  ( .D(n10059), .CP(Clk), .Q(matrixInput[217])
         );
    VMW_FD \matrixInput_reg[127]  ( .D(n10149), .CP(Clk), .Q(matrixInput[127])
         );
    VMW_FD \matrixInput_reg[114]  ( .D(n10162), .CP(Clk), .Q(matrixInput[114])
         );
    VMW_FD \matrixInput_reg[419]  ( .D(n9857), .CP(Clk), .Q(matrixInput[419])
         );
    VMW_FD \matrixInput_reg[400]  ( .D(n9876), .CP(Clk), .Q(matrixInput[400])
         );
    VMW_FD \matrixInput_reg[387]  ( .D(n9889), .CP(Clk), .Q(matrixInput[387])
         );
    VMW_AO22 U400 ( .A(matrixInput[61]), .B(n9707), .C(matrixInput[53]), .D(
        n9697), .Z(n10223) );
    VMW_AO22 U427 ( .A(matrixInput[498]), .B(n9707), .C(matrixInput[490]), .D(
        n9697), .Z(n9786) );
    VMW_AO22 U590 ( .A(matrixInput[351]), .B(n9707), .C(matrixInput[343]), .D(
        n9697), .Z(n9933) );
    VMW_AO22 U687 ( .A(matrixInput[264]), .B(n9707), .C(matrixInput[256]), .D(
        n9697), .Z(n10020) );
    VMW_AO22 U730 ( .A(matrixInput[225]), .B(n9707), .C(matrixInput[217]), .D(
        n9697), .Z(n10059) );
    VMW_AO22 U872 ( .A(cOutput[61]), .B(n9702), .C(cOutput[29]), .D(n9701), 
        .Z(n9719) );
    VMW_FD \matrixInput_reg[34]  ( .D(n10242), .CP(Clk), .Q(matrixInput[34])
         );
    VMW_AO22 U717 ( .A(matrixInput[237]), .B(n9707), .C(matrixInput[229]), .D(
        n9697), .Z(n10047) );
    VMW_AO22 U449 ( .A(matrixInput[478]), .B(n9707), .C(matrixInput[470]), .D(
        n9697), .Z(n9806) );
    VMW_AO22 U779 ( .A(matrixInput[181]), .B(n9707), .C(matrixInput[173]), .D(
        n9697), .Z(n10103) );
    VMW_AO22 U855 ( .A(matrixInput[112]), .B(n9707), .C(matrixInput[104]), .D(
        n9697), .Z(n10172) );
    VMW_PULLDOWN U264 ( .Z(n9762) );
    VMW_AO22 U343 ( .A(vectorInput[22]), .B(n9706), .C(vectorInput[14]), .D(
        n9696), .Z(n10326) );
    VMW_AO22 U662 ( .A(matrixInput[287]), .B(n9707), .C(matrixInput[279]), .D(
        n9697), .Z(n9997) );
    VMW_FD \matrixInput_reg[366]  ( .D(n9910), .CP(Clk), .Q(matrixInput[366])
         );
    VMW_FD \matrixInput_reg[355]  ( .D(n9921), .CP(Clk), .Q(matrixInput[355])
         );
    VMW_AO22 U358 ( .A(matrixInput[99]), .B(n9707), .C(matrixInput[91]), .D(
        n9697), .Z(n10185) );
    VMW_AO22 U364 ( .A(matrixInput[94]), .B(n9707), .C(matrixInput[86]), .D(
        n9697), .Z(n10190) );
    VMW_AO22 U552 ( .A(matrixInput[386]), .B(n9707), .C(matrixInput[378]), .D(
        n9697), .Z(n9898) );
    VMW_AO22 U575 ( .A(matrixInput[365]), .B(n9707), .C(matrixInput[357]), .D(
        n9697), .Z(n9919) );
    VMW_INV U920 ( .A(\holder[2] ), .Z(n9678) );
    VMW_AO22 U645 ( .A(matrixInput[302]), .B(n9707), .C(matrixInput[294]), .D(
        n9697), .Z(n9982) );
    VMW_OAI21 U897 ( .A(n9712), .B(n9713), .C(n9703), .Z(n9692) );
    VMW_OAI21 U907 ( .A(n9732), .B(n9733), .C(n9703), .Z(n9677) );
    VMW_FD \vectorInput_reg[56]  ( .D(n10284), .CP(Clk), .Q(vectorInput[56])
         );
    VMW_FD \matrixInput_reg[376]  ( .D(n9900), .CP(Clk), .Q(matrixInput[376])
         );
    VMW_FD \matrixInput_reg[345]  ( .D(n9931), .CP(Clk), .Q(matrixInput[345])
         );
    VMW_AO22 U549 ( .A(matrixInput[388]), .B(n9707), .C(matrixInput[380]), .D(
        n9697), .Z(n9896) );
    VMW_AO22 U679 ( .A(matrixInput[271]), .B(n9707), .C(matrixInput[263]), .D(
        n9697), .Z(n10013) );
    VMW_AO22 U745 ( .A(matrixInput[211]), .B(n9707), .C(matrixInput[203]), .D(
        n9697), .Z(n10073) );
    VMW_FD \vectorInput_reg[46]  ( .D(n10294), .CP(Clk), .Q(vectorInput[46])
         );
    VMW_AO22 U452 ( .A(matrixInput[476]), .B(n9707), .C(matrixInput[468]), .D(
        n9697), .Z(n9808) );
    VMW_AO22 U475 ( .A(matrixInput[455]), .B(n9707), .C(matrixInput[447]), .D(
        n9697), .Z(n9829) );
    VMW_AO22 U807 ( .A(matrixInput[156]), .B(n9707), .C(matrixInput[148]), .D(
        n9697), .Z(n10128) );
    VMW_FD \matrixInput_reg[5]  ( .D(n10271), .CP(Clk), .Q(matrixInput[5]) );
    VMW_PULLDOWN U251 ( .Z(n9749) );
    VMW_OAI211 U276 ( .A(n9671), .B(n9690), .C(n9691), .D(n9692), .Z(n10342)
         );
    VMW_NOR2 U281 ( .A(n9700), .B(Addr[2]), .Z(n9701) );
    VMW_AO22 U311 ( .A(vectorInput[51]), .B(n9706), .C(vectorInput[43]), .D(
        n9696), .Z(n10297) );
    VMW_AO22 U336 ( .A(vectorInput[28]), .B(n9706), .C(vectorInput[20]), .D(
        n9696), .Z(n10320) );
    VMW_AO22 U527 ( .A(matrixInput[11]), .B(n9707), .C(matrixInput[3]), .D(
        n9697), .Z(n10273) );
    VMW_AO22 U762 ( .A(matrixInput[197]), .B(n9707), .C(matrixInput[189]), .D(
        n9697), .Z(n10087) );
    VMW_AO22 U820 ( .A(matrixInput[144]), .B(n9707), .C(matrixInput[136]), .D(
        n9697), .Z(n10140) );
    VMW_AO22 U869 ( .A(cOutput[37]), .B(n9699), .C(cOutput[5]), .D(n9698), .Z(
        n9716) );
    VMW_FD \matrixInput_reg[423]  ( .D(n9853), .CP(Clk), .Q(matrixInput[423])
         );
    VMW_FD \matrixInput_reg[410]  ( .D(n9866), .CP(Clk), .Q(matrixInput[410])
         );
    VMW_FD \matrixInput_reg[409]  ( .D(n9867), .CP(Clk), .Q(matrixInput[409])
         );
    VMW_FD \matrixInput_reg[397]  ( .D(n9879), .CP(Clk), .Q(matrixInput[397])
         );
    VMW_FD \matrixInput_reg[234]  ( .D(n10042), .CP(Clk), .Q(matrixInput[234])
         );
    VMW_FD \matrixInput_reg[207]  ( .D(n10069), .CP(Clk), .Q(matrixInput[207])
         );
    VMW_FD \vectorInput_reg[3]  ( .D(n10337), .CP(Clk), .Q(vectorInput[3]) );
    VMW_FD \matrixInput_reg[104]  ( .D(n10172), .CP(Clk), .Q(matrixInput[104])
         );
    VMW_FD \matrixInput_reg[137]  ( .D(n10139), .CP(Clk), .Q(matrixInput[137])
         );
    VMW_AO22 U617 ( .A(matrixInput[327]), .B(n9707), .C(matrixInput[319]), .D(
        n9697), .Z(n9957) );
    VMW_BUFIZ U955 ( .A(n9764), .E(RD), .Z(\DataOut[8]1 ) );
    VMW_AO22 U630 ( .A(matrixInput[315]), .B(n9707), .C(matrixInput[307]), .D(
        n9697), .Z(n9969) );
    VMW_AO22 U787 ( .A(matrixInput[174]), .B(n9707), .C(matrixInput[166]), .D(
        n9697), .Z(n10110) );
    VMW_FD \matrixInput_reg[17]  ( .D(n10259), .CP(Clk), .Q(matrixInput[17])
         );
    VMW_AO22 U490 ( .A(matrixInput[441]), .B(n9707), .C(matrixInput[433]), .D(
        n9697), .Z(n9843) );
    VMW_AO22 U293 ( .A(vectorInput[13]), .B(n9706), .C(vectorInput[5]), .D(
        n9696), .Z(n10335) );
    VMW_AO22 U324 ( .A(vectorInput[39]), .B(n9706), .C(vectorInput[31]), .D(
        n9696), .Z(n10309) );
    VMW_AO22 U500 ( .A(matrixInput[432]), .B(n9707), .C(matrixInput[424]), .D(
        n9697), .Z(n9852) );
    VMW_BUFIZ U947 ( .A(\holder[3] ), .E(RD), .Z(\DataOut[3]1 ) );
    VMW_FD \matrixInput_reg[24]  ( .D(n10252), .CP(Clk), .Q(matrixInput[24])
         );
    VMW_AO22 U535 ( .A(matrixInput[401]), .B(n9707), .C(matrixInput[393]), .D(
        n9697), .Z(n9883) );
    VMW_AO22 U605 ( .A(matrixInput[40]), .B(n9707), .C(matrixInput[32]), .D(
        n9697), .Z(n10244) );
    VMW_AO22 U795 ( .A(matrixInput[167]), .B(n9707), .C(matrixInput[159]), .D(
        n9697), .Z(n10117) );
    VMW_FD \vectorInput_reg[61]  ( .D(n10279), .CP(Clk), .Q(vectorInput[61])
         );
    VMW_AO22 U622 ( .A(matrixInput[322]), .B(n9707), .C(matrixInput[314]), .D(
        n9697), .Z(n9962) );
    VMW_FD \vectorInput_reg[52]  ( .D(n10288), .CP(Clk), .Q(vectorInput[52])
         );
    IntMatMul_Control_pVectorSize8_pWordSize8_pScan1_DW01_cmp2_15_0 lt_130 ( 
        .A({Addr[14], Addr[13], Addr[12], Addr[11], Addr[10], Addr[9], Addr[8], 
        Addr[7], Addr[6], Addr[5], Addr[4], Addr[3], UNCONNECTED_1, 
        UNCONNECTED_2, UNCONNECTED_3}), .B({Logic01, Logic01, Logic01, Logic01, 
        Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, Logic11, 
        Logic01, Logic01, Logic01}), .LEQ(n10349), .TC(n10349), .LT_LE(n164)
         );
    VMW_FD \matrixInput_reg[8]  ( .D(n10268), .CP(Clk), .Q(matrixInput[8]) );
    VMW_AO22 U303 ( .A(vectorInput[58]), .B(n9706), .C(vectorInput[50]), .D(
        n9696), .Z(n10290) );
    VMW_AO22 U512 ( .A(matrixInput[421]), .B(n9707), .C(matrixInput[413]), .D(
        n9697), .Z(n9863) );
    VMW_AO22 U388 ( .A(matrixInput[72]), .B(n9707), .C(matrixInput[64]), .D(
        n9697), .Z(n10212) );
    VMW_AO22 U482 ( .A(matrixInput[448]), .B(n9707), .C(matrixInput[440]), .D(
        n9697), .Z(n9836) );
    VMW_AO22 U599 ( .A(matrixInput[343]), .B(n9707), .C(matrixInput[335]), .D(
        n9697), .Z(n9941) );
    VMW_AO22 U739 ( .A(matrixInput[217]), .B(n9707), .C(matrixInput[209]), .D(
        n9697), .Z(n10067) );
    VMW_FD \matrixInput_reg[362]  ( .D(n9914), .CP(Clk), .Q(matrixInput[362])
         );
    VMW_FD \matrixInput_reg[351]  ( .D(n9925), .CP(Clk), .Q(matrixInput[351])
         );
    VMW_FD \matrixInput_reg[348]  ( .D(n9928), .CP(Clk), .Q(matrixInput[348])
         );
    VMW_AO22 U409 ( .A(DataIn[2]), .B(n9707), .C(matrixInput[506]), .D(n9697), 
        .Z(n9770) );
    VMW_AO22 U467 ( .A(matrixInput[462]), .B(n9707), .C(matrixInput[454]), .D(
        n9697), .Z(n9822) );
    VMW_AO22 U757 ( .A(matrixInput[201]), .B(n9707), .C(matrixInput[193]), .D(
        n9697), .Z(n10083) );
    VMW_AO22 U815 ( .A(matrixInput[148]), .B(n9707), .C(matrixInput[140]), .D(
        n9697), .Z(n10136) );
    VMW_AO22 U832 ( .A(matrixInput[133]), .B(n9707), .C(matrixInput[125]), .D(
        n9697), .Z(n10151) );
    VMW_FD \matrixInput_reg[30]  ( .D(n10246), .CP(Clk), .Q(matrixInput[30])
         );
    VMW_FD \matrixInput_reg[29]  ( .D(n10247), .CP(Clk), .Q(matrixInput[29])
         );
    VMW_PULLDOWN U265 ( .Z(n9763) );
    VMW_AND2 U280 ( .A(Addr[2]), .B(n9700), .Z(n9699) );
    VMW_AO22 U288 ( .A(vectorInput[14]), .B(n9706), .C(vectorInput[6]), .D(
        n9696), .Z(n10334) );
    VMW_AO22 U351 ( .A(matrixInput[106]), .B(n9707), .C(matrixInput[98]), .D(
        n9697), .Z(n10178) );
    VMW_AO22 U440 ( .A(matrixInput[487]), .B(n9707), .C(matrixInput[479]), .D(
        n9697), .Z(n9797) );
    VMW_AO22 U540 ( .A(matrixInput[397]), .B(n9707), .C(matrixInput[389]), .D(
        n9697), .Z(n9887) );
    VMW_AO22 U670 ( .A(matrixInput[279]), .B(n9707), .C(matrixInput[271]), .D(
        n9697), .Z(n10005) );
    VMW_AO22 U770 ( .A(matrixInput[189]), .B(n9707), .C(matrixInput[181]), .D(
        n9697), .Z(n10095) );
    VMW_BUFIZ U929 ( .A(n9745), .E(RD), .Z(\DataOut[14]1 ) );
    VMW_FD \matrixInput_reg[437]  ( .D(n9839), .CP(Clk), .Q(matrixInput[437])
         );
    VMW_FD \matrixInput_reg[404]  ( .D(n9872), .CP(Clk), .Q(matrixInput[404])
         );
    VMW_FD \matrixInput_reg[383]  ( .D(n9893), .CP(Clk), .Q(matrixInput[383])
         );
    VMW_FD \matrixInput_reg[123]  ( .D(n10153), .CP(Clk), .Q(matrixInput[123])
         );
    VMW_FD \matrixInput_reg[239]  ( .D(n10037), .CP(Clk), .Q(matrixInput[239])
         );
    VMW_FD \matrixInput_reg[220]  ( .D(n10056), .CP(Clk), .Q(matrixInput[220])
         );
    VMW_FD \matrixInput_reg[213]  ( .D(n10063), .CP(Clk), .Q(matrixInput[213])
         );
    VMW_FD \matrixInput_reg[110]  ( .D(n10166), .CP(Clk), .Q(matrixInput[110])
         );
    VMW_FD \matrixInput_reg[109]  ( .D(n10167), .CP(Clk), .Q(matrixInput[109])
         );
    VMW_BUFIZ U932 ( .A(n9747), .E(RD), .Z(\DataOut[25]1 ) );
    VMW_FD \matrixInput_reg[39]  ( .D(n10237), .CP(Clk), .Q(matrixInput[39])
         );
    VMW_FD \matrixInput_reg[13]  ( .D(n10263), .CP(Clk), .Q(matrixInput[13])
         );
    VMW_FD \matrixInput_reg[20]  ( .D(n10256), .CP(Clk), .Q(matrixInput[20])
         );
    VMW_AO22 U376 ( .A(matrixInput[83]), .B(n9707), .C(matrixInput[75]), .D(
        n9697), .Z(n10201) );
    VMW_AO22 U885 ( .A(cOutput[33]), .B(n9699), .C(cOutput[1]), .D(n9698), .Z(
        n9732) );
    VMW_INV U915 ( .A(Addr[1]), .Z(n9700) );
    VMW_AO22 U393 ( .A(matrixInput[13]), .B(n9707), .C(matrixInput[5]), .D(
        n9697), .Z(n10271) );
    VMW_AO22 U567 ( .A(matrixInput[372]), .B(n9707), .C(matrixInput[364]), .D(
        n9697), .Z(n9912) );
    VMW_AO22 U582 ( .A(matrixInput[358]), .B(n9707), .C(matrixInput[350]), .D(
        n9697), .Z(n9926) );
    VMW_AO22 U657 ( .A(matrixInput[291]), .B(n9707), .C(matrixInput[283]), .D(
        n9697), .Z(n9993) );
    VMW_AO22 U829 ( .A(matrixInput[136]), .B(n9707), .C(matrixInput[128]), .D(
        n9697), .Z(n10148) );
    VMW_FD \matrixInput_reg[203]  ( .D(n10073), .CP(Clk), .Q(matrixInput[203])
         );
    VMW_FD \matrixInput_reg[119]  ( .D(n10157), .CP(Clk), .Q(matrixInput[119])
         );
    VMW_FD \matrixInput_reg[100]  ( .D(n10176), .CP(Clk), .Q(matrixInput[100])
         );
    VMW_FD \matrixInput_reg[133]  ( .D(n10143), .CP(Clk), .Q(matrixInput[133])
         );
    VMW_AO22 U860 ( .A(matrixInput[8]), .B(n9707), .C(matrixInput[0]), .D(
        n9697), .Z(n10276) );
    VMW_FD \matrixInput_reg[427]  ( .D(n9849), .CP(Clk), .Q(matrixInput[427])
         );
    VMW_FD \matrixInput_reg[414]  ( .D(n9862), .CP(Clk), .Q(matrixInput[414])
         );
    VMW_FD \matrixInput_reg[393]  ( .D(n9883), .CP(Clk), .Q(matrixInput[393])
         );
    VMW_FD \matrixInput_reg[230]  ( .D(n10046), .CP(Clk), .Q(matrixInput[230])
         );
    VMW_FD \matrixInput_reg[229]  ( .D(n10047), .CP(Clk), .Q(matrixInput[229])
         );
    VMW_FD \vectorInput_reg[7]  ( .D(n10333), .CP(Clk), .Q(vectorInput[7]) );
    VMW_AO22 U412 ( .A(matrixInput[511]), .B(n9707), .C(matrixInput[503]), .D(
        n9697), .Z(n9773) );
    VMW_AO22 U435 ( .A(matrixInput[491]), .B(n9707), .C(matrixInput[483]), .D(
        n9697), .Z(n9793) );
    VMW_AO22 U695 ( .A(matrixInput[257]), .B(n9707), .C(matrixInput[249]), .D(
        n9697), .Z(n10027) );
    VMW_AO22 U705 ( .A(matrixInput[31]), .B(n9707), .C(matrixInput[23]), .D(
        n9697), .Z(n10253) );
    VMW_AO22 U722 ( .A(matrixInput[232]), .B(n9707), .C(matrixInput[224]), .D(
        n9697), .Z(n10052) );
    VMW_FD \matrixInput_reg[1]  ( .D(n10275), .CP(Clk), .Q(matrixInput[1]) );
    VMW_AO22 U847 ( .A(matrixInput[119]), .B(n9707), .C(matrixInput[111]), .D(
        n9697), .Z(n10165) );
    VMW_FD \vectorInput_reg[42]  ( .D(n10298), .CP(Clk), .Q(vectorInput[42])
         );
    VMW_AO22 U318 ( .A(vectorInput[45]), .B(n9706), .C(vectorInput[37]), .D(
        n9696), .Z(n10303) );
    VMW_AO22 U509 ( .A(matrixInput[424]), .B(n9707), .C(matrixInput[416]), .D(
        n9697), .Z(n9860) );
    VMW_AO22 U337 ( .A(vectorInput[9]), .B(n9706), .C(vectorInput[1]), .D(
        n9696), .Z(n10339) );
    VMW_AO22 U499 ( .A(matrixInput[433]), .B(n9707), .C(matrixInput[425]), .D(
        n9697), .Z(n9851) );
    VMW_AO22 U639 ( .A(matrixInput[37]), .B(n9707), .C(matrixInput[29]), .D(
        n9697), .Z(n10247) );
    VMW_AO22 U868 ( .A(cOutput[62]), .B(n9702), .C(cOutput[30]), .D(n9701), 
        .Z(n9715) );
    VMW_FD \matrixInput_reg[471]  ( .D(n9805), .CP(Clk), .Q(matrixInput[471])
         );
    VMW_FD \matrixInput_reg[468]  ( .D(n9808), .CP(Clk), .Q(matrixInput[468])
         );
    VMW_FD \matrixInput_reg[372]  ( .D(n9904), .CP(Clk), .Q(matrixInput[372])
         );
    VMW_FD \matrixInput_reg[358]  ( .D(n9918), .CP(Clk), .Q(matrixInput[358])
         );
    VMW_FD \matrixInput_reg[341]  ( .D(n9935), .CP(Clk), .Q(matrixInput[341])
         );
    VMW_FD \matrixInput_reg[442]  ( .D(n9834), .CP(Clk), .Q(matrixInput[442])
         );
    VMW_FD \matrixInput_reg[266]  ( .D(n10010), .CP(Clk), .Q(matrixInput[266])
         );
    VMW_FD \matrixInput_reg[165]  ( .D(n10111), .CP(Clk), .Q(matrixInput[165])
         );
    VMW_FD \matrixInput_reg[255]  ( .D(n10021), .CP(Clk), .Q(matrixInput[255])
         );
    VMW_FD \matrixInput_reg[156]  ( .D(n10120), .CP(Clk), .Q(matrixInput[156])
         );
    VMW_AO22 U501 ( .A(matrixInput[431]), .B(n9707), .C(matrixInput[423]), .D(
        n9697), .Z(n9853) );
    VMW_AO22 U526 ( .A(matrixInput[408]), .B(n9707), .C(matrixInput[400]), .D(
        n9697), .Z(n9876) );
    VMW_AO22 U616 ( .A(matrixInput[39]), .B(n9707), .C(matrixInput[31]), .D(
        n9697), .Z(n10245) );
    VMW_AO22 U786 ( .A(matrixInput[175]), .B(n9707), .C(matrixInput[167]), .D(
        n9697), .Z(n10109) );
    VMW_BUFIZ U954 ( .A(\holder[1] ), .E(RD), .Z(\DataOut[1]1 ) );
    VMW_AO22 U631 ( .A(matrixInput[314]), .B(n9707), .C(matrixInput[306]), .D(
        n9697), .Z(n9970) );
    VMW_FD \matrixInput_reg[76]  ( .D(n10200), .CP(Clk), .Q(matrixInput[76])
         );
    VMW_AO22 U310 ( .A(vectorInput[52]), .B(n9706), .C(vectorInput[44]), .D(
        n9696), .Z(n10296) );
    VMW_AO22 U491 ( .A(matrixInput[440]), .B(n9707), .C(matrixInput[432]), .D(
        n9697), .Z(n9844) );
    VMW_AO22 U359 ( .A(matrixInput[98]), .B(n9707), .C(matrixInput[90]), .D(
        n9697), .Z(n10186) );
    VMW_AO22 U548 ( .A(matrixInput[389]), .B(n9707), .C(matrixInput[381]), .D(
        n9697), .Z(n9895) );
    VMW_FD \matrixInput_reg[490]  ( .D(n9786), .CP(Clk), .Q(matrixInput[490])
         );
    VMW_FD \matrixInput_reg[45]  ( .D(n10231), .CP(Clk), .Q(matrixInput[45])
         );
    VMW_FD \matrixInput_reg[489]  ( .D(n9787), .CP(Clk), .Q(matrixInput[489])
         );
    VMW_FD \matrixInput_reg[324]  ( .D(n9952), .CP(Clk), .Q(matrixInput[324])
         );
    VMW_FD \matrixInput_reg[317]  ( .D(n9959), .CP(Clk), .Q(matrixInput[317])
         );
    VMW_FD \matrixInput_reg[287]  ( .D(n9989), .CP(Clk), .Q(matrixInput[287])
         );
    VMW_FD \matrixInput_reg[184]  ( .D(n10092), .CP(Clk), .Q(matrixInput[184])
         );
    VMW_FD \matrixInput_reg[500]  ( .D(n9776), .CP(Clk), .Q(matrixInput[500])
         );
    VMW_AO22 U474 ( .A(matrixInput[456]), .B(n9707), .C(matrixInput[448]), .D(
        n9697), .Z(n9828) );
    VMW_AO22 U678 ( .A(matrixInput[272]), .B(n9707), .C(matrixInput[264]), .D(
        n9697), .Z(n10012) );
    VMW_AO22 U744 ( .A(matrixInput[212]), .B(n9707), .C(matrixInput[204]), .D(
        n9697), .Z(n10072) );
    VMW_FD \vectorInput_reg[27]  ( .D(n10313), .CP(Clk), .Q(vectorInput[27])
         );
    VMW_AO22 U453 ( .A(matrixInput[475]), .B(n9707), .C(matrixInput[467]), .D(
        n9697), .Z(n9809) );
    VMW_AO22 U806 ( .A(matrixInput[157]), .B(n9707), .C(matrixInput[149]), .D(
        n9697), .Z(n10127) );
    VMW_FD \matrixInput_reg[97]  ( .D(n10179), .CP(Clk), .Q(matrixInput[97])
         );
    VMW_FD \vectorInput_reg[14]  ( .D(n10326), .CP(Clk), .Q(vectorInput[14])
         );
    VMW_AO22 U763 ( .A(matrixInput[196]), .B(n9707), .C(matrixInput[188]), .D(
        n9697), .Z(n10088) );
    VMW_AO22 U821 ( .A(matrixInput[143]), .B(n9707), .C(matrixInput[135]), .D(
        n9697), .Z(n10141) );
    VMW_FD \holder_reg[1]  ( .D(n10347), .CP(Clk), .Q(\holder[1] ) );
    VMW_PULLDOWN U245 ( .Z(n9743) );
    VMW_PULLDOWN U250 ( .Z(n9748) );
    VMW_PULLDOWN U259 ( .Z(n9757) );
    VMW_AO22 U778 ( .A(matrixInput[182]), .B(n9707), .C(matrixInput[174]), .D(
        n9697), .Z(n10102) );
    VMW_FD \matrixInput_reg[509]  ( .D(n9767), .CP(Clk), .Q(matrixInput[509])
         );
    VMW_FD \matrixInput_reg[297]  ( .D(n9979), .CP(Clk), .Q(matrixInput[297])
         );
    VMW_FD \matrixInput_reg[194]  ( .D(n10082), .CP(Clk), .Q(matrixInput[194])
         );
    VMW_OAI211 U277 ( .A(n9671), .B(n9693), .C(n9694), .D(n9695), .Z(n10341)
         );
    VMW_AO22 U289 ( .A(DataIn[7]), .B(n9706), .C(vectorInput[63]), .D(n9696), 
        .Z(n10277) );
    VMW_AO22 U319 ( .A(vectorInput[44]), .B(n9706), .C(vectorInput[36]), .D(
        n9696), .Z(n10304) );
    VMW_AO22 U342 ( .A(vectorInput[23]), .B(n9706), .C(vectorInput[15]), .D(
        n9696), .Z(n10325) );
    VMW_AO22 U448 ( .A(matrixInput[479]), .B(n9707), .C(matrixInput[471]), .D(
        n9697), .Z(n9805) );
    VMW_AO22 U553 ( .A(matrixInput[385]), .B(n9707), .C(matrixInput[377]), .D(
        n9697), .Z(n9899) );
    VMW_AO22 U663 ( .A(matrixInput[286]), .B(n9707), .C(matrixInput[278]), .D(
        n9697), .Z(n9998) );
    VMW_FD \matrixInput_reg[510]  ( .D(n9766), .CP(Clk), .Q(matrixInput[510])
         );
    VMW_FD \matrixInput_reg[499]  ( .D(n9777), .CP(Clk), .Q(matrixInput[499])
         );
    VMW_FD \matrixInput_reg[334]  ( .D(n9942), .CP(Clk), .Q(matrixInput[334])
         );
    VMW_FD \matrixInput_reg[480]  ( .D(n9796), .CP(Clk), .Q(matrixInput[480])
         );
    VMW_FD \matrixInput_reg[307]  ( .D(n9969), .CP(Clk), .Q(matrixInput[307])
         );
    VMW_AO22 U365 ( .A(matrixInput[93]), .B(n9707), .C(matrixInput[85]), .D(
        n9697), .Z(n10191) );
    VMW_INV U921 ( .A(\holder[6] ), .Z(n9690) );
    VMW_FD \matrixInput_reg[87]  ( .D(n10189), .CP(Clk), .Q(matrixInput[87])
         );
    VMW_AO22 U380 ( .A(matrixInput[79]), .B(n9707), .C(matrixInput[71]), .D(
        n9697), .Z(n10205) );
    VMW_AO22 U401 ( .A(matrixInput[60]), .B(n9707), .C(matrixInput[52]), .D(
        n9697), .Z(n10224) );
    VMW_AO22 U574 ( .A(matrixInput[366]), .B(n9707), .C(matrixInput[358]), .D(
        n9697), .Z(n9918) );
    VMW_AO22 U591 ( .A(matrixInput[350]), .B(n9707), .C(matrixInput[342]), .D(
        n9697), .Z(n9934) );
    VMW_AO22 U644 ( .A(matrixInput[303]), .B(n9707), .C(matrixInput[295]), .D(
        n9697), .Z(n9981) );
    VMW_OAI21 U896 ( .A(n9710), .B(n9711), .C(n9705), .Z(n9694) );
    VMW_OAI21 U906 ( .A(n9730), .B(n9731), .C(n9705), .Z(n9679) );
    VMW_FD \matrixInput_reg[478]  ( .D(n9798), .CP(Clk), .Q(matrixInput[478])
         );
    VMW_FD \matrixInput_reg[461]  ( .D(n9815), .CP(Clk), .Q(matrixInput[461])
         );
    VMW_FD \matrixInput_reg[452]  ( .D(n9824), .CP(Clk), .Q(matrixInput[452])
         );
    VMW_FD \matrixInput_reg[276]  ( .D(n10000), .CP(Clk), .Q(matrixInput[276])
         );
    VMW_FD \matrixInput_reg[245]  ( .D(n10031), .CP(Clk), .Q(matrixInput[245])
         );
    VMW_FD \matrixInput_reg[146]  ( .D(n10130), .CP(Clk), .Q(matrixInput[146])
         );
    VMW_FD \vectorInput_reg[37]  ( .D(n10303), .CP(Clk), .Q(vectorInput[37])
         );
    VMW_FD \matrixInput_reg[175]  ( .D(n10101), .CP(Clk), .Q(matrixInput[175])
         );
    VMW_AO22 U392 ( .A(matrixInput[68]), .B(n9707), .C(matrixInput[60]), .D(
        n9697), .Z(n10216) );
    VMW_AO22 U413 ( .A(matrixInput[510]), .B(n9707), .C(matrixInput[502]), .D(
        n9697), .Z(n9774) );
    VMW_AO22 U426 ( .A(matrixInput[499]), .B(n9707), .C(matrixInput[491]), .D(
        n9697), .Z(n9785) );
    VMW_AO22 U686 ( .A(matrixInput[265]), .B(n9707), .C(matrixInput[257]), .D(
        n9697), .Z(n10019) );
    VMW_AO22 U716 ( .A(matrixInput[30]), .B(n9707), .C(matrixInput[22]), .D(
        n9697), .Z(n10254) );
    VMW_AO22 U731 ( .A(matrixInput[224]), .B(n9707), .C(matrixInput[216]), .D(
        n9697), .Z(n10060) );
    VMW_AO22 U873 ( .A(cOutput[36]), .B(n9699), .C(cOutput[4]), .D(n9698), .Z(
        n9720) );
    VMW_FD \matrixInput_reg[55]  ( .D(n10221), .CP(Clk), .Q(matrixInput[55])
         );
    VMW_FD \matrixInput_reg[66]  ( .D(n10210), .CP(Clk), .Q(matrixInput[66])
         );
    VMW_AO22 U854 ( .A(matrixInput[113]), .B(n9707), .C(matrixInput[105]), .D(
        n9697), .Z(n10171) );
    VMW_AO22 U861 ( .A(cOutput[39]), .B(n9699), .C(cOutput[7]), .D(n9698), .Z(
        n9708) );
    VMW_AO22 U434 ( .A(matrixInput[492]), .B(n9707), .C(matrixInput[484]), .D(
        n9697), .Z(n9792) );
    VMW_AO22 U583 ( .A(matrixInput[42]), .B(n9707), .C(matrixInput[34]), .D(
        n9697), .Z(n10242) );
    VMW_AO22 U694 ( .A(matrixInput[32]), .B(n9707), .C(matrixInput[24]), .D(
        n9697), .Z(n10252) );
    VMW_AO22 U723 ( .A(matrixInput[231]), .B(n9707), .C(matrixInput[223]), .D(
        n9697), .Z(n10053) );
    VMW_FD \matrixInput_reg[93]  ( .D(n10183), .CP(Clk), .Q(matrixInput[93])
         );
    VMW_FD \vectorInput_reg[23]  ( .D(n10317), .CP(Clk), .Q(vectorInput[23])
         );
    VMW_AO22 U704 ( .A(matrixInput[248]), .B(n9707), .C(matrixInput[240]), .D(
        n9697), .Z(n10036) );
    VMW_AO22 U846 ( .A(matrixInput[120]), .B(n9707), .C(matrixInput[112]), .D(
        n9697), .Z(n10164) );
    VMW_FD \vectorInput_reg[10]  ( .D(n10330), .CP(Clk), .Q(vectorInput[10])
         );
    VMW_AO22 U498 ( .A(matrixInput[434]), .B(n9707), .C(matrixInput[426]), .D(
        n9697), .Z(n9850) );
    VMW_AO22 U508 ( .A(matrixInput[425]), .B(n9707), .C(matrixInput[417]), .D(
        n9697), .Z(n9859) );
    VMW_AO22 U350 ( .A(matrixInput[107]), .B(n9707), .C(matrixInput[99]), .D(
        n9697), .Z(n10177) );
    VMW_AO22 U638 ( .A(matrixInput[10]), .B(n9707), .C(matrixInput[2]), .D(
        n9697), .Z(n10274) );
    VMW_FD \matrixInput_reg[504]  ( .D(n9772), .CP(Clk), .Q(matrixInput[504])
         );
    VMW_FD \matrixInput_reg[283]  ( .D(n9993), .CP(Clk), .Q(matrixInput[283])
         );
    VMW_FD \matrixInput_reg[199]  ( .D(n10077), .CP(Clk), .Q(matrixInput[199])
         );
    VMW_FD \matrixInput_reg[180]  ( .D(n10096), .CP(Clk), .Q(matrixInput[180])
         );
    VMW_AO22 U671 ( .A(matrixInput[278]), .B(n9707), .C(matrixInput[270]), .D(
        n9697), .Z(n10006) );
    VMW_FD \matrixInput_reg[494]  ( .D(n9782), .CP(Clk), .Q(matrixInput[494])
         );
    VMW_FD \matrixInput_reg[313]  ( .D(n9963), .CP(Clk), .Q(matrixInput[313])
         );
    VMW_FD \matrixInput_reg[339]  ( .D(n9937), .CP(Clk), .Q(matrixInput[339])
         );
    VMW_FD \matrixInput_reg[320]  ( .D(n9956), .CP(Clk), .Q(matrixInput[320])
         );
    VMW_BUFIZ U933 ( .A(n9748), .E(RD), .Z(\DataOut[16]1 ) );
    VMW_FD \matrixInput_reg[72]  ( .D(n10204), .CP(Clk), .Q(matrixInput[72])
         );
    VMW_FD \matrixInput_reg[58]  ( .D(n10218), .CP(Clk), .Q(matrixInput[58])
         );
    VMW_FD \matrixInput_reg[41]  ( .D(n10235), .CP(Clk), .Q(matrixInput[41])
         );
    VMW_AO22 U377 ( .A(matrixInput[82]), .B(n9707), .C(matrixInput[74]), .D(
        n9697), .Z(n10202) );
    VMW_AO22 U541 ( .A(matrixInput[396]), .B(n9707), .C(matrixInput[388]), .D(
        n9697), .Z(n9888) );
    VMW_AO22 U566 ( .A(matrixInput[373]), .B(n9707), .C(matrixInput[365]), .D(
        n9697), .Z(n9911) );
    VMW_AO22 U884 ( .A(cOutput[58]), .B(n9702), .C(cOutput[26]), .D(n9701), 
        .Z(n9731) );
    VMW_INV U914 ( .A(WR), .Z(n9740) );
    VMW_AO22 U656 ( .A(matrixInput[292]), .B(n9707), .C(matrixInput[284]), .D(
        n9697), .Z(n9992) );
    VMW_AO22 U756 ( .A(matrixInput[202]), .B(n9707), .C(matrixInput[194]), .D(
        n9697), .Z(n10082) );
    VMW_AO22 U828 ( .A(matrixInput[137]), .B(n9707), .C(matrixInput[129]), .D(
        n9697), .Z(n10147) );
    VMW_FD \matrixInput_reg[262]  ( .D(n10014), .CP(Clk), .Q(matrixInput[262])
         );
    VMW_FD \matrixInput_reg[251]  ( .D(n10025), .CP(Clk), .Q(matrixInput[251])
         );
    VMW_FD \matrixInput_reg[178]  ( .D(n10098), .CP(Clk), .Q(matrixInput[178])
         );
    VMW_FD \matrixInput_reg[161]  ( .D(n10115), .CP(Clk), .Q(matrixInput[161])
         );
    VMW_FD \matrixInput_reg[248]  ( .D(n10028), .CP(Clk), .Q(matrixInput[248])
         );
    VMW_FD \matrixInput_reg[152]  ( .D(n10124), .CP(Clk), .Q(matrixInput[152])
         );
    VMW_FD \matrixInput_reg[475]  ( .D(n9801), .CP(Clk), .Q(matrixInput[475])
         );
    VMW_FD \matrixInput_reg[446]  ( .D(n9830), .CP(Clk), .Q(matrixInput[446])
         );
    VMW_AO22 U814 ( .A(matrixInput[149]), .B(n9707), .C(matrixInput[141]), .D(
        n9697), .Z(n10135) );
    VMW_AO22 U441 ( .A(matrixInput[486]), .B(n9707), .C(matrixInput[478]), .D(
        n9697), .Z(n9798) );
    VMW_AO22 U466 ( .A(matrixInput[463]), .B(n9707), .C(matrixInput[455]), .D(
        n9697), .Z(n9821) );
    VMW_AO22 U833 ( .A(matrixInput[132]), .B(n9707), .C(matrixInput[124]), .D(
        n9697), .Z(n10152) );
    VMW_FD \matrixInput_reg[51]  ( .D(n10225), .CP(Clk), .Q(matrixInput[51])
         );
    VMW_FD \matrixInput_reg[48]  ( .D(n10228), .CP(Clk), .Q(matrixInput[48])
         );
    VMW_PULLDOWN U257 ( .Z(n9755) );
    VMW_AO22 U292 ( .A(DataIn[4]), .B(n9706), .C(vectorInput[60]), .D(n9696), 
        .Z(n10280) );
    VMW_AO22 U302 ( .A(vectorInput[59]), .B(n9706), .C(vectorInput[51]), .D(
        n9696), .Z(n10289) );
    VMW_AO22 U325 ( .A(vectorInput[38]), .B(n9706), .C(vectorInput[30]), .D(
        n9696), .Z(n10310) );
    VMW_AO22 U534 ( .A(matrixInput[402]), .B(n9707), .C(matrixInput[394]), .D(
        n9697), .Z(n9882) );
    VMW_AO22 U771 ( .A(matrixInput[188]), .B(n9707), .C(matrixInput[180]), .D(
        n9697), .Z(n10096) );
    VMW_BUFIZ U928 ( .A(\holder[0] ), .E(RD), .Z(\DataOut[0]1 ) );
    VMW_FD \matrixInput_reg[465]  ( .D(n9811), .CP(Clk), .Q(matrixInput[465])
         );
    VMW_FD \matrixInput_reg[456]  ( .D(n9820), .CP(Clk), .Q(matrixInput[456])
         );
    VMW_FD \matrixInput_reg[62]  ( .D(n10214), .CP(Clk), .Q(matrixInput[62])
         );
    VMW_FD \matrixInput_reg[258]  ( .D(n10018), .CP(Clk), .Q(matrixInput[258])
         );
    VMW_FD \matrixInput_reg[241]  ( .D(n10035), .CP(Clk), .Q(matrixInput[241])
         );
    VMW_FD \matrixInput_reg[142]  ( .D(n10134), .CP(Clk), .Q(matrixInput[142])
         );
    VMW_BUFIZ U946 ( .A(n9759), .E(RD), .Z(\DataOut[17]1 ) );
    VMW_FD \matrixInput_reg[272]  ( .D(n10004), .CP(Clk), .Q(matrixInput[272])
         );
    VMW_FD \matrixInput_reg[171]  ( .D(n10105), .CP(Clk), .Q(matrixInput[171])
         );
    VMW_FD \matrixInput_reg[168]  ( .D(n10108), .CP(Clk), .Q(matrixInput[168])
         );
    VMW_FD \vectorInput_reg[19]  ( .D(n10321), .CP(Clk), .Q(vectorInput[19])
         );
    VMW_AO22 U483 ( .A(matrixInput[51]), .B(n9707), .C(matrixInput[43]), .D(
        n9697), .Z(n10233) );
    VMW_AO22 U604 ( .A(matrixInput[338]), .B(n9707), .C(matrixInput[330]), .D(
        n9697), .Z(n9946) );
    VMW_FD \vectorInput_reg[33]  ( .D(n10307), .CP(Clk), .Q(vectorInput[33])
         );
    VMW_AO22 U623 ( .A(matrixInput[321]), .B(n9707), .C(matrixInput[313]), .D(
        n9697), .Z(n9963) );
    VMW_AO22 U794 ( .A(matrixInput[23]), .B(n9707), .C(matrixInput[15]), .D(
        n9697), .Z(n10261) );
    VMW_FD \matrixInput_reg[83]  ( .D(n10193), .CP(Clk), .Q(matrixInput[83])
         );
    VMW_AO22 U513 ( .A(matrixInput[420]), .B(n9707), .C(matrixInput[412]), .D(
        n9697), .Z(n9864) );
    VMW_AO22 U295 ( .A(DataIn[2]), .B(n9706), .C(vectorInput[58]), .D(n9696), 
        .Z(n10282) );
    VMW_AO22 U389 ( .A(matrixInput[71]), .B(n9707), .C(matrixInput[63]), .D(
        n9697), .Z(n10213) );
    VMW_AO22 U408 ( .A(DataIn[3]), .B(n9707), .C(matrixInput[507]), .D(n9697), 
        .Z(n9769) );
    VMW_AO22 U738 ( .A(matrixInput[28]), .B(n9707), .C(matrixInput[20]), .D(
        n9697), .Z(n10256) );
    VMW_FD \matrixInput_reg[484]  ( .D(n9792), .CP(Clk), .Q(matrixInput[484])
         );
    VMW_FD \matrixInput_reg[330]  ( .D(n9946), .CP(Clk), .Q(matrixInput[330])
         );
    VMW_FD \matrixInput_reg[329]  ( .D(n9947), .CP(Clk), .Q(matrixInput[329])
         );
    VMW_FD \matrixInput_reg[303]  ( .D(n9973), .CP(Clk), .Q(matrixInput[303])
         );
    VMW_FD \holder_reg[5]  ( .D(n10343), .CP(Clk), .Q(\holder[5] ) );
    VMW_AO22 U598 ( .A(matrixInput[344]), .B(n9707), .C(matrixInput[336]), .D(
        n9697), .Z(n9940) );
    VMW_FD \matrixInput_reg[293]  ( .D(n9983), .CP(Clk), .Q(matrixInput[293])
         );
    VMW_FD \matrixInput_reg[190]  ( .D(n10086), .CP(Clk), .Q(matrixInput[190])
         );
    VMW_FD \matrixInput_reg[189]  ( .D(n10087), .CP(Clk), .Q(matrixInput[189])
         );
    VMW_AO22 U305 ( .A(vectorInput[57]), .B(n9706), .C(vectorInput[49]), .D(
        n9696), .Z(n10291) );
    VMW_AO22 U514 ( .A(matrixInput[419]), .B(n9707), .C(matrixInput[411]), .D(
        n9697), .Z(n9865) );
    VMW_AO22 U322 ( .A(vectorInput[41]), .B(n9706), .C(vectorInput[33]), .D(
        n9696), .Z(n10307) );
    VMW_AO22 U484 ( .A(matrixInput[447]), .B(n9707), .C(matrixInput[439]), .D(
        n9697), .Z(n9837) );
    VMW_AO22 U603 ( .A(matrixInput[339]), .B(n9707), .C(matrixInput[331]), .D(
        n9697), .Z(n9945) );
    VMW_AO22 U624 ( .A(matrixInput[320]), .B(n9707), .C(matrixInput[312]), .D(
        n9697), .Z(n9964) );
    VMW_AO22 U793 ( .A(matrixInput[168]), .B(n9707), .C(matrixInput[160]), .D(
        n9697), .Z(n10116) );
    VMW_FD \vectorInput_reg[31]  ( .D(n10309), .CP(Clk), .Q(vectorInput[31])
         );
    VMW_FD \vectorInput_reg[28]  ( .D(n10312), .CP(Clk), .Q(vectorInput[28])
         );
    VMW_AO22 U428 ( .A(matrixInput[56]), .B(n9707), .C(matrixInput[48]), .D(
        n9697), .Z(n10228) );
    VMW_AO22 U533 ( .A(matrixInput[403]), .B(n9707), .C(matrixInput[395]), .D(
        n9697), .Z(n9881) );
    VMW_AO22 U688 ( .A(matrixInput[263]), .B(n9707), .C(matrixInput[255]), .D(
        n9697), .Z(n10021) );
    VMW_AO22 U718 ( .A(matrixInput[236]), .B(n9707), .C(matrixInput[228]), .D(
        n9697), .Z(n10048) );
    VMW_BUFIZ U941 ( .A(n9754), .E(RD), .Z(\DataOut[30]1 ) );
    VMW_FD \matrixInput_reg[98]  ( .D(n10178), .CP(Clk), .Q(matrixInput[98])
         );
    VMW_FD \matrixInput_reg[81]  ( .D(n10195), .CP(Clk), .Q(matrixInput[81])
         );
    VMW_FD \matrixInput_reg[486]  ( .D(n9790), .CP(Clk), .Q(matrixInput[486])
         );
    VMW_FD \matrixInput_reg[332]  ( .D(n9944), .CP(Clk), .Q(matrixInput[332])
         );
    VMW_FD \matrixInput_reg[318]  ( .D(n9958), .CP(Clk), .Q(matrixInput[318])
         );
    VMW_FD \matrixInput_reg[301]  ( .D(n9975), .CP(Clk), .Q(matrixInput[301])
         );
    VMW_FD \holder_reg[7]  ( .D(n10341), .CP(Clk), .Q(\holder[7] ) );
    VMW_FD \matrixInput_reg[291]  ( .D(n9985), .CP(Clk), .Q(matrixInput[291])
         );
    VMW_FD \matrixInput_reg[288]  ( .D(n9988), .CP(Clk), .Q(matrixInput[288])
         );
    VMW_FD \matrixInput_reg[192]  ( .D(n10084), .CP(Clk), .Q(matrixInput[192])
         );
    VMW_AO22 U776 ( .A(matrixInput[184]), .B(n9707), .C(matrixInput[176]), .D(
        n9697), .Z(n10100) );
    VMW_OAI211 U270 ( .A(n9671), .B(n9672), .C(n9673), .D(n9674), .Z(n10348)
         );
    VMW_AO22 U446 ( .A(matrixInput[481]), .B(n9707), .C(matrixInput[473]), .D(
        n9697), .Z(n9803) );
    VMW_AO22 U461 ( .A(matrixInput[53]), .B(n9707), .C(matrixInput[45]), .D(
        n9697), .Z(n10231) );
    VMW_AO22 U834 ( .A(matrixInput[131]), .B(n9707), .C(matrixInput[123]), .D(
        n9697), .Z(n10153) );
    VMW_NOR2 U279 ( .A(Addr[1]), .B(Addr[2]), .Z(n9698) );
    VMW_AO22 U339 ( .A(vectorInput[26]), .B(n9706), .C(vectorInput[18]), .D(
        n9696), .Z(n10322) );
    VMW_AO22 U357 ( .A(matrixInput[100]), .B(n9707), .C(matrixInput[92]), .D(
        n9697), .Z(n10184) );
    VMW_AO22 U370 ( .A(matrixInput[88]), .B(n9707), .C(matrixInput[80]), .D(
        n9697), .Z(n10196) );
    VMW_AO22 U651 ( .A(matrixInput[297]), .B(n9707), .C(matrixInput[289]), .D(
        n9697), .Z(n9987) );
    VMW_AO22 U751 ( .A(matrixInput[207]), .B(n9707), .C(matrixInput[199]), .D(
        n9697), .Z(n10077) );
    VMW_AO22 U813 ( .A(matrixInput[150]), .B(n9707), .C(matrixInput[142]), .D(
        n9697), .Z(n10134) );
    VMW_FD \matrixInput_reg[53]  ( .D(n10223), .CP(Clk), .Q(matrixInput[53])
         );
    VMW_FD \matrixInput_reg[79]  ( .D(n10197), .CP(Clk), .Q(matrixInput[79])
         );
    VMW_FD \matrixInput_reg[60]  ( .D(n10216), .CP(Clk), .Q(matrixInput[60])
         );
    VMW_OAI21 U898 ( .A(n9714), .B(n9715), .C(n9705), .Z(n9691) );
    VMW_FD \matrixInput_reg[467]  ( .D(n9809), .CP(Clk), .Q(matrixInput[467])
         );
    VMW_FD \matrixInput_reg[454]  ( .D(n9822), .CP(Clk), .Q(matrixInput[454])
         );
    VMW_OAI21 U908 ( .A(n9734), .B(n9735), .C(n9705), .Z(n9676) );
    VMW_FD \matrixInput_reg[270]  ( .D(n10006), .CP(Clk), .Q(matrixInput[270])
         );
    VMW_FD \matrixInput_reg[269]  ( .D(n10007), .CP(Clk), .Q(matrixInput[269])
         );
    VMW_FD \matrixInput_reg[243]  ( .D(n10033), .CP(Clk), .Q(matrixInput[243])
         );
    VMW_FD \matrixInput_reg[159]  ( .D(n10117), .CP(Clk), .Q(matrixInput[159])
         );
    VMW_FD \matrixInput_reg[140]  ( .D(n10136), .CP(Clk), .Q(matrixInput[140])
         );
    VMW_FD \matrixInput_reg[173]  ( .D(n10103), .CP(Clk), .Q(matrixInput[173])
         );
    VMW_FD \matrixInput_reg[70]  ( .D(n10206), .CP(Clk), .Q(matrixInput[70])
         );
    VMW_FD \matrixInput_reg[69]  ( .D(n10207), .CP(Clk), .Q(matrixInput[69])
         );
    VMW_AO22 U546 ( .A(matrixInput[391]), .B(n9707), .C(matrixInput[383]), .D(
        n9697), .Z(n9893) );
    VMW_AO22 U561 ( .A(matrixInput[44]), .B(n9707), .C(matrixInput[36]), .D(
        n9697), .Z(n10240) );
    VMW_AO22 U883 ( .A(cOutput[42]), .B(n9699), .C(cOutput[10]), .D(n9698), 
        .Z(n9730) );
    VMW_INV U913 ( .A(Addr[0]), .Z(n9704) );
    VMW_FD \matrixInput_reg[43]  ( .D(n10233), .CP(Clk), .Q(matrixInput[43])
         );
    VMW_AO22 U395 ( .A(matrixInput[66]), .B(n9707), .C(matrixInput[58]), .D(
        n9697), .Z(n10218) );
    VMW_AO22 U433 ( .A(matrixInput[493]), .B(n9707), .C(matrixInput[485]), .D(
        n9697), .Z(n9791) );
    VMW_AO22 U676 ( .A(matrixInput[274]), .B(n9707), .C(matrixInput[266]), .D(
        n9697), .Z(n10010) );
    VMW_BUFIZ U934 ( .A(n9749), .E(RD), .Z(\DataOut[31] ) );
    VMW_AO22 U808 ( .A(matrixInput[155]), .B(n9707), .C(matrixInput[147]), .D(
        n9697), .Z(n10129) );
    VMW_FD \matrixInput_reg[279]  ( .D(n9997), .CP(Clk), .Q(matrixInput[279])
         );
    VMW_FD \matrixInput_reg[260]  ( .D(n10016), .CP(Clk), .Q(matrixInput[260])
         );
    VMW_FD \matrixInput_reg[163]  ( .D(n10113), .CP(Clk), .Q(matrixInput[163])
         );
    VMW_FD \matrixInput_reg[477]  ( .D(n9799), .CP(Clk), .Q(matrixInput[477])
         );
    VMW_FD \matrixInput_reg[253]  ( .D(n10023), .CP(Clk), .Q(matrixInput[253])
         );
    VMW_FD \matrixInput_reg[150]  ( .D(n10126), .CP(Clk), .Q(matrixInput[150])
         );
    VMW_FD \matrixInput_reg[149]  ( .D(n10127), .CP(Clk), .Q(matrixInput[149])
         );
    VMW_FD \matrixInput_reg[444]  ( .D(n9832), .CP(Clk), .Q(matrixInput[444])
         );
    VMW_FD \matrixInput_reg[91]  ( .D(n10185), .CP(Clk), .Q(matrixInput[91])
         );
    VMW_FD \matrixInput_reg[88]  ( .D(n10188), .CP(Clk), .Q(matrixInput[88])
         );
    VMW_AO22 U584 ( .A(matrixInput[357]), .B(n9707), .C(matrixInput[349]), .D(
        n9697), .Z(n9927) );
    VMW_AO22 U693 ( .A(matrixInput[258]), .B(n9707), .C(matrixInput[250]), .D(
        n9697), .Z(n10026) );
    VMW_AO22 U703 ( .A(matrixInput[249]), .B(n9707), .C(matrixInput[241]), .D(
        n9697), .Z(n10035) );
    VMW_AO22 U841 ( .A(matrixInput[125]), .B(n9707), .C(matrixInput[117]), .D(
        n9697), .Z(n10159) );
    VMW_AO22 U724 ( .A(matrixInput[230]), .B(n9707), .C(matrixInput[222]), .D(
        n9697), .Z(n10054) );
    VMW_FD \vectorInput_reg[38]  ( .D(n10302), .CP(Clk), .Q(vectorInput[38])
         );
    VMW_FD \vectorInput_reg[21]  ( .D(n10319), .CP(Clk), .Q(vectorInput[21])
         );
    VMW_AO22 U414 ( .A(matrixInput[509]), .B(n9707), .C(matrixInput[501]), .D(
        n9697), .Z(n9775) );
    VMW_AO22 U866 ( .A(cOutput[54]), .B(n9702), .C(cOutput[22]), .D(n9701), 
        .Z(n9713) );
    VMW_FD \matrixInput_reg[298]  ( .D(n9978), .CP(Clk), .Q(matrixInput[298])
         );
    VMW_FD \vectorInput_reg[12]  ( .D(n10328), .CP(Clk), .Q(vectorInput[12])
         );
    VMW_FD \matrixInput_reg[281]  ( .D(n9995), .CP(Clk), .Q(matrixInput[281])
         );
    VMW_FD \matrixInput_reg[182]  ( .D(n10094), .CP(Clk), .Q(matrixInput[182])
         );
    VMW_AO22 U387 ( .A(matrixInput[73]), .B(n9707), .C(matrixInput[65]), .D(
        n9697), .Z(n10211) );
    VMW_AO22 U421 ( .A(matrixInput[504]), .B(n9707), .C(matrixInput[496]), .D(
        n9697), .Z(n9780) );
    VMW_AO22 U528 ( .A(matrixInput[47]), .B(n9707), .C(matrixInput[39]), .D(
        n9697), .Z(n10237) );
    VMW_FD \matrixInput_reg[506]  ( .D(n9770), .CP(Clk), .Q(matrixInput[506])
         );
    VMW_AO22 U618 ( .A(matrixInput[326]), .B(n9707), .C(matrixInput[318]), .D(
        n9697), .Z(n9958) );
    VMW_AO22 U788 ( .A(matrixInput[173]), .B(n9707), .C(matrixInput[165]), .D(
        n9697), .Z(n10111) );
    VMW_AO22 U853 ( .A(matrixInput[114]), .B(n9707), .C(matrixInput[106]), .D(
        n9697), .Z(n10170) );
    VMW_BUFIZ U948 ( .A(n9760), .E(RD), .Z(\DataOut[15]1 ) );
    VMW_FD \matrixInput_reg[496]  ( .D(n9780), .CP(Clk), .Q(matrixInput[496])
         );
    VMW_FD \matrixInput_reg[322]  ( .D(n9954), .CP(Clk), .Q(matrixInput[322])
         );
    VMW_FD \matrixInput_reg[311]  ( .D(n9965), .CP(Clk), .Q(matrixInput[311])
         );
    VMW_FD \matrixInput_reg[308]  ( .D(n9968), .CP(Clk), .Q(matrixInput[308])
         );
    VMW_FD \matrixInput_reg[247]  ( .D(n10029), .CP(Clk), .Q(matrixInput[247])
         );
    VMW_FD \matrixInput_reg[144]  ( .D(n10132), .CP(Clk), .Q(matrixInput[144])
         );
    VMW_FD \matrixInput_reg[463]  ( .D(n9813), .CP(Clk), .Q(matrixInput[463])
         );
    VMW_FD \matrixInput_reg[450]  ( .D(n9826), .CP(Clk), .Q(matrixInput[450])
         );
    VMW_FD \matrixInput_reg[274]  ( .D(n10002), .CP(Clk), .Q(matrixInput[274])
         );
    VMW_FD \matrixInput_reg[177]  ( .D(n10099), .CP(Clk), .Q(matrixInput[177])
         );
    VMW_FD \matrixInput_reg[449]  ( .D(n9827), .CP(Clk), .Q(matrixInput[449])
         );
    VMW_FD \matrixInput_reg[57]  ( .D(n10219), .CP(Clk), .Q(matrixInput[57])
         );
    VMW_AO22 U681 ( .A(matrixInput[269]), .B(n9707), .C(matrixInput[261]), .D(
        n9697), .Z(n10015) );
    VMW_AO22 U711 ( .A(matrixInput[242]), .B(n9707), .C(matrixInput[234]), .D(
        n9697), .Z(n10042) );
    VMW_AO22 U736 ( .A(matrixInput[219]), .B(n9707), .C(matrixInput[211]), .D(
        n9697), .Z(n10065) );
    VMW_FD \matrixInput_reg[64]  ( .D(n10212), .CP(Clk), .Q(matrixInput[64])
         );
    VMW_AO22 U874 ( .A(cOutput[52]), .B(n9702), .C(cOutput[20]), .D(n9701), 
        .Z(n9721) );
    VMW_AO22 U406 ( .A(DataIn[5]), .B(n9707), .C(matrixInput[509]), .D(n9697), 
        .Z(n9767) );
    VMW_AO22 U596 ( .A(matrixInput[346]), .B(n9707), .C(matrixInput[338]), .D(
        n9697), .Z(n9938) );
    VMW_AO22 U758 ( .A(matrixInput[200]), .B(n9707), .C(matrixInput[192]), .D(
        n9697), .Z(n10084) );
    VMW_FD \holder_reg[3]  ( .D(n10345), .CP(Clk), .Q(\holder[3] ) );
    VMW_AO22 U345 ( .A(vectorInput[20]), .B(n9706), .C(vectorInput[12]), .D(
        n9696), .Z(n10328) );
    VMW_AO22 U362 ( .A(matrixInput[96]), .B(n9707), .C(matrixInput[88]), .D(
        n9697), .Z(n10188) );
    VMW_AO22 U468 ( .A(matrixInput[461]), .B(n9707), .C(matrixInput[453]), .D(
        n9697), .Z(n9823) );
    VMW_AO22 U573 ( .A(matrixInput[367]), .B(n9707), .C(matrixInput[359]), .D(
        n9697), .Z(n9917) );
    VMW_AO22 U643 ( .A(matrixInput[304]), .B(n9707), .C(matrixInput[296]), .D(
        n9697), .Z(n9980) );
    VMW_FD \matrixInput_reg[482]  ( .D(n9794), .CP(Clk), .Q(matrixInput[482])
         );
    VMW_FD \matrixInput_reg[336]  ( .D(n9940), .CP(Clk), .Q(matrixInput[336])
         );
    VMW_FD \matrixInput_reg[295]  ( .D(n9981), .CP(Clk), .Q(matrixInput[295])
         );
    VMW_FD \matrixInput_reg[196]  ( .D(n10080), .CP(Clk), .Q(matrixInput[196])
         );
    VMW_FD \matrixInput_reg[305]  ( .D(n9971), .CP(Clk), .Q(matrixInput[305])
         );
    VMW_AO22 U891 ( .A(cOutput[40]), .B(n9699), .C(cOutput[8]), .D(n9698), .Z(
        n9738) );
    VMW_OAI21 U901 ( .A(n9720), .B(n9721), .C(n9703), .Z(n9686) );
    VMW_FD \matrixInput_reg[85]  ( .D(n10191), .CP(Clk), .Q(matrixInput[85])
         );
    VMW_BUFIZ U926 ( .A(n9743), .E(RD), .Z(\DataOut[19]1 ) );
    VMW_AO22 U379 ( .A(matrixInput[80]), .B(n9707), .C(matrixInput[72]), .D(
        n9697), .Z(n10204) );
    VMW_AO22 U554 ( .A(matrixInput[384]), .B(n9707), .C(matrixInput[376]), .D(
        n9697), .Z(n9900) );
    VMW_AO22 U568 ( .A(matrixInput[371]), .B(n9707), .C(matrixInput[363]), .D(
        n9697), .Z(n9913) );
    VMW_AO22 U664 ( .A(matrixInput[285]), .B(n9707), .C(matrixInput[277]), .D(
        n9697), .Z(n9999) );
    VMW_FD \vectorInput_reg[35]  ( .D(n10305), .CP(Clk), .Q(vectorInput[35])
         );
    VMW_FD \matrixInput_reg[502]  ( .D(n9774), .CP(Clk), .Q(matrixInput[502])
         );
    VMW_FD \matrixInput_reg[492]  ( .D(n9784), .CP(Clk), .Q(matrixInput[492])
         );
    VMW_FD \matrixInput_reg[315]  ( .D(n9961), .CP(Clk), .Q(matrixInput[315])
         );
    VMW_FD \matrixInput_reg[326]  ( .D(n9950), .CP(Clk), .Q(matrixInput[326])
         );
    VMW_AO22 U454 ( .A(matrixInput[474]), .B(n9707), .C(matrixInput[466]), .D(
        n9697), .Z(n9810) );
    VMW_AO22 U658 ( .A(matrixInput[290]), .B(n9707), .C(matrixInput[282]), .D(
        n9697), .Z(n9994) );
    VMW_FD \matrixInput_reg[285]  ( .D(n9991), .CP(Clk), .Q(matrixInput[285])
         );
    VMW_FD \matrixInput_reg[186]  ( .D(n10090), .CP(Clk), .Q(matrixInput[186])
         );
    VMW_AO22 U764 ( .A(matrixInput[195]), .B(n9707), .C(matrixInput[187]), .D(
        n9697), .Z(n10089) );
    VMW_FD \vectorInput_reg[25]  ( .D(n10315), .CP(Clk), .Q(vectorInput[25])
         );
    VMW_AO22 U826 ( .A(matrixInput[138]), .B(n9707), .C(matrixInput[130]), .D(
        n9697), .Z(n10146) );
    VMW_FD \vectorInput_reg[16]  ( .D(n10324), .CP(Clk), .Q(vectorInput[16])
         );
    VMW_PULLDOWN U262 ( .Z(n9760) );
    VMW_AO22 U801 ( .A(matrixInput[161]), .B(n9707), .C(matrixInput[153]), .D(
        n9697), .Z(n10123) );
    VMW_AO22 U473 ( .A(matrixInput[457]), .B(n9707), .C(matrixInput[449]), .D(
        n9697), .Z(n9827) );
    VMW_AO22 U743 ( .A(matrixInput[213]), .B(n9707), .C(matrixInput[205]), .D(
        n9697), .Z(n10071) );
    VMW_FD \matrixInput_reg[95]  ( .D(n10181), .CP(Clk), .Q(matrixInput[95])
         );
    VMW_FD \matrixInput_reg[473]  ( .D(n9803), .CP(Clk), .Q(matrixInput[473])
         );
    VMW_FD \matrixInput_reg[459]  ( .D(n9817), .CP(Clk), .Q(matrixInput[459])
         );
    VMW_FD \matrixInput_reg[440]  ( .D(n9836), .CP(Clk), .Q(matrixInput[440])
         );
    VMW_FD \matrixInput_reg[264]  ( .D(n10012), .CP(Clk), .Q(matrixInput[264])
         );
    VMW_PULLDOWN U246 ( .Z(n9744) );
    VMW_PULLDOWN U247 ( .Z(n9745) );
    VMW_PULLDOWN U255 ( .Z(n9753) );
    VMW_PULLDOWN U269 ( .Z(Logic01) );
    VMW_AO22 U287 ( .A(vectorInput[15]), .B(n9706), .C(vectorInput[7]), .D(
        n9696), .Z(n10333) );
    VMW_AO22 U317 ( .A(vectorInput[46]), .B(n9706), .C(vectorInput[38]), .D(
        n9696), .Z(n10302) );
    VMW_AO22 U848 ( .A(matrixInput[118]), .B(n9707), .C(matrixInput[110]), .D(
        n9697), .Z(n10166) );
    VMW_FD \matrixInput_reg[257]  ( .D(n10019), .CP(Clk), .Q(matrixInput[257])
         );
    VMW_FD \matrixInput_reg[167]  ( .D(n10109), .CP(Clk), .Q(matrixInput[167])
         );
    VMW_FD \matrixInput_reg[154]  ( .D(n10122), .CP(Clk), .Q(matrixInput[154])
         );
    VMW_AO22 U496 ( .A(matrixInput[436]), .B(n9707), .C(matrixInput[428]), .D(
        n9697), .Z(n9848) );
    VMW_AO22 U330 ( .A(vectorInput[34]), .B(n9706), .C(vectorInput[26]), .D(
        n9696), .Z(n10314) );
    VMW_AO22 U506 ( .A(matrixInput[427]), .B(n9707), .C(matrixInput[419]), .D(
        n9697), .Z(n9857) );
    VMW_AO22 U521 ( .A(matrixInput[413]), .B(n9707), .C(matrixInput[405]), .D(
        n9697), .Z(n9871) );
    VMW_AO22 U611 ( .A(matrixInput[332]), .B(n9707), .C(matrixInput[324]), .D(
        n9697), .Z(n9952) );
    VMW_AO22 U636 ( .A(matrixInput[309]), .B(n9707), .C(matrixInput[301]), .D(
        n9697), .Z(n9975) );
    VMW_AO22 U781 ( .A(matrixInput[179]), .B(n9707), .C(matrixInput[171]), .D(
        n9697), .Z(n10105) );
    VMW_BUFIZ U953 ( .A(n9763), .E(RD), .Z(\DataOut[11]1 ) );
    VMW_FD \matrixInput_reg[74]  ( .D(n10202), .CP(Clk), .Q(matrixInput[74])
         );
    VMW_FD \matrixInput_reg[47]  ( .D(n10229), .CP(Clk), .Q(matrixInput[47])
         );
    VMW_AO22 U397 ( .A(matrixInput[64]), .B(n9707), .C(matrixInput[56]), .D(
        n9697), .Z(n10220) );
    VMW_AO22 U586 ( .A(matrixInput[355]), .B(n9707), .C(matrixInput[347]), .D(
        n9697), .Z(n9929) );
    VMW_AO22 U726 ( .A(matrixInput[228]), .B(n9707), .C(matrixInput[220]), .D(
        n9697), .Z(n10056) );
    VMW_FD \matrixInput_reg[462]  ( .D(n9814), .CP(Clk), .Q(matrixInput[462])
         );
    VMW_FD \matrixInput_reg[451]  ( .D(n9825), .CP(Clk), .Q(matrixInput[451])
         );
    VMW_FD \matrixInput_reg[448]  ( .D(n9828), .CP(Clk), .Q(matrixInput[448])
         );
    VMW_FD \matrixInput_reg[275]  ( .D(n10001), .CP(Clk), .Q(matrixInput[275])
         );
    VMW_FD \matrixInput_reg[246]  ( .D(n10030), .CP(Clk), .Q(matrixInput[246])
         );
    VMW_FD \matrixInput_reg[145]  ( .D(n10131), .CP(Clk), .Q(matrixInput[145])
         );
    VMW_FD \matrixInput_reg[176]  ( .D(n10100), .CP(Clk), .Q(matrixInput[176])
         );
    VMW_AO22 U864 ( .A(cOutput[63]), .B(n9702), .C(cOutput[31]), .D(n9701), 
        .Z(n9711) );
    VMW_AO22 U416 ( .A(matrixInput[12]), .B(n9707), .C(matrixInput[4]), .D(
        n9697), .Z(n10272) );
    VMW_AO22 U431 ( .A(matrixInput[495]), .B(n9707), .C(matrixInput[487]), .D(
        n9697), .Z(n9789) );
    VMW_AO22 U843 ( .A(matrixInput[123]), .B(n9707), .C(matrixInput[115]), .D(
        n9697), .Z(n10161) );
    VMW_FD \matrixInput_reg[56]  ( .D(n10220), .CP(Clk), .Q(matrixInput[56])
         );
    VMW_AO22 U478 ( .A(matrixInput[452]), .B(n9707), .C(matrixInput[444]), .D(
        n9697), .Z(n9832) );
    VMW_AO22 U691 ( .A(matrixInput[260]), .B(n9707), .C(matrixInput[252]), .D(
        n9697), .Z(n10024) );
    VMW_AO22 U701 ( .A(matrixInput[251]), .B(n9707), .C(matrixInput[243]), .D(
        n9697), .Z(n10033) );
    VMW_AO22 U748 ( .A(matrixInput[208]), .B(n9707), .C(matrixInput[200]), .D(
        n9697), .Z(n10076) );
    VMW_FD \matrixInput_reg[483]  ( .D(n9793), .CP(Clk), .Q(matrixInput[483])
         );
    VMW_FD \matrixInput_reg[337]  ( .D(n9939), .CP(Clk), .Q(matrixInput[337])
         );
    VMW_FD \matrixInput_reg[65]  ( .D(n10211), .CP(Clk), .Q(matrixInput[65])
         );
    VMW_FD \matrixInput_reg[304]  ( .D(n9972), .CP(Clk), .Q(matrixInput[304])
         );
    VMW_FD \holder_reg[2]  ( .D(n10346), .CP(Clk), .Q(\holder[2] ) );
    VMW_FD \matrixInput_reg[294]  ( .D(n9982), .CP(Clk), .Q(matrixInput[294])
         );
    VMW_OAI211 U272 ( .A(n9671), .B(n9678), .C(n9679), .D(n9680), .Z(n10346)
         );
    VMW_AO22 U355 ( .A(matrixInput[102]), .B(n9707), .C(matrixInput[94]), .D(
        n9697), .Z(n10182) );
    VMW_AO22 U544 ( .A(matrixInput[393]), .B(n9707), .C(matrixInput[385]), .D(
        n9697), .Z(n9891) );
    VMW_BUFIZ U936 ( .A(n9751), .E(RD), .Z(\DataOut[12]1 ) );
    VMW_FD \matrixInput_reg[197]  ( .D(n10079), .CP(Clk), .Q(matrixInput[197])
         );
    VMW_AO22 U369 ( .A(matrixInput[89]), .B(n9707), .C(matrixInput[81]), .D(
        n9697), .Z(n10195) );
    VMW_AO22 U372 ( .A(matrixInput[87]), .B(n9707), .C(matrixInput[79]), .D(
        n9697), .Z(n10197) );
    VMW_AO22 U653 ( .A(matrixInput[295]), .B(n9707), .C(matrixInput[287]), .D(
        n9697), .Z(n9989) );
    VMW_AO22 U674 ( .A(matrixInput[276]), .B(n9707), .C(matrixInput[268]), .D(
        n9697), .Z(n10008) );
    VMW_FD \vectorInput_reg[34]  ( .D(n10306), .CP(Clk), .Q(vectorInput[34])
         );
    VMW_AO22 U881 ( .A(cOutput[34]), .B(n9699), .C(cOutput[2]), .D(n9698), .Z(
        n9728) );
    VMW_INV U911 ( .A(n9696), .Z(n9706) );
    VMW_AO22 U563 ( .A(matrixInput[376]), .B(n9707), .C(matrixInput[368]), .D(
        n9697), .Z(n9908) );
    VMW_FD \matrixInput_reg[284]  ( .D(n9992), .CP(Clk), .Q(matrixInput[284])
         );
    VMW_FD \matrixInput_reg[84]  ( .D(n10192), .CP(Clk), .Q(matrixInput[84])
         );
    VMW_AO22 U463 ( .A(matrixInput[466]), .B(n9707), .C(matrixInput[458]), .D(
        n9697), .Z(n9818) );
    VMW_AO22 U578 ( .A(matrixInput[362]), .B(n9707), .C(matrixInput[354]), .D(
        n9697), .Z(n9922) );
    VMW_FD \matrixInput_reg[503]  ( .D(n9773), .CP(Clk), .Q(matrixInput[503])
         );
    VMW_AO22 U648 ( .A(matrixInput[299]), .B(n9707), .C(matrixInput[291]), .D(
        n9697), .Z(n9985) );
    VMW_FD \matrixInput_reg[187]  ( .D(n10089), .CP(Clk), .Q(matrixInput[187])
         );
    VMW_AO22 U811 ( .A(matrixInput[152]), .B(n9707), .C(matrixInput[144]), .D(
        n9697), .Z(n10132) );
    VMW_FD \matrixInput_reg[493]  ( .D(n9783), .CP(Clk), .Q(matrixInput[493])
         );
    VMW_FD \matrixInput_reg[327]  ( .D(n9949), .CP(Clk), .Q(matrixInput[327])
         );
    VMW_FD \matrixInput_reg[314]  ( .D(n9962), .CP(Clk), .Q(matrixInput[314])
         );
    VMW_FD \matrixInput_reg[94]  ( .D(n10182), .CP(Clk), .Q(matrixInput[94])
         );
    VMW_AO22 U753 ( .A(matrixInput[205]), .B(n9707), .C(matrixInput[197]), .D(
        n9697), .Z(n10079) );
    VMW_AO22 U774 ( .A(matrixInput[186]), .B(n9707), .C(matrixInput[178]), .D(
        n9697), .Z(n10098) );
    VMW_AO22 U836 ( .A(matrixInput[129]), .B(n9707), .C(matrixInput[121]), .D(
        n9697), .Z(n10155) );
    VMW_FD \vectorInput_reg[24]  ( .D(n10316), .CP(Clk), .Q(vectorInput[24])
         );
    VMW_PULLDOWN U260 ( .Z(n9758) );
    VMW_AO22 U285 ( .A(vectorInput[17]), .B(n9706), .C(vectorInput[9]), .D(
        n9696), .Z(n10331) );
    VMW_AO22 U297 ( .A(DataIn[0]), .B(n9706), .C(vectorInput[56]), .D(n9696), 
        .Z(n10284) );
    VMW_AO22 U320 ( .A(vectorInput[43]), .B(n9706), .C(vectorInput[35]), .D(
        n9696), .Z(n10305) );
    VMW_AO22 U444 ( .A(matrixInput[483]), .B(n9707), .C(matrixInput[475]), .D(
        n9697), .Z(n9801) );
    VMW_AO22 U601 ( .A(matrixInput[341]), .B(n9707), .C(matrixInput[333]), .D(
        n9697), .Z(n9943) );
    VMW_AO22 U791 ( .A(matrixInput[170]), .B(n9707), .C(matrixInput[162]), .D(
        n9697), .Z(n10114) );
    VMW_AO22 U858 ( .A(matrixInput[109]), .B(n9707), .C(matrixInput[101]), .D(
        n9697), .Z(n10175) );
    VMW_FD \matrixInput_reg[265]  ( .D(n10011), .CP(Clk), .Q(matrixInput[265])
         );
    VMW_FD \matrixInput_reg[166]  ( .D(n10110), .CP(Clk), .Q(matrixInput[166])
         );
    VMW_FD \vectorInput_reg[17]  ( .D(n10323), .CP(Clk), .Q(vectorInput[17])
         );
    VMW_FD \matrixInput_reg[155]  ( .D(n10121), .CP(Clk), .Q(matrixInput[155])
         );
    VMW_FD \matrixInput_reg[472]  ( .D(n9804), .CP(Clk), .Q(matrixInput[472])
         );
    VMW_FD \matrixInput_reg[256]  ( .D(n10020), .CP(Clk), .Q(matrixInput[256])
         );
    VMW_FD \matrixInput_reg[458]  ( .D(n9818), .CP(Clk), .Q(matrixInput[458])
         );
    VMW_FD \matrixInput_reg[441]  ( .D(n9835), .CP(Clk), .Q(matrixInput[441])
         );
    VMW_BUFIZ U943 ( .A(n9756), .E(RD), .Z(\DataOut[20]1 ) );
    VMW_FD \matrixInput_reg[75]  ( .D(n10201), .CP(Clk), .Q(matrixInput[75])
         );
    VMW_FD \matrixInput_reg[46]  ( .D(n10230), .CP(Clk), .Q(matrixInput[46])
         );
    VMW_AO22 U531 ( .A(matrixInput[405]), .B(n9707), .C(matrixInput[397]), .D(
        n9697), .Z(n9879) );
    VMW_AO22 U307 ( .A(vectorInput[55]), .B(n9706), .C(vectorInput[47]), .D(
        n9696), .Z(n10293) );
    VMW_AO22 U516 ( .A(matrixInput[48]), .B(n9707), .C(matrixInput[40]), .D(
        n9697), .Z(n10236) );
    VMW_AO22 U315 ( .A(vectorInput[11]), .B(n9706), .C(vectorInput[3]), .D(
        n9696), .Z(n10337) );
    VMW_AO22 U332 ( .A(vectorInput[32]), .B(n9706), .C(vectorInput[24]), .D(
        n9696), .Z(n10316) );
    VMW_AO22 U486 ( .A(matrixInput[445]), .B(n9707), .C(matrixInput[437]), .D(
        n9697), .Z(n9839) );
    VMW_AO22 U523 ( .A(matrixInput[411]), .B(n9707), .C(matrixInput[403]), .D(
        n9697), .Z(n9873) );
    VMW_AO22 U613 ( .A(matrixInput[330]), .B(n9707), .C(matrixInput[322]), .D(
        n9697), .Z(n9954) );
    VMW_AO22 U626 ( .A(matrixInput[318]), .B(n9707), .C(matrixInput[310]), .D(
        n9697), .Z(n9966) );
    VMW_AO22 U783 ( .A(matrixInput[24]), .B(n9707), .C(matrixInput[16]), .D(
        n9697), .Z(n10260) );
    VMW_FD \matrixInput_reg[99]  ( .D(n10177), .CP(Clk), .Q(matrixInput[99])
         );
    VMW_FD \matrixInput_reg[80]  ( .D(n10196), .CP(Clk), .Q(matrixInput[80])
         );
    VMW_BUFIZ U951 ( .A(n9761), .E(RD), .Z(\DataOut[22]1 ) );
    VMW_AO22 U494 ( .A(matrixInput[50]), .B(n9707), .C(matrixInput[42]), .D(
        n9697), .Z(n10234) );
    VMW_AO22 U438 ( .A(matrixInput[488]), .B(n9707), .C(matrixInput[480]), .D(
        n9697), .Z(n9796) );
    VMW_AO22 U504 ( .A(matrixInput[428]), .B(n9707), .C(matrixInput[420]), .D(
        n9697), .Z(n9856) );
    VMW_AO22 U634 ( .A(matrixInput[311]), .B(n9707), .C(matrixInput[303]), .D(
        n9697), .Z(n9973) );
    VMW_FD \vectorInput_reg[30]  ( .D(n10310), .CP(Clk), .Q(vectorInput[30])
         );
    VMW_FD \vectorInput_reg[29]  ( .D(n10311), .CP(Clk), .Q(vectorInput[29])
         );
    VMW_AO22 U698 ( .A(matrixInput[254]), .B(n9707), .C(matrixInput[246]), .D(
        n9697), .Z(n10030) );
    VMW_AO22 U708 ( .A(matrixInput[245]), .B(n9707), .C(matrixInput[237]), .D(
        n9697), .Z(n10039) );
    VMW_FD \matrixInput_reg[193]  ( .D(n10083), .CP(Clk), .Q(matrixInput[193])
         );
    VMW_FD \holder_reg[6]  ( .D(n10342), .CP(Clk), .Q(\holder[6] ) );
    VMW_FD \matrixInput_reg[487]  ( .D(n9789), .CP(Clk), .Q(matrixInput[487])
         );
    VMW_FD \matrixInput_reg[333]  ( .D(n9943), .CP(Clk), .Q(matrixInput[333])
         );
    VMW_FD \matrixInput_reg[290]  ( .D(n9986), .CP(Clk), .Q(matrixInput[290])
         );
    VMW_FD \matrixInput_reg[289]  ( .D(n9987), .CP(Clk), .Q(matrixInput[289])
         );
    VMW_FD \matrixInput_reg[319]  ( .D(n9957), .CP(Clk), .Q(matrixInput[319])
         );
    VMW_FD \matrixInput_reg[300]  ( .D(n9976), .CP(Clk), .Q(matrixInput[300])
         );
    VMW_AO22 U456 ( .A(matrixInput[472]), .B(n9707), .C(matrixInput[464]), .D(
        n9697), .Z(n9812) );
    VMW_AO22 U471 ( .A(matrixInput[458]), .B(n9707), .C(matrixInput[450]), .D(
        n9697), .Z(n9826) );
    VMW_AO22 U741 ( .A(matrixInput[215]), .B(n9707), .C(matrixInput[207]), .D(
        n9697), .Z(n10069) );
    VMW_AO22 U803 ( .A(matrixInput[159]), .B(n9707), .C(matrixInput[151]), .D(
        n9697), .Z(n10125) );
    VMW_FD \matrixInput_reg[78]  ( .D(n10198), .CP(Clk), .Q(matrixInput[78])
         );
    VMW_FD \matrixInput_reg[52]  ( .D(n10224), .CP(Clk), .Q(matrixInput[52])
         );
    VMW_FD \matrixInput_reg[61]  ( .D(n10215), .CP(Clk), .Q(matrixInput[61])
         );
    VMW_AO22 U766 ( .A(matrixInput[193]), .B(n9707), .C(matrixInput[185]), .D(
        n9697), .Z(n10091) );
    VMW_PULLDOWN U248 ( .Z(n9746) );
    VMW_PULLDOWN U249 ( .Z(n9747) );
    VMW_PULLDOWN U252 ( .Z(n9750) );
    VMW_PULLDOWN U267 ( .Z(n10349) );
    VMW_AO22 U299 ( .A(vectorInput[62]), .B(n9706), .C(vectorInput[54]), .D(
        n9696), .Z(n10286) );
    VMW_AO22 U329 ( .A(vectorInput[35]), .B(n9706), .C(vectorInput[27]), .D(
        n9696), .Z(n10313) );
    VMW_AO22 U347 ( .A(vectorInput[18]), .B(n9706), .C(vectorInput[10]), .D(
        n9696), .Z(n10330) );
    VMW_AO22 U824 ( .A(matrixInput[140]), .B(n9707), .C(matrixInput[132]), .D(
        n9697), .Z(n10144) );
    VMW_AO22 U888 ( .A(cOutput[57]), .B(n9702), .C(cOutput[25]), .D(n9701), 
        .Z(n9735) );
    VMW_INV U918 ( .A(\holder[7] ), .Z(n9693) );
    VMW_FD \matrixInput_reg[242]  ( .D(n10034), .CP(Clk), .Q(matrixInput[242])
         );
    VMW_FD \matrixInput_reg[466]  ( .D(n9810), .CP(Clk), .Q(matrixInput[466])
         );
    VMW_FD \matrixInput_reg[455]  ( .D(n9821), .CP(Clk), .Q(matrixInput[455])
         );
    VMW_FD \matrixInput_reg[271]  ( .D(n10005), .CP(Clk), .Q(matrixInput[271])
         );
    VMW_FD \matrixInput_reg[158]  ( .D(n10118), .CP(Clk), .Q(matrixInput[158])
         );
    VMW_FD \matrixInput_reg[141]  ( .D(n10135), .CP(Clk), .Q(matrixInput[141])
         );
    VMW_FD \matrixInput_reg[268]  ( .D(n10008), .CP(Clk), .Q(matrixInput[268])
         );
    VMW_FD \matrixInput_reg[172]  ( .D(n10104), .CP(Clk), .Q(matrixInput[172])
         );
    VMW_AO22 U360 ( .A(matrixInput[16]), .B(n9707), .C(matrixInput[8]), .D(
        n9697), .Z(n10268) );
    VMW_AO22 U556 ( .A(matrixInput[382]), .B(n9707), .C(matrixInput[374]), .D(
        n9697), .Z(n9902) );
    VMW_AO22 U571 ( .A(matrixInput[368]), .B(n9707), .C(matrixInput[360]), .D(
        n9697), .Z(n9916) );
    VMW_AO22 U641 ( .A(matrixInput[306]), .B(n9707), .C(matrixInput[298]), .D(
        n9697), .Z(n9978) );
    VMW_AO22 U666 ( .A(matrixInput[283]), .B(n9707), .C(matrixInput[275]), .D(
        n9697), .Z(n10001) );
    VMW_BUFIZ U924 ( .A(n9741), .E(RD), .Z(\DataOut[27]1 ) );
    VMW_FD \matrixInput_reg[71]  ( .D(n10205), .CP(Clk), .Q(matrixInput[71])
         );
    VMW_FD \matrixInput_reg[68]  ( .D(n10208), .CP(Clk), .Q(matrixInput[68])
         );
    VMW_AO22 U385 ( .A(matrixInput[75]), .B(n9707), .C(matrixInput[67]), .D(
        n9697), .Z(n10209) );
    VMW_AO22 U734 ( .A(matrixInput[221]), .B(n9707), .C(matrixInput[213]), .D(
        n9697), .Z(n10063) );
    VMW_AO22 U818 ( .A(matrixInput[146]), .B(n9707), .C(matrixInput[138]), .D(
        n9697), .Z(n10138) );
    VMW_OR3 U893 ( .A(Addr[1]), .B(Addr[0]), .C(n9740), .Z(n9697) );
    VMW_OAI21 U903 ( .A(n9724), .B(n9725), .C(n9703), .Z(n9683) );
    VMW_FD \matrixInput_reg[42]  ( .D(n10234), .CP(Clk), .Q(matrixInput[42])
         );
    VMW_FD \matrixInput_reg[476]  ( .D(n9800), .CP(Clk), .Q(matrixInput[476])
         );
    VMW_FD \matrixInput_reg[445]  ( .D(n9831), .CP(Clk), .Q(matrixInput[445])
         );
    VMW_FD \matrixInput_reg[278]  ( .D(n9998), .CP(Clk), .Q(matrixInput[278])
         );
    VMW_FD \matrixInput_reg[261]  ( .D(n10015), .CP(Clk), .Q(matrixInput[261])
         );
    VMW_FD \matrixInput_reg[252]  ( .D(n10024), .CP(Clk), .Q(matrixInput[252])
         );
    VMW_FD \matrixInput_reg[162]  ( .D(n10114), .CP(Clk), .Q(matrixInput[162])
         );
    VMW_FD \matrixInput_reg[151]  ( .D(n10125), .CP(Clk), .Q(matrixInput[151])
         );
    VMW_FD \matrixInput_reg[148]  ( .D(n10128), .CP(Clk), .Q(matrixInput[148])
         );
    VMW_FD \vectorInput_reg[39]  ( .D(n10301), .CP(Clk), .Q(vectorInput[39])
         );
    VMW_FD \vectorInput_reg[20]  ( .D(n10320), .CP(Clk), .Q(vectorInput[20])
         );
    VMW_FD \vectorInput_reg[13]  ( .D(n10327), .CP(Clk), .Q(vectorInput[13])
         );
    VMW_AO22 U404 ( .A(DataIn[6]), .B(n9707), .C(matrixInput[510]), .D(n9697), 
        .Z(n9766) );
    VMW_AO22 U423 ( .A(matrixInput[502]), .B(n9707), .C(matrixInput[494]), .D(
        n9697), .Z(n9782) );
    VMW_AO22 U594 ( .A(matrixInput[41]), .B(n9707), .C(matrixInput[33]), .D(
        n9697), .Z(n10243) );
    VMW_AO22 U876 ( .A(cOutput[60]), .B(n9702), .C(cOutput[28]), .D(n9701), 
        .Z(n9723) );
    VMW_AO22 U538 ( .A(matrixInput[398]), .B(n9707), .C(matrixInput[390]), .D(
        n9697), .Z(n9886) );
    VMW_AO22 U683 ( .A(matrixInput[33]), .B(n9707), .C(matrixInput[25]), .D(
        n9697), .Z(n10251) );
    VMW_AO22 U851 ( .A(matrixInput[116]), .B(n9707), .C(matrixInput[108]), .D(
        n9697), .Z(n10168) );
    VMW_FD \matrixInput_reg[90]  ( .D(n10186), .CP(Clk), .Q(matrixInput[90])
         );
    VMW_FD \matrixInput_reg[89]  ( .D(n10187), .CP(Clk), .Q(matrixInput[89])
         );
    VMW_AO22 U713 ( .A(matrixInput[240]), .B(n9707), .C(matrixInput[232]), .D(
        n9697), .Z(n10044) );
    VMW_FD \matrixInput_reg[507]  ( .D(n9769), .CP(Clk), .Q(matrixInput[507])
         );
    VMW_FD \matrixInput_reg[497]  ( .D(n9779), .CP(Clk), .Q(matrixInput[497])
         );
    VMW_FD \matrixInput_reg[310]  ( .D(n9966), .CP(Clk), .Q(matrixInput[310])
         );
    VMW_FD \matrixInput_reg[309]  ( .D(n9967), .CP(Clk), .Q(matrixInput[309])
         );
    VMW_FD \matrixInput_reg[323]  ( .D(n9953), .CP(Clk), .Q(matrixInput[323])
         );
    VMW_FD \matrixInput_reg[183]  ( .D(n10093), .CP(Clk), .Q(matrixInput[183])
         );
    VMW_AO22 U382 ( .A(matrixInput[14]), .B(n9707), .C(matrixInput[6]), .D(
        n9697), .Z(n10270) );
    VMW_AO22 U403 ( .A(DataIn[7]), .B(n9707), .C(matrixInput[511]), .D(n9697), 
        .Z(n9765) );
    VMW_AO22 U424 ( .A(matrixInput[501]), .B(n9707), .C(matrixInput[493]), .D(
        n9697), .Z(n9783) );
    VMW_AO22 U608 ( .A(matrixInput[335]), .B(n9707), .C(matrixInput[327]), .D(
        n9697), .Z(n9949) );
    VMW_FD \matrixInput_reg[299]  ( .D(n9977), .CP(Clk), .Q(matrixInput[299])
         );
    VMW_FD \matrixInput_reg[280]  ( .D(n9996), .CP(Clk), .Q(matrixInput[280])
         );
    VMW_AO22 U684 ( .A(matrixInput[267]), .B(n9707), .C(matrixInput[259]), .D(
        n9697), .Z(n10017) );
    VMW_AO22 U714 ( .A(matrixInput[239]), .B(n9707), .C(matrixInput[231]), .D(
        n9697), .Z(n10045) );
    VMW_AO22 U798 ( .A(matrixInput[164]), .B(n9707), .C(matrixInput[156]), .D(
        n9697), .Z(n10120) );
    VMW_AO22 U856 ( .A(matrixInput[111]), .B(n9707), .C(matrixInput[103]), .D(
        n9697), .Z(n10173) );
    VMW_FD \vectorInput_reg[22]  ( .D(n10318), .CP(Clk), .Q(vectorInput[22])
         );
    VMW_AO22 U593 ( .A(matrixInput[348]), .B(n9707), .C(matrixInput[340]), .D(
        n9697), .Z(n9936) );
    VMW_AO22 U871 ( .A(cOutput[45]), .B(n9699), .C(cOutput[13]), .D(n9698), 
        .Z(n9718) );
    VMW_FD \vectorInput_reg[11]  ( .D(n10329), .CP(Clk), .Q(vectorInput[11])
         );
    VMW_FD \matrixInput_reg[92]  ( .D(n10184), .CP(Clk), .Q(matrixInput[92])
         );
    VMW_AO22 U518 ( .A(matrixInput[416]), .B(n9707), .C(matrixInput[408]), .D(
        n9697), .Z(n9868) );
    VMW_AO22 U733 ( .A(matrixInput[222]), .B(n9707), .C(matrixInput[214]), .D(
        n9697), .Z(n10062) );
    VMW_FD \matrixInput_reg[495]  ( .D(n9781), .CP(Clk), .Q(matrixInput[495])
         );
    VMW_FD \matrixInput_reg[338]  ( .D(n9938), .CP(Clk), .Q(matrixInput[338])
         );
    VMW_FD \matrixInput_reg[321]  ( .D(n9955), .CP(Clk), .Q(matrixInput[321])
         );
    VMW_FD \matrixInput_reg[312]  ( .D(n9964), .CP(Clk), .Q(matrixInput[312])
         );
    VMW_FD \matrixInput_reg[282]  ( .D(n9994), .CP(Clk), .Q(matrixInput[282])
         );
    VMW_AO22 U309 ( .A(vectorInput[53]), .B(n9706), .C(vectorInput[45]), .D(
        n9696), .Z(n10295) );
    VMW_AO22 U488 ( .A(matrixInput[443]), .B(n9707), .C(matrixInput[435]), .D(
        n9697), .Z(n9841) );
    VMW_FD \matrixInput_reg[505]  ( .D(n9771), .CP(Clk), .Q(matrixInput[505])
         );
    VMW_AO22 U340 ( .A(vectorInput[25]), .B(n9706), .C(vectorInput[17]), .D(
        n9696), .Z(n10323) );
    VMW_AO22 U367 ( .A(matrixInput[91]), .B(n9707), .C(matrixInput[83]), .D(
        n9697), .Z(n10193) );
    VMW_AO22 U628 ( .A(matrixInput[317]), .B(n9707), .C(matrixInput[309]), .D(
        n9697), .Z(n9967) );
    VMW_FD \matrixInput_reg[198]  ( .D(n10078), .CP(Clk), .Q(matrixInput[198])
         );
    VMW_FD \matrixInput_reg[181]  ( .D(n10095), .CP(Clk), .Q(matrixInput[181])
         );
    VMW_OR3 U894 ( .A(n9740), .B(Addr[1]), .C(n9704), .Z(n9696) );
    VMW_OAI21 U904 ( .A(n9726), .B(n9727), .C(n9705), .Z(n9682) );
    VMW_AO22 U551 ( .A(matrixInput[387]), .B(n9707), .C(matrixInput[379]), .D(
        n9697), .Z(n9897) );
    VMW_AO22 U576 ( .A(matrixInput[364]), .B(n9707), .C(matrixInput[356]), .D(
        n9697), .Z(n9920) );
    VMW_AO22 U646 ( .A(matrixInput[301]), .B(n9707), .C(matrixInput[293]), .D(
        n9697), .Z(n9983) );
    VMW_AO22 U661 ( .A(matrixInput[35]), .B(n9707), .C(matrixInput[27]), .D(
        n9697), .Z(n10249) );
    VMW_INV U923 ( .A(\holder[0] ), .Z(n9672) );
    VMW_FD \matrixInput_reg[73]  ( .D(n10203), .CP(Clk), .Q(matrixInput[73])
         );
    VMW_FD \matrixInput_reg[59]  ( .D(n10217), .CP(Clk), .Q(matrixInput[59])
         );
    VMW_FD \matrixInput_reg[40]  ( .D(n10236), .CP(Clk), .Q(matrixInput[40])
         );
    VMW_AO22 U451 ( .A(matrixInput[477]), .B(n9707), .C(matrixInput[469]), .D(
        n9697), .Z(n9807) );
    VMW_AO22 U823 ( .A(matrixInput[141]), .B(n9707), .C(matrixInput[133]), .D(
        n9697), .Z(n10143) );
    VMW_AO22 U838 ( .A(matrixInput[19]), .B(n9707), .C(matrixInput[11]), .D(
        n9697), .Z(n10265) );
    VMW_FD \matrixInput_reg[474]  ( .D(n9802), .CP(Clk), .Q(matrixInput[474])
         );
    VMW_FD \matrixInput_reg[447]  ( .D(n9829), .CP(Clk), .Q(matrixInput[447])
         );
    VMW_FD \matrixInput_reg[263]  ( .D(n10013), .CP(Clk), .Q(matrixInput[263])
         );
    VMW_FD \matrixInput_reg[179]  ( .D(n10097), .CP(Clk), .Q(matrixInput[179])
         );
    VMW_FD \matrixInput_reg[160]  ( .D(n10116), .CP(Clk), .Q(matrixInput[160])
         );
    VMW_FD \matrixInput_reg[153]  ( .D(n10123), .CP(Clk), .Q(matrixInput[153])
         );
    VMW_FD \matrixInput_reg[250]  ( .D(n10026), .CP(Clk), .Q(matrixInput[250])
         );
    VMW_FD \matrixInput_reg[249]  ( .D(n10027), .CP(Clk), .Q(matrixInput[249])
         );
    VMW_FD \matrixInput_reg[50]  ( .D(n10226), .CP(Clk), .Q(matrixInput[50])
         );
    VMW_FD \matrixInput_reg[49]  ( .D(n10227), .CP(Clk), .Q(matrixInput[49])
         );
    VMW_AO22 U476 ( .A(matrixInput[454]), .B(n9707), .C(matrixInput[446]), .D(
        n9697), .Z(n9830) );
    VMW_AO22 U746 ( .A(matrixInput[210]), .B(n9707), .C(matrixInput[202]), .D(
        n9697), .Z(n10074) );
    VMW_AO22 U761 ( .A(matrixInput[26]), .B(n9707), .C(matrixInput[18]), .D(
        n9697), .Z(n10258) );
    VMW_FD \matrixInput_reg[63]  ( .D(n10213), .CP(Clk), .Q(matrixInput[63])
         );
    VMW_AO22 U804 ( .A(matrixInput[158]), .B(n9707), .C(matrixInput[150]), .D(
        n9697), .Z(n10126) );
    VMW_AND2 U282 ( .A(Addr[1]), .B(Addr[2]), .Z(n9702) );
    VMW_AO22 U503 ( .A(matrixInput[429]), .B(n9707), .C(matrixInput[421]), .D(
        n9697), .Z(n9855) );
    VMW_AO22 U633 ( .A(matrixInput[312]), .B(n9707), .C(matrixInput[304]), .D(
        n9697), .Z(n9972) );
    VMW_BUFIZ U938 ( .A(n9752), .E(RD), .Z(\DataOut[28]1 ) );
    VMW_FD \matrixInput_reg[143]  ( .D(n10133), .CP(Clk), .Q(matrixInput[143])
         );
    VMW_FD \matrixInput_reg[464]  ( .D(n9812), .CP(Clk), .Q(matrixInput[464])
         );
    VMW_FD \matrixInput_reg[457]  ( .D(n9819), .CP(Clk), .Q(matrixInput[457])
         );
    VMW_FD \matrixInput_reg[273]  ( .D(n10003), .CP(Clk), .Q(matrixInput[273])
         );
    VMW_FD \matrixInput_reg[259]  ( .D(n10017), .CP(Clk), .Q(matrixInput[259])
         );
    VMW_FD \matrixInput_reg[240]  ( .D(n10036), .CP(Clk), .Q(matrixInput[240])
         );
    VMW_FD \matrixInput_reg[170]  ( .D(n10106), .CP(Clk), .Q(matrixInput[170])
         );
    VMW_FD \matrixInput_reg[169]  ( .D(n10107), .CP(Clk), .Q(matrixInput[169])
         );
    VMW_AO22 U290 ( .A(DataIn[6]), .B(n9706), .C(vectorInput[62]), .D(n9696), 
        .Z(n10278) );
    VMW_AO22 U300 ( .A(vectorInput[61]), .B(n9706), .C(vectorInput[53]), .D(
        n9696), .Z(n10287) );
    VMW_AO22 U312 ( .A(vectorInput[50]), .B(n9706), .C(vectorInput[42]), .D(
        n9696), .Z(n10298) );
    VMW_AO22 U493 ( .A(matrixInput[438]), .B(n9707), .C(matrixInput[430]), .D(
        n9697), .Z(n9846) );
    VMW_AO22 U335 ( .A(vectorInput[29]), .B(n9706), .C(vectorInput[21]), .D(
        n9696), .Z(n10319) );
    VMW_FD \matrixInput_reg[82]  ( .D(n10194), .CP(Clk), .Q(matrixInput[82])
         );
    VMW_AO22 U399 ( .A(matrixInput[62]), .B(n9707), .C(matrixInput[54]), .D(
        n9697), .Z(n10222) );
    VMW_AO22 U418 ( .A(matrixInput[507]), .B(n9707), .C(matrixInput[499]), .D(
        n9697), .Z(n9777) );
    VMW_AO22 U524 ( .A(matrixInput[410]), .B(n9707), .C(matrixInput[402]), .D(
        n9697), .Z(n9874) );
    VMW_AO22 U588 ( .A(matrixInput[353]), .B(n9707), .C(matrixInput[345]), .D(
        n9697), .Z(n9931) );
    VMW_AO22 U614 ( .A(matrixInput[329]), .B(n9707), .C(matrixInput[321]), .D(
        n9697), .Z(n9955) );
    VMW_AO22 U784 ( .A(matrixInput[177]), .B(n9707), .C(matrixInput[169]), .D(
        n9697), .Z(n10107) );
    VMW_FD \vectorInput_reg[18]  ( .D(n10322), .CP(Clk), .Q(vectorInput[18])
         );
    VMW_AO22 U728 ( .A(matrixInput[227]), .B(n9707), .C(matrixInput[219]), .D(
        n9697), .Z(n10057) );
    VMW_FD \vectorInput_reg[32]  ( .D(n10308), .CP(Clk), .Q(vectorInput[32])
         );
    VMW_FD \holder_reg[4]  ( .D(n10344), .CP(Clk), .Q(\holder[4] ) );
    VMW_FD \matrixInput_reg[292]  ( .D(n9984), .CP(Clk), .Q(matrixInput[292])
         );
    VMW_AO22 U481 ( .A(matrixInput[449]), .B(n9707), .C(matrixInput[441]), .D(
        n9697), .Z(n9835) );
    VMW_AO22 U621 ( .A(matrixInput[323]), .B(n9707), .C(matrixInput[315]), .D(
        n9697), .Z(n9961) );
    VMW_AO22 U878 ( .A(cOutput[51]), .B(n9702), .C(cOutput[19]), .D(n9701), 
        .Z(n9725) );
    VMW_FD \matrixInput_reg[485]  ( .D(n9791), .CP(Clk), .Q(matrixInput[485])
         );
    VMW_FD \matrixInput_reg[331]  ( .D(n9945), .CP(Clk), .Q(matrixInput[331])
         );
    VMW_FD \matrixInput_reg[328]  ( .D(n9948), .CP(Clk), .Q(matrixInput[328])
         );
    VMW_FD \matrixInput_reg[191]  ( .D(n10085), .CP(Clk), .Q(matrixInput[191])
         );
    VMW_FD \matrixInput_reg[188]  ( .D(n10088), .CP(Clk), .Q(matrixInput[188])
         );
    VMW_FD \matrixInput_reg[302]  ( .D(n9974), .CP(Clk), .Q(matrixInput[302])
         );
    VMW_FD \matrixInput_reg[267]  ( .D(n10009), .CP(Clk), .Q(matrixInput[267])
         );
    VMW_FD \matrixInput_reg[254]  ( .D(n10022), .CP(Clk), .Q(matrixInput[254])
         );
    VMW_FD \matrixInput_reg[164]  ( .D(n10112), .CP(Clk), .Q(matrixInput[164])
         );
    VMW_FD \matrixInput_reg[470]  ( .D(n9806), .CP(Clk), .Q(matrixInput[470])
         );
    VMW_FD \matrixInput_reg[157]  ( .D(n10119), .CP(Clk), .Q(matrixInput[157])
         );
    VMW_FD \matrixInput_reg[469]  ( .D(n9807), .CP(Clk), .Q(matrixInput[469])
         );
    VMW_FD \matrixInput_reg[443]  ( .D(n9833), .CP(Clk), .Q(matrixInput[443])
         );
    VMW_FD \matrixInput_reg[77]  ( .D(n10199), .CP(Clk), .Q(matrixInput[77])
         );
    VMW_AO22 U511 ( .A(matrixInput[422]), .B(n9707), .C(matrixInput[414]), .D(
        n9697), .Z(n9862) );
    VMW_AO22 U327 ( .A(vectorInput[37]), .B(n9706), .C(vectorInput[29]), .D(
        n9696), .Z(n10311) );
    VMW_AO22 U536 ( .A(matrixInput[400]), .B(n9707), .C(matrixInput[392]), .D(
        n9697), .Z(n9884) );
    VMW_FD \matrixInput_reg[44]  ( .D(n10232), .CP(Clk), .Q(matrixInput[44])
         );
    VMW_AO22 U349 ( .A(matrixInput[17]), .B(n9707), .C(matrixInput[9]), .D(
        n9697), .Z(n10267) );
    VMW_AO22 U606 ( .A(matrixInput[337]), .B(n9707), .C(matrixInput[329]), .D(
        n9697), .Z(n9947) );
    VMW_BUFIZ U944 ( .A(n9757), .E(RD), .Z(\DataOut[26]1 ) );
    VMW_AO22 U796 ( .A(matrixInput[166]), .B(n9707), .C(matrixInput[158]), .D(
        n9697), .Z(n10118) );
    VMW_FD \matrixInput_reg[185]  ( .D(n10091), .CP(Clk), .Q(matrixInput[185])
         );
    VMW_AO22 U443 ( .A(matrixInput[484]), .B(n9707), .C(matrixInput[476]), .D(
        n9697), .Z(n9800) );
    VMW_AO22 U558 ( .A(matrixInput[380]), .B(n9707), .C(matrixInput[372]), .D(
        n9697), .Z(n9904) );
    VMW_AO22 U668 ( .A(matrixInput[281]), .B(n9707), .C(matrixInput[273]), .D(
        n9697), .Z(n10003) );
    VMW_FD \matrixInput_reg[501]  ( .D(n9775), .CP(Clk), .Q(matrixInput[501])
         );
    VMW_FD \matrixInput_reg[286]  ( .D(n9990), .CP(Clk), .Q(matrixInput[286])
         );
    VMW_FD \matrixInput_reg[491]  ( .D(n9785), .CP(Clk), .Q(matrixInput[491])
         );
    VMW_FD \matrixInput_reg[488]  ( .D(n9788), .CP(Clk), .Q(matrixInput[488])
         );
    VMW_FD \matrixInput_reg[316]  ( .D(n9960), .CP(Clk), .Q(matrixInput[316])
         );
    VMW_FD \matrixInput_reg[325]  ( .D(n9951), .CP(Clk), .Q(matrixInput[325])
         );
    VMW_OAI211 U275 ( .A(n9671), .B(n9687), .C(n9688), .D(n9689), .Z(n10343)
         );
    VMW_AO22 U754 ( .A(matrixInput[204]), .B(n9707), .C(matrixInput[196]), .D(
        n9697), .Z(n10080) );
    VMW_AO22 U773 ( .A(matrixInput[187]), .B(n9707), .C(matrixInput[179]), .D(
        n9697), .Z(n10097) );
    VMW_AO22 U831 ( .A(matrixInput[134]), .B(n9707), .C(matrixInput[126]), .D(
        n9697), .Z(n10150) );
    VMW_FD \matrixInput_reg[96]  ( .D(n10180), .CP(Clk), .Q(matrixInput[96])
         );
    VMW_FD \vectorInput_reg[26]  ( .D(n10314), .CP(Clk), .Q(vectorInput[26])
         );
    VMW_FD \vectorInput_reg[15]  ( .D(n10325), .CP(Clk), .Q(vectorInput[15])
         );
    VMW_AO22 U458 ( .A(matrixInput[470]), .B(n9707), .C(matrixInput[462]), .D(
        n9697), .Z(n9814) );
    VMW_AO22 U464 ( .A(matrixInput[465]), .B(n9707), .C(matrixInput[457]), .D(
        n9697), .Z(n9819) );
    VMW_AO22 U768 ( .A(matrixInput[191]), .B(n9707), .C(matrixInput[183]), .D(
        n9697), .Z(n10093) );
    VMW_AO22 U816 ( .A(matrixInput[21]), .B(n9707), .C(matrixInput[13]), .D(
        n9697), .Z(n10263) );
    VMW_FD \matrixInput_reg[498]  ( .D(n9778), .CP(Clk), .Q(matrixInput[498])
         );
    VMW_FD \matrixInput_reg[481]  ( .D(n9795), .CP(Clk), .Q(matrixInput[481])
         );
    VMW_FD \matrixInput_reg[335]  ( .D(n9941), .CP(Clk), .Q(matrixInput[335])
         );
    VMW_FD \matrixInput_reg[306]  ( .D(n9970), .CP(Clk), .Q(matrixInput[306])
         );
    VMW_FD \matrixInput_reg[195]  ( .D(n10081), .CP(Clk), .Q(matrixInput[195])
         );
    VMW_FD \holder_reg[0]  ( .D(n10348), .CP(Clk), .Q(\holder[0] ) );
    VMW_FD \matrixInput_reg[511]  ( .D(n9765), .CP(Clk), .Q(matrixInput[511])
         );
    VMW_FD \matrixInput_reg[508]  ( .D(n9768), .CP(Clk), .Q(matrixInput[508])
         );
    VMW_PULLDOWN U266 ( .Z(n9764) );
    VMW_AND2 U283 ( .A(n9704), .B(n9671), .Z(n9703) );
    VMW_AO22 U313 ( .A(vectorInput[49]), .B(n9706), .C(vectorInput[41]), .D(
        n9696), .Z(n10299) );
    VMW_AO22 U352 ( .A(matrixInput[105]), .B(n9707), .C(matrixInput[97]), .D(
        n9697), .Z(n10179) );
    VMW_AO22 U375 ( .A(matrixInput[84]), .B(n9707), .C(matrixInput[76]), .D(
        n9697), .Z(n10200) );
    VMW_AO22 U564 ( .A(matrixInput[375]), .B(n9707), .C(matrixInput[367]), .D(
        n9697), .Z(n9909) );
    VMW_FD \matrixInput_reg[296]  ( .D(n9980), .CP(Clk), .Q(matrixInput[296])
         );
    VMW_AO22 U654 ( .A(matrixInput[294]), .B(n9707), .C(matrixInput[286]), .D(
        n9697), .Z(n9990) );
    VMW_AO22 U886 ( .A(cOutput[49]), .B(n9702), .C(cOutput[17]), .D(n9701), 
        .Z(n9733) );
    VMW_INV U916 ( .A(\holder[1] ), .Z(n9675) );
    VMW_FD \vectorInput_reg[36]  ( .D(n10304), .CP(Clk), .Q(vectorInput[36])
         );
    VMW_AO22 U673 ( .A(matrixInput[277]), .B(n9707), .C(matrixInput[269]), .D(
        n9697), .Z(n10007) );
    VMW_FD \matrixInput_reg[86]  ( .D(n10190), .CP(Clk), .Q(matrixInput[86])
         );
    VMW_AO22 U390 ( .A(matrixInput[70]), .B(n9707), .C(matrixInput[62]), .D(
        n9697), .Z(n10214) );
    VMW_AO22 U411 ( .A(DataIn[0]), .B(n9707), .C(matrixInput[504]), .D(n9697), 
        .Z(n9772) );
    VMW_AO22 U436 ( .A(matrixInput[490]), .B(n9707), .C(matrixInput[482]), .D(
        n9697), .Z(n9794) );
    VMW_AO22 U543 ( .A(matrixInput[394]), .B(n9707), .C(matrixInput[386]), .D(
        n9697), .Z(n9890) );
    VMW_AO22 U696 ( .A(matrixInput[256]), .B(n9707), .C(matrixInput[248]), .D(
        n9697), .Z(n10028) );
    VMW_BUFIZ U931 ( .A(\holder[4] ), .E(RD), .Z(\DataOut[4]1 ) );
    VMW_FD \matrixInput_reg[479]  ( .D(n9797), .CP(Clk), .Q(matrixInput[479])
         );
    VMW_FD \matrixInput_reg[453]  ( .D(n9823), .CP(Clk), .Q(matrixInput[453])
         );
    VMW_FD \matrixInput_reg[460]  ( .D(n9816), .CP(Clk), .Q(matrixInput[460])
         );
    VMW_FD \matrixInput_reg[277]  ( .D(n9999), .CP(Clk), .Q(matrixInput[277])
         );
    VMW_FD \matrixInput_reg[244]  ( .D(n10032), .CP(Clk), .Q(matrixInput[244])
         );
    VMW_FD \matrixInput_reg[147]  ( .D(n10129), .CP(Clk), .Q(matrixInput[147])
         );
    VMW_FD \matrixInput_reg[174]  ( .D(n10102), .CP(Clk), .Q(matrixInput[174])
         );
    VMW_AO22 U706 ( .A(matrixInput[247]), .B(n9707), .C(matrixInput[239]), .D(
        n9697), .Z(n10037) );
    VMW_AO22 U844 ( .A(matrixInput[122]), .B(n9707), .C(matrixInput[114]), .D(
        n9697), .Z(n10162) );
    VMW_AO22 U581 ( .A(matrixInput[359]), .B(n9707), .C(matrixInput[351]), .D(
        n9697), .Z(n9925) );
    VMW_AO22 U632 ( .A(matrixInput[313]), .B(n9707), .C(matrixInput[305]), .D(
        n9697), .Z(n9971) );
    VMW_AO22 U721 ( .A(matrixInput[233]), .B(n9707), .C(matrixInput[225]), .D(
        n9697), .Z(n10051) );
    VMW_AO22 U863 ( .A(cOutput[47]), .B(n9699), .C(cOutput[15]), .D(n9698), 
        .Z(n9710) );
    VMW_FD \matrixInput_reg[67]  ( .D(n10209), .CP(Clk), .Q(matrixInput[67])
         );
    VMW_FD \matrixInput_reg[54]  ( .D(n10222), .CP(Clk), .Q(matrixInput[54])
         );
    VMW_AO22 U492 ( .A(matrixInput[439]), .B(n9707), .C(matrixInput[431]), .D(
        n9697), .Z(n9845) );
    VMW_AO22 U334 ( .A(vectorInput[30]), .B(n9706), .C(vectorInput[22]), .D(
        n9696), .Z(n10318) );
    VMW_AO22 U502 ( .A(matrixInput[430]), .B(n9707), .C(matrixInput[422]), .D(
        n9697), .Z(n9854) );
    VMW_AO22 U525 ( .A(matrixInput[409]), .B(n9707), .C(matrixInput[401]), .D(
        n9697), .Z(n9875) );
    VMW_FD \matrixInput_reg[9]  ( .D(n10267), .CP(Clk), .Q(matrixInput[9]) );
    VMW_FD \vectorInput_reg[60]  ( .D(n10280), .CP(Clk), .Q(vectorInput[60])
         );
    VMW_AO22 U398 ( .A(matrixInput[63]), .B(n9707), .C(matrixInput[55]), .D(
        n9697), .Z(n10221) );
    VMW_AO22 U615 ( .A(matrixInput[328]), .B(n9707), .C(matrixInput[320]), .D(
        n9697), .Z(n9956) );
    VMW_FD \vectorInput_reg[53]  ( .D(n10287), .CP(Clk), .Q(vectorInput[53])
         );
    VMW_AO22 U729 ( .A(matrixInput[226]), .B(n9707), .C(matrixInput[218]), .D(
        n9697), .Z(n10058) );
    VMW_AO22 U785 ( .A(matrixInput[176]), .B(n9707), .C(matrixInput[168]), .D(
        n9697), .Z(n10108) );
    VMW_AO22 U419 ( .A(matrixInput[506]), .B(n9707), .C(matrixInput[498]), .D(
        n9697), .Z(n9778) );
    VMW_AO22 U450 ( .A(matrixInput[54]), .B(n9707), .C(matrixInput[46]), .D(
        n9697), .Z(n10230) );
    VMW_AO22 U589 ( .A(matrixInput[352]), .B(n9707), .C(matrixInput[344]), .D(
        n9697), .Z(n9932) );
    VMW_AO22 U822 ( .A(matrixInput[142]), .B(n9707), .C(matrixInput[134]), .D(
        n9697), .Z(n10142) );
    VMW_FD \matrixInput_reg[363]  ( .D(n9913), .CP(Clk), .Q(matrixInput[363])
         );
    VMW_FD \matrixInput_reg[350]  ( .D(n9926), .CP(Clk), .Q(matrixInput[350])
         );
    VMW_FD \matrixInput_reg[349]  ( .D(n9927), .CP(Clk), .Q(matrixInput[349])
         );
    VMW_FD \matrixInput_reg[31]  ( .D(n10245), .CP(Clk), .Q(matrixInput[31])
         );
    VMW_FD \matrixInput_reg[28]  ( .D(n10248), .CP(Clk), .Q(matrixInput[28])
         );
    VMW_AO22 U747 ( .A(matrixInput[209]), .B(n9707), .C(matrixInput[201]), .D(
        n9697), .Z(n10075) );
    VMW_AO22 U760 ( .A(matrixInput[198]), .B(n9707), .C(matrixInput[190]), .D(
        n9697), .Z(n10086) );
    VMW_AO22 U805 ( .A(matrixInput[22]), .B(n9707), .C(matrixInput[14]), .D(
        n9697), .Z(n10262) );
    VMW_AO22 U298 ( .A(vectorInput[63]), .B(n9706), .C(vectorInput[55]), .D(
        n9696), .Z(n10285) );
    VMW_AO22 U308 ( .A(vectorInput[54]), .B(n9706), .C(vectorInput[46]), .D(
        n9696), .Z(n10294) );
    VMW_AO22 U341 ( .A(vectorInput[24]), .B(n9706), .C(vectorInput[16]), .D(
        n9696), .Z(n10324) );
    VMW_AO22 U366 ( .A(matrixInput[92]), .B(n9707), .C(matrixInput[84]), .D(
        n9697), .Z(n10192) );
    VMW_AO22 U477 ( .A(matrixInput[453]), .B(n9707), .C(matrixInput[445]), .D(
        n9697), .Z(n9831) );
    VMW_AO22 U577 ( .A(matrixInput[363]), .B(n9707), .C(matrixInput[355]), .D(
        n9697), .Z(n9921) );
    VMW_OAI21 U895 ( .A(n9708), .B(n9709), .C(n9703), .Z(n9695) );
    VMW_OAI21 U905 ( .A(n9728), .B(n9729), .C(n9703), .Z(n9680) );
    VMW_BUFIZ U939 ( .A(\holder[2] ), .E(RD), .Z(\DataOut[2]1 ) );
    VMW_FD \matrixInput_reg[238]  ( .D(n10038), .CP(Clk), .Q(matrixInput[238])
         );
    VMW_FD \matrixInput_reg[221]  ( .D(n10055), .CP(Clk), .Q(matrixInput[221])
         );
    VMW_FD \matrixInput_reg[122]  ( .D(n10154), .CP(Clk), .Q(matrixInput[122])
         );
    VMW_FD \matrixInput_reg[436]  ( .D(n9840), .CP(Clk), .Q(matrixInput[436])
         );
    VMW_FD \matrixInput_reg[212]  ( .D(n10064), .CP(Clk), .Q(matrixInput[212])
         );
    VMW_FD \matrixInput_reg[111]  ( .D(n10165), .CP(Clk), .Q(matrixInput[111])
         );
    VMW_FD \matrixInput_reg[108]  ( .D(n10168), .CP(Clk), .Q(matrixInput[108])
         );
    VMW_FD \matrixInput_reg[405]  ( .D(n9871), .CP(Clk), .Q(matrixInput[405])
         );
    VMW_FD \matrixInput_reg[382]  ( .D(n9894), .CP(Clk), .Q(matrixInput[382])
         );
    VMW_AO22 U647 ( .A(matrixInput[300]), .B(n9707), .C(matrixInput[292]), .D(
        n9697), .Z(n9984) );
    VMW_AO22 U660 ( .A(matrixInput[288]), .B(n9707), .C(matrixInput[280]), .D(
        n9697), .Z(n9996) );
    VMW_INV U922 ( .A(\holder[4] ), .Z(n9684) );
    VMW_FD \matrixInput_reg[12]  ( .D(n10264), .CP(Clk), .Q(matrixInput[12])
         );
    VMW_FD \matrixInput_reg[38]  ( .D(n10238), .CP(Clk), .Q(matrixInput[38])
         );
    VMW_FD \matrixInput_reg[21]  ( .D(n10255), .CP(Clk), .Q(matrixInput[21])
         );
    VMW_AO22 U383 ( .A(matrixInput[77]), .B(n9707), .C(matrixInput[69]), .D(
        n9697), .Z(n10207) );
    VMW_AO22 U425 ( .A(matrixInput[500]), .B(n9707), .C(matrixInput[492]), .D(
        n9697), .Z(n9784) );
    VMW_AO22 U550 ( .A(matrixInput[45]), .B(n9707), .C(matrixInput[37]), .D(
        n9697), .Z(n10239) );
    VMW_AO22 U685 ( .A(matrixInput[266]), .B(n9707), .C(matrixInput[258]), .D(
        n9697), .Z(n10018) );
    VMW_AO22 U839 ( .A(matrixInput[127]), .B(n9707), .C(matrixInput[119]), .D(
        n9697), .Z(n10157) );
    VMW_FD \matrixInput_reg[426]  ( .D(n9850), .CP(Clk), .Q(matrixInput[426])
         );
    VMW_FD \matrixInput_reg[415]  ( .D(n9861), .CP(Clk), .Q(matrixInput[415])
         );
    VMW_FD \matrixInput_reg[392]  ( .D(n9884), .CP(Clk), .Q(matrixInput[392])
         );
    VMW_FD \matrixInput_reg[231]  ( .D(n10045), .CP(Clk), .Q(matrixInput[231])
         );
    VMW_FD \matrixInput_reg[228]  ( .D(n10048), .CP(Clk), .Q(matrixInput[228])
         );
    VMW_FD \matrixInput_reg[202]  ( .D(n10074), .CP(Clk), .Q(matrixInput[202])
         );
    VMW_FD \vectorInput_reg[6]  ( .D(n10334), .CP(Clk), .Q(vectorInput[6]) );
    VMW_FD \matrixInput_reg[118]  ( .D(n10158), .CP(Clk), .Q(matrixInput[118])
         );
    VMW_FD \matrixInput_reg[101]  ( .D(n10175), .CP(Clk), .Q(matrixInput[101])
         );
    VMW_FD \matrixInput_reg[132]  ( .D(n10144), .CP(Clk), .Q(matrixInput[132])
         );
    VMW_FD \vectorInput_reg[43]  ( .D(n10297), .CP(Clk), .Q(vectorInput[43])
         );
    VMW_AO22 U715 ( .A(matrixInput[238]), .B(n9707), .C(matrixInput[230]), .D(
        n9697), .Z(n10046) );
    VMW_AO22 U857 ( .A(matrixInput[110]), .B(n9707), .C(matrixInput[102]), .D(
        n9697), .Z(n10174) );
    VMW_AO22 U870 ( .A(cOutput[53]), .B(n9702), .C(cOutput[21]), .D(n9701), 
        .Z(n9717) );
    VMW_FD \matrixInput_reg[0]  ( .D(n10276), .CP(Clk), .Q(matrixInput[0]) );
    VMW_AO22 U402 ( .A(matrixInput[59]), .B(n9707), .C(matrixInput[51]), .D(
        n9697), .Z(n10225) );
    VMW_AO22 U592 ( .A(matrixInput[349]), .B(n9707), .C(matrixInput[341]), .D(
        n9697), .Z(n9935) );
    VMW_AO22 U732 ( .A(matrixInput[223]), .B(n9707), .C(matrixInput[215]), .D(
        n9697), .Z(n10061) );
    VMW_FD \matrixInput_reg[373]  ( .D(n9903), .CP(Clk), .Q(matrixInput[373])
         );
    VMW_FD \matrixInput_reg[359]  ( .D(n9917), .CP(Clk), .Q(matrixInput[359])
         );
    VMW_FD \matrixInput_reg[340]  ( .D(n9936), .CP(Clk), .Q(matrixInput[340])
         );
    VMW_AO22 U489 ( .A(matrixInput[442]), .B(n9707), .C(matrixInput[434]), .D(
        n9697), .Z(n9842) );
    VMW_AO22 U391 ( .A(matrixInput[69]), .B(n9707), .C(matrixInput[61]), .D(
        n9697), .Z(n10215) );
    VMW_AO22 U437 ( .A(matrixInput[489]), .B(n9707), .C(matrixInput[481]), .D(
        n9697), .Z(n9795) );
    VMW_AO22 U519 ( .A(matrixInput[415]), .B(n9707), .C(matrixInput[407]), .D(
        n9697), .Z(n9869) );
    VMW_AO22 U629 ( .A(matrixInput[316]), .B(n9707), .C(matrixInput[308]), .D(
        n9697), .Z(n9968) );
    VMW_AO22 U697 ( .A(matrixInput[255]), .B(n9707), .C(matrixInput[247]), .D(
        n9697), .Z(n10029) );
    VMW_AO22 U707 ( .A(matrixInput[246]), .B(n9707), .C(matrixInput[238]), .D(
        n9697), .Z(n10038) );
    VMW_FD \matrixInput_reg[432]  ( .D(n9844), .CP(Clk), .Q(matrixInput[432])
         );
    VMW_FD \matrixInput_reg[418]  ( .D(n9858), .CP(Clk), .Q(matrixInput[418])
         );
    VMW_FD \matrixInput_reg[386]  ( .D(n9890), .CP(Clk), .Q(matrixInput[386])
         );
    VMW_FD \matrixInput_reg[401]  ( .D(n9875), .CP(Clk), .Q(matrixInput[401])
         );
    VMW_FD \matrixInput_reg[225]  ( .D(n10051), .CP(Clk), .Q(matrixInput[225])
         );
    VMW_FD \matrixInput_reg[126]  ( .D(n10150), .CP(Clk), .Q(matrixInput[126])
         );
    VMW_FD \matrixInput_reg[216]  ( .D(n10060), .CP(Clk), .Q(matrixInput[216])
         );
    VMW_FD \matrixInput_reg[115]  ( .D(n10161), .CP(Clk), .Q(matrixInput[115])
         );
    VMW_AO22 U580 ( .A(matrixInput[360]), .B(n9707), .C(matrixInput[352]), .D(
        n9697), .Z(n9924) );
    VMW_AO22 U845 ( .A(matrixInput[121]), .B(n9707), .C(matrixInput[113]), .D(
        n9697), .Z(n10163) );
    VMW_AO22 U410 ( .A(DataIn[1]), .B(n9707), .C(matrixInput[505]), .D(n9697), 
        .Z(n9771) );
    VMW_AO22 U720 ( .A(matrixInput[234]), .B(n9707), .C(matrixInput[226]), .D(
        n9697), .Z(n10050) );
    VMW_AO22 U862 ( .A(cOutput[55]), .B(n9702), .C(cOutput[23]), .D(n9701), 
        .Z(n9709) );
    VMW_FD \matrixInput_reg[35]  ( .D(n10241), .CP(Clk), .Q(matrixInput[35])
         );
    VMW_AO22 U769 ( .A(matrixInput[190]), .B(n9707), .C(matrixInput[182]), .D(
        n9697), .Z(n10094) );
    VMW_FD \matrixInput_reg[367]  ( .D(n9909), .CP(Clk), .Q(matrixInput[367])
         );
    VMW_FD \matrixInput_reg[354]  ( .D(n9922), .CP(Clk), .Q(matrixInput[354])
         );
    VMW_PULLDOWN U253 ( .Z(n9751) );
    VMW_AO22 U348 ( .A(vectorInput[8]), .B(n9706), .C(vectorInput[0]), .D(
        n9696), .Z(n10340) );
    VMW_AO22 U353 ( .A(matrixInput[104]), .B(n9707), .C(matrixInput[96]), .D(
        n9697), .Z(n10180) );
    VMW_AO22 U374 ( .A(matrixInput[85]), .B(n9707), .C(matrixInput[77]), .D(
        n9697), .Z(n10199) );
    VMW_AO22 U459 ( .A(matrixInput[469]), .B(n9707), .C(matrixInput[461]), .D(
        n9697), .Z(n9815) );
    VMW_AO22 U542 ( .A(matrixInput[395]), .B(n9707), .C(matrixInput[387]), .D(
        n9697), .Z(n9889) );
    VMW_AO22 U565 ( .A(matrixInput[374]), .B(n9707), .C(matrixInput[366]), .D(
        n9697), .Z(n9910) );
    VMW_AO22 U655 ( .A(matrixInput[293]), .B(n9707), .C(matrixInput[285]), .D(
        n9697), .Z(n9991) );
    VMW_AO22 U887 ( .A(cOutput[41]), .B(n9699), .C(cOutput[9]), .D(n9698), .Z(
        n9734) );
    VMW_INV U917 ( .A(\holder[5] ), .Z(n9687) );
    VMW_AO22 U672 ( .A(matrixInput[34]), .B(n9707), .C(matrixInput[26]), .D(
        n9697), .Z(n10250) );
    VMW_FD \vectorInput_reg[57]  ( .D(n10283), .CP(Clk), .Q(vectorInput[57])
         );
    VMW_AO22 U559 ( .A(matrixInput[379]), .B(n9707), .C(matrixInput[371]), .D(
        n9697), .Z(n9905) );
    VMW_BUFIZ U930 ( .A(n9746), .E(RD), .Z(\DataOut[9]1 ) );
    VMW_AO22 U669 ( .A(matrixInput[280]), .B(n9707), .C(matrixInput[272]), .D(
        n9697), .Z(n10004) );
    VMW_FD \matrixInput_reg[377]  ( .D(n9899), .CP(Clk), .Q(matrixInput[377])
         );
    VMW_FD \matrixInput_reg[344]  ( .D(n9932), .CP(Clk), .Q(matrixInput[344])
         );
    VMW_PULLDOWN U254 ( .Z(n9752) );
    VMW_OAI211 U273 ( .A(n9671), .B(n9681), .C(n9682), .D(n9683), .Z(n10345)
         );
    VMW_OAI211 U274 ( .A(n9671), .B(n9684), .C(n9685), .D(n9686), .Z(n10344)
         );
    VMW_AO22 U442 ( .A(matrixInput[485]), .B(n9707), .C(matrixInput[477]), .D(
        n9697), .Z(n9799) );
    VMW_AO22 U465 ( .A(matrixInput[464]), .B(n9707), .C(matrixInput[456]), .D(
        n9697), .Z(n9820) );
    VMW_AO22 U755 ( .A(matrixInput[203]), .B(n9707), .C(matrixInput[195]), .D(
        n9697), .Z(n10081) );
    VMW_AO22 U772 ( .A(matrixInput[25]), .B(n9707), .C(matrixInput[17]), .D(
        n9697), .Z(n10259) );
    VMW_AO22 U830 ( .A(matrixInput[135]), .B(n9707), .C(matrixInput[127]), .D(
        n9697), .Z(n10149) );
    VMW_FD \matrixInput_reg[4]  ( .D(n10272), .CP(Clk), .Q(matrixInput[4]) );
    VMW_FD \vectorInput_reg[47]  ( .D(n10293), .CP(Clk), .Q(vectorInput[47])
         );
    VMW_AO22 U291 ( .A(DataIn[5]), .B(n9706), .C(vectorInput[61]), .D(n9696), 
        .Z(n10279) );
    VMW_AO22 U620 ( .A(matrixInput[324]), .B(n9707), .C(matrixInput[316]), .D(
        n9697), .Z(n9960) );
    VMW_AO22 U817 ( .A(matrixInput[147]), .B(n9707), .C(matrixInput[139]), .D(
        n9697), .Z(n10137) );
    VMW_AO22 U879 ( .A(cOutput[43]), .B(n9699), .C(cOutput[11]), .D(n9698), 
        .Z(n9726) );
    VMW_FD \matrixInput_reg[206]  ( .D(n10070), .CP(Clk), .Q(matrixInput[206])
         );
    VMW_FD \matrixInput_reg[105]  ( .D(n10171), .CP(Clk), .Q(matrixInput[105])
         );
    VMW_FD \matrixInput_reg[422]  ( .D(n9854), .CP(Clk), .Q(matrixInput[422])
         );
    VMW_FD \matrixInput_reg[411]  ( .D(n9865), .CP(Clk), .Q(matrixInput[411])
         );
    VMW_FD \matrixInput_reg[396]  ( .D(n9880), .CP(Clk), .Q(matrixInput[396])
         );
    VMW_FD \matrixInput_reg[235]  ( .D(n10041), .CP(Clk), .Q(matrixInput[235])
         );
    VMW_FD \matrixInput_reg[136]  ( .D(n10140), .CP(Clk), .Q(matrixInput[136])
         );
    VMW_FD \matrixInput_reg[408]  ( .D(n9868), .CP(Clk), .Q(matrixInput[408])
         );
    VMW_FD \vectorInput_reg[2]  ( .D(n10338), .CP(Clk), .Q(vectorInput[2]) );
    VMW_FD \matrixInput_reg[16]  ( .D(n10260), .CP(Clk), .Q(matrixInput[16])
         );
    VMW_AO22 U296 ( .A(DataIn[1]), .B(n9706), .C(vectorInput[57]), .D(n9696), 
        .Z(n10283) );
    VMW_AO22 U301 ( .A(vectorInput[60]), .B(n9706), .C(vectorInput[52]), .D(
        n9696), .Z(n10288) );
    VMW_AO22 U510 ( .A(matrixInput[423]), .B(n9707), .C(matrixInput[415]), .D(
        n9697), .Z(n9861) );
    VMW_AO22 U306 ( .A(vectorInput[56]), .B(n9706), .C(vectorInput[48]), .D(
        n9696), .Z(n10292) );
    VMW_AO22 U321 ( .A(vectorInput[42]), .B(n9706), .C(vectorInput[34]), .D(
        n9696), .Z(n10306) );
    VMW_AO22 U326 ( .A(vectorInput[10]), .B(n9706), .C(vectorInput[2]), .D(
        n9696), .Z(n10338) );
    VMW_AO22 U480 ( .A(matrixInput[450]), .B(n9707), .C(matrixInput[442]), .D(
        n9697), .Z(n9834) );
    VMW_FD \matrixInput_reg[25]  ( .D(n10251), .CP(Clk), .Q(matrixInput[25])
         );
    VMW_AO22 U530 ( .A(matrixInput[406]), .B(n9707), .C(matrixInput[398]), .D(
        n9697), .Z(n9878) );
    VMW_AO22 U537 ( .A(matrixInput[399]), .B(n9707), .C(matrixInput[391]), .D(
        n9697), .Z(n9885) );
    VMW_AO22 U600 ( .A(matrixInput[342]), .B(n9707), .C(matrixInput[334]), .D(
        n9697), .Z(n9942) );
    VMW_AO22 U607 ( .A(matrixInput[336]), .B(n9707), .C(matrixInput[328]), .D(
        n9697), .Z(n9948) );
    VMW_AO22 U797 ( .A(matrixInput[165]), .B(n9707), .C(matrixInput[157]), .D(
        n9697), .Z(n10119) );
    VMW_BUFIZ U945 ( .A(n9758), .E(RD), .Z(\DataOut[24]1 ) );
    VMW_AO22 U859 ( .A(matrixInput[108]), .B(n9707), .C(matrixInput[100]), .D(
        n9697), .Z(n10176) );
    VMW_FD \matrixInput_reg[237]  ( .D(n10039), .CP(Clk), .Q(matrixInput[237])
         );
    VMW_FD \matrixInput_reg[204]  ( .D(n10072), .CP(Clk), .Q(matrixInput[204])
         );
    VMW_FD \matrixInput_reg[107]  ( .D(n10169), .CP(Clk), .Q(matrixInput[107])
         );
    VMW_FD \matrixInput_reg[134]  ( .D(n10142), .CP(Clk), .Q(matrixInput[134])
         );
    VMW_FD \matrixInput_reg[439]  ( .D(n9837), .CP(Clk), .Q(matrixInput[439])
         );
    VMW_FD \matrixInput_reg[420]  ( .D(n9856), .CP(Clk), .Q(matrixInput[420])
         );
    VMW_FD \matrixInput_reg[413]  ( .D(n9863), .CP(Clk), .Q(matrixInput[413])
         );
    VMW_FD \matrixInput_reg[394]  ( .D(n9882), .CP(Clk), .Q(matrixInput[394])
         );
    VMW_FD \vectorInput_reg[0]  ( .D(n10340), .CP(Clk), .Q(vectorInput[0]) );
    VMW_AO22 U790 ( .A(matrixInput[171]), .B(n9707), .C(matrixInput[163]), .D(
        n9697), .Z(n10113) );
    VMW_BUFIZ U942 ( .A(n9755), .E(RD), .Z(\DataOut[29]1 ) );
    VMW_FD \matrixInput_reg[14]  ( .D(n10262), .CP(Clk), .Q(matrixInput[14])
         );
    VMW_FD \matrixInput_reg[27]  ( .D(n10249), .CP(Clk), .Q(matrixInput[27])
         );
    VMW_AO22 U487 ( .A(matrixInput[444]), .B(n9707), .C(matrixInput[436]), .D(
        n9697), .Z(n9840) );
    VMW_AO22 U517 ( .A(matrixInput[417]), .B(n9707), .C(matrixInput[409]), .D(
        n9697), .Z(n9867) );
    VMW_AO22 U368 ( .A(matrixInput[90]), .B(n9707), .C(matrixInput[82]), .D(
        n9697), .Z(n10194) );
    VMW_AO22 U579 ( .A(matrixInput[361]), .B(n9707), .C(matrixInput[353]), .D(
        n9697), .Z(n9923) );
    VMW_AO22 U627 ( .A(matrixInput[38]), .B(n9707), .C(matrixInput[30]), .D(
        n9697), .Z(n10246) );
    VMW_AO22 U649 ( .A(matrixInput[298]), .B(n9707), .C(matrixInput[290]), .D(
        n9697), .Z(n9986) );
    VMW_AO22 U810 ( .A(matrixInput[153]), .B(n9707), .C(matrixInput[145]), .D(
        n9697), .Z(n10131) );
    VMW_FD \matrixInput_reg[375]  ( .D(n9901), .CP(Clk), .Q(matrixInput[375])
         );
    VMW_FD \matrixInput_reg[346]  ( .D(n9930), .CP(Clk), .Q(matrixInput[346])
         );
    VMW_FD \matrixInput_reg[6]  ( .D(n10270), .CP(Clk), .Q(matrixInput[6]) );
    VMW_AO22 U445 ( .A(matrixInput[482]), .B(n9707), .C(matrixInput[474]), .D(
        n9697), .Z(n9802) );
    VMW_AO22 U462 ( .A(matrixInput[467]), .B(n9707), .C(matrixInput[459]), .D(
        n9697), .Z(n9817) );
    VMW_AO22 U752 ( .A(matrixInput[206]), .B(n9707), .C(matrixInput[198]), .D(
        n9697), .Z(n10078) );
    VMW_AO22 U775 ( .A(matrixInput[185]), .B(n9707), .C(matrixInput[177]), .D(
        n9697), .Z(n10099) );
    VMW_FD \vectorInput_reg[45]  ( .D(n10295), .CP(Clk), .Q(vectorInput[45])
         );
    VMW_AO22 U837 ( .A(matrixInput[128]), .B(n9707), .C(matrixInput[120]), .D(
        n9697), .Z(n10156) );
    VMW_PULLDOWN U261 ( .Z(n9759) );
    VMW_PULLUP U268 ( .Z(Logic11) );
    VMW_AO22 U749 ( .A(matrixInput[9]), .B(n9707), .C(matrixInput[1]), .D(
        n9697), .Z(n10275) );
    VMW_FD \matrixInput_reg[365]  ( .D(n9911), .CP(Clk), .Q(matrixInput[365])
         );
    VMW_FD \matrixInput_reg[356]  ( .D(n9920), .CP(Clk), .Q(matrixInput[356])
         );
    VMW_AO22 U328 ( .A(vectorInput[36]), .B(n9706), .C(vectorInput[28]), .D(
        n9696), .Z(n10312) );
    VMW_AO22 U354 ( .A(matrixInput[103]), .B(n9707), .C(matrixInput[95]), .D(
        n9697), .Z(n10181) );
    VMW_AO22 U479 ( .A(matrixInput[451]), .B(n9707), .C(matrixInput[443]), .D(
        n9697), .Z(n9833) );
    VMW_BUFIZ U937 ( .A(\holder[6] ), .E(RD), .Z(\DataOut[6]1 ) );
    VMW_AO22 U373 ( .A(matrixInput[86]), .B(n9707), .C(matrixInput[78]), .D(
        n9697), .Z(n10198) );
    VMW_AO22 U545 ( .A(matrixInput[392]), .B(n9707), .C(matrixInput[384]), .D(
        n9697), .Z(n9892) );
    VMW_AO22 U562 ( .A(matrixInput[377]), .B(n9707), .C(matrixInput[369]), .D(
        n9697), .Z(n9907) );
    VMW_AO22 U652 ( .A(matrixInput[296]), .B(n9707), .C(matrixInput[288]), .D(
        n9697), .Z(n9988) );
    VMW_AO22 U675 ( .A(matrixInput[275]), .B(n9707), .C(matrixInput[267]), .D(
        n9697), .Z(n10009) );
    VMW_FD \vectorInput_reg[55]  ( .D(n10285), .CP(Clk), .Q(vectorInput[55])
         );
    VMW_AO22 U880 ( .A(cOutput[59]), .B(n9702), .C(cOutput[27]), .D(n9701), 
        .Z(n9727) );
    VMW_OAI21 U910 ( .A(n9738), .B(n9739), .C(n9705), .Z(n9673) );
    VMW_AO22 U384 ( .A(matrixInput[76]), .B(n9707), .C(matrixInput[68]), .D(
        n9697), .Z(n10208) );
    VMW_AO22 U396 ( .A(matrixInput[65]), .B(n9707), .C(matrixInput[57]), .D(
        n9697), .Z(n10219) );
    VMW_AO22 U417 ( .A(matrixInput[57]), .B(n9707), .C(matrixInput[49]), .D(
        n9697), .Z(n10227) );
    VMW_AO22 U727 ( .A(matrixInput[29]), .B(n9707), .C(matrixInput[21]), .D(
        n9697), .Z(n10255) );
    VMW_FD \matrixInput_reg[430]  ( .D(n9846), .CP(Clk), .Q(matrixInput[430])
         );
    VMW_FD \matrixInput_reg[429]  ( .D(n9847), .CP(Clk), .Q(matrixInput[429])
         );
    VMW_FD \matrixInput_reg[403]  ( .D(n9873), .CP(Clk), .Q(matrixInput[403])
         );
    VMW_FD \vectorInput_reg[9]  ( .D(n10331), .CP(Clk), .Q(vectorInput[9]) );
    VMW_FD \matrixInput_reg[384]  ( .D(n9892), .CP(Clk), .Q(matrixInput[384])
         );
    VMW_FD \matrixInput_reg[227]  ( .D(n10049), .CP(Clk), .Q(matrixInput[227])
         );
    VMW_FD \matrixInput_reg[214]  ( .D(n10062), .CP(Clk), .Q(matrixInput[214])
         );
    VMW_FD \matrixInput_reg[124]  ( .D(n10152), .CP(Clk), .Q(matrixInput[124])
         );
    VMW_FD \matrixInput_reg[117]  ( .D(n10159), .CP(Clk), .Q(matrixInput[117])
         );
    VMW_AO22 U865 ( .A(cOutput[38]), .B(n9699), .C(cOutput[6]), .D(n9698), .Z(
        n9712) );
    VMW_AO22 U405 ( .A(matrixInput[58]), .B(n9707), .C(matrixInput[50]), .D(
        n9697), .Z(n10226) );
    VMW_AO22 U430 ( .A(matrixInput[496]), .B(n9707), .C(matrixInput[488]), .D(
        n9697), .Z(n9788) );
    VMW_AO22 U587 ( .A(matrixInput[354]), .B(n9707), .C(matrixInput[346]), .D(
        n9697), .Z(n9930) );
    VMW_AO22 U842 ( .A(matrixInput[124]), .B(n9707), .C(matrixInput[116]), .D(
        n9697), .Z(n10160) );
    VMW_FD \matrixInput_reg[37]  ( .D(n10239), .CP(Clk), .Q(matrixInput[37])
         );
    VMW_AO22 U595 ( .A(matrixInput[347]), .B(n9707), .C(matrixInput[339]), .D(
        n9697), .Z(n9937) );
    VMW_AO22 U690 ( .A(matrixInput[261]), .B(n9707), .C(matrixInput[253]), .D(
        n9697), .Z(n10023) );
    VMW_AO22 U700 ( .A(matrixInput[252]), .B(n9707), .C(matrixInput[244]), .D(
        n9697), .Z(n10032) );
    VMW_AO22 U735 ( .A(matrixInput[220]), .B(n9707), .C(matrixInput[212]), .D(
        n9697), .Z(n10064) );
    VMW_FD \vectorInput_reg[58]  ( .D(n10282), .CP(Clk), .Q(vectorInput[58])
         );
    VMW_FD \vectorInput_reg[41]  ( .D(n10299), .CP(Clk), .Q(vectorInput[41])
         );
    VMW_AO22 U422 ( .A(matrixInput[503]), .B(n9707), .C(matrixInput[495]), .D(
        n9697), .Z(n9781) );
    VMW_AO22 U877 ( .A(cOutput[35]), .B(n9699), .C(cOutput[3]), .D(n9698), .Z(
        n9724) );
    VMW_AO22 U682 ( .A(matrixInput[268]), .B(n9707), .C(matrixInput[260]), .D(
        n9697), .Z(n10016) );
    VMW_AO22 U712 ( .A(matrixInput[241]), .B(n9707), .C(matrixInput[233]), .D(
        n9697), .Z(n10043) );
    VMW_AO22 U850 ( .A(matrixInput[117]), .B(n9707), .C(matrixInput[109]), .D(
        n9697), .Z(n10167) );
    VMW_FD \matrixInput_reg[2]  ( .D(n10274), .CP(Clk), .Q(matrixInput[2]) );
    VMW_FD \matrixInput_reg[371]  ( .D(n9905), .CP(Clk), .Q(matrixInput[371])
         );
    VMW_FD \matrixInput_reg[368]  ( .D(n9908), .CP(Clk), .Q(matrixInput[368])
         );
    VMW_FD \matrixInput_reg[342]  ( .D(n9934), .CP(Clk), .Q(matrixInput[342])
         );
    VMW_AO22 U346 ( .A(vectorInput[19]), .B(n9706), .C(vectorInput[11]), .D(
        n9696), .Z(n10329) );
    VMW_AO22 U539 ( .A(matrixInput[46]), .B(n9707), .C(matrixInput[38]), .D(
        n9697), .Z(n10238) );
    VMW_AO22 U557 ( .A(matrixInput[381]), .B(n9707), .C(matrixInput[373]), .D(
        n9697), .Z(n9903) );
    VMW_AO22 U609 ( .A(matrixInput[334]), .B(n9707), .C(matrixInput[326]), .D(
        n9697), .Z(n9950) );
    VMW_AO22 U799 ( .A(matrixInput[163]), .B(n9707), .C(matrixInput[155]), .D(
        n9697), .Z(n10121) );
    VMW_AO22 U361 ( .A(matrixInput[97]), .B(n9707), .C(matrixInput[89]), .D(
        n9697), .Z(n10187) );
    VMW_AO22 U640 ( .A(matrixInput[307]), .B(n9707), .C(matrixInput[299]), .D(
        n9697), .Z(n9977) );
    VMW_AO22 U667 ( .A(matrixInput[282]), .B(n9707), .C(matrixInput[274]), .D(
        n9697), .Z(n10002) );
    VMW_BUFIZ U925 ( .A(n9742), .E(RD), .Z(\DataOut[23]1 ) );
    VMW_FD \matrixInput_reg[10]  ( .D(n10266), .CP(Clk), .Q(matrixInput[10])
         );
    VMW_AO22 U470 ( .A(matrixInput[459]), .B(n9707), .C(matrixInput[451]), .D(
        n9697), .Z(n9825) );
    VMW_AO22 U570 ( .A(matrixInput[369]), .B(n9707), .C(matrixInput[361]), .D(
        n9697), .Z(n9915) );
    VMW_AO22 U819 ( .A(matrixInput[145]), .B(n9707), .C(matrixInput[137]), .D(
        n9697), .Z(n10139) );
    VMW_AO22 U892 ( .A(cOutput[56]), .B(n9702), .C(cOutput[24]), .D(n9701), 
        .Z(n9739) );
    VMW_FD \matrixInput_reg[23]  ( .D(n10253), .CP(Clk), .Q(matrixInput[23])
         );
    VMW_OAI21 U902 ( .A(n9722), .B(n9723), .C(n9705), .Z(n9685) );
    VMW_FD \matrixInput_reg[424]  ( .D(n9852), .CP(Clk), .Q(matrixInput[424])
         );
    VMW_FD \matrixInput_reg[417]  ( .D(n9859), .CP(Clk), .Q(matrixInput[417])
         );
    VMW_FD \matrixInput_reg[390]  ( .D(n9886), .CP(Clk), .Q(matrixInput[390])
         );
    VMW_FD \matrixInput_reg[389]  ( .D(n9887), .CP(Clk), .Q(matrixInput[389])
         );
    VMW_FD \vectorInput_reg[4]  ( .D(n10336), .CP(Clk), .Q(vectorInput[4]) );
    VMW_FD \matrixInput_reg[219]  ( .D(n10057), .CP(Clk), .Q(matrixInput[219])
         );
    VMW_FD \matrixInput_reg[103]  ( .D(n10173), .CP(Clk), .Q(matrixInput[103])
         );
    VMW_FD \matrixInput_reg[200]  ( .D(n10076), .CP(Clk), .Q(matrixInput[200])
         );
    VMW_FD \matrixInput_reg[233]  ( .D(n10043), .CP(Clk), .Q(matrixInput[233])
         );
    VMW_FD \matrixInput_reg[130]  ( .D(n10146), .CP(Clk), .Q(matrixInput[130])
         );
    VMW_FD \matrixInput_reg[129]  ( .D(n10147), .CP(Clk), .Q(matrixInput[129])
         );
    VMW_AO22 U740 ( .A(matrixInput[216]), .B(n9707), .C(matrixInput[208]), .D(
        n9697), .Z(n10068) );
    VMW_AO22 U802 ( .A(matrixInput[160]), .B(n9707), .C(matrixInput[152]), .D(
        n9697), .Z(n10124) );
    VMW_FD \matrixInput_reg[33]  ( .D(n10243), .CP(Clk), .Q(matrixInput[33])
         );
    VMW_FD \matrixInput_reg[19]  ( .D(n10257), .CP(Clk), .Q(matrixInput[19])
         );
    VMW_AO22 U767 ( .A(matrixInput[192]), .B(n9707), .C(matrixInput[184]), .D(
        n9697), .Z(n10092) );
    VMW_AND2 U284 ( .A(Addr[0]), .B(n9671), .Z(n9705) );
    VMW_AO22 U333 ( .A(vectorInput[31]), .B(n9706), .C(vectorInput[23]), .D(
        n9696), .Z(n10317) );
    VMW_AO22 U457 ( .A(matrixInput[471]), .B(n9707), .C(matrixInput[463]), .D(
        n9697), .Z(n9813) );
    VMW_AO22 U612 ( .A(matrixInput[331]), .B(n9707), .C(matrixInput[323]), .D(
        n9697), .Z(n9953) );
    VMW_AO22 U782 ( .A(matrixInput[178]), .B(n9707), .C(matrixInput[170]), .D(
        n9697), .Z(n10106) );
    VMW_AO22 U825 ( .A(matrixInput[139]), .B(n9707), .C(matrixInput[131]), .D(
        n9697), .Z(n10145) );
    VMW_AO22 U889 ( .A(cOutput[32]), .B(n9699), .C(cOutput[0]), .D(n9698), .Z(
        n9736) );
    VMW_INV U919 ( .A(\holder[3] ), .Z(n9681) );
    VMW_FD \matrixInput_reg[434]  ( .D(n9842), .CP(Clk), .Q(matrixInput[434])
         );
    VMW_FD \matrixInput_reg[223]  ( .D(n10053), .CP(Clk), .Q(matrixInput[223])
         );
    VMW_FD \matrixInput_reg[139]  ( .D(n10137), .CP(Clk), .Q(matrixInput[139])
         );
    VMW_FD \matrixInput_reg[120]  ( .D(n10156), .CP(Clk), .Q(matrixInput[120])
         );
    VMW_FD \matrixInput_reg[210]  ( .D(n10066), .CP(Clk), .Q(matrixInput[210])
         );
    VMW_FD \matrixInput_reg[113]  ( .D(n10163), .CP(Clk), .Q(matrixInput[113])
         );
    VMW_FD \matrixInput_reg[209]  ( .D(n10067), .CP(Clk), .Q(matrixInput[209])
         );
    VMW_FD \matrixInput_reg[407]  ( .D(n9869), .CP(Clk), .Q(matrixInput[407])
         );
    VMW_FD \matrixInput_reg[399]  ( .D(n9877), .CP(Clk), .Q(matrixInput[399])
         );
    VMW_FD \matrixInput_reg[380]  ( .D(n9896), .CP(Clk), .Q(matrixInput[380])
         );
    VMW_AO22 U505 ( .A(matrixInput[49]), .B(n9707), .C(matrixInput[41]), .D(
        n9697), .Z(n10235) );
    VMW_AO22 U522 ( .A(matrixInput[412]), .B(n9707), .C(matrixInput[404]), .D(
        n9697), .Z(n9872) );
    VMW_BUFIZ U950 ( .A(\holder[5] ), .E(RD), .Z(\DataOut[5]1 ) );
    VMW_AO22 U314 ( .A(vectorInput[48]), .B(n9706), .C(vectorInput[40]), .D(
        n9696), .Z(n10300) );
    VMW_AO22 U495 ( .A(matrixInput[437]), .B(n9707), .C(matrixInput[429]), .D(
        n9697), .Z(n9847) );
    VMW_AO22 U439 ( .A(matrixInput[55]), .B(n9707), .C(matrixInput[47]), .D(
        n9697), .Z(n10229) );
    VMW_AO22 U635 ( .A(matrixInput[310]), .B(n9707), .C(matrixInput[302]), .D(
        n9697), .Z(n9974) );
    VMW_FD \vectorInput_reg[62]  ( .D(n10278), .CP(Clk), .Q(vectorInput[62])
         );
    VMW_AO22 U699 ( .A(matrixInput[253]), .B(n9707), .C(matrixInput[245]), .D(
        n9697), .Z(n10031) );
    VMW_AO22 U709 ( .A(matrixInput[244]), .B(n9707), .C(matrixInput[236]), .D(
        n9697), .Z(n10040) );
    VMW_FD \vectorInput_reg[51]  ( .D(n10289), .CP(Clk), .Q(vectorInput[51])
         );
    VMW_FD \vectorInput_reg[48]  ( .D(n10292), .CP(Clk), .Q(vectorInput[48])
         );
    VMW_FD \matrixInput_reg[378]  ( .D(n9898), .CP(Clk), .Q(matrixInput[378])
         );
    VMW_FD \matrixInput_reg[352]  ( .D(n9924), .CP(Clk), .Q(matrixInput[352])
         );
    VMW_FD \matrixInput_reg[361]  ( .D(n9915), .CP(Clk), .Q(matrixInput[361])
         );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_6 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n1, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_5 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n2, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n2) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n2), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_4 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n3, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n3) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n3), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_7 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_7 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n31, n32, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , \CARRYB[2][1] , 
        \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , \ab[3][3] , 
        \A1[2] , n33, n34, n35, \A2[3] , \ab[2][0] , \ab[6][0] , \ab[2][2] , 
        \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , 
        \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[5][1] , 
        \SUMB[3][4] , lsb_0, \ab[4][2] , \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , \ab[4][0] , 
        \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , \ab[1][1] , \ab[0][7] , 
        \CARRYB[1][5] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , n36, \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , \SUMB[3][3] , 
        \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , \A2[4] , 
        \A2[2] , \A2[6] , \SUMB[1][3] , \CARRYB[1][3] , \CARRYB[5][1] , 
        \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , \A1[1] , 
        \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , \ab[3][2] , 
        \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n31) );
    VMW_PULLDOWN U5 ( .Z(n33) );
    VMW_PULLDOWN U6 ( .Z(n34) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n32), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n35) );
    VMW_PULLDOWN U8 ( .Z(n36) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n33), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n34), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n31), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_7 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n36), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n32) );
    VMW_FADD S0_1 ( .CI(n35), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_6 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_6 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n37, n38, n40, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , n41, \A2[3] , \ab[6][0] , \ab[2][2] , 
        \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , 
        \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[4][2] , 
        \ab[5][1] , \SUMB[3][4] , lsb_0, \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[0][7] , 
        \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , \ab[0][1] , 
        \ab[4][3] , \ab[5][0] , \SUMB[4][2] , \CARRYB[3][1] , n39, n42, 
        \SUMB[1][3] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , \CARRYB[2][2] , 
        \A2[2] , \A2[6] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , 
        \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , 
        \ab[3][2] , \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , 
        \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n37) );
    VMW_PULLDOWN U5 ( .Z(n39) );
    VMW_PULLDOWN U6 ( .Z(n40) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n38), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n41) );
    VMW_PULLDOWN U8 ( .Z(n42) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n39), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n40), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n37), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_6 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n42), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n38) );
    VMW_FADD S0_1 ( .CI(n41), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_5 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_5 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n43, n44, n46, n47, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , n48, lsb_0, \A2[3] , \ab[6][0] , 
        \ab[2][2] , \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , 
        \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , 
        \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[0][6] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , \ab[4][0] , 
        \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , \ab[0][7] , \CARRYB[1][5] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \CARRYB[1][1] , \SUMB[3][3] , \ab[1][4] , \CARRYB[4][0] , 
        n45, \A2[2] , \A2[6] , \ab[1][6] , \SUMB[3][1] , \ab[0][5] , 
        \CARRYB[4][2] , \SUMB[1][3] , \CARRYB[1][3] , \CARRYB[5][1] , 
        \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , \A1[1] , 
        \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , \ab[3][2] , 
        \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , 
        \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n43) );
    VMW_PULLDOWN U5 ( .Z(n45) );
    VMW_PULLDOWN U6 ( .Z(n46) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n44), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n47) );
    VMW_PULLDOWN U8 ( .Z(n48) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n45), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n46), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n43), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_5 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n48), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n44) );
    VMW_FADD S0_1 ( .CI(n47), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_3 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n4, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n4) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n4), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_4 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_4 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n49, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , n50, n51, n52, 
        \SUMB[1][2] , \CARRYB[2][3] , n53, \ab[1][3] , \A1[4] , \ab[4][2] , 
        \ab[5][1] , \SUMB[3][4] , n54, lsb_0, \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , 
        \CARRYB[1][0] , \SUMB[2][1] , \ab[0][7] , \ab[1][5] , \SUMB[3][2] , 
        \CARRYB[1][5] , \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , 
        \SUMB[2][5] , \ab[0][2] , \ab[1][1] , \ab[4][1] , \ab[0][3] , 
        \SUMB[2][4] , \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , 
        \CARRYB[1][1] , \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , 
        \CARRYB[4][2] , \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , 
        \SUMB[2][2] , \ab[4][3] , \ab[5][0] , \A2[6] , \SUMB[1][3] , 
        \ab[0][1] , \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , 
        \CARRYB[6][0] , \CARRYB[2][2] , \A1[5] , \A2[4] , \A2[2] , \ab[6][1] , 
        \ab[2][3] , \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , 
        \ab[7][0] , \ab[2][1] , \ab[3][2] , \A1[3] , \SUMB[1][1] , 
        \CARRYB[2][0] , \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n49) );
    VMW_PULLDOWN U5 ( .Z(n51) );
    VMW_PULLDOWN U6 ( .Z(n52) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n50), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n53) );
    VMW_PULLDOWN U8 ( .Z(n54) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n51), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n52), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n49), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_4 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n54), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n50) );
    VMW_FADD S0_1 ( .CI(n53), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_3 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_3 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n55, n56, n60, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , lsb_0, \A2[3] , \ab[6][0] , 
        \ab[2][2] , \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , 
        \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , 
        \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , n57, n58, \ab[0][7] , 
        \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \SUMB[2][2] , n59, \ab[1][2] , 
        \ab[0][1] , \ab[4][3] , \ab[5][0] , \SUMB[4][2] , \CARRYB[3][1] , 
        \A2[2] , \A2[6] , \SUMB[1][3] , \ab[3][4] , \SUMB[5][1] , 
        \CARRYB[6][0] , \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n55) );
    VMW_PULLDOWN U5 ( .Z(n57) );
    VMW_PULLDOWN U6 ( .Z(n58) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n56), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n59) );
    VMW_PULLDOWN U8 ( .Z(n60) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n57), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n58), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n55), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_3 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n60), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n56) );
    VMW_FADD S0_1 ( .CI(n59), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_2 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_2 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n61, n66, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , \CARRYB[3][0] , 
        \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[4][2] , \ab[5][1] , 
        \SUMB[3][4] , lsb_0, \ab[0][6] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , \CARRYB[1][0] , 
        \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , 
        \SUMB[2][5] , \ab[0][2] , n62, n63, \ab[0][7] , \CARRYB[1][5] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \CARRYB[1][1] , n64, \ab[1][4] , \SUMB[3][3] , 
        \SUMB[3][1] , \CARRYB[4][0] , n65, \ab[1][6] , \ab[0][5] , 
        \CARRYB[4][2] , \SUMB[1][3] , \CARRYB[1][3] , \CARRYB[5][1] , 
        \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A2[2] , \A2[6] , \A1[5] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n61) );
    VMW_PULLDOWN U5 ( .Z(n63) );
    VMW_PULLDOWN U6 ( .Z(n64) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n62), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n65) );
    VMW_PULLDOWN U8 ( .Z(n66) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n63), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n64), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n61), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_2 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n66), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n62) );
    VMW_FADD S0_1 ( .CI(n65), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_2 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n5, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n5) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n5), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_1 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_1 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n67, n69, n72, \A1[13] , \A2[5] , \CARRYB[2][1] , \SUMB[5][2] , 
        \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , \A2[1] , \SUMB[1][4] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , n68, lsb_0, \A2[3] , \ab[6][0] , 
        \ab[2][2] , \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , 
        \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , 
        \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , n70, n71, \ab[0][6] , 
        \ab[1][5] , \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \SUMB[2][4] , \A2[2] , \A2[6] , \ab[0][7] , 
        \ab[0][3] , \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , 
        \CARRYB[1][1] , \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , 
        \CARRYB[4][2] , \SUMB[1][3] , \CARRYB[1][3] , \CARRYB[5][1] , 
        \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , \A1[1] , 
        \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , \ab[3][2] , 
        \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , 
        \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n67) );
    VMW_PULLDOWN U5 ( .Z(n69) );
    VMW_PULLDOWN U6 ( .Z(n70) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n68), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n71) );
    VMW_PULLDOWN U8 ( .Z(n72) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n69), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n70), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n67), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_1 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n72), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n68) );
    VMW_FADD S0_1 ( .CI(n71), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_1 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n6, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n6) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n6), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_0 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_0 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n73, n74, n75, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \SUMB[1][2] , \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , 
        \CARRYB[2][3] , \ab[1][3] , \A1[4] , \ab[4][2] , \ab[5][1] , 
        \SUMB[3][4] , lsb_0, \ab[0][6] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \CARRYB[1][0] , 
        \SUMB[2][1] , n76, n78, \ab[1][5] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \ab[0][7] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , \ab[0][1] , 
        \ab[4][3] , \ab[5][0] , n77, \A2[6] , \SUMB[1][3] , \SUMB[4][2] , 
        \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \A2[4] , \A2[2] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n73) );
    VMW_PULLDOWN U5 ( .Z(n75) );
    VMW_PULLDOWN U6 ( .Z(n76) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n74), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n77) );
    VMW_PULLDOWN U8 ( .Z(n78) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n75), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n76), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n73), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_14_0 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n78), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n74) );
    VMW_FADD S0_1 ( .CI(n77), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_0 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n7, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n7) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n7), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize8_pWordSize8 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, vectorAInput, vectorBInput, cOutput );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [63:0] vectorAInput;
output [7:0] cOutput;
input  [63:0] vectorBInput;
input  Clk, Reset, RD, WR;
    wire n832, n834, n826, \result60[1] , \n642[8] , \n730[7] , \result463[5] , 
        \result552[2] , \n553[7] , \n464[7] , \n642[1] , \result60[5] , 
        \result285[2] , \result463[1] , \n730[3] , n829, n828, n833, \n642[5] , 
        \result285[6] , \result552[6] , \result552[4] , \n553[3] , \n464[3] , 
        \n642[7] , \n553[1] , \n464[1] , \result60[7] , \result285[4] , 
        \n730[8] , n821, \n642[3] , \n730[1] , \result463[3] , \n553[8] , 
        \n464[8] , \result285[0] , \result552[0] , \n464[5] , \n553[5] , 
        \result463[7] , \result60[3] , \result641[1] , \n730[5] , \n286[2] , 
        \n197[4] , \result196[1] , \n106[3] , \result374[5] , n823, n825, n820, 
        \result641[5] , \result196[5] , \n106[7] , \n375[4] , \result374[1] , 
        \n286[6] , n827, \result641[7] , \n286[4] , \result641[3] , 
        \result196[7] , \result196[3] , \n106[5] , \result374[3] , \n375[6] , 
        \n197[2] , \n106[8] , \n375[2] , \n197[6] , \n106[1] , \result374[7] , 
        \n286[8] , n822, n830, \result641[6] , \result641[2] , \result196[2] , 
        \n375[3] , \n197[7] , \result374[6] , \n286[1] , \result641[4] , 
        \result196[6] , \n286[5] , \result196[4] , \n106[4] , \result374[2] , 
        \n375[7] , \n197[3] , \n106[6] , \result374[0] , \n375[5] , \n197[1] , 
        \n286[7] , \result641[0] , \n197[8] , \result196[0] , \n286[3] , 
        \n375[1] , \n197[5] , \n106[2] , \result374[4] , n831, \n642[2] , 
        \n375[8] , \result285[1] , \result552[1] , \n553[4] , \n464[4] , 
        \result60[2] , \result463[6] , \result552[5] , \n730[4] , \n642[6] , 
        \result285[5] , n824, \result60[6] , \result60[4] , \result463[2] , 
        \result463[0] , \n642[4] , \n730[2] , \result285[7] , \result60[0] , 
        \result552[7] , \n553[2] , \n464[2] , \result552[3] , \n730[6] , 
        \n464[6] , \result463[4] , \n553[6] , \result285[3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 , UNCONNECTED_23 , UNCONNECTED_24 , 
	UNCONNECTED_25 , UNCONNECTED_26 , UNCONNECTED_27 , UNCONNECTED_28 , 
	UNCONNECTED_29 , UNCONNECTED_30 , UNCONNECTED_31 , UNCONNECTED_32 , 
	UNCONNECTED_33 , UNCONNECTED_34 , UNCONNECTED_35 , UNCONNECTED_36 , 
	UNCONNECTED_37 , UNCONNECTED_38 , UNCONNECTED_39 , UNCONNECTED_40 , 
	UNCONNECTED_41 , UNCONNECTED_42 , UNCONNECTED_43 , UNCONNECTED_44 , 
	UNCONNECTED_45 , UNCONNECTED_46 , UNCONNECTED_47 , UNCONNECTED_48 , 
	UNCONNECTED_49 , UNCONNECTED_50 , UNCONNECTED_51 , UNCONNECTED_52 , 
	UNCONNECTED_53 , UNCONNECTED_54 , UNCONNECTED_55 , UNCONNECTED_56 , 
	UNCONNECTED_57 , UNCONNECTED_58 , UNCONNECTED_59 , UNCONNECTED_60 , 
	UNCONNECTED_61 , UNCONNECTED_62 , UNCONNECTED_63 , UNCONNECTED_64 ;
    VMW_PULLDOWN U20 ( .Z(n832) );
    VMW_PULLDOWN U21 ( .Z(n823) );
    VMW_FD \cOutput_reg[2]  ( .D(\result60[2] ), .CP(Clk), .Q(cOutput[2]) );
    VMW_PULLDOWN U26 ( .Z(n820) );
    VMW_PULLDOWN U28 ( .Z(n828) );
    VMW_PULLDOWN U33 ( .Z(n827) );
    VMW_FD \cOutput_reg[6]  ( .D(\result60[6] ), .CP(Clk), .Q(cOutput[6]) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_2 mul_48_6 ( .A(
        vectorAInput[55:48]), .B(vectorBInput[55:48]), .TC(n825), .PRODUCT({
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, UNCONNECTED_8, \n642[1] , 
        \n642[2] , \n642[3] , \n642[4] , \n642[5] , \n642[6] , \n642[7] , 
        \n642[8] }) );
    VMW_PULLDOWN U34 ( .Z(n831) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_6 add_48_6 ( .A({
        \result552[7] , \result552[6] , \result552[5] , \result552[4] , 
        \result552[3] , \result552[2] , \result552[1] , \result552[0] }), .B({
        \n642[1] , \n642[2] , \n642[3] , \n642[4] , \n642[5] , \n642[6] , 
        \n642[7] , \n642[8] }), .CI(n834), .SUM({\result641[7] , 
        \result641[6] , \result641[5] , \result641[4] , \result641[3] , 
        \result641[2] , \result641[1] , \result641[0] }) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_2 add_48_1 ( .A({
        \n106[1] , \n106[2] , \n106[3] , \n106[4] , \n106[5] , \n106[6] , 
        \n106[7] , \n106[8] }), .B({\n197[1] , \n197[2] , \n197[3] , \n197[4] , 
        \n197[5] , \n197[6] , \n197[7] , \n197[8] }), .CI(n824), .SUM({
        \result196[7] , \result196[6] , \result196[5] , \result196[4] , 
        \result196[3] , \result196[2] , \result196[1] , \result196[0] }) );
    VMW_FD \cOutput_reg[4]  ( .D(\result60[4] ), .CP(Clk), .Q(cOutput[4]) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_4 mul_48_1 ( .A(
        vectorAInput[15:8]), .B(vectorBInput[15:8]), .TC(n827), .PRODUCT({
        UNCONNECTED_9, UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, 
        UNCONNECTED_13, UNCONNECTED_14, UNCONNECTED_15, UNCONNECTED_16, 
        \n197[1] , \n197[2] , \n197[3] , \n197[4] , \n197[5] , \n197[6] , 
        \n197[7] , \n197[8] }) );
    VMW_PULLDOWN U27 ( .Z(n829) );
    VMW_FD \cOutput_reg[0]  ( .D(\result60[0] ), .CP(Clk), .Q(cOutput[0]) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_4 add_48_7 ( .A({
        \result641[7] , \result641[6] , \result641[5] , \result641[4] , 
        \result641[3] , \result641[2] , \result641[1] , \result641[0] }), .B({
        \n730[1] , \n730[2] , \n730[3] , \n730[4] , \n730[5] , \n730[6] , 
        \n730[7] , \n730[8] }), .CI(n832), .SUM({\result60[7] , \result60[6] , 
        \result60[5] , \result60[4] , \result60[3] , \result60[2] , 
        \result60[1] , \result60[0] }) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_7 mul_48 ( .A(
        vectorAInput[7:0]), .B(vectorBInput[7:0]), .TC(n831), .PRODUCT({
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, UNCONNECTED_23, UNCONNECTED_24, 
        \n106[1] , \n106[2] , \n106[3] , \n106[4] , \n106[5] , \n106[6] , 
        \n106[7] , \n106[8] }) );
    VMW_PULLDOWN U22 ( .Z(n834) );
    VMW_PULLDOWN U29 ( .Z(n826) );
    VMW_PULLDOWN U32 ( .Z(n824) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_1 mul_48_7 ( .A(
        vectorAInput[63:56]), .B(vectorBInput[63:56]), .TC(n823), .PRODUCT({
        UNCONNECTED_25, UNCONNECTED_26, UNCONNECTED_27, UNCONNECTED_28, 
        UNCONNECTED_29, UNCONNECTED_30, UNCONNECTED_31, UNCONNECTED_32, 
        \n730[1] , \n730[2] , \n730[3] , \n730[4] , \n730[5] , \n730[6] , 
        \n730[7] , \n730[8] }) );
    VMW_PULLDOWN U23 ( .Z(n825) );
    VMW_PULLDOWN U24 ( .Z(n822) );
    VMW_PULLDOWN U25 ( .Z(n830) );
    VMW_PULLDOWN U30 ( .Z(n833) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_6 mul_48_5 ( .A(
        vectorAInput[47:40]), .B(vectorBInput[47:40]), .TC(n830), .PRODUCT({
        UNCONNECTED_33, UNCONNECTED_34, UNCONNECTED_35, UNCONNECTED_36, 
        UNCONNECTED_37, UNCONNECTED_38, UNCONNECTED_39, UNCONNECTED_40, 
        \n553[1] , \n553[2] , \n553[3] , \n553[4] , \n553[5] , \n553[6] , 
        \n553[7] , \n553[8] }) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_5 add_48_2 ( .A({
        \result196[7] , \result196[6] , \result196[5] , \result196[4] , 
        \result196[3] , \result196[2] , \result196[1] , \result196[0] }), .B({
        \n286[1] , \n286[2] , \n286[3] , \n286[4] , \n286[5] , \n286[6] , 
        \n286[7] , \n286[8] }), .CI(n833), .SUM({\result285[7] , 
        \result285[6] , \result285[5] , \result285[4] , \result285[3] , 
        \result285[2] , \result285[1] , \result285[0] }) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_1 add_48_5 ( .A({
        \result463[7] , \result463[6] , \result463[5] , \result463[4] , 
        \result463[3] , \result463[2] , \result463[1] , \result463[0] }), .B({
        \n553[1] , \n553[2] , \n553[3] , \n553[4] , \n553[5] , \n553[6] , 
        \n553[7] , \n553[8] }), .CI(n822), .SUM({\result552[7] , 
        \result552[6] , \result552[5] , \result552[4] , \result552[3] , 
        \result552[2] , \result552[1] , \result552[0] }) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_0 mul_48_2 ( .A(
        vectorAInput[23:16]), .B(vectorBInput[23:16]), .TC(n821), .PRODUCT({
        UNCONNECTED_41, UNCONNECTED_42, UNCONNECTED_43, UNCONNECTED_44, 
        UNCONNECTED_45, UNCONNECTED_46, UNCONNECTED_47, UNCONNECTED_48, 
        \n286[1] , \n286[2] , \n286[3] , \n286[4] , \n286[5] , \n286[6] , 
        \n286[7] , \n286[8] }) );
    VMW_FD \cOutput_reg[1]  ( .D(\result60[1] ), .CP(Clk), .Q(cOutput[1]) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_3 mul_48_3 ( .A(
        vectorAInput[31:24]), .B(vectorBInput[31:24]), .TC(n826), .PRODUCT({
        UNCONNECTED_49, UNCONNECTED_50, UNCONNECTED_51, UNCONNECTED_52, 
        UNCONNECTED_53, UNCONNECTED_54, UNCONNECTED_55, UNCONNECTED_56, 
        \n375[1] , \n375[2] , \n375[3] , \n375[4] , \n375[5] , \n375[6] , 
        \n375[7] , \n375[8] }) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_0 add_48_4 ( .A({
        \result374[7] , \result374[6] , \result374[5] , \result374[4] , 
        \result374[3] , \result374[2] , \result374[1] , \result374[0] }), .B({
        \n464[1] , \n464[2] , \n464[3] , \n464[4] , \n464[5] , \n464[6] , 
        \n464[7] , \n464[8] }), .CI(n820), .SUM({\result463[7] , 
        \result463[6] , \result463[5] , \result463[4] , \result463[3] , 
        \result463[2] , \result463[1] , \result463[0] }) );
    VMW_FD \cOutput_reg[7]  ( .D(\result60[7] ), .CP(Clk), .Q(cOutput[7]) );
    VMW_FD \cOutput_reg[5]  ( .D(\result60[5] ), .CP(Clk), .Q(cOutput[5]) );
    VMW_PULLDOWN U31 ( .Z(n821) );
    VMW_FD \cOutput_reg[3]  ( .D(\result60[3] ), .CP(Clk), .Q(cOutput[3]) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW01_add_8_3 add_48_3 ( .A({
        \result285[7] , \result285[6] , \result285[5] , \result285[4] , 
        \result285[3] , \result285[2] , \result285[1] , \result285[0] }), .B({
        \n375[1] , \n375[2] , \n375[3] , \n375[4] , \n375[5] , \n375[6] , 
        \n375[7] , \n375[8] }), .CI(n828), .SUM({\result374[7] , 
        \result374[6] , \result374[5] , \result374[4] , \result374[3] , 
        \result374[2] , \result374[1] , \result374[0] }) );
    VectorDotProduct_pVectorSize8_pWordSize8_DW02_mult_8_8_5 mul_48_4 ( .A(
        vectorAInput[39:32]), .B(vectorBInput[39:32]), .TC(n829), .PRODUCT({
        UNCONNECTED_57, UNCONNECTED_58, UNCONNECTED_59, UNCONNECTED_60, 
        UNCONNECTED_61, UNCONNECTED_62, UNCONNECTED_63, UNCONNECTED_64, 
        \n464[1] , \n464[2] , \n464[3] , \n464[4] , \n464[5] , \n464[6] , 
        \n464[7] , \n464[8] }) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \matrixInput[53] , \vectorInput[51] , \matrixInput[483] , 
        \matrixInput[79] , \matrixInput[60] , \cOutput[54] , 
        \matrixInput[462] , \matrixInput[337] , \matrixInput[304] , 
        \matrixInput[294] , \matrixInput[197] , \matrixInput[98] , 
        \matrixInput[81] , \matrixInput[451] , \matrixInput[448] , 
        \matrixInput[176] , \vectorInput[48] , \matrixInput[275] , 
        \matrixInput[145] , \vectorInput[62] , \matrixInput[246] , 
        \vectorInput[58] , \matrixInput[256] , \matrixInput[155] , 
        \matrixInput[91] , \matrixInput[88] , \matrixInput[166] , 
        \vectorInput[41] , \matrixInput[472] , \matrixInput[458] , 
        \matrixInput[441] , \matrixInput[265] , \matrixInput[70] , 
        \matrixInput[69] , \cOutput[44] , \matrixInput[43] , \cOutput[6] , 
        \vectorInput[55] , \matrixInput[503] , \matrixInput[284] , 
        \matrixInput[187] , \matrixInput[493] , \matrixInput[327] , 
        \matrixInput[314] , \matrixInput[271] , \matrixInput[268] , 
        \matrixInput[242] , \matrixInput[172] , \matrixInput[487] , 
        \matrixInput[466] , \matrixInput[158] , \matrixInput[141] , 
        \matrixInput[455] , \matrixInput[319] , \matrixInput[290] , 
        \matrixInput[289] , \matrixInput[193] , \matrixInput[85] , 
        \matrixInput[300] , \matrixInput[333] , \matrixInput[57] , 
        \cOutput[63] , \cOutput[50] , \cOutput[49] , \matrixInput[64] , 
        \matrixInput[507] , \matrixInput[497] , \matrixInput[323] , 
        \matrixInput[310] , \matrixInput[309] , \matrixInput[299] , 
        \matrixInput[280] , \matrixInput[183] , \matrixInput[74] , 
        \cOutput[2] , \matrixInput[476] , \matrixInput[445] , 
        \matrixInput[47] , \cOutput[59] , \cOutput[40] , \matrixInput[252] , 
        \vectorInput[47] , \vectorInput[45] , \matrixInput[278] , 
        \matrixInput[151] , \matrixInput[148] , \matrixInput[261] , 
        \matrixInput[474] , \matrixInput[447] , \matrixInput[162] , 
        \matrixInput[95] , \matrixInput[250] , \matrixInput[249] , 
        \matrixInput[153] , \matrixInput[179] , \matrixInput[160] , 
        \matrixInput[505] , \matrixInput[495] , \matrixInput[338] , 
        \matrixInput[321] , \matrixInput[263] , \matrixInput[97] , 
        \matrixInput[312] , \matrixInput[282] , \cOutput[0] , 
        \matrixInput[198] , \matrixInput[181] , \matrixInput[76] , 
        \matrixInput[485] , \matrixInput[292] , \matrixInput[45] , 
        \cOutput[42] , \cOutput[9] , \matrixInput[191] , \matrixInput[188] , 
        \matrixInput[331] , \matrixInput[328] , \matrixInput[302] , 
        \cOutput[61] , \cOutput[52] , \matrixInput[55] , \vectorInput[57] , 
        \matrixInput[170] , \matrixInput[169] , \matrixInput[66] , 
        \matrixInput[273] , \matrixInput[501] , \matrixInput[464] , 
        \matrixInput[259] , \matrixInput[240] , \matrixInput[143] , 
        \matrixInput[457] , \matrixInput[87] , \matrixInput[72] , 
        \cOutput[46] , \matrixInput[58] , \matrixInput[41] , 
        \matrixInput[185] , \vectorInput[60] , \vectorInput[53] , 
        \vectorInput[43] , \matrixInput[491] , \matrixInput[488] , 
        \matrixInput[325] , \matrixInput[286] , \cOutput[4] , 
        \matrixInput[316] , \matrixInput[267] , \matrixInput[254] , 
        \matrixInput[93] , \matrixInput[157] , \matrixInput[479] , 
        \matrixInput[470] , \matrixInput[443] , \matrixInput[164] , 
        \matrixInput[469] , \matrixInput[83] , \matrixInput[460] , 
        \matrixInput[453] , \matrixInput[277] , \matrixInput[174] , 
        \matrixInput[244] , \matrixInput[147] , \matrixInput[51] , 
        \matrixInput[48] , \matrixInput[62] , \vectorInput[36] , 
        \matrixInput[511] , \matrixInput[498] , \matrixInput[481] , 
        \matrixInput[306] , \cOutput[56] , \matrixInput[335] , 
        \matrixInput[508] , \matrixInput[296] , \matrixInput[195] , 
        \matrixInput[436] , \matrixInput[405] , \matrixInput[238] , 
        \matrixInput[221] , \matrixInput[212] , \matrixInput[111] , 
        \matrixInput[108] , \matrixInput[122] , \matrixInput[382] , 
        \matrixInput[363] , \matrixInput[350] , \matrixInput[349] , 
        \cOutput[19] , \vectorInput[3] , \matrixInput[373] , 
        \matrixInput[359] , \matrixInput[340] , \matrixInput[34] , 
        \matrixInput[7] , \cOutput[33] , \matrixInput[24] , \matrixInput[17] , 
        \cOutput[23] , \cOutput[10] , \vectorInput[26] , \vectorInput[15] , 
        \matrixInput[426] , \matrixInput[415] , \matrixInput[392] , 
        \matrixInput[231] , \matrixInput[228] , \matrixInput[132] , 
        \matrixInput[202] , \matrixInput[118] , \matrixInput[101] , 
        \matrixInput[30] , \matrixInput[29] , \matrixInput[3] , \cOutput[37] , 
        \matrixInput[367] , \matrixInput[354] , \vectorInput[32] , 
        \matrixInput[432] , \matrixInput[418] , \matrixInput[386] , 
        \matrixInput[401] , \matrixInput[216] , \matrixInput[115] , 
        \vectorInput[22] , \vectorInput[18] , \matrixInput[126] , 
        \vectorInput[11] , \matrixInput[225] , \matrixInput[136] , 
        \matrixInput[235] , \matrixInput[206] , \matrixInput[105] , 
        \matrixInput[422] , \matrixInput[411] , \matrixInput[396] , 
        \matrixInput[408] , \cOutput[27] , \vectorInput[7] , \matrixInput[13] , 
        \cOutput[14] , \matrixInput[39] , \matrixInput[20] , 
        \matrixInput[377] , \matrixInput[344] , \cOutput[25] , 
        \vectorInput[5] , \matrixInput[22] , \matrixInput[11] , \cOutput[16] , 
        \matrixInput[8] , \matrixInput[375] , \matrixInput[346] , 
        \vectorInput[39] , \vectorInput[13] , \matrixInput[237] , 
        \matrixInput[134] , \vectorInput[20] , \matrixInput[439] , 
        \matrixInput[420] , \matrixInput[204] , \matrixInput[107] , 
        \matrixInput[413] , \matrixInput[394] , \vectorInput[30] , 
        \matrixInput[430] , \matrixInput[429] , \matrixInput[403] , 
        \matrixInput[384] , \vectorInput[29] , \matrixInput[227] , 
        \matrixInput[214] , \matrixInput[117] , \matrixInput[124] , 
        \matrixInput[32] , \matrixInput[1] , \matrixInput[18] , 
        \vectorInput[24] , \vectorInput[17] , \matrixInput[424] , 
        \matrixInput[365] , \cOutput[35] , \matrixInput[356] , 
        \matrixInput[417] , \matrixInput[390] , \matrixInput[389] , 
        \matrixInput[130] , \matrixInput[129] , \matrixInput[233] , 
        \matrixInput[219] , \matrixInput[103] , \matrixInput[200] , 
        \vectorInput[1] , \matrixInput[371] , \matrixInput[342] , 
        \matrixInput[368] , \matrixInput[15] , \matrixInput[26] , 
        \cOutput[38] , \cOutput[21] , \cOutput[12] , \matrixInput[378] , 
        \matrixInput[361] , \matrixInput[352] , \cOutput[31] , \cOutput[28] , 
        \vectorInput[34] , \vectorInput[8] , \matrixInput[210] , 
        \matrixInput[113] , \matrixInput[36] , \matrixInput[5] , 
        \matrixInput[209] , \matrixInput[434] , \matrixInput[407] , 
        \matrixInput[399] , \matrixInput[380] , \matrixInput[223] , 
        \matrixInput[139] , \matrixInput[120] , \vectorInput[25] , 
        \vectorInput[16] , \matrixInput[232] , \matrixInput[218] , 
        \matrixInput[201] , \matrixInput[131] , \matrixInput[128] , 
        \matrixInput[425] , \matrixInput[102] , \matrixInput[416] , 
        \matrixInput[391] , \matrixInput[388] , \matrixInput[370] , 
        \matrixInput[369] , \matrixInput[343] , \cOutput[39] , \cOutput[20] , 
        \vectorInput[9] , \vectorInput[0] , \matrixInput[27] , 
        \matrixInput[14] , \cOutput[13] , \matrixInput[379] , 
        \matrixInput[360] , \matrixInput[353] , \matrixInput[37] , 
        \matrixInput[4] , \vectorInput[35] , \matrixInput[435] , 
        \matrixInput[406] , \cOutput[30] , \cOutput[29] , \matrixInput[398] , 
        \matrixInput[381] , \matrixInput[211] , \matrixInput[208] , 
        \matrixInput[222] , \matrixInput[112] , \matrixInput[138] , 
        \matrixInput[121] , \vectorInput[4] , \matrixInput[10] , 
        \matrixInput[23] , \matrixInput[9] , \cOutput[24] , \cOutput[17] , 
        \matrixInput[374] , \matrixInput[347] , \vectorInput[38] , 
        \vectorInput[21] , \vectorInput[12] , \matrixInput[438] , 
        \matrixInput[421] , \matrixInput[412] , \matrixInput[395] , 
        \matrixInput[236] , \matrixInput[135] , \matrixInput[106] , 
        \matrixInput[205] , \vectorInput[31] , \vectorInput[28] , 
        \matrixInput[116] , \matrixInput[431] , \matrixInput[402] , 
        \matrixInput[385] , \matrixInput[226] , \matrixInput[215] , 
        \matrixInput[125] , \matrixInput[428] , \cOutput[34] , 
        \matrixInput[364] , \matrixInput[33] , \matrixInput[0] , 
        \matrixInput[19] , \matrixInput[357] , \matrixInput[366] , 
        \matrixInput[31] , \matrixInput[28] , \cOutput[36] , \matrixInput[2] , 
        \matrixInput[355] , \vectorInput[33] , \matrixInput[217] , 
        \vectorInput[23] , \vectorInput[19] , \matrixInput[114] , 
        \vectorInput[10] , \matrixInput[433] , \matrixInput[419] , 
        \matrixInput[400] , \matrixInput[224] , \matrixInput[127] , 
        \matrixInput[387] , \matrixInput[423] , \matrixInput[410] , 
        \matrixInput[409] , \matrixInput[397] , \matrixInput[234] , 
        \matrixInput[207] , \matrixInput[137] , \matrixInput[104] , 
        \matrixInput[12] , \vectorInput[6] , \matrixInput[38] , 
        \matrixInput[21] , \cOutput[26] , \cOutput[15] , \vectorInput[37] , 
        \matrixInput[437] , \matrixInput[404] , \matrixInput[383] , 
        \matrixInput[376] , \matrixInput[345] , \matrixInput[110] , 
        \matrixInput[109] , \matrixInput[239] , \matrixInput[213] , 
        \matrixInput[123] , \matrixInput[220] , \matrixInput[362] , 
        \matrixInput[351] , \matrixInput[348] , \matrixInput[35] , 
        \matrixInput[6] , \cOutput[18] , \cOutput[32] , \matrixInput[372] , 
        \matrixInput[358] , \matrixInput[341] , \cOutput[22] , 
        \vectorInput[27] , \vectorInput[14] , \vectorInput[2] , 
        \matrixInput[16] , \cOutput[11] , \matrixInput[230] , 
        \matrixInput[133] , \matrixInput[25] , \matrixInput[229] , 
        \matrixInput[119] , \matrixInput[100] , \matrixInput[490] , 
        \matrixInput[427] , \matrixInput[203] , \matrixInput[414] , 
        \matrixInput[393] , \matrixInput[324] , \matrixInput[73] , 
        \matrixInput[59] , \matrixInput[40] , \cOutput[47] , 
        \matrixInput[489] , \matrixInput[317] , \matrixInput[287] , 
        \vectorInput[52] , \vectorInput[42] , \matrixInput[500] , \cOutput[5] , 
        \matrixInput[471] , \matrixInput[468] , \matrixInput[442] , 
        \matrixInput[184] , \matrixInput[92] , \matrixInput[266] , 
        \matrixInput[255] , \matrixInput[156] , \matrixInput[165] , 
        \matrixInput[276] , \matrixInput[175] , \matrixInput[82] , 
        \vectorInput[61] , \matrixInput[146] , \matrixInput[478] , 
        \matrixInput[461] , \matrixInput[245] , \matrixInput[452] , 
        \cOutput[57] , \matrixInput[50] , \matrixInput[49] , \vectorInput[46] , 
        \matrixInput[510] , \matrixInput[509] , \matrixInput[297] , 
        \matrixInput[63] , \matrixInput[499] , \matrixInput[194] , 
        \matrixInput[480] , \matrixInput[334] , \matrixInput[307] , 
        \matrixInput[251] , \matrixInput[248] , \matrixInput[152] , 
        \matrixInput[504] , \matrixInput[475] , \matrixInput[446] , 
        \matrixInput[262] , \matrixInput[178] , \matrixInput[161] , 
        \matrixInput[199] , \matrixInput[180] , \matrixInput[96] , 
        \cOutput[1] , \matrixInput[494] , \matrixInput[339] , 
        \matrixInput[283] , \matrixInput[320] , \matrixInput[313] , 
        \matrixInput[77] , \cOutput[43] , \matrixInput[44] , 
        \matrixInput[484] , \matrixInput[303] , \matrixInput[330] , 
        \matrixInput[329] , \matrixInput[293] , \matrixInput[190] , 
        \matrixInput[189] , \cOutput[8] , \matrixInput[54] , \matrixInput[67] , 
        \vectorInput[56] , \matrixInput[465] , \cOutput[60] , \cOutput[53] , 
        \matrixInput[456] , \matrixInput[272] , \matrixInput[258] , 
        \matrixInput[171] , \matrixInput[168] , \matrixInput[241] , 
        \matrixInput[142] , \vectorInput[54] , \matrixInput[467] , 
        \matrixInput[86] , \matrixInput[454] , \matrixInput[270] , 
        \matrixInput[269] , \matrixInput[173] , \matrixInput[140] , 
        \matrixInput[486] , \matrixInput[243] , \matrixInput[159] , 
        \matrixInput[84] , \matrixInput[332] , \matrixInput[318] , 
        \matrixInput[301] , \matrixInput[291] , \matrixInput[288] , 
        \matrixInput[192] , \matrixInput[56] , \matrixInput[506] , 
        \matrixInput[298] , \matrixInput[65] , \cOutput[62] , \cOutput[51] , 
        \cOutput[48] , \matrixInput[281] , \cOutput[3] , \matrixInput[496] , 
        \matrixInput[322] , \matrixInput[182] , \matrixInput[311] , 
        \matrixInput[308] , \cOutput[58] , \cOutput[41] , \matrixInput[149] , 
        \matrixInput[75] , \matrixInput[46] , \vectorInput[44] , 
        \matrixInput[279] , \matrixInput[260] , \matrixInput[253] , 
        \matrixInput[150] , \matrixInput[163] , \matrixInput[477] , 
        \matrixInput[444] , \matrixInput[94] , \matrixInput[52] , 
        \cOutput[55] , \matrixInput[78] , \matrixInput[61] , \vectorInput[63] , 
        \vectorInput[50] , \vectorInput[49] , \matrixInput[482] , 
        \matrixInput[305] , \matrixInput[295] , \matrixInput[196] , 
        \matrixInput[336] , \matrixInput[99] , \matrixInput[80] , 
        \matrixInput[274] , \matrixInput[247] , \matrixInput[177] , 
        \vectorInput[59] , \vectorInput[40] , \matrixInput[473] , 
        \matrixInput[463] , \matrixInput[144] , \matrixInput[459] , 
        \matrixInput[450] , \matrixInput[449] , \matrixInput[90] , 
        \matrixInput[89] , \matrixInput[440] , \matrixInput[257] , 
        \matrixInput[154] , \matrixInput[502] , \matrixInput[492] , 
        \matrixInput[326] , \matrixInput[264] , \matrixInput[167] , 
        \matrixInput[71] , \matrixInput[68] , \matrixInput[42] , \cOutput[45] , 
        \matrixInput[315] , \matrixInput[186] , \matrixInput[285] , 
        \cOutput[7] ;
    IntMatMul_Control_pVectorSize8_pWordSize8_pScan1 U_IntMatMul_Control ( 
        .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(
        DataIn), .DataOut(DataOut), .vectorInput({\vectorInput[63] , 
        \vectorInput[62] , \vectorInput[61] , \vectorInput[60] , 
        \vectorInput[59] , \vectorInput[58] , \vectorInput[57] , 
        \vectorInput[56] , \vectorInput[55] , \vectorInput[54] , 
        \vectorInput[53] , \vectorInput[52] , \vectorInput[51] , 
        \vectorInput[50] , \vectorInput[49] , \vectorInput[48] , 
        \vectorInput[47] , \vectorInput[46] , \vectorInput[45] , 
        \vectorInput[44] , \vectorInput[43] , \vectorInput[42] , 
        \vectorInput[41] , \vectorInput[40] , \vectorInput[39] , 
        \vectorInput[38] , \vectorInput[37] , \vectorInput[36] , 
        \vectorInput[35] , \vectorInput[34] , \vectorInput[33] , 
        \vectorInput[32] , \vectorInput[31] , \vectorInput[30] , 
        \vectorInput[29] , \vectorInput[28] , \vectorInput[27] , 
        \vectorInput[26] , \vectorInput[25] , \vectorInput[24] , 
        \vectorInput[23] , \vectorInput[22] , \vectorInput[21] , 
        \vectorInput[20] , \vectorInput[19] , \vectorInput[18] , 
        \vectorInput[17] , \vectorInput[16] , \vectorInput[15] , 
        \vectorInput[14] , \vectorInput[13] , \vectorInput[12] , 
        \vectorInput[11] , \vectorInput[10] , \vectorInput[9] , 
        \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , 
        \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , 
        \vectorInput[0] }), .matrixInput({\matrixInput[511] , 
        \matrixInput[510] , \matrixInput[509] , \matrixInput[508] , 
        \matrixInput[507] , \matrixInput[506] , \matrixInput[505] , 
        \matrixInput[504] , \matrixInput[503] , \matrixInput[502] , 
        \matrixInput[501] , \matrixInput[500] , \matrixInput[499] , 
        \matrixInput[498] , \matrixInput[497] , \matrixInput[496] , 
        \matrixInput[495] , \matrixInput[494] , \matrixInput[493] , 
        \matrixInput[492] , \matrixInput[491] , \matrixInput[490] , 
        \matrixInput[489] , \matrixInput[488] , \matrixInput[487] , 
        \matrixInput[486] , \matrixInput[485] , \matrixInput[484] , 
        \matrixInput[483] , \matrixInput[482] , \matrixInput[481] , 
        \matrixInput[480] , \matrixInput[479] , \matrixInput[478] , 
        \matrixInput[477] , \matrixInput[476] , \matrixInput[475] , 
        \matrixInput[474] , \matrixInput[473] , \matrixInput[472] , 
        \matrixInput[471] , \matrixInput[470] , \matrixInput[469] , 
        \matrixInput[468] , \matrixInput[467] , \matrixInput[466] , 
        \matrixInput[465] , \matrixInput[464] , \matrixInput[463] , 
        \matrixInput[462] , \matrixInput[461] , \matrixInput[460] , 
        \matrixInput[459] , \matrixInput[458] , \matrixInput[457] , 
        \matrixInput[456] , \matrixInput[455] , \matrixInput[454] , 
        \matrixInput[453] , \matrixInput[452] , \matrixInput[451] , 
        \matrixInput[450] , \matrixInput[449] , \matrixInput[448] , 
        \matrixInput[447] , \matrixInput[446] , \matrixInput[445] , 
        \matrixInput[444] , \matrixInput[443] , \matrixInput[442] , 
        \matrixInput[441] , \matrixInput[440] , \matrixInput[439] , 
        \matrixInput[438] , \matrixInput[437] , \matrixInput[436] , 
        \matrixInput[435] , \matrixInput[434] , \matrixInput[433] , 
        \matrixInput[432] , \matrixInput[431] , \matrixInput[430] , 
        \matrixInput[429] , \matrixInput[428] , \matrixInput[427] , 
        \matrixInput[426] , \matrixInput[425] , \matrixInput[424] , 
        \matrixInput[423] , \matrixInput[422] , \matrixInput[421] , 
        \matrixInput[420] , \matrixInput[419] , \matrixInput[418] , 
        \matrixInput[417] , \matrixInput[416] , \matrixInput[415] , 
        \matrixInput[414] , \matrixInput[413] , \matrixInput[412] , 
        \matrixInput[411] , \matrixInput[410] , \matrixInput[409] , 
        \matrixInput[408] , \matrixInput[407] , \matrixInput[406] , 
        \matrixInput[405] , \matrixInput[404] , \matrixInput[403] , 
        \matrixInput[402] , \matrixInput[401] , \matrixInput[400] , 
        \matrixInput[399] , \matrixInput[398] , \matrixInput[397] , 
        \matrixInput[396] , \matrixInput[395] , \matrixInput[394] , 
        \matrixInput[393] , \matrixInput[392] , \matrixInput[391] , 
        \matrixInput[390] , \matrixInput[389] , \matrixInput[388] , 
        \matrixInput[387] , \matrixInput[386] , \matrixInput[385] , 
        \matrixInput[384] , \matrixInput[383] , \matrixInput[382] , 
        \matrixInput[381] , \matrixInput[380] , \matrixInput[379] , 
        \matrixInput[378] , \matrixInput[377] , \matrixInput[376] , 
        \matrixInput[375] , \matrixInput[374] , \matrixInput[373] , 
        \matrixInput[372] , \matrixInput[371] , \matrixInput[370] , 
        \matrixInput[369] , \matrixInput[368] , \matrixInput[367] , 
        \matrixInput[366] , \matrixInput[365] , \matrixInput[364] , 
        \matrixInput[363] , \matrixInput[362] , \matrixInput[361] , 
        \matrixInput[360] , \matrixInput[359] , \matrixInput[358] , 
        \matrixInput[357] , \matrixInput[356] , \matrixInput[355] , 
        \matrixInput[354] , \matrixInput[353] , \matrixInput[352] , 
        \matrixInput[351] , \matrixInput[350] , \matrixInput[349] , 
        \matrixInput[348] , \matrixInput[347] , \matrixInput[346] , 
        \matrixInput[345] , \matrixInput[344] , \matrixInput[343] , 
        \matrixInput[342] , \matrixInput[341] , \matrixInput[340] , 
        \matrixInput[339] , \matrixInput[338] , \matrixInput[337] , 
        \matrixInput[336] , \matrixInput[335] , \matrixInput[334] , 
        \matrixInput[333] , \matrixInput[332] , \matrixInput[331] , 
        \matrixInput[330] , \matrixInput[329] , \matrixInput[328] , 
        \matrixInput[327] , \matrixInput[326] , \matrixInput[325] , 
        \matrixInput[324] , \matrixInput[323] , \matrixInput[322] , 
        \matrixInput[321] , \matrixInput[320] , \matrixInput[319] , 
        \matrixInput[318] , \matrixInput[317] , \matrixInput[316] , 
        \matrixInput[315] , \matrixInput[314] , \matrixInput[313] , 
        \matrixInput[312] , \matrixInput[311] , \matrixInput[310] , 
        \matrixInput[309] , \matrixInput[308] , \matrixInput[307] , 
        \matrixInput[306] , \matrixInput[305] , \matrixInput[304] , 
        \matrixInput[303] , \matrixInput[302] , \matrixInput[301] , 
        \matrixInput[300] , \matrixInput[299] , \matrixInput[298] , 
        \matrixInput[297] , \matrixInput[296] , \matrixInput[295] , 
        \matrixInput[294] , \matrixInput[293] , \matrixInput[292] , 
        \matrixInput[291] , \matrixInput[290] , \matrixInput[289] , 
        \matrixInput[288] , \matrixInput[287] , \matrixInput[286] , 
        \matrixInput[285] , \matrixInput[284] , \matrixInput[283] , 
        \matrixInput[282] , \matrixInput[281] , \matrixInput[280] , 
        \matrixInput[279] , \matrixInput[278] , \matrixInput[277] , 
        \matrixInput[276] , \matrixInput[275] , \matrixInput[274] , 
        \matrixInput[273] , \matrixInput[272] , \matrixInput[271] , 
        \matrixInput[270] , \matrixInput[269] , \matrixInput[268] , 
        \matrixInput[267] , \matrixInput[266] , \matrixInput[265] , 
        \matrixInput[264] , \matrixInput[263] , \matrixInput[262] , 
        \matrixInput[261] , \matrixInput[260] , \matrixInput[259] , 
        \matrixInput[258] , \matrixInput[257] , \matrixInput[256] , 
        \matrixInput[255] , \matrixInput[254] , \matrixInput[253] , 
        \matrixInput[252] , \matrixInput[251] , \matrixInput[250] , 
        \matrixInput[249] , \matrixInput[248] , \matrixInput[247] , 
        \matrixInput[246] , \matrixInput[245] , \matrixInput[244] , 
        \matrixInput[243] , \matrixInput[242] , \matrixInput[241] , 
        \matrixInput[240] , \matrixInput[239] , \matrixInput[238] , 
        \matrixInput[237] , \matrixInput[236] , \matrixInput[235] , 
        \matrixInput[234] , \matrixInput[233] , \matrixInput[232] , 
        \matrixInput[231] , \matrixInput[230] , \matrixInput[229] , 
        \matrixInput[228] , \matrixInput[227] , \matrixInput[226] , 
        \matrixInput[225] , \matrixInput[224] , \matrixInput[223] , 
        \matrixInput[222] , \matrixInput[221] , \matrixInput[220] , 
        \matrixInput[219] , \matrixInput[218] , \matrixInput[217] , 
        \matrixInput[216] , \matrixInput[215] , \matrixInput[214] , 
        \matrixInput[213] , \matrixInput[212] , \matrixInput[211] , 
        \matrixInput[210] , \matrixInput[209] , \matrixInput[208] , 
        \matrixInput[207] , \matrixInput[206] , \matrixInput[205] , 
        \matrixInput[204] , \matrixInput[203] , \matrixInput[202] , 
        \matrixInput[201] , \matrixInput[200] , \matrixInput[199] , 
        \matrixInput[198] , \matrixInput[197] , \matrixInput[196] , 
        \matrixInput[195] , \matrixInput[194] , \matrixInput[193] , 
        \matrixInput[192] , \matrixInput[191] , \matrixInput[190] , 
        \matrixInput[189] , \matrixInput[188] , \matrixInput[187] , 
        \matrixInput[186] , \matrixInput[185] , \matrixInput[184] , 
        \matrixInput[183] , \matrixInput[182] , \matrixInput[181] , 
        \matrixInput[180] , \matrixInput[179] , \matrixInput[178] , 
        \matrixInput[177] , \matrixInput[176] , \matrixInput[175] , 
        \matrixInput[174] , \matrixInput[173] , \matrixInput[172] , 
        \matrixInput[171] , \matrixInput[170] , \matrixInput[169] , 
        \matrixInput[168] , \matrixInput[167] , \matrixInput[166] , 
        \matrixInput[165] , \matrixInput[164] , \matrixInput[163] , 
        \matrixInput[162] , \matrixInput[161] , \matrixInput[160] , 
        \matrixInput[159] , \matrixInput[158] , \matrixInput[157] , 
        \matrixInput[156] , \matrixInput[155] , \matrixInput[154] , 
        \matrixInput[153] , \matrixInput[152] , \matrixInput[151] , 
        \matrixInput[150] , \matrixInput[149] , \matrixInput[148] , 
        \matrixInput[147] , \matrixInput[146] , \matrixInput[145] , 
        \matrixInput[144] , \matrixInput[143] , \matrixInput[142] , 
        \matrixInput[141] , \matrixInput[140] , \matrixInput[139] , 
        \matrixInput[138] , \matrixInput[137] , \matrixInput[136] , 
        \matrixInput[135] , \matrixInput[134] , \matrixInput[133] , 
        \matrixInput[132] , \matrixInput[131] , \matrixInput[130] , 
        \matrixInput[129] , \matrixInput[128] , \matrixInput[127] , 
        \matrixInput[126] , \matrixInput[125] , \matrixInput[124] , 
        \matrixInput[123] , \matrixInput[122] , \matrixInput[121] , 
        \matrixInput[120] , \matrixInput[119] , \matrixInput[118] , 
        \matrixInput[117] , \matrixInput[116] , \matrixInput[115] , 
        \matrixInput[114] , \matrixInput[113] , \matrixInput[112] , 
        \matrixInput[111] , \matrixInput[110] , \matrixInput[109] , 
        \matrixInput[108] , \matrixInput[107] , \matrixInput[106] , 
        \matrixInput[105] , \matrixInput[104] , \matrixInput[103] , 
        \matrixInput[102] , \matrixInput[101] , \matrixInput[100] , 
        \matrixInput[99] , \matrixInput[98] , \matrixInput[97] , 
        \matrixInput[96] , \matrixInput[95] , \matrixInput[94] , 
        \matrixInput[93] , \matrixInput[92] , \matrixInput[91] , 
        \matrixInput[90] , \matrixInput[89] , \matrixInput[88] , 
        \matrixInput[87] , \matrixInput[86] , \matrixInput[85] , 
        \matrixInput[84] , \matrixInput[83] , \matrixInput[82] , 
        \matrixInput[81] , \matrixInput[80] , \matrixInput[79] , 
        \matrixInput[78] , \matrixInput[77] , \matrixInput[76] , 
        \matrixInput[75] , \matrixInput[74] , \matrixInput[73] , 
        \matrixInput[72] , \matrixInput[71] , \matrixInput[70] , 
        \matrixInput[69] , \matrixInput[68] , \matrixInput[67] , 
        \matrixInput[66] , \matrixInput[65] , \matrixInput[64] , 
        \matrixInput[63] , \matrixInput[62] , \matrixInput[61] , 
        \matrixInput[60] , \matrixInput[59] , \matrixInput[58] , 
        \matrixInput[57] , \matrixInput[56] , \matrixInput[55] , 
        \matrixInput[54] , \matrixInput[53] , \matrixInput[52] , 
        \matrixInput[51] , \matrixInput[50] , \matrixInput[49] , 
        \matrixInput[48] , \matrixInput[47] , \matrixInput[46] , 
        \matrixInput[45] , \matrixInput[44] , \matrixInput[43] , 
        \matrixInput[42] , \matrixInput[41] , \matrixInput[40] , 
        \matrixInput[39] , \matrixInput[38] , \matrixInput[37] , 
        \matrixInput[36] , \matrixInput[35] , \matrixInput[34] , 
        \matrixInput[33] , \matrixInput[32] , \matrixInput[31] , 
        \matrixInput[30] , \matrixInput[29] , \matrixInput[28] , 
        \matrixInput[27] , \matrixInput[26] , \matrixInput[25] , 
        \matrixInput[24] , \matrixInput[23] , \matrixInput[22] , 
        \matrixInput[21] , \matrixInput[20] , \matrixInput[19] , 
        \matrixInput[18] , \matrixInput[17] , \matrixInput[16] , 
        \matrixInput[15] , \matrixInput[14] , \matrixInput[13] , 
        \matrixInput[12] , \matrixInput[11] , \matrixInput[10] , 
        \matrixInput[9] , \matrixInput[8] , \matrixInput[7] , \matrixInput[6] , 
        \matrixInput[5] , \matrixInput[4] , \matrixInput[3] , \matrixInput[2] , 
        \matrixInput[1] , \matrixInput[0] }), .cOutput({\cOutput[63] , 
        \cOutput[62] , \cOutput[61] , \cOutput[60] , \cOutput[59] , 
        \cOutput[58] , \cOutput[57] , \cOutput[56] , \cOutput[55] , 
        \cOutput[54] , \cOutput[53] , \cOutput[52] , \cOutput[51] , 
        \cOutput[50] , \cOutput[49] , \cOutput[48] , \cOutput[47] , 
        \cOutput[46] , \cOutput[45] , \cOutput[44] , \cOutput[43] , 
        \cOutput[42] , \cOutput[41] , \cOutput[40] , \cOutput[39] , 
        \cOutput[38] , \cOutput[37] , \cOutput[36] , \cOutput[35] , 
        \cOutput[34] , \cOutput[33] , \cOutput[32] , \cOutput[31] , 
        \cOutput[30] , \cOutput[29] , \cOutput[28] , \cOutput[27] , 
        \cOutput[26] , \cOutput[25] , \cOutput[24] , \cOutput[23] , 
        \cOutput[22] , \cOutput[21] , \cOutput[20] , \cOutput[19] , 
        \cOutput[18] , \cOutput[17] , \cOutput[16] , \cOutput[15] , 
        \cOutput[14] , \cOutput[13] , \cOutput[12] , \cOutput[11] , 
        \cOutput[10] , \cOutput[9] , \cOutput[8] , \cOutput[7] , \cOutput[6] , 
        \cOutput[5] , \cOutput[4] , \cOutput[3] , \cOutput[2] , \cOutput[1] , 
        \cOutput[0] }) );
    VectorDotProduct_pVectorSize8_pWordSize8 VectorDotProduct_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[63] , \vectorInput[62] , 
        \vectorInput[61] , \vectorInput[60] , \vectorInput[59] , 
        \vectorInput[58] , \vectorInput[57] , \vectorInput[56] , 
        \vectorInput[55] , \vectorInput[54] , \vectorInput[53] , 
        \vectorInput[52] , \vectorInput[51] , \vectorInput[50] , 
        \vectorInput[49] , \vectorInput[48] , \vectorInput[47] , 
        \vectorInput[46] , \vectorInput[45] , \vectorInput[44] , 
        \vectorInput[43] , \vectorInput[42] , \vectorInput[41] , 
        \vectorInput[40] , \vectorInput[39] , \vectorInput[38] , 
        \vectorInput[37] , \vectorInput[36] , \vectorInput[35] , 
        \vectorInput[34] , \vectorInput[33] , \vectorInput[32] , 
        \vectorInput[31] , \vectorInput[30] , \vectorInput[29] , 
        \vectorInput[28] , \vectorInput[27] , \vectorInput[26] , 
        \vectorInput[25] , \vectorInput[24] , \vectorInput[23] , 
        \vectorInput[22] , \vectorInput[21] , \vectorInput[20] , 
        \vectorInput[19] , \vectorInput[18] , \vectorInput[17] , 
        \vectorInput[16] , \vectorInput[15] , \vectorInput[14] , 
        \vectorInput[13] , \vectorInput[12] , \vectorInput[11] , 
        \vectorInput[10] , \vectorInput[9] , \vectorInput[8] , 
        \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , \vectorInput[4] , 
        \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , \vectorInput[0] 
        }), .vectorBInput({\matrixInput[127] , \matrixInput[126] , 
        \matrixInput[125] , \matrixInput[124] , \matrixInput[123] , 
        \matrixInput[122] , \matrixInput[121] , \matrixInput[120] , 
        \matrixInput[119] , \matrixInput[118] , \matrixInput[117] , 
        \matrixInput[116] , \matrixInput[115] , \matrixInput[114] , 
        \matrixInput[113] , \matrixInput[112] , \matrixInput[111] , 
        \matrixInput[110] , \matrixInput[109] , \matrixInput[108] , 
        \matrixInput[107] , \matrixInput[106] , \matrixInput[105] , 
        \matrixInput[104] , \matrixInput[103] , \matrixInput[102] , 
        \matrixInput[101] , \matrixInput[100] , \matrixInput[99] , 
        \matrixInput[98] , \matrixInput[97] , \matrixInput[96] , 
        \matrixInput[95] , \matrixInput[94] , \matrixInput[93] , 
        \matrixInput[92] , \matrixInput[91] , \matrixInput[90] , 
        \matrixInput[89] , \matrixInput[88] , \matrixInput[87] , 
        \matrixInput[86] , \matrixInput[85] , \matrixInput[84] , 
        \matrixInput[83] , \matrixInput[82] , \matrixInput[81] , 
        \matrixInput[80] , \matrixInput[79] , \matrixInput[78] , 
        \matrixInput[77] , \matrixInput[76] , \matrixInput[75] , 
        \matrixInput[74] , \matrixInput[73] , \matrixInput[72] , 
        \matrixInput[71] , \matrixInput[70] , \matrixInput[69] , 
        \matrixInput[68] , \matrixInput[67] , \matrixInput[66] , 
        \matrixInput[65] , \matrixInput[64] }), .cOutput({\cOutput[15] , 
        \cOutput[14] , \cOutput[13] , \cOutput[12] , \cOutput[11] , 
        \cOutput[10] , \cOutput[9] , \cOutput[8] }) );
    VectorDotProduct_pVectorSize8_pWordSize8 VectorDotProduct_2 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[63] , \vectorInput[62] , 
        \vectorInput[61] , \vectorInput[60] , \vectorInput[59] , 
        \vectorInput[58] , \vectorInput[57] , \vectorInput[56] , 
        \vectorInput[55] , \vectorInput[54] , \vectorInput[53] , 
        \vectorInput[52] , \vectorInput[51] , \vectorInput[50] , 
        \vectorInput[49] , \vectorInput[48] , \vectorInput[47] , 
        \vectorInput[46] , \vectorInput[45] , \vectorInput[44] , 
        \vectorInput[43] , \vectorInput[42] , \vectorInput[41] , 
        \vectorInput[40] , \vectorInput[39] , \vectorInput[38] , 
        \vectorInput[37] , \vectorInput[36] , \vectorInput[35] , 
        \vectorInput[34] , \vectorInput[33] , \vectorInput[32] , 
        \vectorInput[31] , \vectorInput[30] , \vectorInput[29] , 
        \vectorInput[28] , \vectorInput[27] , \vectorInput[26] , 
        \vectorInput[25] , \vectorInput[24] , \vectorInput[23] , 
        \vectorInput[22] , \vectorInput[21] , \vectorInput[20] , 
        \vectorInput[19] , \vectorInput[18] , \vectorInput[17] , 
        \vectorInput[16] , \vectorInput[15] , \vectorInput[14] , 
        \vectorInput[13] , \vectorInput[12] , \vectorInput[11] , 
        \vectorInput[10] , \vectorInput[9] , \vectorInput[8] , 
        \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , \vectorInput[4] , 
        \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , \vectorInput[0] 
        }), .vectorBInput({\matrixInput[191] , \matrixInput[190] , 
        \matrixInput[189] , \matrixInput[188] , \matrixInput[187] , 
        \matrixInput[186] , \matrixInput[185] , \matrixInput[184] , 
        \matrixInput[183] , \matrixInput[182] , \matrixInput[181] , 
        \matrixInput[180] , \matrixInput[179] , \matrixInput[178] , 
        \matrixInput[177] , \matrixInput[176] , \matrixInput[175] , 
        \matrixInput[174] , \matrixInput[173] , \matrixInput[172] , 
        \matrixInput[171] , \matrixInput[170] , \matrixInput[169] , 
        \matrixInput[168] , \matrixInput[167] , \matrixInput[166] , 
        \matrixInput[165] , \matrixInput[164] , \matrixInput[163] , 
        \matrixInput[162] , \matrixInput[161] , \matrixInput[160] , 
        \matrixInput[159] , \matrixInput[158] , \matrixInput[157] , 
        \matrixInput[156] , \matrixInput[155] , \matrixInput[154] , 
        \matrixInput[153] , \matrixInput[152] , \matrixInput[151] , 
        \matrixInput[150] , \matrixInput[149] , \matrixInput[148] , 
        \matrixInput[147] , \matrixInput[146] , \matrixInput[145] , 
        \matrixInput[144] , \matrixInput[143] , \matrixInput[142] , 
        \matrixInput[141] , \matrixInput[140] , \matrixInput[139] , 
        \matrixInput[138] , \matrixInput[137] , \matrixInput[136] , 
        \matrixInput[135] , \matrixInput[134] , \matrixInput[133] , 
        \matrixInput[132] , \matrixInput[131] , \matrixInput[130] , 
        \matrixInput[129] , \matrixInput[128] }), .cOutput({\cOutput[23] , 
        \cOutput[22] , \cOutput[21] , \cOutput[20] , \cOutput[19] , 
        \cOutput[18] , \cOutput[17] , \cOutput[16] }) );
    VectorDotProduct_pVectorSize8_pWordSize8 VectorDotProduct_3 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[63] , \vectorInput[62] , 
        \vectorInput[61] , \vectorInput[60] , \vectorInput[59] , 
        \vectorInput[58] , \vectorInput[57] , \vectorInput[56] , 
        \vectorInput[55] , \vectorInput[54] , \vectorInput[53] , 
        \vectorInput[52] , \vectorInput[51] , \vectorInput[50] , 
        \vectorInput[49] , \vectorInput[48] , \vectorInput[47] , 
        \vectorInput[46] , \vectorInput[45] , \vectorInput[44] , 
        \vectorInput[43] , \vectorInput[42] , \vectorInput[41] , 
        \vectorInput[40] , \vectorInput[39] , \vectorInput[38] , 
        \vectorInput[37] , \vectorInput[36] , \vectorInput[35] , 
        \vectorInput[34] , \vectorInput[33] , \vectorInput[32] , 
        \vectorInput[31] , \vectorInput[30] , \vectorInput[29] , 
        \vectorInput[28] , \vectorInput[27] , \vectorInput[26] , 
        \vectorInput[25] , \vectorInput[24] , \vectorInput[23] , 
        \vectorInput[22] , \vectorInput[21] , \vectorInput[20] , 
        \vectorInput[19] , \vectorInput[18] , \vectorInput[17] , 
        \vectorInput[16] , \vectorInput[15] , \vectorInput[14] , 
        \vectorInput[13] , \vectorInput[12] , \vectorInput[11] , 
        \vectorInput[10] , \vectorInput[9] , \vectorInput[8] , 
        \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , \vectorInput[4] , 
        \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , \vectorInput[0] 
        }), .vectorBInput({\matrixInput[255] , \matrixInput[254] , 
        \matrixInput[253] , \matrixInput[252] , \matrixInput[251] , 
        \matrixInput[250] , \matrixInput[249] , \matrixInput[248] , 
        \matrixInput[247] , \matrixInput[246] , \matrixInput[245] , 
        \matrixInput[244] , \matrixInput[243] , \matrixInput[242] , 
        \matrixInput[241] , \matrixInput[240] , \matrixInput[239] , 
        \matrixInput[238] , \matrixInput[237] , \matrixInput[236] , 
        \matrixInput[235] , \matrixInput[234] , \matrixInput[233] , 
        \matrixInput[232] , \matrixInput[231] , \matrixInput[230] , 
        \matrixInput[229] , \matrixInput[228] , \matrixInput[227] , 
        \matrixInput[226] , \matrixInput[225] , \matrixInput[224] , 
        \matrixInput[223] , \matrixInput[222] , \matrixInput[221] , 
        \matrixInput[220] , \matrixInput[219] , \matrixInput[218] , 
        \matrixInput[217] , \matrixInput[216] , \matrixInput[215] , 
        \matrixInput[214] , \matrixInput[213] , \matrixInput[212] , 
        \matrixInput[211] , \matrixInput[210] , \matrixInput[209] , 
        \matrixInput[208] , \matrixInput[207] , \matrixInput[206] , 
        \matrixInput[205] , \matrixInput[204] , \matrixInput[203] , 
        \matrixInput[202] , \matrixInput[201] , \matrixInput[200] , 
        \matrixInput[199] , \matrixInput[198] , \matrixInput[197] , 
        \matrixInput[196] , \matrixInput[195] , \matrixInput[194] , 
        \matrixInput[193] , \matrixInput[192] }), .cOutput({\cOutput[31] , 
        \cOutput[30] , \cOutput[29] , \cOutput[28] , \cOutput[27] , 
        \cOutput[26] , \cOutput[25] , \cOutput[24] }) );
    VectorDotProduct_pVectorSize8_pWordSize8 VectorDotProduct_4 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[63] , \vectorInput[62] , 
        \vectorInput[61] , \vectorInput[60] , \vectorInput[59] , 
        \vectorInput[58] , \vectorInput[57] , \vectorInput[56] , 
        \vectorInput[55] , \vectorInput[54] , \vectorInput[53] , 
        \vectorInput[52] , \vectorInput[51] , \vectorInput[50] , 
        \vectorInput[49] , \vectorInput[48] , \vectorInput[47] , 
        \vectorInput[46] , \vectorInput[45] , \vectorInput[44] , 
        \vectorInput[43] , \vectorInput[42] , \vectorInput[41] , 
        \vectorInput[40] , \vectorInput[39] , \vectorInput[38] , 
        \vectorInput[37] , \vectorInput[36] , \vectorInput[35] , 
        \vectorInput[34] , \vectorInput[33] , \vectorInput[32] , 
        \vectorInput[31] , \vectorInput[30] , \vectorInput[29] , 
        \vectorInput[28] , \vectorInput[27] , \vectorInput[26] , 
        \vectorInput[25] , \vectorInput[24] , \vectorInput[23] , 
        \vectorInput[22] , \vectorInput[21] , \vectorInput[20] , 
        \vectorInput[19] , \vectorInput[18] , \vectorInput[17] , 
        \vectorInput[16] , \vectorInput[15] , \vectorInput[14] , 
        \vectorInput[13] , \vectorInput[12] , \vectorInput[11] , 
        \vectorInput[10] , \vectorInput[9] , \vectorInput[8] , 
        \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , \vectorInput[4] , 
        \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , \vectorInput[0] 
        }), .vectorBInput({\matrixInput[319] , \matrixInput[318] , 
        \matrixInput[317] , \matrixInput[316] , \matrixInput[315] , 
        \matrixInput[314] , \matrixInput[313] , \matrixInput[312] , 
        \matrixInput[311] , \matrixInput[310] , \matrixInput[309] , 
        \matrixInput[308] , \matrixInput[307] , \matrixInput[306] , 
        \matrixInput[305] , \matrixInput[304] , \matrixInput[303] , 
        \matrixInput[302] , \matrixInput[301] , \matrixInput[300] , 
        \matrixInput[299] , \matrixInput[298] , \matrixInput[297] , 
        \matrixInput[296] , \matrixInput[295] , \matrixInput[294] , 
        \matrixInput[293] , \matrixInput[292] , \matrixInput[291] , 
        \matrixInput[290] , \matrixInput[289] , \matrixInput[288] , 
        \matrixInput[287] , \matrixInput[286] , \matrixInput[285] , 
        \matrixInput[284] , \matrixInput[283] , \matrixInput[282] , 
        \matrixInput[281] , \matrixInput[280] , \matrixInput[279] , 
        \matrixInput[278] , \matrixInput[277] , \matrixInput[276] , 
        \matrixInput[275] , \matrixInput[274] , \matrixInput[273] , 
        \matrixInput[272] , \matrixInput[271] , \matrixInput[270] , 
        \matrixInput[269] , \matrixInput[268] , \matrixInput[267] , 
        \matrixInput[266] , \matrixInput[265] , \matrixInput[264] , 
        \matrixInput[263] , \matrixInput[262] , \matrixInput[261] , 
        \matrixInput[260] , \matrixInput[259] , \matrixInput[258] , 
        \matrixInput[257] , \matrixInput[256] }), .cOutput({\cOutput[39] , 
        \cOutput[38] , \cOutput[37] , \cOutput[36] , \cOutput[35] , 
        \cOutput[34] , \cOutput[33] , \cOutput[32] }) );
    VectorDotProduct_pVectorSize8_pWordSize8 VectorDotProduct_5 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[63] , \vectorInput[62] , 
        \vectorInput[61] , \vectorInput[60] , \vectorInput[59] , 
        \vectorInput[58] , \vectorInput[57] , \vectorInput[56] , 
        \vectorInput[55] , \vectorInput[54] , \vectorInput[53] , 
        \vectorInput[52] , \vectorInput[51] , \vectorInput[50] , 
        \vectorInput[49] , \vectorInput[48] , \vectorInput[47] , 
        \vectorInput[46] , \vectorInput[45] , \vectorInput[44] , 
        \vectorInput[43] , \vectorInput[42] , \vectorInput[41] , 
        \vectorInput[40] , \vectorInput[39] , \vectorInput[38] , 
        \vectorInput[37] , \vectorInput[36] , \vectorInput[35] , 
        \vectorInput[34] , \vectorInput[33] , \vectorInput[32] , 
        \vectorInput[31] , \vectorInput[30] , \vectorInput[29] , 
        \vectorInput[28] , \vectorInput[27] , \vectorInput[26] , 
        \vectorInput[25] , \vectorInput[24] , \vectorInput[23] , 
        \vectorInput[22] , \vectorInput[21] , \vectorInput[20] , 
        \vectorInput[19] , \vectorInput[18] , \vectorInput[17] , 
        \vectorInput[16] , \vectorInput[15] , \vectorInput[14] , 
        \vectorInput[13] , \vectorInput[12] , \vectorInput[11] , 
        \vectorInput[10] , \vectorInput[9] , \vectorInput[8] , 
        \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , \vectorInput[4] , 
        \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , \vectorInput[0] 
        }), .vectorBInput({\matrixInput[383] , \matrixInput[382] , 
        \matrixInput[381] , \matrixInput[380] , \matrixInput[379] , 
        \matrixInput[378] , \matrixInput[377] , \matrixInput[376] , 
        \matrixInput[375] , \matrixInput[374] , \matrixInput[373] , 
        \matrixInput[372] , \matrixInput[371] , \matrixInput[370] , 
        \matrixInput[369] , \matrixInput[368] , \matrixInput[367] , 
        \matrixInput[366] , \matrixInput[365] , \matrixInput[364] , 
        \matrixInput[363] , \matrixInput[362] , \matrixInput[361] , 
        \matrixInput[360] , \matrixInput[359] , \matrixInput[358] , 
        \matrixInput[357] , \matrixInput[356] , \matrixInput[355] , 
        \matrixInput[354] , \matrixInput[353] , \matrixInput[352] , 
        \matrixInput[351] , \matrixInput[350] , \matrixInput[349] , 
        \matrixInput[348] , \matrixInput[347] , \matrixInput[346] , 
        \matrixInput[345] , \matrixInput[344] , \matrixInput[343] , 
        \matrixInput[342] , \matrixInput[341] , \matrixInput[340] , 
        \matrixInput[339] , \matrixInput[338] , \matrixInput[337] , 
        \matrixInput[336] , \matrixInput[335] , \matrixInput[334] , 
        \matrixInput[333] , \matrixInput[332] , \matrixInput[331] , 
        \matrixInput[330] , \matrixInput[329] , \matrixInput[328] , 
        \matrixInput[327] , \matrixInput[326] , \matrixInput[325] , 
        \matrixInput[324] , \matrixInput[323] , \matrixInput[322] , 
        \matrixInput[321] , \matrixInput[320] }), .cOutput({\cOutput[47] , 
        \cOutput[46] , \cOutput[45] , \cOutput[44] , \cOutput[43] , 
        \cOutput[42] , \cOutput[41] , \cOutput[40] }) );
    VectorDotProduct_pVectorSize8_pWordSize8 VectorDotProduct_6 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[63] , \vectorInput[62] , 
        \vectorInput[61] , \vectorInput[60] , \vectorInput[59] , 
        \vectorInput[58] , \vectorInput[57] , \vectorInput[56] , 
        \vectorInput[55] , \vectorInput[54] , \vectorInput[53] , 
        \vectorInput[52] , \vectorInput[51] , \vectorInput[50] , 
        \vectorInput[49] , \vectorInput[48] , \vectorInput[47] , 
        \vectorInput[46] , \vectorInput[45] , \vectorInput[44] , 
        \vectorInput[43] , \vectorInput[42] , \vectorInput[41] , 
        \vectorInput[40] , \vectorInput[39] , \vectorInput[38] , 
        \vectorInput[37] , \vectorInput[36] , \vectorInput[35] , 
        \vectorInput[34] , \vectorInput[33] , \vectorInput[32] , 
        \vectorInput[31] , \vectorInput[30] , \vectorInput[29] , 
        \vectorInput[28] , \vectorInput[27] , \vectorInput[26] , 
        \vectorInput[25] , \vectorInput[24] , \vectorInput[23] , 
        \vectorInput[22] , \vectorInput[21] , \vectorInput[20] , 
        \vectorInput[19] , \vectorInput[18] , \vectorInput[17] , 
        \vectorInput[16] , \vectorInput[15] , \vectorInput[14] , 
        \vectorInput[13] , \vectorInput[12] , \vectorInput[11] , 
        \vectorInput[10] , \vectorInput[9] , \vectorInput[8] , 
        \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , \vectorInput[4] , 
        \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , \vectorInput[0] 
        }), .vectorBInput({\matrixInput[447] , \matrixInput[446] , 
        \matrixInput[445] , \matrixInput[444] , \matrixInput[443] , 
        \matrixInput[442] , \matrixInput[441] , \matrixInput[440] , 
        \matrixInput[439] , \matrixInput[438] , \matrixInput[437] , 
        \matrixInput[436] , \matrixInput[435] , \matrixInput[434] , 
        \matrixInput[433] , \matrixInput[432] , \matrixInput[431] , 
        \matrixInput[430] , \matrixInput[429] , \matrixInput[428] , 
        \matrixInput[427] , \matrixInput[426] , \matrixInput[425] , 
        \matrixInput[424] , \matrixInput[423] , \matrixInput[422] , 
        \matrixInput[421] , \matrixInput[420] , \matrixInput[419] , 
        \matrixInput[418] , \matrixInput[417] , \matrixInput[416] , 
        \matrixInput[415] , \matrixInput[414] , \matrixInput[413] , 
        \matrixInput[412] , \matrixInput[411] , \matrixInput[410] , 
        \matrixInput[409] , \matrixInput[408] , \matrixInput[407] , 
        \matrixInput[406] , \matrixInput[405] , \matrixInput[404] , 
        \matrixInput[403] , \matrixInput[402] , \matrixInput[401] , 
        \matrixInput[400] , \matrixInput[399] , \matrixInput[398] , 
        \matrixInput[397] , \matrixInput[396] , \matrixInput[395] , 
        \matrixInput[394] , \matrixInput[393] , \matrixInput[392] , 
        \matrixInput[391] , \matrixInput[390] , \matrixInput[389] , 
        \matrixInput[388] , \matrixInput[387] , \matrixInput[386] , 
        \matrixInput[385] , \matrixInput[384] }), .cOutput({\cOutput[55] , 
        \cOutput[54] , \cOutput[53] , \cOutput[52] , \cOutput[51] , 
        \cOutput[50] , \cOutput[49] , \cOutput[48] }) );
    VectorDotProduct_pVectorSize8_pWordSize8 VectorDotProduct_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[63] , \vectorInput[62] , 
        \vectorInput[61] , \vectorInput[60] , \vectorInput[59] , 
        \vectorInput[58] , \vectorInput[57] , \vectorInput[56] , 
        \vectorInput[55] , \vectorInput[54] , \vectorInput[53] , 
        \vectorInput[52] , \vectorInput[51] , \vectorInput[50] , 
        \vectorInput[49] , \vectorInput[48] , \vectorInput[47] , 
        \vectorInput[46] , \vectorInput[45] , \vectorInput[44] , 
        \vectorInput[43] , \vectorInput[42] , \vectorInput[41] , 
        \vectorInput[40] , \vectorInput[39] , \vectorInput[38] , 
        \vectorInput[37] , \vectorInput[36] , \vectorInput[35] , 
        \vectorInput[34] , \vectorInput[33] , \vectorInput[32] , 
        \vectorInput[31] , \vectorInput[30] , \vectorInput[29] , 
        \vectorInput[28] , \vectorInput[27] , \vectorInput[26] , 
        \vectorInput[25] , \vectorInput[24] , \vectorInput[23] , 
        \vectorInput[22] , \vectorInput[21] , \vectorInput[20] , 
        \vectorInput[19] , \vectorInput[18] , \vectorInput[17] , 
        \vectorInput[16] , \vectorInput[15] , \vectorInput[14] , 
        \vectorInput[13] , \vectorInput[12] , \vectorInput[11] , 
        \vectorInput[10] , \vectorInput[9] , \vectorInput[8] , 
        \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , \vectorInput[4] , 
        \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , \vectorInput[0] 
        }), .vectorBInput({\matrixInput[63] , \matrixInput[62] , 
        \matrixInput[61] , \matrixInput[60] , \matrixInput[59] , 
        \matrixInput[58] , \matrixInput[57] , \matrixInput[56] , 
        \matrixInput[55] , \matrixInput[54] , \matrixInput[53] , 
        \matrixInput[52] , \matrixInput[51] , \matrixInput[50] , 
        \matrixInput[49] , \matrixInput[48] , \matrixInput[47] , 
        \matrixInput[46] , \matrixInput[45] , \matrixInput[44] , 
        \matrixInput[43] , \matrixInput[42] , \matrixInput[41] , 
        \matrixInput[40] , \matrixInput[39] , \matrixInput[38] , 
        \matrixInput[37] , \matrixInput[36] , \matrixInput[35] , 
        \matrixInput[34] , \matrixInput[33] , \matrixInput[32] , 
        \matrixInput[31] , \matrixInput[30] , \matrixInput[29] , 
        \matrixInput[28] , \matrixInput[27] , \matrixInput[26] , 
        \matrixInput[25] , \matrixInput[24] , \matrixInput[23] , 
        \matrixInput[22] , \matrixInput[21] , \matrixInput[20] , 
        \matrixInput[19] , \matrixInput[18] , \matrixInput[17] , 
        \matrixInput[16] , \matrixInput[15] , \matrixInput[14] , 
        \matrixInput[13] , \matrixInput[12] , \matrixInput[11] , 
        \matrixInput[10] , \matrixInput[9] , \matrixInput[8] , 
        \matrixInput[7] , \matrixInput[6] , \matrixInput[5] , \matrixInput[4] , 
        \matrixInput[3] , \matrixInput[2] , \matrixInput[1] , \matrixInput[0] 
        }), .cOutput({\cOutput[7] , \cOutput[6] , \cOutput[5] , \cOutput[4] , 
        \cOutput[3] , \cOutput[2] , \cOutput[1] , \cOutput[0] }) );
    VectorDotProduct_pVectorSize8_pWordSize8 VectorDotProduct_7 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[63] , \vectorInput[62] , 
        \vectorInput[61] , \vectorInput[60] , \vectorInput[59] , 
        \vectorInput[58] , \vectorInput[57] , \vectorInput[56] , 
        \vectorInput[55] , \vectorInput[54] , \vectorInput[53] , 
        \vectorInput[52] , \vectorInput[51] , \vectorInput[50] , 
        \vectorInput[49] , \vectorInput[48] , \vectorInput[47] , 
        \vectorInput[46] , \vectorInput[45] , \vectorInput[44] , 
        \vectorInput[43] , \vectorInput[42] , \vectorInput[41] , 
        \vectorInput[40] , \vectorInput[39] , \vectorInput[38] , 
        \vectorInput[37] , \vectorInput[36] , \vectorInput[35] , 
        \vectorInput[34] , \vectorInput[33] , \vectorInput[32] , 
        \vectorInput[31] , \vectorInput[30] , \vectorInput[29] , 
        \vectorInput[28] , \vectorInput[27] , \vectorInput[26] , 
        \vectorInput[25] , \vectorInput[24] , \vectorInput[23] , 
        \vectorInput[22] , \vectorInput[21] , \vectorInput[20] , 
        \vectorInput[19] , \vectorInput[18] , \vectorInput[17] , 
        \vectorInput[16] , \vectorInput[15] , \vectorInput[14] , 
        \vectorInput[13] , \vectorInput[12] , \vectorInput[11] , 
        \vectorInput[10] , \vectorInput[9] , \vectorInput[8] , 
        \vectorInput[7] , \vectorInput[6] , \vectorInput[5] , \vectorInput[4] , 
        \vectorInput[3] , \vectorInput[2] , \vectorInput[1] , \vectorInput[0] 
        }), .vectorBInput({\matrixInput[511] , \matrixInput[510] , 
        \matrixInput[509] , \matrixInput[508] , \matrixInput[507] , 
        \matrixInput[506] , \matrixInput[505] , \matrixInput[504] , 
        \matrixInput[503] , \matrixInput[502] , \matrixInput[501] , 
        \matrixInput[500] , \matrixInput[499] , \matrixInput[498] , 
        \matrixInput[497] , \matrixInput[496] , \matrixInput[495] , 
        \matrixInput[494] , \matrixInput[493] , \matrixInput[492] , 
        \matrixInput[491] , \matrixInput[490] , \matrixInput[489] , 
        \matrixInput[488] , \matrixInput[487] , \matrixInput[486] , 
        \matrixInput[485] , \matrixInput[484] , \matrixInput[483] , 
        \matrixInput[482] , \matrixInput[481] , \matrixInput[480] , 
        \matrixInput[479] , \matrixInput[478] , \matrixInput[477] , 
        \matrixInput[476] , \matrixInput[475] , \matrixInput[474] , 
        \matrixInput[473] , \matrixInput[472] , \matrixInput[471] , 
        \matrixInput[470] , \matrixInput[469] , \matrixInput[468] , 
        \matrixInput[467] , \matrixInput[466] , \matrixInput[465] , 
        \matrixInput[464] , \matrixInput[463] , \matrixInput[462] , 
        \matrixInput[461] , \matrixInput[460] , \matrixInput[459] , 
        \matrixInput[458] , \matrixInput[457] , \matrixInput[456] , 
        \matrixInput[455] , \matrixInput[454] , \matrixInput[453] , 
        \matrixInput[452] , \matrixInput[451] , \matrixInput[450] , 
        \matrixInput[449] , \matrixInput[448] }), .cOutput({\cOutput[63] , 
        \cOutput[62] , \cOutput[61] , \cOutput[60] , \cOutput[59] , 
        \cOutput[58] , \cOutput[57] , \cOutput[56] }) );
endmodule

