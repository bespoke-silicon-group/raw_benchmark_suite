
module DES_Control_WIDTH64_MEMSPACE2_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, key, start, rdy
     );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
output [63:0] key;
input  Clk, Reset, RD, WR, rdy;
output ScanEnable, start;
    wire n379, n454, n468, n421, n406, n387, n433, n395, n414, n370, n461, 
        n446, n428, n408, n389, n466, n441, n377, n392, n413, n434, n401, n380, 
        n426, n448, n453, n393, n412, n435, n376, \ScanReg[15] , n467, 
        \ScanReg[26] , n440, \ScanReg[2] , n388, n409, \ScanReg[18] , n449, 
        n452, \ScanReg[11] , \ScanReg[6] , \ScanReg[22] , n400, n381, n427, 
        n407, \ScanReg[20] , \ScanReg[13] , \ScanReg[4] , n420, n386, n469, 
        n378, n455, n472, \ScanReg[29] , \ScanReg[30] , n429, \ScanReg[17] , 
        n447, \ScanReg[24] , n460, \ScanReg[0] , n371, \ScanReg[9] , n432, 
        n394, n415, n439, \ScanReg[16] , \ScanReg[25] , n470, n457, 
        \ScanReg[8] , \ScanReg[1] , \ScanReg[7] , n405, n384, n422, 
        \ScanReg[5] , n396, n417, \ScanReg[21] , \ScanReg[12] , n430, n373, 
        n368, n445, n462, \ScanReg[28] , \ScanReg[31] , \ScanReg[19] , n374, 
        n465, n442, n459, n402, n391, \ScanReg[10] , n437, n383, \ScanReg[23] , 
        n410, n425, \ScanReg[14] , \ScanReg[27] , n450, n398, \ScanReg[3] , 
        n419, n436, n390, n411, n464, n458, n375, n443, n399, n418, n451, n438, 
        n367, n403, n424, n382, n404, n385, n423, n471, n456, n369, n463, n444, 
        n372, n397, n416, n431;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U54 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_AND2 U73 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_AO22 U113 ( .A(key[63]), .B(n373), .C(DataIn[31]), .D(n374), .Z(n409)
         );
    VMW_AO22 U134 ( .A(key[44]), .B(n373), .C(DataIn[12]), .D(n374), .Z(n428)
         );
    VMW_AND2 U68 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_AND2 U96 ( .A(\ScanReg[6] ), .B(n369), .Z(n388) );
    VMW_BUFIZ U198 ( .A(n392), .E(n381), .Z(\arr[2] ) );
    VMW_BUFIZ U204 ( .A(n398), .E(n381), .Z(\arr[24] ) );
    VMW_FD \key_reg[36]  ( .D(n436), .CP(Clk), .Q(key[36]) );
    VMW_OAI21 U108 ( .A(RD), .B(WR), .C(n372), .Z(n371) );
    VMW_AO22 U141 ( .A(key[38]), .B(n373), .C(DataIn[6]), .D(n374), .Z(n434)
         );
    VMW_AO22 U166 ( .A(key[15]), .B(n373), .C(key[47]), .D(n374), .Z(n457) );
    VMW_FD \key_reg[15]  ( .D(n457), .CP(Clk), .Q(key[15]) );
    VMW_BUFIZ U183 ( .A(n376), .E(n381), .Z(\arr[19] ) );
    VMW_FD \key_reg[26]  ( .D(n446), .CP(Clk), .Q(key[26]) );
    VMW_FD \key_reg[7]  ( .D(n465), .CP(Clk), .Q(key[7]) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AND2 U46 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U61 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U84 ( .A(\ScanReg[7] ), .B(n369), .Z(n400) );
    VMW_AO22 U148 ( .A(key[31]), .B(n373), .C(key[63]), .D(n374), .Z(n441) );
    VMW_AO22 U153 ( .A(key[27]), .B(n373), .C(key[59]), .D(n374), .Z(n445) );
    VMW_AND3 U174 ( .A(n367), .B(Addr[1]), .C(Addr[0]), .Z(n370) );
    VMW_BUFIZ U191 ( .A(n385), .E(n381), .Z(\arr[25] ) );
    VMW_FD \key_reg[32]  ( .D(n440), .CP(Clk), .Q(key[32]) );
    VMW_FD \key_reg[18]  ( .D(n454), .CP(Clk), .Q(key[18]) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_FD \key_reg[3]  ( .D(n469), .CP(Clk), .Q(key[3]) );
    VMW_AND2 U101 ( .A(\ScanReg[27] ), .B(n369), .Z(n383) );
    VMW_FD \key_reg[22]  ( .D(n450), .CP(Clk), .Q(key[22]) );
    VMW_FD \key_reg[11]  ( .D(n461), .CP(Clk), .Q(key[11]) );
    VMW_AO22 U126 ( .A(key[51]), .B(n373), .C(DataIn[19]), .D(n374), .Z(n421)
         );
    VMW_AND2 U48 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U66 ( .A(DataIn[9]), .B(WR), .Z(ScanOut[9]) );
    VMW_AO21 U106 ( .A(RD), .B(ScanEnable), .C(n370), .Z(n381) );
    VMW_AO22 U121 ( .A(key[56]), .B(n373), .C(DataIn[24]), .D(n374), .Z(n416)
         );
    VMW_BUFIZ U211 ( .A(n405), .E(n381), .Z(\arr[22] ) );
    VMW_FD \key_reg[13]  ( .D(n459), .CP(Clk), .Q(key[13]) );
    VMW_FD \key_reg[1]  ( .D(n471), .CP(Clk), .Q(key[1]) );
    VMW_FD \key_reg[39]  ( .D(n433), .CP(Clk), .Q(key[39]) );
    VMW_FD \key_reg[20]  ( .D(n452), .CP(Clk), .Q(key[20]) );
    VMW_AND2 U83 ( .A(\ScanReg[5] ), .B(n369), .Z(n401) );
    VMW_AO22 U168 ( .A(key[13]), .B(n373), .C(key[45]), .D(n374), .Z(n459) );
    VMW_AND2 U98 ( .A(\ScanReg[16] ), .B(n369), .Z(n386) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(key[4]), .B(n373), .C(key[36]), .D(n374), .Z(n468) );
    VMW_AO22 U154 ( .A(key[26]), .B(n373), .C(key[58]), .D(n374), .Z(n446) );
    VMW_AO22 U173 ( .A(\ScanReg[0] ), .B(n369), .C(rdy), .D(n370), .Z(n377) );
    VMW_BUFIZ U184 ( .A(n377), .E(n381), .Z(\arr[0] ) );
    VMW_BUFIZ U196 ( .A(n390), .E(n381), .Z(\arr[21] ) );
    VMW_FD \key_reg[8]  ( .D(n464), .CP(Clk), .Q(key[8]) );
    VMW_FD \key_reg[30]  ( .D(n442), .CP(Clk), .Q(key[30]) );
    VMW_FD \key_reg[29]  ( .D(n443), .CP(Clk), .Q(key[29]) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AND2 U53 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_AND2 U91 ( .A(\ScanReg[13] ), .B(n369), .Z(n393) );
    VMW_AO22 U146 ( .A(key[33]), .B(n373), .C(DataIn[1]), .D(n374), .Z(n439)
         );
    VMW_AO22 U161 ( .A(key[1]), .B(n373), .C(key[33]), .D(n374), .Z(n471) );
    VMW_FD \key_reg[24]  ( .D(n448), .CP(Clk), .Q(key[24]) );
    VMW_FD \key_reg[17]  ( .D(n455), .CP(Clk), .Q(key[17]) );
    VMW_FD \key_reg[34]  ( .D(n438), .CP(Clk), .Q(key[34]) );
    VMW_FD \key_reg[5]  ( .D(n467), .CP(Clk), .Q(key[5]) );
    VMW_BUFIZ U203 ( .A(n397), .E(n381), .Z(\arr[3] ) );
    VMW_AND2 U74 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_AO22 U114 ( .A(key[62]), .B(n373), .C(DataIn[30]), .D(n374), .Z(n410)
         );
    VMW_AO22 U133 ( .A(key[45]), .B(n373), .C(DataIn[13]), .D(n374), .Z(n427)
         );
    VMW_AND2 U99 ( .A(\ScanReg[25] ), .B(n369), .Z(n385) );
    VMW_BUFIZ U197 ( .A(n391), .E(n381), .Z(\arr[28] ) );
    VMW_FD \key_reg[62]  ( .D(n410), .CP(Clk), .Q(key[62]) );
    VMW_FD \key_reg[51]  ( .D(n421), .CP(Clk), .Q(key[51]) );
    VMW_FD \key_reg[48]  ( .D(n424), .CP(Clk), .Q(key[48]) );
    VMW_AO22 U155 ( .A(key[25]), .B(n373), .C(key[57]), .D(n374), .Z(n447) );
    VMW_AO22 U172 ( .A(key[0]), .B(n373), .C(key[32]), .D(n374), .Z(n472) );
    VMW_AND2 U47 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U49 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_AND2 U52 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U67 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U82 ( .A(\ScanReg[26] ), .B(n369), .Z(n402) );
    VMW_AO22 U169 ( .A(key[12]), .B(n373), .C(key[44]), .D(n374), .Z(n460) );
    VMW_AND2 U107 ( .A(\ScanReg[19] ), .B(n369), .Z(n376) );
    VMW_AO22 U120 ( .A(key[57]), .B(n373), .C(DataIn[25]), .D(n374), .Z(n415)
         );
    VMW_BUFIZ U210 ( .A(n404), .E(n381), .Z(\arr[18] ) );
    VMW_FD \key_reg[58]  ( .D(n414), .CP(Clk), .Q(key[58]) );
    VMW_FD \key_reg[41]  ( .D(n431), .CP(Clk), .Q(key[41]) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U75 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_AO22 U115 ( .A(key[61]), .B(n373), .C(DataIn[29]), .D(n374), .Z(n411)
         );
    VMW_AO22 U132 ( .A(key[46]), .B(n373), .C(DataIn[14]), .D(n374), .Z(n426)
         );
    VMW_BUFIZ U202 ( .A(n396), .E(n381), .Z(\arr[20] ) );
    VMW_AND2 U90 ( .A(\ScanReg[30] ), .B(n369), .Z(n394) );
    VMW_FD \key_reg[55]  ( .D(n417), .CP(Clk), .Q(key[55]) );
    VMW_AO22 U129 ( .A(key[49]), .B(n373), .C(DataIn[17]), .D(n374), .Z(n423)
         );
    VMW_AO22 U147 ( .A(key[32]), .B(n373), .C(DataIn[0]), .D(n374), .Z(n440)
         );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_AO22 U160 ( .A(key[20]), .B(n373), .C(key[52]), .D(n374), .Z(n452) );
    VMW_FD \key_reg[45]  ( .D(n427), .CP(Clk), .Q(key[45]) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_BUFIZ U185 ( .A(n378), .E(n381), .Z(\arr[23] ) );
    VMW_AND2 U55 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U69 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_AO22 U109 ( .A(key[9]), .B(n373), .C(key[41]), .D(n374), .Z(n463) );
    VMW_INV U182 ( .A(n370), .Z(n369) );
    VMW_AND2 U72 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_AND2 U97 ( .A(\ScanReg[12] ), .B(n369), .Z(n387) );
    VMW_AO22 U140 ( .A(key[39]), .B(n373), .C(DataIn[7]), .D(n374), .Z(n433)
         );
    VMW_AO22 U167 ( .A(key[14]), .B(n373), .C(key[46]), .D(n374), .Z(n458) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD \key_reg[57]  ( .D(n415), .CP(Clk), .Q(key[57]) );
    VMW_FD \key_reg[47]  ( .D(n425), .CP(Clk), .Q(key[47]) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_AO22 U112 ( .A(key[6]), .B(n373), .C(key[38]), .D(n374), .Z(n466) );
    VMW_AO22 U135 ( .A(key[43]), .B(n373), .C(DataIn[11]), .D(n374), .Z(n429)
         );
    VMW_BUFIZ U205 ( .A(n399), .E(n381), .Z(\arr[17] ) );
    VMW_AND2 U60 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_BUFIZ U199 ( .A(n393), .E(n381), .Z(\arr[13] ) );
    VMW_AND2 U100 ( .A(\ScanReg[14] ), .B(n369), .Z(n384) );
    VMW_FD \key_reg[43]  ( .D(n429), .CP(Clk), .Q(key[43]) );
    VMW_AO22 U127 ( .A(key[50]), .B(n373), .C(DataIn[18]), .D(n374), .Z(n422)
         );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_AND2 U85 ( .A(\ScanReg[17] ), .B(n369), .Z(n399) );
    VMW_AO22 U149 ( .A(key[30]), .B(n373), .C(key[62]), .D(n374), .Z(n442) );
    VMW_AO22 U152 ( .A(key[28]), .B(n373), .C(key[60]), .D(n374), .Z(n444) );
    VMW_AND4 U175 ( .A(Addr[0]), .B(WR), .C(n367), .D(n375), .Z(n374) );
    VMW_AND4 U43 ( .A(WR), .B(Addr[1]), .C(n367), .D(n368), .Z(start) );
    VMW_AND2 U45 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U57 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AO22 U137 ( .A(key[41]), .B(n373), .C(DataIn[9]), .D(n374), .Z(n431)
         );
    VMW_BUFIZ U190 ( .A(n384), .E(n381), .Z(\arr[14] ) );
    VMW_FD \key_reg[60]  ( .D(n412), .CP(Clk), .Q(key[60]) );
    VMW_FD \key_reg[53]  ( .D(n419), .CP(Clk), .Q(key[53]) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_AND2 U70 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_BUFIZ U207 ( .A(n401), .E(n381), .Z(\arr[5] ) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AND2 U79 ( .A(\ScanReg[22] ), .B(n369), .Z(n405) );
    VMW_AND2 U95 ( .A(\ScanReg[31] ), .B(n369), .Z(n389) );
    VMW_AO22 U110 ( .A(key[8]), .B(n373), .C(key[40]), .D(n374), .Z(n464) );
    VMW_AO22 U159 ( .A(key[21]), .B(n373), .C(key[53]), .D(n374), .Z(n451) );
    VMW_FD \key_reg[42]  ( .D(n430), .CP(Clk), .Q(key[42]) );
    VMW_AO22 U119 ( .A(key[58]), .B(n373), .C(DataIn[26]), .D(n374), .Z(n414)
         );
    VMW_AO22 U142 ( .A(key[37]), .B(n373), .C(DataIn[5]), .D(n374), .Z(n435)
         );
    VMW_AO22 U165 ( .A(key[16]), .B(n373), .C(key[48]), .D(n374), .Z(n456) );
    VMW_INV U180 ( .A(Addr[0]), .Z(n368) );
    VMW_FD \key_reg[52]  ( .D(n420), .CP(Clk), .Q(key[52]) );
    VMW_BUFIZ U192 ( .A(n386), .E(n381), .Z(\arr[16] ) );
    VMW_FD \key_reg[61]  ( .D(n411), .CP(Clk), .Q(key[61]) );
    VMW_AND2 U87 ( .A(\ScanReg[3] ), .B(n369), .Z(n397) );
    VMW_AO22 U150 ( .A(key[2]), .B(n373), .C(key[34]), .D(n374), .Z(n470) );
    VMW_FD \key_reg[46]  ( .D(n426), .CP(Clk), .Q(key[46]) );
    VMW_XNOR2 U177 ( .A(Addr[2]), .B(ScanId), .Z(n372) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(key[52]), .B(n373), .C(DataIn[20]), .D(n374), .Z(n420)
         );
    VMW_FD \key_reg[56]  ( .D(n416), .CP(Clk), .Q(key[56]) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U50 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U59 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_AND2 U62 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_AND2 U65 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_AND2 U102 ( .A(\ScanReg[4] ), .B(n369), .Z(n382) );
    VMW_AND2 U105 ( .A(\ScanReg[23] ), .B(n369), .Z(n378) );
    VMW_BUFIZ U189 ( .A(n383), .E(n381), .Z(\arr[27] ) );
    VMW_AND2 U80 ( .A(\ScanReg[18] ), .B(n369), .Z(n404) );
    VMW_AO22 U122 ( .A(key[55]), .B(n373), .C(DataIn[23]), .D(n374), .Z(n417)
         );
    VMW_BUFIZ U212 ( .A(n406), .E(n381), .Z(\arr[11] ) );
    VMW_FD \key_reg[54]  ( .D(n418), .CP(Clk), .Q(key[54]) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_AO22 U139 ( .A(key[3]), .B(n373), .C(key[35]), .D(n374), .Z(n469) );
    VMW_AO22 U157 ( .A(key[23]), .B(n373), .C(key[55]), .D(n374), .Z(n449) );
    VMW_AO22 U170 ( .A(key[11]), .B(n373), .C(key[43]), .D(n374), .Z(n461) );
    VMW_FD \key_reg[44]  ( .D(n428), .CP(Clk), .Q(key[44]) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_BUFIZ U195 ( .A(n389), .E(n381), .Z(\arr[31] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AND2 U77 ( .A(\ScanReg[1] ), .B(n369), .Z(n407) );
    VMW_AND2 U89 ( .A(\ScanReg[29] ), .B(n369), .Z(n395) );
    VMW_BUFIZ U187 ( .A(n380), .E(n381), .Z(\arr[9] ) );
    VMW_BUFIZ U209 ( .A(n403), .E(n381), .Z(\arr[15] ) );
    VMW_FD \key_reg[63]  ( .D(n409), .CP(Clk), .Q(key[63]) );
    VMW_FD \key_reg[50]  ( .D(n422), .CP(Clk), .Q(key[50]) );
    VMW_FD \key_reg[49]  ( .D(n423), .CP(Clk), .Q(key[49]) );
    VMW_AND2 U92 ( .A(\ScanReg[2] ), .B(n369), .Z(n392) );
    VMW_AO22 U145 ( .A(key[34]), .B(n373), .C(DataIn[2]), .D(n374), .Z(n438)
         );
    VMW_AO22 U162 ( .A(key[19]), .B(n373), .C(key[51]), .D(n374), .Z(n453) );
    VMW_INV U179 ( .A(Addr[1]), .Z(n375) );
    VMW_AO22 U117 ( .A(key[5]), .B(n373), .C(key[37]), .D(n374), .Z(n467) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_BUFIZ U200 ( .A(n394), .E(n381), .Z(\arr[30] ) );
    VMW_AND2 U58 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AO22 U130 ( .A(key[48]), .B(n373), .C(DataIn[16]), .D(n374), .Z(n424)
         );
    VMW_FD \key_reg[59]  ( .D(n413), .CP(Clk), .Q(key[59]) );
    VMW_FD \key_reg[40]  ( .D(n432), .CP(Clk), .Q(key[40]) );
    VMW_AO22 U138 ( .A(key[40]), .B(n373), .C(DataIn[8]), .D(n374), .Z(n432)
         );
    VMW_BUFIZ U194 ( .A(n388), .E(n381), .Z(\arr[6] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_BUFIZ U208 ( .A(n402), .E(n381), .Z(\arr[26] ) );
    VMW_AND2 U64 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_AND2 U81 ( .A(\ScanReg[15] ), .B(n369), .Z(n403) );
    VMW_AO22 U156 ( .A(key[24]), .B(n373), .C(key[56]), .D(n374), .Z(n448) );
    VMW_AO22 U171 ( .A(key[10]), .B(n373), .C(key[42]), .D(n374), .Z(n462) );
    VMW_FD \key_reg[16]  ( .D(n456), .CP(Clk), .Q(key[16]) );
    VMW_FD \key_reg[25]  ( .D(n447), .CP(Clk), .Q(key[25]) );
    VMW_FD \key_reg[35]  ( .D(n437), .CP(Clk), .Q(key[35]) );
    VMW_FD \key_reg[4]  ( .D(n468), .CP(Clk), .Q(key[4]) );
    VMW_AND2 U104 ( .A(\ScanReg[10] ), .B(n369), .Z(n379) );
    VMW_AND2 U44 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U51 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_AND2 U76 ( .A(\ScanReg[8] ), .B(n369), .Z(n408) );
    VMW_AO22 U116 ( .A(key[60]), .B(n373), .C(DataIn[28]), .D(n374), .Z(n412)
         );
    VMW_AO22 U123 ( .A(key[54]), .B(n373), .C(DataIn[22]), .D(n374), .Z(n418)
         );
    VMW_BUFIZ U213 ( .A(n407), .E(n381), .Z(\arr[1] ) );
    VMW_FD \key_reg[0]  ( .D(n472), .CP(Clk), .Q(key[0]) );
    VMW_AND2 U56 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AND2 U88 ( .A(\ScanReg[20] ), .B(n369), .Z(n396) );
    VMW_AND2 U93 ( .A(\ScanReg[28] ), .B(n369), .Z(n391) );
    VMW_AO22 U131 ( .A(key[47]), .B(n373), .C(DataIn[15]), .D(n374), .Z(n425)
         );
    VMW_BUFIZ U201 ( .A(n395), .E(n381), .Z(\arr[29] ) );
    VMW_FD \key_reg[38]  ( .D(n434), .CP(Clk), .Q(key[38]) );
    VMW_FD \key_reg[12]  ( .D(n460), .CP(Clk), .Q(key[12]) );
    VMW_FD \key_reg[21]  ( .D(n451), .CP(Clk), .Q(key[21]) );
    VMW_INV U178 ( .A(n374), .Z(n373) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(\ScanReg[21] ), .B(n369), .Z(n390) );
    VMW_AO22 U143 ( .A(key[36]), .B(n373), .C(DataIn[4]), .D(n374), .Z(n436)
         );
    VMW_AO22 U144 ( .A(key[35]), .B(n373), .C(DataIn[3]), .D(n374), .Z(n437)
         );
    VMW_AO22 U163 ( .A(key[18]), .B(n373), .C(key[50]), .D(n374), .Z(n454) );
    VMW_INV U181 ( .A(n371), .Z(ScanEnable) );
    VMW_BUFIZ U186 ( .A(n379), .E(n381), .Z(\arr[10] ) );
    VMW_FD \key_reg[31]  ( .D(n441), .CP(Clk), .Q(key[31]) );
    VMW_FD \key_reg[9]  ( .D(n463), .CP(Clk), .Q(key[9]) );
    VMW_FD \key_reg[28]  ( .D(n444), .CP(Clk), .Q(key[28]) );
    VMW_FD \key_reg[33]  ( .D(n439), .CP(Clk), .Q(key[33]) );
    VMW_FD \key_reg[19]  ( .D(n453), .CP(Clk), .Q(key[19]) );
    VMW_AO22 U158 ( .A(key[22]), .B(n373), .C(key[54]), .D(n374), .Z(n450) );
    VMW_AO22 U164 ( .A(key[17]), .B(n373), .C(key[49]), .D(n374), .Z(n455) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_AO22 U136 ( .A(key[42]), .B(n373), .C(DataIn[10]), .D(n374), .Z(n430)
         );
    VMW_FD \key_reg[2]  ( .D(n470), .CP(Clk), .Q(key[2]) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_BUFIZ U206 ( .A(n400), .E(n381), .Z(\arr[7] ) );
    VMW_AND2 U71 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_FD \key_reg[10]  ( .D(n462), .CP(Clk), .Q(key[10]) );
    VMW_AO22 U111 ( .A(key[7]), .B(n373), .C(key[39]), .D(n374), .Z(n465) );
    VMW_AO22 U124 ( .A(key[53]), .B(n373), .C(DataIn[21]), .D(n374), .Z(n419)
         );
    VMW_FD \key_reg[23]  ( .D(n449), .CP(Clk), .Q(key[23]) );
    VMW_BUFIZ U214 ( .A(n408), .E(n381), .Z(\arr[8] ) );
    VMW_AND2 U63 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_AND2 U78 ( .A(\ScanReg[11] ), .B(n369), .Z(n406) );
    VMW_AND2 U86 ( .A(\ScanReg[24] ), .B(n369), .Z(n398) );
    VMW_AND2 U103 ( .A(\ScanReg[9] ), .B(n369), .Z(n380) );
    VMW_BUFIZ U188 ( .A(n382), .E(n381), .Z(\arr[4] ) );
    VMW_AO22 U118 ( .A(key[59]), .B(n373), .C(DataIn[27]), .D(n374), .Z(n413)
         );
    VMW_AO22 U151 ( .A(key[29]), .B(n373), .C(key[61]), .D(n374), .Z(n443) );
    VMW_FD \key_reg[37]  ( .D(n435), .CP(Clk), .Q(key[37]) );
    VMW_FD \key_reg[27]  ( .D(n445), .CP(Clk), .Q(key[27]) );
    VMW_FD \key_reg[14]  ( .D(n458), .CP(Clk), .Q(key[14]) );
    VMW_XNOR2 U176 ( .A(Addr[2]), .B(Id), .Z(n367) );
    VMW_BUFIZ U193 ( .A(n387), .E(n381), .Z(\arr[12] ) );
    VMW_FD \key_reg[6]  ( .D(n466), .CP(Clk), .Q(key[6]) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module DES_ECB_dummy1_DW01_inc_6_0 ( A, SUM );
input  [5:0] A;
output [5:0] SUM;
    wire \carry[4] , \carry[2] , \carry[3] , \carry[5] ;
    VMW_INV U3 ( .A(A[0]), .Z(SUM[0]) );
    VMW_HADD U1_1 ( .A(A[1]), .B(A[0]), .S(SUM[1]), .CO(\carry[2] ) );
    VMW_HADD U1_2 ( .A(A[2]), .B(\carry[2] ), .S(SUM[2]), .CO(\carry[3] ) );
    VMW_HADD U1_5 ( .A(A[5]), .B(\carry[5] ), .S(SUM[5]) );
    VMW_HADD U1_3 ( .A(A[3]), .B(\carry[3] ), .S(SUM[3]), .CO(\carry[4] ) );
    VMW_HADD U1_4 ( .A(A[4]), .B(\carry[4] ), .S(SUM[4]), .CO(\carry[5] ) );
endmodule


module DES_ECB_dummy1 ( Clk, Reset, Start, X, KEY, OUT, RDY );
input  [63:0] X;
input  [63:0] KEY;
output [63:0] OUT;
input  Clk, Reset, Start;
output RDY;
    wire \temp[63] , \temp[59] , \temp[54] , n13015, \temp[44] , \temp[2] , 
        n13928, n14268, n14479, n14158, n14373, n13032, n13129, n13147, n13160, 
        n13771, n13250, n13441, n14043, n13277, n13833, n14064, n13466, n13814, 
        n13984, n14354, n13219, n13389, n13756, n13408, n13598, n13738, n13292, 
        n13302, n13483, n13513, n13961, n14081, n14111, n13185, n13604, n13623, 
        n14221, n14430, n13794, n13029, n13325, n13534, n14206, n14396, n14417, 
        \arr12639[31] , \arr12639[28] , n13946, n14136, \arr12639[38] , n13085, 
        n13115, n13225, n13289, n13319, n13638, n13498, n13508, n13434, n13694, 
        n13846, n14036, \arr12639[12] , n13704, n13047, n13132, n13723, n14296, 
        \arr12639[21] , n14306, n14487, n13202, n13392, n14321, n13413, n13583, 
        n13656, n13828, n13861, n14011, n14181, \arr12639[3] , n14058, n14254, 
        n14368, n14445, n13350, n13377, n13566, n14164, n13884, n13914, n14143, 
        n13541, n13933, \temp[40] , \arr12639[35] , n13060, n14273, n14462, 
        n13671, n13055, n14246, n14457, n13072, n13342, n13365, \i[2] , n13644, 
        n13896, n14176, n13906, n13553, n13574, n13921, n14151, n13663, n14261, 
        n14470, n13097, n13169, n13259, n13448, n13237, n13426, n13778, n13854, 
        n13716, n14024, n13107, n13686, n13120, n14284, n14314, n14495, n14505, 
        n13731, n13210, n13873, n14333, n13280, n13380, n13591, n13401, 
        \temp[6] , n14003, n14193, n13968, n14088, n14118, n14228, n14439, 
        n13973, n13310, n13501, n13491, n13005, n13006, \arr12639[63] , n13007, 
        \temp[50] , \temp[49] , n13020, n13631, n14093, n14103, n14233, n14422, 
        n13786, \temp[61] , n13049, n13069, n13155, n13172, n13197, n13616, 
        n13337, n13954, n14214, n14384, n14405, n13526, n13868, n14018, n14124, 
        n14188, n14328, n14361, \arr12639[7] , n13242, n13763, n13821, n14051, 
        n13265, n13453, n13474, n13806, n14076, \arr12639[16] , n13996, n13744, 
        n14346, \arr12639[25] , n13678, n13152, n13359, n13548, \i6749[2] , 
        n13175, n13245, n13262, n13743, n14341, n13454, n13473, n13801, n13991, 
        n14071, n13764, n13826, n14056, \arr12639[14] , n13658, n14366, 
        \arr12639[27] , n13379, \i6749[0] , n13568, n14123, n13008, 
        \arr12639[61] , n13009, \temp[56] , \temp[52] , n13330, n13521, n13953, 
        \temp[42] , n13027, n13190, n14213, n14383, n14402, n13611, n13781, 
        n14234, n14425, n13127, n13217, n13287, n13317, n13496, n13636, n14094, 
        n14104, n13506, n13387, n13406, n13848, n13974, n14004, n14038, n14298, 
        n14308, \arr12639[5] , n14489, n14194, n13596, n13736, n13874, n14334, 
        n14283, n14313, n14502, n14492, \arr12639[37] , n13075, n13090, n13100, 
        n13681, n13230, n13711, n14023, n13421, \temp[4] , n13853, \i[0] , 
        n13948, n14208, n14398, n14419, n14138, n13664, n14266, n14477, n13040, 
        n13052, n13345, n13362, n13554, n13573, n13926, n14156, n13891, n13901, 
        n14171, n13643, n13067, n13149, n13279, n14241, n14450, n13468, 
        \temp[9] , n13758, \arr12639[1] , n13676, n13808, n14078, n13998, 
        n14348, n13357, n13546, n13934, n14274, n14465, n13370, n13883, n14144, 
        n13913, n13561, n14163, n13651, n14253, n14442, n13012, n13082, n13135, 
        n13199, n13788, n13205, n13339, n13618, \i6749[4] , n13528, n13584, 
        n13866, n14016, n14186, \arr12639[10] , n13395, n13414, n14326, 
        \arr12639[23] , n13724, n14291, n14301, n14480, n13099, n13112, n13703, 
        n13222, n13433, n13693, n13841, n14031, n13239, n13428, n13109, n13718, 
        n13322, n13688, n13941, n14131, n13533, n14201, n14391, n14410, n13013, 
        \arr12639[56] , \temp[46] , n13035, \arr12639[33] , n13182, n13793, 
        n13603, n13624, n14226, n14437, n13140, n13295, n13514, n13966, n14086, 
        n14116, \i[4] , \arr12639[19] , n13305, n13484, \temp[0] , n13898, 
        n14178, n14248, n14459, n13908, n13751, \arr12639[8] , n13167, n13257, 
        n13270, n13461, n13813, n14353, n13983, n13834, n14063, n13446, n14044, 
        n13776, n14267, n14374, n14476, \arr12639[46] , n13026, \temp[33] , 
        n13053, n13074, n13665, n13344, n13555, n14157, n13363, n13927, n14170, 
        n13572, n13890, n13900, n14240, n14451, n13091, n13126, n13148, n13278, 
        n13469, n13642, n13759, n13216, n13386, n13597, n13407, n13875, n14005, 
        n14195, n13710, n13737, n14335, n13101, n13680, n13191, n13231, n13420, 
        \temp[23] , n14282, n14312, n14493, n14503, n13331, \temp[10] , n13852, 
        n13949, n14022, n14139, n14209, n14399, n14418, \temp[19] , n13520, 
        n13952, n14122, n13610, n13780, n13637, n14212, n14382, n14403, n13153, 
        n13286, n14235, n14424, n13316, n13507, n13497, n13742, n13849, n13975, 
        n14039, n14095, n14105, n14299, n14309, n14488, n14340, n13244, n13263, 
        n13472, n14070, n13800, n13990, n14057, n13455, n13827, n13048, n13174, 
        n14367, n13765, n13098, n13108, n13141, n13378, n13659, \temp[27] , 
        n13569, n13899, n13909, n14249, n14458, n14179, n14352, n13166, n13256, 
        n13271, \temp[14] , n13750, n14062, n13812, n13982, n13447, n13460, 
        n13835, n14045, n13777, n14375, n13238, n13429, n13689, n13719, n13183, 
        n13323, n13532, n13940, n13602, n14130, n13792, \arr12639[52] , n13034, 
        n14200, n14390, n14411, n13625, n13294, n13304, n13967, n14227, n14436, 
        n13485, n13515, n14087, n14117, n13198, n13619, n13789, \arr12639[59] , 
        \arr12639[42] , n13134, n13204, n13338, n13529, n13394, n13867, n13415, 
        n13585, n13725, n14017, n14187, n14327, n13028, \temp[37] , n13066, 
        n13083, n13113, n13692, n13702, n13223, n13840, n14290, n14300, n14481, 
        n13432, n13809, n13999, n14030, n14079, n14275, n14349, n14464, n13356, 
        n13677, n13935, n14145, n13371, n13547, n13560, n13882, n13912, n14162, 
        n14252, n14443, \temp[35] , n13041, n13650, n13046, n13829, n14059, 
        n14369, n13061, n13351, n13376, n13657, n14255, n14444, n13540, n13567, 
        n13885, n13915, n14165, n13932, n14142, n13670, n13639, n14272, n14463, 
        n13224, n13288, n13509, n13318, n13499, n13435, n14037, n13847, n13014, 
        \arr12639[50] , \arr12639[40] , n13033, n13084, n14297, n14307, n14486, 
        n13114, n13705, n13128, n13133, n13695, n14320, n13203, n13582, n13722, 
        n14010, n14180, n13218, n13393, n13412, n13599, n13860, n13388, n13409, 
        n13293, n13739, n13512, n14080, n14110, n13303, n13482, n13622, n13960, 
        n14220, n14431, n14207, n14397, n14416, \arr12639[49] , n13184, n13795, 
        n13605, n13021, \arr12639[44] , n13146, n13161, n13324, n14137, n13535, 
        n13929, n13947, n14159, n14269, n14478, n13251, \temp[25] , n13770, 
        n14372, n13276, n13440, n13467, \temp[16] , n13832, n14042, n13757, 
        n13815, n13985, n14065, n13154, n13173, n13762, n14355, n13243, n13452, 
        n13820, n14360, n13264, n13807, n13997, n14050, n13475, n14077, n13745, 
        n14347, n13068, n13281, n13311, n13358, n13679, n13490, n13549, n13972, 
        n14092, n14102, n13500, \temp[28] , n14232, n14423, \temp[31] , n13196, 
        n13630, n14215, n14385, n14404, n13617, \temp[62] , \arr12639[62] , 
        \arr12639[58] , \arr12639[55] , \arr12639[54] , \temp[38] , n13096, 
        n13106, n13236, n13336, n13527, n13787, n13955, n14125, n13855, n13869, 
        n14019, n14025, n14189, n14329, n13427, n14504, n14285, n14315, n14494, 
        n13687, \temp[21] , n13717, n13054, n13121, n14332, n13730, n13211, 
        n13381, n13400, \temp[12] , n14002, n14192, n13872, n13590, n13645, 
        n13969, n14229, n14438, n14089, n14119, n13016, \arr12639[45] , n13073, 
        n13343, n13364, n13575, n13897, n13907, n14247, n14456, n13920, n14177, 
        n13552, n14150, n13168, n13258, n13449, n13662, n14260, n14471, n13779, 
        n13274, n13465, n13817, n14067, n13987, n13078, n13144, n13755, n14357, 
        n13163, n14370, n13253, n13772, n13830, n14040, n13442, n13669, n13348, 
        n13559, \temp[39] , n13031, n13186, n13797, n13291, n13326, n13607, 
        n13945, n14205, n14395, n14414, n13510, n13537, n13962, n14135, n13301, 
        n13480, n14082, n14112, n13620, n13131, \temp[29] , \temp[30] , n13879, 
        n14009, n14199, n14222, n14433, n14339, n13720, n14322, n13063, n13086, 
        n13201, \temp[20] , n13580, n13862, n13226, n13391, n13410, n13437, 
        \temp[13] , n13845, n14012, n14182, n14035, n13116, n13707, n13353, 
        n13542, n13697, n13930, n13979, n14099, n14109, n14239, n14295, n14305, 
        n14484, n14428, n14140, n13672, n14270, n14461, n14257, n14446, 
        \arr12639[41] , \temp[34] , n13044, n13178, n13248, n13374, n13655, 
        n13887, n14167, n13917, n13565, n13459, n13341, n13769, n13839, n14049, 
        n14152, n14379, n13550, n13922, n14262, n14473, n13038, n13056, n13071, 
        n13660, n13647, n14245, n14454, n13366, n13577, n14175, n13895, n13905, 
        n13094, n13104, n13123, n13298, n13308, n13489, n13629, n13519, n13732, 
        n13213, n13383, n13402, n14330, n13592, n13234, n13870, n14000, n14190, 
        n13425, n13857, n14027, n13685, n14506, n13715, n14287, n14317, n14496, 
        \arr12639[51] , \arr12639[48] , n13138, n13208, n13398, n13419, n13589, 
        n13729, n13194, n13615, n13785, n13334, n13525, n14217, n14387, n14406, 
        n13957, n14127, \temp[60] , \arr12639[60] , \arr12639[53] , n13023, 
        n13283, n13313, n13492, n13502, n13970, n14090, n14100, n13088, n13151, 
        n13156, n13266, n13632, n13939, n14230, n14421, n14279, n14468, n14075, 
        n14149, n13477, n13805, n13995, n14345, n13171, \temp[24] , n13747, 
        n14362, n13760, n13176, n13241, n13450, \temp[17] , n14052, n13246, 
        n13822, n13825, n13889, n14169, n14259, n14448, n13919, n13457, n14055, 
        n13740, n13767, n14365, n13228, n13261, n13470, \temp[26] , n14342, 
        n13802, n13992, n13439, \temp[15] , n14072, n13709, n13118, n13699, 
        n14237, n14426, n13024, n13635, n13011, \arr12639[57] , n13018, n13193, 
        n13284, n13977, n14097, n14107, n13314, n13505, n13333, n13495, n13950, 
        n14120, n13522, n13612, n13782, n14210, n14380, n14401, n13799, 
        \arr12639[43] , n13093, n13188, n13609, n13328, n13539, n13712, n14280, 
        n14310, n14491, n14501, n13103, n13682, n13214, n13233, n13422, n13850, 
        n14020, n13877, n14007, n14197, n13384, n13595, n13405, \temp[36] , 
        n13051, n13124, n14337, n13361, n13735, n13819, n14069, n13892, n13989, 
        n14359, n13902, n13570, n14172, n13640, n13043, n13076, n13667, n14242, 
        n14453, n13346, n13557, n13925, n14265, n14474, n13373, n13562, n14155, 
        n13652, n13880, n13910, n14160, n13064, n14250, n14441, n13675, n13036, 
        n13081, n13111, n13158, n13268, n13354, n14277, n14466, n13545, n13937, 
        n14147, n13479, \temp[22] , n13749, n13690, n14292, n14302, n14483, 
        n13700, n13136, n13206, n13221, \temp[11] , n14032, n13396, n13430, 
        n13842, n14015, n14185, n13417, n13587, n13727, n13865, n14325, n13959, 
        n14219, n14389, n14408, n14129, n14225, n14434, \temp[32] , n13296, 
        n13306, n13627, n14085, n14115, n13487, n13321, \temp[18] , n13517, 
        n13965, n13530, n14132, n13942, n14202, n14392, n14413, n13181, n13600, 
        n13790, \temp[57] , \arr12639[47] , n13164, n13254, n13445, n14508, 
        n13859, n14029, n14289, n14319, n14498, n13775, n13837, n14047, n14377, 
        n13058, n13143, n13273, n13752, n14350, n13462, n13649, n13810, n13980, 
        n14060, n13360, n13368, n13579, n13571, \temp[8] , n13818, n13988, 
        n14068, n14358, \arr12639[0] , n13893, n13903, n14173, n13019, n13050, 
        n13641, n14243, n14452, n13077, n14264, n14475, n13189, n13347, n13666, 
        n13924, n14154, n13556, n13608, \temp[47] , n13025, n13089, n13092, 
        n13102, n13329, n13538, n13798, \i6749[5] , n13683, n13119, n13125, 
        n13215, n13232, n13713, n13851, n14281, n14311, n14500, n14490, n13385, 
        n13404, n13423, n13876, n14021, n13594, n13734, n14006, n14196, 
        \arr12639[11] , n13229, n14336, \arr12639[22] , n13438, n13698, n13708, 
        \arr12639[32] , \i[5] , n13634, n14236, n14427, n13177, n13192, n13285, 
        n13315, n13494, n13976, n13504, n13332, n13523, n13951, n14096, 
        \arr12639[18] , n14106, n14121, n13247, n13456, \temp[1] , n13613, 
        n13783, n14211, n14381, n14400, n13824, n13888, n13918, n14258, 
        \arr12639[9] , n14449, n14054, n14168, n13766, n14364, n14343, n13037, 
        n13059, n13142, n13150, n13165, n13255, n13260, n13741, n13803, n13993, 
        n14073, n13471, n14046, \arr12639[15] , n13444, n13836, n14376, 
        \arr12639[26] , n13774, n14351, n13753, n13272, n13463, n14061, n13811, 
        n13981, n13369, \i6749[1] , n13648, n13578, n13626, n13297, n13516, 
        n14224, n14435, n13307, n13486, n13320, n13964, n14084, n14114, n13531, 
        n13943, n13010, n14133, \temp[58] , \temp[53] , n13180, n13791, n13601, 
        n14203, n14393, n14412, \temp[43] , n13080, n14509, n13858, n14028, 
        \arr12639[4] , n14288, n14318, n14499, n13110, n13701, n13691, 
        \arr12639[36] , n13042, n13137, n13207, n13220, n13431, n14293, n14303, 
        n14482, n13586, n13843, n14033, n13397, n13416, n13864, n14014, n14184, 
        n13372, \temp[5] , n13726, n13958, n14128, n14218, n14324, n14388, 
        n14409, n14161, n13563, n13881, n13911, n14251, n14440, n13653, 
        \arr12639[34] , n13045, n13062, n13065, \i[1] , n14276, n14467, n13674, 
        n13159, n13269, n13355, n13544, n14146, n13478, n13936, n13748, n13352, 
        n13931, n13543, n14141, n13673, n13654, n14271, n14460, \i[3] , n14256, 
        n14447, n13179, n13249, n13375, n13564, n13886, n13916, n13458, n14166, 
        n13768, n14323, n13017, \temp[41] , n13087, n13117, n13130, n13721, 
        n13200, n13390, n13863, n14013, n14183, n13411, n13227, n13581, n13844, 
        n14034, n13436, n13696, n14294, n14304, n14485, n13706, n13187, 
        \temp[7] , n13978, n14238, n14429, n14098, n14108, n13606, n14204, 
        n14394, n14415, n13796, n13327, n13536, n13944, n14134, n14083, n14113, 
        \temp[51] , n13290, n13300, n13963, n13481, n13511, \temp[48] , 
        \temp[45] , n13030, n14223, n14432, n13079, n13145, n13275, n13621, 
        n13816, n13878, \arr12639[6] , n13986, n14008, n14198, n14338, n13464, 
        n14066, \arr12639[17] , n13162, n13754, n13773, n14356, \arr12639[24] , 
        n13252, n13443, n13831, n14371, n14041, n13157, n13267, n13349, n13668, 
        \i6749[3] , n13558, n13476, \temp[3] , n13938, n14148, n14278, n14469, 
        n13746, n13804, n13994, n14074, n13170, n14344, n13761, n13139, n13209, 
        n13240, n14363, n13451, n13823, n14053, n13399, n13588, n13418, n13728, 
        n13784, n14216, n14386, n14407, \arr12639[30] , \arr12639[29] , 
        \temp[55] , n13022, n13195, n13614, n13282, n13335, n14126, n13524, 
        n13956, n14091, n14101, n13312, n13503, n13493, n13971, n14231, n14420, 
        n13633, \arr12639[39] , n13039, n13628, n13122, n13299, n13309, n13518, 
        n13488, n14331, n13212, n13733, n14001, n14191, n13235, n13382, n13593, 
        n13403, n13424, n13871, n14026, \arr12639[13] , n14507, n13856, n14316, 
        n14497, n14286, \arr12639[20] , n13070, n13095, n13714, n13105, n13684, 
        n13340, n13551, n13838, n14048, n14378, \arr12639[2] , n13661, n13923, 
        n14153, n14263, n14472, n13057, n13367, n13646, n14244, n14455, n13576, 
        n13894, n13904, n14174;
    VMW_AO21 U3925 ( .A(\temp[63] ), .B(n13005), .C(n13006), .Z(\arr12639[63] 
        ) );
    VMW_AO21 U3950 ( .A(\temp[38] ), .B(n13005), .C(n13031), .Z(\arr12639[38] 
        ) );
    VMW_AO22 U4120 ( .A(n13593), .B(n13594), .C(\temp[6] ), .D(n13370), .Z(
        n13396) );
    VMW_AND3 U4210 ( .A(n13688), .B(n13681), .C(n13478), .Z(n13104) );
    VMW_AOI211 U4968 ( .A(n13653), .B(n14367), .C(n13669), .D(n13932), .Z(
        n14366) );
    VMW_NAND3 U5068 ( .A(n13586), .B(n13606), .C(n13337), .Z(n13853) );
    VMW_INV U5358 ( .A(n13212), .Z(n13539) );
    VMW_AND2 U4380 ( .A(n13596), .B(n13440), .Z(n13902) );
    VMW_OR4 U4591 ( .A(n14148), .B(n14149), .C(n14146), .D(n14147), .Z(n13083)
         );
    VMW_AO21 U4401 ( .A(n13651), .B(n13932), .C(n13934), .Z(n13933) );
    VMW_OAI22 U4873 ( .A(n13643), .B(n14172), .C(n13642), .D(n14155), .Z(
        n14299) );
    VMW_AO22 U5264 ( .A(n14056), .B(n13451), .C(X[21]), .D(Start), .Z(n14488)
         );
    VMW_INV U5475 ( .A(n14366), .Z(n14458) );
    VMW_OAI22 U4731 ( .A(n13635), .B(n14163), .C(n13616), .D(n14164), .Z(
        n14233) );
    VMW_NOR4 U3977 ( .A(n13134), .B(n13135), .C(n13136), .D(n13137), .Z(n13133
        ) );
    VMW_AO22 U4097 ( .A(n13538), .B(n13539), .C(\temp[2] ), .D(n13212), .Z(
        n13537) );
    VMW_OAI22 U4716 ( .A(n13642), .B(n13714), .C(n13628), .D(n13713), .Z(
        n14226) );
    VMW_OAI21 U5154 ( .A(n13548), .B(n13780), .C(n13355), .Z(n13964) );
    VMW_AO22 U4107 ( .A(n13457), .B(n13563), .C(\temp[28] ), .D(n13261), .Z(
        n13562) );
    VMW_OAI22 U4686 ( .A(n13616), .B(n13618), .C(n13615), .D(n13644), .Z(
        n14211) );
    VMW_NOR4 U3989 ( .A(n13180), .B(n13181), .C(n13182), .D(n13183), .Z(n13179
        ) );
    VMW_NOR4 U3992 ( .A(n13195), .B(n13196), .C(n13197), .D(n13198), .Z(n13194
        ) );
    VMW_INV U4169 ( .A(KEY[46]), .Z(n13649) );
    VMW_INV U4237 ( .A(KEY[35]), .Z(n13725) );
    VMW_NAND2 U4426 ( .A(n13732), .B(n13493), .Z(n13986) );
    VMW_INV U5173 ( .A(n13453), .Z(n13659) );
    VMW_OAI22 U4854 ( .A(n13644), .B(n14159), .C(n13637), .D(n13717), .Z(
        n13307) );
    VMW_MUX2 U5243 ( .A(n14481), .B(\temp[28] ), .S(n13005), .Z(\arr12639[28] 
        ) );
    VMW_INV U5452 ( .A(n13898), .Z(n13911) );
    VMW_AOI211 U4259 ( .A(n13149), .B(n13736), .C(n13740), .D(n13741), .Z(
        n13739) );
    VMW_OAI22 U4778 ( .A(n13637), .B(n14103), .C(n13635), .D(n14112), .Z(
        n14254) );
    VMW_FD \OUT_reg[55]  ( .D(\arr12639[57] ), .CP(Clk), .Q(OUT[55]) );
    VMW_AO21 U4448 ( .A(n13530), .B(n13757), .C(n14009), .Z(n14008) );
    VMW_AO22 U5196 ( .A(n13578), .B(n13329), .C(n13322), .D(n13835), .Z(n14425
        ) );
    VMW_FD \temp_reg[59]  ( .D(\arr12639[59] ), .CP(Clk), .Q(\temp[59] ) );
    VMW_FD \temp_reg[40]  ( .D(\arr12639[40] ), .CP(Clk), .Q(\temp[40] ) );
    VMW_AND2 U4055 ( .A(\i6749[3] ), .B(n13445), .Z(n14506) );
    VMW_AO22 U4072 ( .A(n13479), .B(n13480), .C(\temp[19] ), .D(n13092), .Z(
        n13478) );
    VMW_OAI22 U4663 ( .A(n13626), .B(n14097), .C(n13624), .D(n14102), .Z(
        n14200) );
    VMW_AND3 U5006 ( .A(n13456), .B(n13659), .C(n13652), .Z(n14411) );
    VMW_NOR2 U4342 ( .A(n13329), .B(n13575), .Z(n13837) );
    VMW_OAI22 U4553 ( .A(n13626), .B(n14092), .C(n13624), .D(n14089), .Z(
        n13081) );
    VMW_INV U5336 ( .A(n13133), .Z(n13495) );
    VMW_OAI211 U4365 ( .A(n13749), .B(n13875), .C(n13876), .D(n13877), .Z(
        n13874) );
    VMW_OAI2222 U4921 ( .A(n13640), .B(n13718), .C(n13631), .D(n13721), .E(
        n13628), .F(n13720), .G(n13626), .H(n13719), .Z(n13392) );
    VMW_OAI22 U5281 ( .A(n14072), .B(n13804), .C(n13344), .D(n13569), .Z(
        n14497) );
    VMW_INV U5311 ( .A(n13266), .Z(n13566) );
    VMW_INV U5490 ( .A(n14474), .Z(n14427) );
    VMW_OR4 U4574 ( .A(n14138), .B(n14139), .C(n14136), .D(n14137), .Z(n13093)
         );
    VMW_AND2 U4896 ( .A(n13686), .B(n13680), .Z(n13866) );
    VMW_AO22 U4906 ( .A(n13353), .B(n13894), .C(n13424), .D(n13692), .Z(n13895
        ) );
    VMW_OAI21 U5021 ( .A(n13102), .B(n13894), .C(n13475), .Z(n14416) );
    VMW_AO22 U4069 ( .A(n13470), .B(n13464), .C(n13467), .D(n13471), .Z(n13070
        ) );
    VMW_AO21 U4359 ( .A(n13273), .B(n13863), .C(n13349), .Z(n13435) );
    VMW_OAI22 U4548 ( .A(n13620), .B(n13635), .C(n13618), .D(n13633), .Z(
        n14126) );
    VMW_OR4 U4644 ( .A(n14188), .B(n14189), .C(n14186), .D(n14187), .Z(n13129)
         );
    VMW_OAI22 U4678 ( .A(n13616), .B(n14096), .C(n13644), .D(n14097), .Z(
        n14207) );
    VMW_FD \temp_reg[50]  ( .D(\arr12639[50] ), .CP(Clk), .Q(\temp[50] ) );
    VMW_FD \temp_reg[49]  ( .D(\arr12639[49] ), .CP(Clk), .Q(\temp[49] ) );
    VMW_NAND5 U5121 ( .A(n13897), .B(n13401), .C(n13904), .D(n13396), .E(
        n13603), .Z(n14037) );
    VMW_FD \temp_reg[63]  ( .D(\arr12639[63] ), .CP(Clk), .Q(\temp[63] ) );
    VMW_FD \OUT_reg[45]  ( .D(\arr12639[50] ), .CP(Clk), .Q(OUT[45]) );
    VMW_AO21 U3926 ( .A(\temp[62] ), .B(n13005), .C(n13007), .Z(\arr12639[62] 
        ) );
    VMW_AO21 U3930 ( .A(\temp[58] ), .B(n13005), .C(n13011), .Z(\arr12639[58] 
        ) );
    VMW_AO21 U3937 ( .A(\temp[51] ), .B(n13005), .C(n13018), .Z(\arr12639[51] 
        ) );
    VMW_NOR4 U3959 ( .A(n13049), .B(n13050), .C(n13051), .D(n13052), .Z(n13048
        ) );
    VMW_NOR4 U4007 ( .A(n13267), .B(n13268), .C(n13269), .D(n13270), .Z(n13266
        ) );
    VMW_OR2 U4155 ( .A(n13629), .B(n13607), .Z(n13637) );
    VMW_OAI2222 U4744 ( .A(n13635), .B(n13715), .C(n13619), .D(n13714), .E(
        n13637), .F(n13713), .G(n13626), .H(n13712), .Z(n13234) );
    VMW_AND2 U4172 ( .A(n13453), .B(n13651), .Z(n13650) );
    VMW_INV U4242 ( .A(\temp[12] ), .Z(n13502) );
    VMW_INV U4265 ( .A(\temp[7] ), .Z(n13582) );
    VMW_AND2 U4474 ( .A(n13653), .B(n13664), .Z(n14049) );
    VMW_AO22 U5211 ( .A(n13107), .B(n13682), .C(n13680), .D(n13478), .Z(n14419
        ) );
    VMW_INV U5381 ( .A(KEY[43]), .Z(n14166) );
    VMW_INV U5400 ( .A(n13438), .Z(n13776) );
    VMW_OAI2222 U4806 ( .A(n13641), .B(n13645), .C(n13640), .D(n13648), .E(
        n13637), .F(n13647), .G(n13635), .H(n13646), .Z(n13248) );
    VMW_AO21 U4996 ( .A(n13068), .B(n13971), .C(n13659), .Z(n13672) );
    VMW_MUX2 U5236 ( .A(n14477), .B(\temp[30] ), .S(n13005), .Z(\arr12639[30] 
        ) );
    VMW_INV U5427 ( .A(n13730), .Z(n14359) );
    VMW_AO22 U4453 ( .A(n13684), .B(n13362), .C(n13691), .D(n13688), .Z(n13870
        ) );
    VMW_AOI211 U4821 ( .A(n13273), .B(n14277), .C(n13825), .D(n13286), .Z(
        n14276) );
    VMW_OAI211 U5096 ( .A(n14359), .B(n13875), .C(n14433), .D(n14432), .Z(
        n14396) );
    VMW_NAND3 U5106 ( .A(n13832), .B(n13321), .C(n13327), .Z(n14320) );
    VMW_AND2 U4337 ( .A(n13328), .B(n13320), .Z(n13833) );
    VMW_AO22 U4763 ( .A(X[4]), .B(n13774), .C(n13773), .D(\temp[23] ), .Z(
        n13014) );
    VMW_OR4 U4868 ( .A(n14296), .B(n14297), .C(n14294), .D(n14295), .Z(n13295)
         );
    VMW_OR4 U5168 ( .A(n13924), .B(n13950), .C(n13965), .D(n14390), .Z(n14081)
         );
    VMW_AO22 U5258 ( .A(n14050), .B(n13453), .C(n14049), .D(n13659), .Z(n13934
        ) );
    VMW_INV U5449 ( .A(n13864), .Z(n14440) );
    VMW_OAI2222 U4526 ( .A(n13621), .B(n13639), .C(n13619), .D(n13636), .E(
        n13616), .F(n13634), .G(n13632), .H(n13644), .Z(n13045) );
    VMW_OAI22 U4786 ( .A(n13624), .B(n14119), .C(n13643), .D(n14102), .Z(
        n14258) );
    VMW_OAI22 U4954 ( .A(n13628), .B(n13724), .C(n13626), .D(n13726), .Z(
        n13388) );
    VMW_INV U5343 ( .A(\temp[9] ), .Z(n13576) );
    DES_ECB_dummy1_DW01_inc_6_0 add_260 ( .A({\i[5] , \i[4] , \i[3] , \i[2] , 
        \i[1] , \i[0] }), .SUM({\i6749[5] , \i6749[4] , \i6749[3] , \i6749[2] , 
        \i6749[1] , \i6749[0] }) );
    VMW_FD \i_reg[3]  ( .D(n14506), .CP(Clk), .Q(\i[3] ) );
    VMW_NOR4 U4015 ( .A(n13300), .B(n13301), .C(n13302), .D(n13303), .Z(n13299
        ) );
    VMW_AND2 U4020 ( .A(n13324), .B(n13325), .Z(n13323) );
    VMW_NOR2 U4197 ( .A(n13353), .B(n13472), .Z(n13680) );
    VMW_OAI22 U4616 ( .A(n13641), .B(n14166), .C(n13631), .D(n14167), .Z(
        n14174) );
    VMW_OAI22 U4631 ( .A(n13637), .B(n14173), .C(n13631), .D(n14159), .Z(
        n13127) );
    VMW_OAI211 U5073 ( .A(n13319), .B(n13323), .C(n13328), .D(n13575), .Z(
        n13844) );
    VMW_AO21 U4185 ( .A(n13657), .B(n13662), .C(n13666), .Z(n13665) );
    VMW_AOI21 U4280 ( .A(n13339), .B(n13756), .C(n13770), .Z(n13769) );
    VMW_NAND3 U5054 ( .A(n13540), .B(n14401), .C(n13357), .Z(n13789) );
    VMW_OR2 U4310 ( .A(n13559), .B(n13557), .Z(n13806) );
    VMW_OR4 U4501 ( .A(n14087), .B(n14088), .C(n14084), .D(n14086), .Z(n13054)
         );
    VMW_AND2 U4325 ( .A(n13280), .B(n13808), .Z(n13815) );
    VMW_XNOR2 U4491 ( .A(\temp[46] ), .B(n13431), .Z(n14073) );
    VMW_OAI2222 U4534 ( .A(n13615), .B(n13628), .C(n13621), .D(n13645), .E(
        n13619), .F(n13648), .G(n13616), .H(n13647), .Z(n13060) );
    VMW_OAI22 U4946 ( .A(n13642), .B(n14161), .C(n13641), .D(n14159), .Z(
        n13378) );
    VMW_NAND2 U4973 ( .A(n13537), .B(n13239), .Z(n14375) );
    VMW_INV U5364 ( .A(KEY[29]), .Z(n14090) );
    VMW_OR4 U4604 ( .A(n14157), .B(n14158), .C(n14154), .D(n14156), .Z(n13134)
         );
    VMW_INV U5351 ( .A(\temp[5] ), .Z(n13599) );
    VMW_OAI22 U4794 ( .A(n13631), .B(n14097), .C(n13628), .D(n14102), .Z(
        n14262) );
    VMW_AND3 U4032 ( .A(n13351), .B(n13359), .C(n13360), .Z(n13358) );
    VMW_AO21 U5061 ( .A(n13564), .B(n13562), .C(n13809), .Z(n13288) );
    VMW_AND2 U4292 ( .A(n13437), .B(n13531), .Z(n13778) );
    VMW_AND2 U4302 ( .A(n13779), .B(n13421), .Z(n13787) );
    VMW_OAI22 U4623 ( .A(n13616), .B(n14160), .C(n13644), .D(n14161), .Z(
        n13112) );
    VMW_OAI21 U4961 ( .A(n13875), .B(n14359), .C(n13739), .Z(n13405) );
    VMW_AND3 U5046 ( .A(n13754), .B(n13514), .C(n13759), .Z(n13762) );
    VMW_OR2 U4483 ( .A(n13459), .B(n13470), .Z(n14061) );
    VMW_OAI22 U4513 ( .A(n13640), .B(n14094), .C(n14085), .D(n13624), .Z(
        n14100) );
    VMW_INV U5376 ( .A(KEY[19]), .Z(n14159) );
    VMW_FD \OUT_reg[51]  ( .D(\arr12639[41] ), .CP(Clk), .Q(OUT[51]) );
    VMW_FD \OUT_reg[48]  ( .D(\arr12639[1] ), .CP(Clk), .Q(OUT[48]) );
    VMW_OR2 U4129 ( .A(n13607), .B(n13608), .Z(n13609) );
    VMW_OAI22 U4738 ( .A(n13619), .B(n14173), .C(n13643), .D(n14159), .Z(
        n13226) );
    VMW_AND2 U4219 ( .A(n13688), .B(n13363), .Z(n13703) );
    VMW_AND2 U4389 ( .A(n13603), .B(n13907), .Z(n13909) );
    VMW_FD \temp_reg[44]  ( .D(\arr12639[44] ), .CP(Clk), .Q(\temp[44] ) );
    VMW_FD \OUT_reg[62]  ( .D(\arr12639[24] ), .CP(Clk), .Q(OUT[62]) );
    VMW_AO22 U4408 ( .A(n13398), .B(n13955), .C(n13956), .D(n13902), .Z(n13954
        ) );
    VMW_AO22 U4598 ( .A(n13685), .B(n13692), .C(n13680), .D(n13703), .Z(n14151
        ) );
    VMW_AO21 U3942 ( .A(\temp[46] ), .B(n13005), .C(n13023), .Z(\arr12639[46] 
        ) );
    VMW_AND3 U3980 ( .A(n13147), .B(n13148), .C(n13149), .Z(n13146) );
    VMW_NAND2 U4147 ( .A(\i[3] ), .B(\i[2] ), .Z(n13629) );
    VMW_AOI21 U5133 ( .A(n13456), .B(n14446), .C(n14412), .Z(n14362) );
    VMW_OR2 U4160 ( .A(n13617), .B(n13638), .Z(n13642) );
    VMW_AND2 U4250 ( .A(n13496), .B(n13729), .Z(n13140) );
    VMW_AOI21 U4277 ( .A(n13520), .B(n13204), .C(n13762), .Z(n13761) );
    VMW_AOI211 U4756 ( .A(n13787), .B(n13543), .C(n13788), .D(n14246), .Z(
        n13794) );
    VMW_OAI2222 U4814 ( .A(n13636), .B(n13644), .C(n13630), .D(n13641), .E(
        n13627), .F(n13640), .G(n13625), .H(n13637), .Z(n13243) );
    VMW_NAND4 U4984 ( .A(n14393), .B(n14036), .C(n14394), .D(n14395), .Z(
        n14392) );
    VMW_NAND2 U5203 ( .A(n13661), .B(n13655), .Z(n13973) );
    VMW_INV U5393 ( .A(n14479), .Z(n14397) );
    VMW_INV U5412 ( .A(n13661), .Z(n13677) );
    VMW_XOR2 U4441 ( .A(n14000), .B(\temp[36] ), .Z(n13999) );
    VMW_AND2 U4466 ( .A(n13410), .B(n13908), .Z(n14038) );
    VMW_OAI22 U4833 ( .A(n13619), .B(n13727), .C(n13609), .D(n14167), .Z(
        n14279) );
    VMW_MUX2 U5224 ( .A(n14471), .B(\temp[5] ), .S(n13005), .Z(\arr12639[5] )
         );
    VMW_INV U5435 ( .A(n13786), .Z(n13792) );
    VMW_OAI22 U4771 ( .A(n13620), .B(n13624), .C(n13618), .D(n13621), .Z(
        n14251) );
    VMW_OAI211 U5084 ( .A(n13344), .B(n13346), .C(n13569), .D(n13564), .Z(
        n14429) );
    VMW_NAND2 U5114 ( .A(n13693), .B(n13351), .Z(n14325) );
    VMW_OR4 U4928 ( .A(n14338), .B(n14339), .C(n14336), .D(n14337), .Z(n13371)
         );
    VMW_AO22 U5028 ( .A(n13352), .B(n13353), .C(n13478), .D(n13691), .Z(n14406
        ) );
    VMW_MUX2 U5288 ( .A(n14500), .B(\temp[12] ), .S(n13005), .Z(\arr12639[12] 
        ) );
    VMW_INV U5318 ( .A(n13077), .Z(n13483) );
    VMW_AND3 U5014 ( .A(n13467), .B(n13653), .C(n13071), .Z(n13666) );
    VMW_AO21 U4047 ( .A(n13421), .B(n13357), .C(n13422), .Z(n13420) );
    VMW_AND2 U4060 ( .A(n13401), .B(n13409), .Z(n13448) );
    VMW_INV U5184 ( .A(n13512), .Z(n13516) );
    VMW_AND2 U4350 ( .A(n13329), .B(n13606), .Z(n13842) );
    VMW_OAI22 U4671 ( .A(n13644), .B(n13648), .C(n13635), .D(n14096), .Z(
        n14204) );
    VMW_OAI22 U4933 ( .A(n13635), .B(n14166), .C(n13624), .D(n14167), .Z(
        n14341) );
    VMW_INV U5324 ( .A(n13169), .Z(n13508) );
    VMW_AND2 U4377 ( .A(n13899), .B(n13401), .Z(n13898) );
    VMW_OR4 U4541 ( .A(n14117), .B(n14118), .C(n14115), .D(n14116), .Z(n13049)
         );
    VMW_OR4 U4566 ( .A(n14134), .B(n14135), .C(n14132), .D(n14133), .Z(n13088)
         );
    VMW_AO22 U4884 ( .A(X[16]), .B(n13774), .C(\temp[5] ), .D(n13773), .Z(
        n13032) );
    VMW_OAI22 U4914 ( .A(n13616), .B(n13717), .C(n13644), .D(n13723), .Z(
        n13368) );
    VMW_AO22 U5293 ( .A(n14082), .B(n13451), .C(X[57]), .D(Start), .Z(n14503)
         );
    VMW_INV U5303 ( .A(n13058), .Z(n13469) );
    VMW_INV U5482 ( .A(n14152), .Z(n14421) );
    VMW_OAI22 U4656 ( .A(n13644), .B(n14119), .C(n13641), .D(n14096), .Z(
        n14197) );
    VMW_OAI211 U5033 ( .A(n13155), .B(n13147), .C(n13144), .D(n13731), .Z(
        n13745) );
    VMW_NAND2 U4132 ( .A(\i[2] ), .B(n13614), .Z(n13613) );
    VMW_AO21 U4202 ( .A(n13472), .B(n13475), .C(n13364), .Z(n13107) );
    VMW_AND2 U4392 ( .A(n13603), .B(n13903), .Z(n13913) );
    VMW_AO22 U4828 ( .A(X[34]), .B(n13774), .C(n13773), .D(\temp[11] ), .Z(
        n13026) );
    VMW_OAI2222 U4861 ( .A(n13644), .B(n13715), .C(n13633), .D(n13714), .E(
        n13616), .F(n13713), .G(n13640), .H(n13712), .Z(n13291) );
    VMW_AND3 U5128 ( .A(n13459), .B(n13456), .C(n13653), .Z(n14444) );
    VMW_AO22 U5218 ( .A(n13991), .B(n13451), .C(X[9]), .D(Start), .Z(n14470)
         );
    VMW_INV U5388 ( .A(n13069), .Z(n13654) );
    VMW_INV U5409 ( .A(n13602), .Z(n13397) );
    VMW_NOR3 U4413 ( .A(Start), .B(Reset), .C(n13452), .Z(n13445) );
    VMW_OAI2222 U4583 ( .A(n13616), .B(n13627), .C(n13625), .D(n13644), .E(
        n13637), .F(n13649), .G(n13631), .H(n13645), .Z(n13074) );
    VMW_OAI22 U4723 ( .A(n13628), .B(n14170), .C(n13626), .D(n14166), .Z(
        n14229) );
    VMW_MUX2 U5276 ( .A(n14494), .B(\temp[17] ), .S(n13005), .Z(\arr12639[17] 
        ) );
    VMW_INV U5467 ( .A(n13984), .Z(n13743) );
    VMW_NAND3 U5146 ( .A(n14048), .B(n13662), .C(n13668), .Z(n13959) );
    VMW_AO21 U3945 ( .A(\temp[43] ), .B(n13005), .C(n13026), .Z(\arr12639[43] 
        ) );
    VMW_NOR4 U3962 ( .A(n13064), .B(n13065), .C(n13066), .D(n13067), .Z(n13063
        ) );
    VMW_NOR4 U3965 ( .A(n13078), .B(n13079), .C(n13080), .D(n13081), .Z(n13077
        ) );
    VMW_AO22 U4085 ( .A(n13510), .B(n13511), .C(\temp[18] ), .D(n13179), .Z(
        n13509) );
    VMW_AO22 U4115 ( .A(n13582), .B(n13583), .C(\temp[7] ), .D(n13314), .Z(
        n13581) );
    VMW_OAI22 U4694 ( .A(n13618), .B(n13637), .C(n13615), .D(n13635), .Z(
        n14215) );
    VMW_AO22 U4704 ( .A(X[14]), .B(n13774), .C(n13773), .D(\temp[30] ), .Z(
        n13007) );
    VMW_NAND3 U5161 ( .A(n13837), .B(n13322), .C(n13572), .Z(n14459) );
    VMW_AND3 U4029 ( .A(n13287), .B(n13288), .C(n13282), .Z(n13349) );
    VMW_INV U4225 ( .A(KEY[18]), .Z(n13714) );
    VMW_OAI22 U4846 ( .A(n13628), .B(n14159), .C(n13626), .D(n13725), .Z(
        n13302) );
    VMW_INV U4289 ( .A(\temp[3] ), .Z(n13544) );
    VMW_OR2 U4319 ( .A(n13569), .B(n13810), .Z(n13285) );
    VMW_XOR2 U4434 ( .A(n13992), .B(\temp[38] ), .Z(n13991) );
    VMW_AO22 U5251 ( .A(n14039), .B(n13444), .C(n14038), .D(n13897), .Z(n13915
        ) );
    VMW_INV U5440 ( .A(n13811), .Z(n14274) );
    VMW_FD \temp_reg[54]  ( .D(\arr12639[54] ), .CP(Clk), .Q(\temp[54] ) );
    VMW_OAI22 U4498 ( .A(n13620), .B(n13621), .C(n13618), .D(n13619), .Z(
        n14086) );
    VMW_OAI22 U4508 ( .A(n13620), .B(n13626), .C(n13618), .D(n13624), .Z(
        n14099) );
    VMW_FD \OUT_reg[58]  ( .D(\arr12639[8] ), .CP(Clk), .Q(OUT[58]) );
    VMW_FD \OUT_reg[41]  ( .D(\arr12639[34] ), .CP(Clk), .Q(OUT[41]) );
    VMW_INV U4222 ( .A(\temp[8] ), .Z(n13573) );
    VMW_AND2 U4433 ( .A(n13525), .B(n13202), .Z(n13529) );
    VMW_OAI22 U4638 ( .A(n13637), .B(n14159), .C(n13635), .D(n13725), .Z(
        n13116) );
    VMW_MUX2 U5256 ( .A(n14485), .B(\temp[24] ), .S(n13005), .Z(\arr12639[24] 
        ) );
    VMW_INV U5447 ( .A(n13327), .Z(n13883) );
    VMW_OAI22 U4841 ( .A(n13609), .B(n14169), .C(n13644), .D(n14167), .Z(
        n14283) );
    VMW_AO22 U5166 ( .A(n13906), .B(n13396), .C(n13409), .D(n13900), .Z(n13966
        ) );
    VMW_AO22 U4082 ( .A(n13497), .B(n13504), .C(\temp[15] ), .D(n13194), .Z(
        n13200) );
    VMW_AO22 U4112 ( .A(n13573), .B(n13574), .C(\temp[8] ), .D(n13304), .Z(
        n13572) );
    VMW_AO22 U4703 ( .A(X[6]), .B(n13774), .C(n13773), .D(\temp[31] ), .Z(
        n13006) );
    VMW_OAI22 U4693 ( .A(n13609), .B(n14094), .C(n14085), .D(n13644), .Z(
        n14214) );
    VMW_NOR5 U5141 ( .A(n14302), .B(n14450), .C(n13855), .D(n14451), .E(n13886
        ), .Z(n14057) );
    VMW_NOR4 U3987 ( .A(n13170), .B(n13171), .C(n13172), .D(n13173), .Z(n13169
        ) );
    VMW_AOI211 U4009 ( .A(n13276), .B(n13277), .C(n13278), .D(n13271), .Z(
        n13275) );
    VMW_OR2 U4135 ( .A(n13612), .B(\i[1] ), .Z(n13617) );
    VMW_AND2 U4205 ( .A(n13683), .B(n13478), .Z(n13359) );
    VMW_OAI22 U4584 ( .A(n13609), .B(n14090), .C(n13619), .D(n13630), .Z(
        n13075) );
    VMW_OAI22 U4724 ( .A(n13641), .B(n14155), .C(n13631), .D(n14169), .Z(
        n14230) );
    VMW_AO22 U5271 ( .A(n14064), .B(n13451), .C(X[37]), .D(Start), .Z(n14492)
         );
    VMW_INV U5460 ( .A(n13944), .Z(n14449) );
    VMW_AND2 U4339 ( .A(n13584), .B(n13320), .Z(n13337) );
    VMW_AOI21 U4395 ( .A(n13901), .B(n13400), .C(n13917), .Z(n13916) );
    VMW_AO22 U4414 ( .A(n13969), .B(n13456), .C(n13970), .D(n13651), .Z(n13968
        ) );
    VMW_OAI22 U4866 ( .A(n13637), .B(n14169), .C(n13635), .D(n14170), .Z(
        n14296) );
    VMW_OAI22 U4528 ( .A(n13609), .B(n14091), .C(n13628), .D(n14092), .Z(
        n13047) );
    VMW_FD \temp_reg[56]  ( .D(\arr12639[56] ), .CP(Clk), .Q(\temp[56] ) );
    VMW_NAND3 U4040 ( .A(n13396), .B(n13397), .C(n13398), .Z(n13395) );
    VMW_AND2 U4199 ( .A(n13472), .B(n13481), .Z(n13683) );
    VMW_OAI22 U4788 ( .A(n13640), .B(n13649), .C(n13631), .D(n13648), .Z(
        n14260) );
    VMW_OAI22 U4618 ( .A(n13626), .B(n14172), .C(n13624), .D(n14155), .Z(
        n14176) );
    VMW_FD \OUT_reg[43]  ( .D(\arr12639[42] ), .CP(Clk), .Q(OUT[43]) );
    VMW_AO22 U4067 ( .A(n13465), .B(n13466), .C(\temp[0] ), .D(n13043), .Z(
        n13464) );
    VMW_AND2 U4357 ( .A(n13807), .B(n13277), .Z(n13346) );
    VMW_NAND3 U4370 ( .A(n13421), .B(n13356), .C(n13238), .Z(n13888) );
    VMW_AND2 U4651 ( .A(n13496), .B(n13488), .Z(n13751) );
    VMW_AND3 U5034 ( .A(n13447), .B(n13152), .C(n13163), .Z(n13740) );
    VMW_OAI22 U4546 ( .A(n13643), .B(n14119), .C(n13631), .D(n14112), .Z(
        n14124) );
    VMW_OAI22 U4561 ( .A(n13640), .B(n14092), .C(n13637), .D(n14089), .Z(
        n13101) );
    VMW_AO22 U4883 ( .A(X[8]), .B(n13774), .C(n13773), .D(\temp[6] ), .Z(
        n13031) );
    VMW_OAI2222 U4913 ( .A(n13635), .B(n13716), .C(n13619), .D(n13715), .E(
        n13637), .F(n13714), .G(n13621), .H(n13713), .Z(n13367) );
    VMW_MUX2 U5294 ( .A(n14503), .B(\temp[0] ), .S(n13005), .Z(\arr12639[0] )
         );
    VMW_INV U5304 ( .A(\temp[29] ), .Z(n13454) );
    VMW_INV U5485 ( .A(n14416), .Z(n13710) );
    VMW_OAI22 U4676 ( .A(n13621), .B(n14091), .C(n13639), .D(n13643), .Z(
        n13173) );
    VMW_OAI22 U4934 ( .A(n13640), .B(n14169), .C(n13637), .D(n14170), .Z(
        n14342) );
    VMW_INV U5323 ( .A(n13092), .Z(n13480) );
    VMW_FD \i_reg[5]  ( .D(n14504), .CP(Clk), .Q(\i[5] ) );
    VMW_NAND2 U4140 ( .A(\i[0] ), .B(\i[1] ), .Z(n13622) );
    VMW_INV U4167 ( .A(KEY[53]), .Z(n13647) );
    VMW_OAI22 U4808 ( .A(n13643), .B(n14091), .C(n13631), .D(n13632), .Z(
        n13250) );
    VMW_NAND3 U5013 ( .A(n13453), .B(n13656), .C(n13657), .Z(n13678) );
    VMW_INV U5183 ( .A(n13200), .Z(n13760) );
    VMW_OAI21 U4998 ( .A(n14404), .B(n14405), .C(n13351), .Z(n14381) );
    VMW_NAND2 U5098 ( .A(n13873), .B(n14190), .Z(n14434) );
    VMW_NOR2 U5108 ( .A(n13888), .B(n13550), .Z(n13892) );
    VMW_MUX2 U5238 ( .A(n14478), .B(\temp[2] ), .S(n13005), .Z(\arr12639[2] )
         );
    VMW_INV U5429 ( .A(n13589), .Z(n13555) );
    VMW_AND2 U4257 ( .A(n13143), .B(n13161), .Z(n13736) );
    VMW_OAI22 U4776 ( .A(n13616), .B(n14091), .C(n14089), .D(n13643), .Z(
        n13265) );
    VMW_NAND3 U5083 ( .A(n13272), .B(n13288), .C(n13412), .Z(n14428) );
    VMW_NAND3 U5113 ( .A(n13686), .B(n13107), .C(n13690), .Z(n14326) );
    VMW_AND2 U4270 ( .A(n13507), .B(n13200), .Z(n13756) );
    VMW_XOR2 U4446 ( .A(n14006), .B(\temp[35] ), .Z(n14005) );
    VMW_XOR2 U4461 ( .A(n14028), .B(\temp[59] ), .Z(n14027) );
    VMW_OAI22 U4834 ( .A(n13624), .B(n13720), .C(n13621), .D(n13719), .Z(
        n14280) );
    VMW_AO22 U5223 ( .A(n13997), .B(n13451), .C(X[17]), .D(Start), .Z(n14471)
         );
    VMW_INV U5432 ( .A(n13779), .Z(n14377) );
    VMW_OR4 U4751 ( .A(n14243), .B(n14244), .C(n14241), .D(n14242), .Z(n13208)
         );
    VMW_OR4 U4813 ( .A(n14271), .B(n14272), .C(n14269), .D(n14270), .Z(n13242)
         );
    VMW_OAI211 U4983 ( .A(n13911), .B(n13921), .C(n14391), .D(n13916), .Z(
        n14390) );
    VMW_NAND2 U5204 ( .A(n13653), .B(n13663), .Z(n13972) );
    VMW_INV U5394 ( .A(n13139), .Z(n13156) );
    VMW_INV U5415 ( .A(n13684), .Z(n14153) );
    VMW_AO21 U3931 ( .A(\temp[57] ), .B(n13005), .C(n13012), .Z(\arr12639[57] 
        ) );
    VMW_AO21 U3939 ( .A(\temp[49] ), .B(n13005), .C(n13020), .Z(\arr12639[49] 
        ) );
    VMW_AOI211 U3979 ( .A(n13143), .B(n13144), .C(n13145), .D(n13138), .Z(
        n13142) );
    VMW_AND3 U4012 ( .A(n13287), .B(n13288), .C(n13272), .Z(n13286) );
    VMW_NOR4 U4035 ( .A(n13371), .B(n13372), .C(n13373), .D(n13374), .Z(n13370
        ) );
    VMW_AND2 U4295 ( .A(n13543), .B(n13540), .Z(n13781) );
    VMW_OAI22 U4514 ( .A(n13616), .B(n14102), .C(n13644), .D(n14103), .Z(
        n14101) );
    VMW_AOI211 U4898 ( .A(n13684), .B(n13104), .C(n13700), .D(n13864), .Z(
        n14311) );
    VMW_AND2 U5008 ( .A(n13151), .B(n13141), .Z(n13159) );
    VMW_OR3 U5134 ( .A(n13940), .B(n13935), .C(n14361), .Z(n14052) );
    VMW_INV U5198 ( .A(n13440), .Z(n13603) );
    VMW_INV U5338 ( .A(n13309), .Z(n13571) );
    VMW_OAI22 U4908 ( .A(n13643), .B(n14167), .C(n13631), .D(n14164), .Z(
        n14328) );
    VMW_INV U5371 ( .A(KEY[5]), .Z(n14094) );
    VMW_OR2 U4305 ( .A(n13796), .B(n13797), .Z(n13795) );
    VMW_XOR2 U4484 ( .A(n14063), .B(\temp[33] ), .Z(n14062) );
    VMW_OAI22 U4624 ( .A(n13619), .B(n14163), .C(n13635), .D(n14164), .Z(
        n14178) );
    VMW_AOI211 U4966 ( .A(n13913), .B(n13901), .C(n14365), .D(n13407), .Z(
        n14364) );
    VMW_AND3 U5041 ( .A(n13755), .B(n13514), .C(n13205), .Z(n13772) );
    VMW_OR4 U5066 ( .A(n13417), .B(n13434), .C(n13829), .D(n14424), .Z(n14000)
         );
    VMW_AO22 U4099 ( .A(n13544), .B(n13545), .C(\temp[3] ), .D(n13207), .Z(
        n13543) );
    VMW_OR2 U4182 ( .A(n13663), .B(n13652), .Z(n13660) );
    VMW_OAI22 U4793 ( .A(n13626), .B(n14103), .C(n13624), .D(n14112), .Z(
        n14261) );
    VMW_AND2 U4322 ( .A(n13280), .B(n13812), .Z(n13276) );
    VMW_OAI22 U4603 ( .A(n13635), .B(n13721), .C(n13633), .D(n13720), .Z(
        n14158) );
    VMW_INV U5356 ( .A(n13380), .Z(n13595) );
    VMW_OR4 U4533 ( .A(n14113), .B(n14114), .C(n14110), .D(n14111), .Z(n13059)
         );
    VMW_OAI22 U4941 ( .A(n13621), .B(n13720), .C(n13619), .D(n13719), .Z(
        n14345) );
    VMW_AO22 U4109 ( .A(n13460), .B(n13568), .C(\temp[27] ), .D(n13246), .Z(
        n13567) );
    VMW_OAI22 U4718 ( .A(n13616), .B(n13721), .C(n13644), .D(n13720), .Z(
        n14228) );
    VMW_OAI22 U4688 ( .A(n13626), .B(n13627), .C(n13624), .D(n13625), .Z(
        n14213) );
    VMW_NOR4 U4000 ( .A(n13233), .B(n13234), .C(n13235), .D(n13236), .Z(n13232
        ) );
    VMW_AND3 U4027 ( .A(n13273), .B(n13280), .C(n13344), .Z(n13343) );
    VMW_INV U4239 ( .A(\temp[15] ), .Z(n13497) );
    VMW_AND2 U4428 ( .A(n13525), .B(n13342), .Z(n13521) );
    VMW_FD \OUT_reg[53]  ( .D(\arr12639[49] ), .CP(Clk), .Q(OUT[53]) );
    VMW_OR2 U4287 ( .A(n13535), .B(n13777), .Z(n13589) );
    VMW_NOR2 U4317 ( .A(n13562), .B(n13808), .Z(n13274) );
    VMW_XOR2 U4496 ( .A(n14083), .B(\temp[32] ), .Z(n14082) );
    VMW_OAI22 U4848 ( .A(n13643), .B(n14170), .C(n13642), .D(n14166), .Z(
        n14286) );
    VMW_AO21 U5148 ( .A(n13650), .B(n13663), .C(n14411), .Z(n14367) );
    VMW_MUX2 U5278 ( .A(n14495), .B(\temp[16] ), .S(n13005), .Z(\arr12639[16] 
        ) );
    VMW_INV U5469 ( .A(n14042), .Z(n13925) );
    VMW_FD \temp_reg[46]  ( .D(\arr12639[46] ), .CP(Clk), .Q(\temp[46] ) );
    VMW_FD \OUT_reg[60]  ( .D(\arr12639[16] ), .CP(Clk), .Q(OUT[60]) );
    VMW_OR2 U4974 ( .A(n13537), .B(n13589), .Z(n13963) );
    VMW_INV U5363 ( .A(KEY[13]), .Z(n14089) );
    VMW_FD \i_reg[1]  ( .D(n14508), .CP(Clk), .Q(\i[1] ) );
    VMW_OAI22 U4506 ( .A(n13633), .B(n14096), .C(n13609), .D(n14097), .Z(
        n14095) );
    VMW_NAND3 U5053 ( .A(n13543), .B(n13551), .C(n13238), .Z(n13790) );
    VMW_OAI211 U4190 ( .A(n13658), .B(n13677), .C(n13678), .D(n13679), .Z(
        n13676) );
    VMW_OR4 U4636 ( .A(n14184), .B(n14185), .C(n14182), .D(n14183), .Z(n13114)
         );
    VMW_NAND4 U5074 ( .A(n14425), .B(n13572), .C(n13320), .D(n13606), .Z(
        n14426) );
    VMW_OAI22 U4611 ( .A(n13621), .B(n14172), .C(n13619), .D(n14155), .Z(
        n14171) );
    VMW_AND4 U4049 ( .A(n13427), .B(n13428), .C(n13429), .D(n13430), .Z(n13426
        ) );
    VMW_AO22 U4330 ( .A(n13272), .B(n13819), .C(n13809), .D(n13820), .Z(n13432
        ) );
    VMW_OAI22 U4521 ( .A(n13615), .B(n13633), .C(n13631), .D(n13649), .Z(
        n14106) );
    VMW_OR4 U4781 ( .A(n14255), .B(n14256), .C(n14253), .D(n14254), .Z(n13267)
         );
    VMW_OAI2222 U4953 ( .A(n13624), .B(n13718), .C(n13643), .D(n13720), .E(
        n13642), .F(n13719), .G(n13641), .H(n13727), .Z(n13387) );
    VMW_INV U5344 ( .A(n13299), .Z(n13577) );
    VMW_AND2 U4379 ( .A(n13900), .B(n13444), .Z(n13901) );
    VMW_OAI22 U4568 ( .A(n13628), .B(n13632), .C(n13615), .D(n13643), .Z(
        n13090) );
    VMW_FD \temp_reg[52]  ( .D(\arr12639[52] ), .CP(Clk), .Q(\temp[52] ) );
    VMW_OAI2222 U4658 ( .A(n13624), .B(n13645), .C(n13621), .D(n13648), .E(
        n13619), .F(n13647), .G(n13616), .H(n13646), .Z(n13191) );
    VMW_FD \temp_reg[61]  ( .D(\arr12639[61] ), .CP(Clk), .Q(\temp[61] ) );
    VMW_FD \OUT_reg[47]  ( .D(\arr12639[58] ), .CP(Clk), .Q(OUT[47]) );
    VMW_INV U4152 ( .A(KEY[12]), .Z(n13634) );
    VMW_AND2 U4175 ( .A(n13459), .B(n13470), .Z(n13655) );
    VMW_AO22 U4764 ( .A(X[12]), .B(n13774), .C(n13773), .D(\temp[22] ), .Z(
        n13015) );
    VMW_AND2 U4245 ( .A(n13148), .B(n13157), .Z(n13730) );
    VMW_XOR2 U4454 ( .A(n14018), .B(\temp[34] ), .Z(n14017) );
    VMW_AO22 U4826 ( .A(X[18]), .B(n13774), .C(n13773), .D(\temp[13] ), .Z(
        n13024) );
    VMW_NAND4 U5091 ( .A(n13427), .B(n13709), .C(n13869), .D(n14312), .Z(
        n14018) );
    VMW_NAND3 U5101 ( .A(n13320), .B(n13322), .C(n13842), .Z(n14436) );
    VMW_OAI22 U4262 ( .A(n13153), .B(n13161), .C(n13749), .D(n13735), .Z(
        n13166) );
    VMW_OAI22 U4801 ( .A(n13642), .B(n14094), .C(n14085), .D(n13628), .Z(
        n14265) );
    VMW_AO21 U4991 ( .A(n13395), .B(n14031), .C(n13904), .Z(n14357) );
    VMW_AO22 U5231 ( .A(n14007), .B(n13200), .C(n14008), .D(n13760), .Z(n14474
        ) );
    VMW_INV U5420 ( .A(n13700), .Z(n13708) );
    VMW_OR2 U4473 ( .A(n14048), .B(n13659), .Z(n14047) );
    VMW_MUX2 U5216 ( .A(n14468), .B(\temp[7] ), .S(n13005), .Z(\arr12639[7] )
         );
    VMW_INV U5386 ( .A(n13345), .Z(n13960) );
    VMW_INV U5407 ( .A(n13396), .Z(n13899) );
    VMW_OR4 U4743 ( .A(n14239), .B(n14240), .C(n14237), .D(n14238), .Z(n13233)
         );
    VMW_NOR4 U5126 ( .A(n14443), .B(n13148), .C(n13139), .D(n13447), .Z(n13929
        ) );
    VMW_FD \OUT_reg[57]  ( .D(\arr12639[32] ), .CP(Clk), .Q(OUT[57]) );
    VMW_NOR4 U3957 ( .A(n13039), .B(n13040), .C(n13041), .D(n13042), .Z(n13038
        ) );
    VMW_AND2 U3970 ( .A(n13103), .B(n13104), .Z(n13102) );
    VMW_NOR4 U3995 ( .A(n13208), .B(n13209), .C(n13210), .D(n13211), .Z(n13207
        ) );
    VMW_AND3 U4052 ( .A(n13440), .B(n13441), .C(n13408), .Z(n13439) );
    VMW_OR2 U4149 ( .A(n13629), .B(n13622), .Z(n13631) );
    VMW_AND3 U4279 ( .A(n13767), .B(n13761), .C(n13768), .Z(n13766) );
    VMW_AOI211 U4758 ( .A(n13357), .B(n13551), .C(n14248), .D(n13237), .Z(
        n14247) );
    VMW_FD \temp_reg[42]  ( .D(\arr12639[42] ), .CP(Clk), .Q(\temp[42] ) );
    VMW_AO22 U4468 ( .A(n13910), .B(n13441), .C(n14041), .D(n13401), .Z(n14040
        ) );
    VMW_OAI22 U4643 ( .A(n13643), .B(n13717), .C(n13642), .D(n13723), .Z(
        n14189) );
    VMW_AO22 U4075 ( .A(n13486), .B(n13487), .C(\temp[21] ), .D(n13082), .Z(
        n13362) );
    VMW_AND2 U4345 ( .A(n13581), .B(n13322), .Z(n13333) );
    VMW_AOI211 U4362 ( .A(n13424), .B(n13870), .C(n13871), .D(n13872), .Z(
        n13869) );
    VMW_OAI22 U4573 ( .A(n13609), .B(n13620), .C(n13624), .D(n13649), .Z(
        n14139) );
    VMW_AOI211 U4891 ( .A(n13202), .B(n13526), .C(n14218), .D(n13340), .Z(
        n14305) );
    VMW_NAND2 U4901 ( .A(n13321), .B(n13337), .Z(n13884) );
    VMW_AO21 U5026 ( .A(n13481), .B(n14418), .C(n13103), .Z(n14417) );
    VMW_OAI22 U4926 ( .A(n13635), .B(n13720), .C(n13633), .D(n13719), .Z(
        n14338) );
    VMW_OAI22 U5286 ( .A(n13342), .B(n13760), .C(n13528), .D(n13200), .Z(
        n14462) );
    VMW_INV U5316 ( .A(n13241), .Z(n13570) );
    VMW_OAI22 U4554 ( .A(n13643), .B(n14103), .C(n13642), .D(n14112), .Z(
        n14128) );
    VMW_INV U5331 ( .A(n13113), .Z(n13498) );
    VMW_OAI22 U4664 ( .A(n13635), .B(n14119), .C(n13628), .D(n14096), .Z(
        n14201) );
    VMW_AND2 U5001 ( .A(n13880), .B(n13337), .Z(n14407) );
    VMW_INV U5191 ( .A(n13569), .Z(n13804) );
    VMW_INV U4230 ( .A(\temp[11] ), .Z(n13489) );
    VMW_OAI2222 U4853 ( .A(n13635), .B(n13723), .C(n13633), .D(n13722), .E(
        n13609), .F(n13721), .G(n13621), .H(n13716), .Z(n13306) );
    VMW_OAI22 U4948 ( .A(n13621), .B(n14163), .C(n13637), .D(n14164), .Z(
        n14348) );
    VMW_NAND3 U5048 ( .A(n13555), .B(n13550), .C(n13421), .Z(n13802) );
    VMW_AO22 U5244 ( .A(n14026), .B(n13543), .C(n14025), .D(n13550), .Z(n14379
        ) );
    VMW_INV U5378 ( .A(KEY[2]), .Z(n14155) );
    VMW_INV U5455 ( .A(n13910), .Z(n13921) );
    VMW_AND2 U4421 ( .A(n13425), .B(n13107), .Z(n13980) );
    VMW_AO22 U4090 ( .A(n13523), .B(n13505), .C(n13524), .D(n13525), .Z(n13201
        ) );
    VMW_OAI22 U4100 ( .A(n13531), .B(n13546), .C(n13547), .D(n13537), .Z(
        n13438) );
    VMW_INV U5174 ( .A(n13464), .Z(n13471) );
    VMW_OR4 U4681 ( .A(n14208), .B(n14209), .C(n14206), .D(n14207), .Z(n13185)
         );
    VMW_OR4 U4711 ( .A(n14223), .B(n14224), .C(n14221), .D(n14222), .Z(n13218)
         );
    VMW_AND3 U3978 ( .A(n13139), .B(n13140), .C(n13141), .Z(n13138) );
    VMW_NOR4 U4013 ( .A(n13290), .B(n13291), .C(n13292), .D(n13293), .Z(n13289
        ) );
    VMW_NOR4 U4034 ( .A(n13366), .B(n13367), .C(n13368), .D(n13369), .Z(n13365
        ) );
    VMW_OR2 U4127 ( .A(\i[1] ), .B(\i[0] ), .Z(n13607) );
    VMW_OAI2222 U4736 ( .A(n13640), .B(n13726), .C(n13637), .D(n13718), .E(
        n13631), .F(n13722), .G(n13628), .H(n13721), .Z(n13224) );
    VMW_OR4 U5153 ( .A(n13874), .B(n13165), .C(n13406), .D(n14371), .Z(n14066)
         );
    VMW_OAI22 U4217 ( .A(n13697), .B(n13698), .C(n13694), .D(n13699), .Z(
        n13696) );
    VMW_AND2 U4387 ( .A(n13904), .B(n13598), .Z(n13907) );
    VMW_NOR5 U4406 ( .A(n13843), .B(n13948), .C(n13852), .D(n13949), .E(n13882
        ), .Z(n13947) );
    VMW_OAI22 U4874 ( .A(n13641), .B(n13714), .C(n13626), .D(n13713), .Z(
        n14300) );
    VMW_AO22 U5263 ( .A(n14407), .B(n13322), .C(n14055), .D(n13578), .Z(n13949
        ) );
    VMW_INV U5472 ( .A(n14276), .Z(n14424) );
    VMW_OR2 U4596 ( .A(n13472), .B(n13481), .Z(n13698) );
    VMW_AND2 U4294 ( .A(n13779), .B(n13543), .Z(n13780) );
    VMW_OAI211 U4304 ( .A(n13540), .B(n13792), .C(n13793), .D(n13794), .Z(
        n13791) );
    VMW_XNOR2 U4485 ( .A(\temp[51] ), .B(n13415), .Z(n14064) );
    VMW_OAI22 U4515 ( .A(n13621), .B(n14096), .C(n13619), .D(n14097), .Z(
        n14104) );
    VMW_NOR2 U4967 ( .A(n13410), .B(n13896), .Z(n13956) );
    VMW_INV U5370 ( .A(KEY[30]), .Z(n14112) );
    VMW_AND2 U4183 ( .A(n13467), .B(n13459), .Z(n13663) );
    VMW_OAI22 U4602 ( .A(n13609), .B(n13719), .C(n13626), .D(n13716), .Z(
        n14157) );
    VMW_OAI22 U4625 ( .A(n13609), .B(n14170), .C(n13616), .D(n14167), .Z(
        n14179) );
    VMW_AO21 U5040 ( .A(n13525), .B(n13200), .C(n13943), .Z(n14363) );
    VMW_OAI22 U4792 ( .A(n13637), .B(n14092), .C(n13635), .D(n14089), .Z(
        n13260) );
    VMW_AND2 U4323 ( .A(n13562), .B(n13812), .Z(n13813) );
    VMW_OAI22 U4532 ( .A(n13644), .B(n13646), .C(n13640), .D(n14096), .Z(
        n14114) );
    VMW_NAND4 U5067 ( .A(n14425), .B(n13832), .C(n13606), .D(n13334), .Z(
        n13857) );
    VMW_OAI22 U4940 ( .A(n13616), .B(n13727), .C(n13609), .D(n14163), .Z(
        n14344) );
    VMW_INV U5357 ( .A(\temp[2] ), .Z(n13538) );
    VMW_AO22 U4098 ( .A(n13541), .B(n13542), .C(\temp[1] ), .D(n13217), .Z(
        n13540) );
    VMW_AO22 U4108 ( .A(n13565), .B(n13566), .C(\temp[26] ), .D(n13266), .Z(
        n13564) );
    VMW_OR4 U4689 ( .A(n14212), .B(n14213), .C(n14210), .D(n14211), .Z(n13180)
         );
    VMW_FD \temp_reg[14]  ( .D(\arr12639[14] ), .CP(Clk), .Q(\temp[14] ) );
    VMW_FD \OUT_reg[32]  ( .D(\arr12639[3] ), .CP(Clk), .Q(OUT[32]) );
    VMW_OR4 U4719 ( .A(n14227), .B(n14228), .C(n14225), .D(n14226), .Z(n13213)
         );
    VMW_INV U4166 ( .A(KEY[4]), .Z(n13646) );
    VMW_INV U4238 ( .A(KEY[36]), .Z(n13726) );
    VMW_FD \temp_reg[27]  ( .D(\arr12639[27] ), .CP(Clk), .Q(\temp[27] ) );
    VMW_FD \OUT_reg[18]  ( .D(\arr12639[13] ), .CP(Clk), .Q(OUT[18]) );
    VMW_AND2 U4429 ( .A(n13505), .B(n13528), .Z(n13522) );
    VMW_OAI22 U4777 ( .A(n13628), .B(n14094), .C(n14085), .D(n13643), .Z(
        n14253) );
    VMW_AO22 U5082 ( .A(n13273), .B(n13282), .C(n13272), .D(n13803), .Z(n13861
        ) );
    VMW_NAND3 U5112 ( .A(n13103), .B(n13353), .C(n13104), .Z(n14327) );
    VMW_AND2 U4256 ( .A(n13156), .B(n13140), .Z(n13151) );
    VMW_AND2 U4447 ( .A(n13758), .B(n13520), .Z(n14007) );
    VMW_OAI22 U5222 ( .A(n13778), .B(n13546), .C(n13994), .D(n13537), .Z(
        n14422) );
    VMW_INV U5433 ( .A(n13780), .Z(n13799) );
    VMW_NOR2 U4271 ( .A(n13507), .B(n13516), .Z(n13524) );
    VMW_OAI22 U4835 ( .A(n13628), .B(n13722), .C(n13626), .D(n13721), .Z(
        n14281) );
    VMW_AO22 U5205 ( .A(n13974), .B(n13453), .C(n13975), .D(n13659), .Z(n14415
        ) );
    VMW_INV U5395 ( .A(n13507), .Z(n13758) );
    VMW_INV U5414 ( .A(n13472), .Z(n14418) );
    VMW_AND2 U4460 ( .A(n13553), .B(n13546), .Z(n14026) );
    VMW_OAI22 U4812 ( .A(n13623), .B(n13635), .C(n13620), .D(n13633), .Z(
        n14272) );
    VMW_AND2 U4982 ( .A(n13907), .B(n13602), .Z(n13967) );
    VMW_AO22 U5135 ( .A(n13200), .B(n13530), .C(n13342), .D(n13943), .Z(n13945
        ) );
    VMW_AO21 U3936 ( .A(\temp[52] ), .B(n13005), .C(n13017), .Z(\arr12639[52] 
        ) );
    VMW_AO21 U3938 ( .A(\temp[50] ), .B(n13005), .C(n13019), .Z(\arr12639[50] 
        ) );
    VMW_AO21 U3944 ( .A(\temp[44] ), .B(n13005), .C(n13025), .Z(\arr12639[44] 
        ) );
    VMW_NAND3 U3963 ( .A(n13069), .B(n13070), .C(n13071), .Z(n13068) );
    VMW_NOR4 U3986 ( .A(n13165), .B(n13166), .C(n13167), .D(n13168), .Z(n13164
        ) );
    VMW_AND3 U4041 ( .A(n13400), .B(n13401), .C(n13402), .Z(n13399) );
    VMW_INV U4141 ( .A(KEY[55]), .Z(n13623) );
    VMW_AND2 U4650 ( .A(n14192), .B(n13447), .Z(n13753) );
    VMW_OAI22 U4750 ( .A(n13640), .B(n14172), .C(n13637), .D(n14155), .Z(
        n14244) );
    VMW_AOI211 U4899 ( .A(n13703), .B(n13364), .C(n14313), .D(n13350), .Z(
        n14312) );
    VMW_OAI22 U4909 ( .A(n13626), .B(n14170), .C(n13624), .D(n14166), .Z(
        n14329) );
    VMW_NAND3 U5009 ( .A(n13444), .B(n13401), .C(n13909), .Z(n14356) );
    VMW_INV U5199 ( .A(n13444), .Z(n13897) );
    VMW_INV U5339 ( .A(n13118), .Z(n13490) );
    VMW_AND2 U5035 ( .A(n14192), .B(n13733), .Z(n13741) );
    VMW_FD \OUT_reg[3]  ( .D(\arr12639[47] ), .CP(Clk), .Q(OUT[3]) );
    VMW_AND3 U4356 ( .A(n13859), .B(n13761), .C(n13860), .Z(n13858) );
    VMW_AO21 U4371 ( .A(n13787), .B(n13550), .C(n13890), .Z(n13889) );
    VMW_OAI22 U4560 ( .A(n13635), .B(n14090), .C(n13633), .D(n13639), .Z(
        n13100) );
    VMW_INV U5295 ( .A(\i[4] ), .Z(n13610) );
    VMW_INV U5305 ( .A(n13038), .Z(n13455) );
    VMW_INV U5484 ( .A(n13952), .Z(n14035) );
    VMW_AO22 U4882 ( .A(X[0]), .B(n13774), .C(n13773), .D(\temp[7] ), .Z(
        n13030) );
    VMW_OR4 U4912 ( .A(n14330), .B(n14331), .C(n14328), .D(n14329), .Z(n13366)
         );
    VMW_INV U5322 ( .A(n13174), .Z(n13513) );
    VMW_OAI22 U4547 ( .A(n13609), .B(n13615), .C(n13628), .D(n13649), .Z(
        n14125) );
    VMW_OAI22 U4935 ( .A(n13619), .B(n14172), .C(n13616), .D(n14155), .Z(
        n14343) );
    VMW_NAND3 U5012 ( .A(n13652), .B(n13650), .C(n13653), .Z(n13679) );
    VMW_INV U5182 ( .A(n13505), .Z(n13525) );
    VMW_AO22 U4066 ( .A(n13462), .B(n13463), .C(\temp[31] ), .D(n13048), .Z(
        n13069) );
    VMW_AO22 U4083 ( .A(n13500), .B(n13506), .C(\temp[16] ), .D(n13189), .Z(
        n13505) );
    VMW_AO22 U4113 ( .A(n13576), .B(n13577), .C(\temp[9] ), .D(n13299), .Z(
        n13575) );
    VMW_INV U4223 ( .A(KEY[33]), .Z(n13712) );
    VMW_OAI22 U4677 ( .A(n13635), .B(n14094), .C(n14085), .D(n13619), .Z(
        n14206) );
    VMW_OAI22 U4809 ( .A(n13631), .B(n14103), .C(n13628), .D(n14112), .Z(
        n14269) );
    VMW_NAND3 U4999 ( .A(n13688), .B(n14406), .C(n13351), .Z(n13706) );
    VMW_FD \temp_reg[3]  ( .D(\arr12639[3] ), .CP(Clk), .Q(\temp[3] ) );
    VMW_NAND4 U5099 ( .A(n13746), .B(n14434), .C(n14435), .D(n14314), .Z(
        n14022) );
    VMW_AO22 U5239 ( .A(n14019), .B(n13447), .C(n14020), .D(n13161), .Z(n14479
        ) );
    VMW_INV U5428 ( .A(n13763), .Z(n13767) );
    VMW_NAND2 U5109 ( .A(n13238), .B(n13535), .Z(n13590) );
    VMW_AND2 U4432 ( .A(n13989), .B(n13990), .Z(n13764) );
    VMW_OAI22 U4692 ( .A(n13642), .B(n14092), .C(n13641), .D(n14089), .Z(
        n13183) );
    VMW_OAI22 U4840 ( .A(n13616), .B(n14163), .C(n13633), .D(n14164), .Z(
        n14282) );
    VMW_AO22 U5257 ( .A(n14046), .B(n13464), .C(n14047), .D(n13471), .Z(n14445
        ) );
    VMW_INV U5446 ( .A(n14436), .Z(n14438) );
    VMW_AOI211 U4702 ( .A(n13759), .B(n14011), .C(n14220), .D(n13203), .Z(
        n14219) );
    VMW_OR2 U4134 ( .A(n13611), .B(n13613), .Z(n13616) );
    VMW_OAI22 U4725 ( .A(n13643), .B(n13712), .C(n13642), .D(n14172), .Z(
        n14231) );
    VMW_OAI211 U5167 ( .A(n13439), .B(n13442), .C(n13396), .D(n13596), .Z(
        n14391) );
    VMW_AO21 U3956 ( .A(\temp[32] ), .B(n13005), .C(n13037), .Z(\arr12639[32] 
        ) );
    VMW_NOR2 U3971 ( .A(n13106), .B(n13107), .Z(n13105) );
    VMW_AND3 U4008 ( .A(n13272), .B(n13273), .C(n13274), .Z(n13271) );
    VMW_AND2 U4198 ( .A(n13681), .B(n13682), .Z(n13424) );
    VMW_NOR2 U4204 ( .A(n13353), .B(n13688), .Z(n13687) );
    VMW_AOI21 U4394 ( .A(n13901), .B(n13909), .C(n13915), .Z(n13914) );
    VMW_AND3 U5140 ( .A(n13328), .B(n13321), .C(n13604), .Z(n14450) );
    VMW_AO22 U4415 ( .A(n13972), .B(n13456), .C(n13973), .D(n13651), .Z(n13971
        ) );
    VMW_NAND3 U4338 ( .A(n13334), .B(n13835), .C(n13575), .Z(n13834) );
    VMW_OAI22 U4529 ( .A(n13624), .B(n14094), .C(n14085), .D(n13641), .Z(
        n14110) );
    VMW_OAI22 U4585 ( .A(n13635), .B(n14092), .C(n13633), .D(n14089), .Z(
        n13076) );
    VMW_OAI22 U4867 ( .A(n13616), .B(n14172), .C(n13644), .D(n14155), .Z(
        n14297) );
    VMW_MUX2 U5270 ( .A(n14491), .B(\temp[1] ), .S(n13005), .Z(\arr12639[1] )
         );
    VMW_INV U5461 ( .A(n13947), .Z(n14451) );
    VMW_FD \temp_reg[37]  ( .D(\arr12639[37] ), .CP(Clk), .Q(\temp[37] ) );
    VMW_FD \OUT_reg[11]  ( .D(\arr12639[46] ), .CP(Clk), .Q(OUT[11]) );
    VMW_OAI22 U4619 ( .A(n13640), .B(n13713), .C(n13628), .D(n13712), .Z(
        n14177) );
    VMW_FD \OUT_reg[22]  ( .D(\arr12639[29] ), .CP(Clk), .Q(OUT[22]) );
    VMW_OR4 U4789 ( .A(n14259), .B(n14260), .C(n14257), .D(n14258), .Z(n13257)
         );
    VMW_AO22 U4091 ( .A(n13523), .B(n13525), .C(n13524), .D(n13505), .Z(n13526
        ) );
    VMW_INV U4231 ( .A(KEY[10]), .Z(n13719) );
    VMW_XOR2 U4420 ( .A(n13979), .B(\temp[41] ), .Z(n13978) );
    VMW_OR4 U4852 ( .A(n14288), .B(n14289), .C(n14286), .D(n14287), .Z(n13305)
         );
    VMW_OAI22 U4949 ( .A(n13609), .B(n14166), .C(n13619), .D(n14167), .Z(
        n14349) );
    VMW_OR3 U5049 ( .A(n13356), .B(n13591), .C(n14422), .Z(n13801) );
    VMW_INV U5379 ( .A(KEY[11]), .Z(n14169) );
    VMW_OAI22 U4710 ( .A(n13633), .B(n14172), .C(n13609), .D(n14155), .Z(
        n14224) );
    VMW_AO22 U5245 ( .A(n14027), .B(n13451), .C(X[39]), .D(Start), .Z(n14482)
         );
    VMW_INV U5454 ( .A(n13905), .Z(n13912) );
    VMW_AO22 U4101 ( .A(n13549), .B(n13543), .C(n13238), .D(n13550), .Z(n13548
        ) );
    VMW_OAI22 U4680 ( .A(n13618), .B(n13641), .C(n13615), .D(n13640), .Z(
        n14209) );
    VMW_INV U5175 ( .A(n13475), .Z(n13353) );
    VMW_AO22 U4126 ( .A(n13333), .B(n13575), .C(n13605), .D(n13606), .Z(n13604
        ) );
    VMW_OAI22 U4737 ( .A(n13642), .B(n13725), .C(n13641), .D(n13724), .Z(
        n13225) );
    VMW_NAND2 U5152 ( .A(n13163), .B(n14190), .Z(n14372) );
    VMW_INV U4148 ( .A(KEY[7]), .Z(n13630) );
    VMW_NAND2 U4216 ( .A(n13695), .B(n13681), .Z(n13694) );
    VMW_OAI22 U4875 ( .A(n13640), .B(n13716), .C(n13624), .D(n13715), .Z(
        n14301) );
    VMW_AND2 U4386 ( .A(n13401), .B(n13902), .Z(n13906) );
    VMW_AND2 U4597 ( .A(n13362), .B(n14150), .Z(n13702) );
    VMW_OR4 U4407 ( .A(n13951), .B(n13952), .C(n13920), .D(n13953), .Z(n13950)
         );
    VMW_AO22 U4759 ( .A(X[38]), .B(n13774), .C(n13773), .D(\temp[27] ), .Z(
        n13010) );
    VMW_MUX2 U5262 ( .A(n14487), .B(\temp[22] ), .S(n13005), .Z(\arr12639[22] 
        ) );
    VMW_INV U5473 ( .A(n14321), .Z(n13893) );
    VMW_FD \temp_reg[10]  ( .D(\arr12639[10] ), .CP(Clk), .Q(\temp[10] ) );
    VMW_FD \OUT_reg[36]  ( .D(\arr12639[19] ), .CP(Clk), .Q(OUT[36]) );
    VMW_AO21 U3943 ( .A(\temp[45] ), .B(n13005), .C(n13024), .Z(\arr12639[45] 
        ) );
    VMW_AO21 U3951 ( .A(\temp[37] ), .B(n13005), .C(n13032), .Z(\arr12639[37] 
        ) );
    VMW_NOR4 U3988 ( .A(n13175), .B(n13176), .C(n13177), .D(n13178), .Z(n13174
        ) );
    VMW_AND3 U3994 ( .A(n13204), .B(n13205), .C(n13206), .Z(n13203) );
    VMW_AND3 U4053 ( .A(n13397), .B(n13443), .C(n13444), .Z(n13442) );
    VMW_OAI21 U4278 ( .A(n13764), .B(n13200), .C(n13765), .Z(n13763) );
    VMW_AO22 U4469 ( .A(n13906), .B(n13444), .C(n13448), .D(n13897), .Z(n14042
        ) );
    VMW_AO21 U5027 ( .A(n13682), .B(n14417), .C(n13359), .Z(n13352) );
    VMW_FD \temp_reg[23]  ( .D(\arr12639[23] ), .CP(Clk), .Q(\temp[23] ) );
    VMW_NAND3 U4344 ( .A(n13581), .B(n13334), .C(n13331), .Z(n13838) );
    VMW_OR2 U4363 ( .A(n13141), .B(n13730), .Z(n13162) );
    VMW_OAI22 U4642 ( .A(n13641), .B(n13722), .C(n13640), .D(n13721), .Z(
        n14188) );
    VMW_AOI211 U4890 ( .A(n13200), .B(n14008), .C(n14220), .D(n13338), .Z(
        n13860) );
    VMW_AO22 U5287 ( .A(n14076), .B(n13451), .C(X[27]), .D(Start), .Z(n14500)
         );
    VMW_INV U5317 ( .A(\temp[22] ), .Z(n13482) );
    VMW_AOI211 U4900 ( .A(n13144), .B(n14315), .C(n13930), .D(n14316), .Z(
        n14314) );
    VMW_OAI22 U4555 ( .A(n13628), .B(n13646), .C(n13626), .D(n14119), .Z(
        n14129) );
    VMW_OAI22 U4572 ( .A(n13643), .B(n13647), .C(n13642), .D(n13646), .Z(
        n14138) );
    VMW_OAI22 U4927 ( .A(n13640), .B(n13722), .C(n13637), .D(n13721), .Z(
        n14339) );
    VMW_INV U5330 ( .A(n13189), .Z(n13506) );
    VMW_AND3 U4001 ( .A(n13238), .B(n13239), .C(n13240), .Z(n13237) );
    VMW_AND3 U4026 ( .A(n13341), .B(n13342), .C(n13204), .Z(n13340) );
    VMW_AND2 U4048 ( .A(n13424), .B(n13425), .Z(n13423) );
    VMW_AO22 U4074 ( .A(n13484), .B(n13485), .C(\temp[23] ), .D(n13072), .Z(
        n13351) );
    VMW_OR4 U4665 ( .A(n14200), .B(n14201), .C(n14198), .D(n14199), .Z(n13195)
         );
    VMW_AND3 U5000 ( .A(n13730), .B(n13156), .C(n13154), .Z(n13145) );
    VMW_INV U5190 ( .A(n13543), .Z(n13550) );
    VMW_NOR2 U4378 ( .A(n13396), .B(n13401), .Z(n13900) );
    VMW_OAI22 U4569 ( .A(n13642), .B(n14091), .C(n13631), .D(n13634), .Z(
        n13091) );
    VMW_FD \temp_reg[33]  ( .D(\arr12639[33] ), .CP(Clk), .Q(\temp[33] ) );
    VMW_FD \OUT_reg[15]  ( .D(\arr12639[62] ), .CP(Clk), .Q(OUT[15]) );
    VMW_OR2 U4153 ( .A(n13617), .B(n13629), .Z(n13635) );
    VMW_AND2 U4174 ( .A(n13464), .B(n13654), .Z(n13653) );
    VMW_OAI22 U4659 ( .A(n13615), .B(n13631), .C(n13609), .D(n13649), .Z(
        n13192) );
    VMW_NAND3 U5090 ( .A(n13103), .B(n13424), .C(n13360), .Z(n14309) );
    VMW_AND2 U5100 ( .A(n13856), .B(n13838), .Z(n13887) );
    VMW_FD \temp_reg[19]  ( .D(\arr12639[19] ), .CP(Clk), .Q(\temp[19] ) );
    VMW_FD \OUT_reg[26]  ( .D(\arr12639[12] ), .CP(Clk), .Q(OUT[26]) );
    VMW_OR2 U4244 ( .A(n13729), .B(n13496), .Z(n13728) );
    VMW_AO22 U4765 ( .A(X[20]), .B(n13774), .C(n13773), .D(\temp[21] ), .Z(
        n13016) );
    VMW_AO22 U4827 ( .A(X[26]), .B(n13774), .C(n13773), .D(\temp[12] ), .Z(
        n13025) );
    VMW_MUX2 U5230 ( .A(n14473), .B(\temp[3] ), .S(n13005), .Z(\arr12639[3] )
         );
    VMW_INV U5421 ( .A(n13728), .Z(n13149) );
    VMW_AO22 U4263 ( .A(n13750), .B(n13447), .C(n13154), .D(n13733), .Z(n13165
        ) );
    VMW_OR2 U4455 ( .A(n13162), .B(n13499), .Z(n14019) );
    VMW_NAND2 U4472 ( .A(n13071), .B(n13659), .Z(n14046) );
    VMW_OAI22 U4800 ( .A(n13619), .B(n14092), .C(n13616), .D(n14089), .Z(
        n13255) );
    VMW_AO22 U5217 ( .A(n13988), .B(n13760), .C(n13764), .D(n13200), .Z(n14469
        ) );
    VMW_INV U5387 ( .A(n13450), .Z(n14505) );
    VMW_INV U5406 ( .A(n13584), .Z(n13328) );
    VMW_NAND2 U4990 ( .A(n14400), .B(n14058), .Z(n14395) );
    VMW_OAI22 U4742 ( .A(n13624), .B(n14172), .C(n13621), .D(n14155), .Z(
        n14240) );
    VMW_AND3 U5127 ( .A(n13144), .B(n13162), .C(n13732), .Z(n13931) );
    VMW_OR2 U4286 ( .A(n13437), .B(n13531), .Z(n13777) );
    VMW_OAI22 U4849 ( .A(n13628), .B(n14172), .C(n13626), .D(n14155), .Z(
        n14287) );
    VMW_OR4 U5149 ( .A(n13940), .B(n13933), .C(n13957), .D(n14458), .Z(n14063)
         );
    VMW_AO22 U5279 ( .A(n14070), .B(n13451), .C(X[3]), .D(Start), .Z(n14496)
         );
    VMW_INV U5468 ( .A(n14040), .Z(n14442) );
    VMW_FD \temp_reg[7]  ( .D(\arr12639[7] ), .CP(Clk), .Q(\temp[7] ) );
    VMW_OAI22 U4975 ( .A(n13543), .B(n13888), .C(n14377), .D(n14375), .Z(
        n14376) );
    VMW_NOR2 U4316 ( .A(n13564), .B(n13562), .Z(n13809) );
    VMW_OAI22 U4507 ( .A(n13615), .B(n13621), .C(n13644), .D(n13645), .Z(
        n14098) );
    VMW_OAI22 U4497 ( .A(n13615), .B(n13616), .C(n13609), .D(n14085), .Z(
        n14084) );
    VMW_OAI2222 U4637 ( .A(n13633), .B(n13724), .C(n13609), .D(n13726), .E(
        n13626), .F(n13717), .G(n13624), .H(n13723), .Z(n13115) );
    VMW_INV U5362 ( .A(KEY[62]), .Z(n14092) );
    VMW_OAI22 U4780 ( .A(n13616), .B(n14119), .C(n13642), .D(n14096), .Z(
        n14256) );
    VMW_AND3 U5052 ( .A(n13537), .B(n13555), .C(n13781), .Z(n13797) );
    VMW_NOR4 U4006 ( .A(n13262), .B(n13263), .C(n13264), .D(n13265), .Z(n13261
        ) );
    VMW_INV U4191 ( .A(Start), .Z(n13451) );
    VMW_OAI22 U4610 ( .A(n13641), .B(n14169), .C(n13640), .D(n14170), .Z(
        n14168) );
    VMW_INV U4196 ( .A(\temp[20] ), .Z(n13476) );
    VMW_AO21 U4331 ( .A(n13813), .B(n13272), .C(n13822), .Z(n13821) );
    VMW_OR4 U4952 ( .A(n14350), .B(n14351), .C(n14348), .D(n14349), .Z(n13386)
         );
    VMW_OAI211 U5075 ( .A(n13834), .B(n13840), .C(n14426), .D(n13881), .Z(
        n14399) );
    VMW_FD \OUT_reg[7]  ( .D(\arr12639[63] ), .CP(Clk), .Q(OUT[7]) );
    VMW_AND2 U4336 ( .A(n13581), .B(n13584), .Z(n13832) );
    VMW_OAI22 U4520 ( .A(n13641), .B(n14091), .C(n13631), .D(n13636), .Z(
        n13042) );
    VMW_OAI22 U4527 ( .A(n13626), .B(n14089), .C(n13624), .D(n14090), .Z(
        n13046) );
    VMW_OAI2222 U4869 ( .A(n13643), .B(n13719), .C(n13642), .D(n13727), .E(
        n13609), .F(n13713), .G(n13619), .H(n13712), .Z(n13296) );
    VMW_OAI211 U5169 ( .A(n13910), .B(n14409), .C(n13401), .D(n13396), .Z(
        n14394) );
    VMW_AO22 U5259 ( .A(n14051), .B(n13451), .C(X[5]), .D(Start), .Z(n14486)
         );
    VMW_INV U5345 ( .A(n13304), .Z(n13574) );
    VMW_INV U5448 ( .A(n13849), .Z(n14304) );
    VMW_FD \temp_reg[5]  ( .D(\arr12639[5] ), .CP(Clk), .Q(\temp[5] ) );
    VMW_INV U5342 ( .A(n13294), .Z(n13580) );
    VMW_OAI22 U4955 ( .A(n13640), .B(n14173), .C(n13631), .D(n13725), .Z(
        n13389) );
    VMW_AO21 U5072 ( .A(n13572), .B(n13835), .C(n13324), .Z(n13321) );
    VMW_OAI22 U4617 ( .A(n13643), .B(n14169), .C(n13642), .D(n14170), .Z(
        n14175) );
    VMW_AND3 U4021 ( .A(n13327), .B(n13328), .C(n13329), .Z(n13326) );
    VMW_OAI22 U4787 ( .A(n13628), .B(n13647), .C(n13626), .D(n13646), .Z(
        n14259) );
    VMW_AND3 U5055 ( .A(n13537), .B(n13781), .C(n13238), .Z(n13422) );
    VMW_FD \OUT_reg[5]  ( .D(\arr12639[55] ), .CP(Clk), .Q(OUT[5]) );
    VMW_AOI21 U4281 ( .A(n13520), .B(n13756), .C(n13772), .Z(n13771) );
    VMW_AND2 U4311 ( .A(n13562), .B(n13808), .Z(n13807) );
    VMW_NOR2 U4490 ( .A(n13806), .B(n13808), .Z(n14072) );
    VMW_OAI22 U4630 ( .A(n13628), .B(n13725), .C(n13626), .D(n13724), .Z(
        n13126) );
    VMW_INV U5365 ( .A(KEY[20]), .Z(n14119) );
    VMW_OAI22 U4500 ( .A(n13630), .B(n13631), .C(n13627), .D(n13628), .Z(
        n14088) );
    VMW_AO22 U4358 ( .A(n13807), .B(n13861), .C(n13862), .D(n13274), .Z(n13416
        ) );
    VMW_NAND4 U4972 ( .A(n13747), .B(n14372), .C(n14373), .D(n14374), .Z(
        n14371) );
    VMW_FD \temp_reg[31]  ( .D(\arr12639[31] ), .CP(Clk), .Q(\temp[31] ) );
    VMW_FD \temp_reg[28]  ( .D(\arr12639[28] ), .CP(Clk), .Q(\temp[28] ) );
    VMW_FD \OUT_reg[17]  ( .D(\arr12639[37] ), .CP(Clk), .Q(OUT[17]) );
    VMW_OAI22 U4549 ( .A(n13625), .B(n13640), .C(n13623), .D(n13637), .Z(
        n14127) );
    VMW_AND3 U3993 ( .A(n13200), .B(n13201), .C(n13202), .Z(n13199) );
    VMW_AO22 U4068 ( .A(n13468), .B(n13469), .C(\temp[30] ), .D(n13058), .Z(
        n13467) );
    VMW_FD \OUT_reg[24]  ( .D(\arr12639[4] ), .CP(Clk), .Q(OUT[24]) );
    VMW_AO22 U4073 ( .A(n13482), .B(n13483), .C(\temp[22] ), .D(n13077), .Z(
        n13481) );
    VMW_INV U4154 ( .A(KEY[61]), .Z(n13636) );
    VMW_OAI22 U4679 ( .A(n13633), .B(n13645), .C(n13609), .D(n13648), .Z(
        n14208) );
    VMW_INV U4168 ( .A(KEY[37]), .Z(n13648) );
    VMW_NOR2 U4173 ( .A(n13467), .B(n13459), .Z(n13652) );
    VMW_NOR2 U4243 ( .A(n13499), .B(n13496), .Z(n13144) );
    VMW_AO22 U4264 ( .A(n13751), .B(n13752), .C(n13753), .D(n13730), .Z(n13167
        ) );
    VMW_OAI22 U4745 ( .A(n13609), .B(n13723), .C(n13616), .D(n13716), .Z(
        n13235) );
    VMW_AOI21 U5120 ( .A(n14356), .B(n14442), .C(n13396), .Z(n13917) );
    VMW_XOR2 U4452 ( .A(n14016), .B(\temp[62] ), .Z(n14015) );
    VMW_AND3 U4475 ( .A(n13456), .B(n13656), .C(n13663), .Z(n14050) );
    VMW_OAI22 U4807 ( .A(n13609), .B(n13630), .C(n13644), .D(n13649), .Z(
        n13249) );
    VMW_OAI21 U4997 ( .A(n13105), .B(n14144), .C(n13362), .Z(n14310) );
    VMW_AO22 U5210 ( .A(n13689), .B(n13478), .C(n13980), .D(n13682), .Z(n14404
        ) );
    VMW_INV U5380 ( .A(KEY[27]), .Z(n14170) );
    VMW_INV U5401 ( .A(n13240), .Z(n14401) );
    VMW_AO22 U4762 ( .A(X[62]), .B(n13774), .C(n13773), .D(\temp[24] ), .Z(
        n13013) );
    VMW_AO22 U4820 ( .A(n14275), .B(n13282), .C(n13813), .D(n13414), .Z(n13278
        ) );
    VMW_AO22 U5237 ( .A(n14017), .B(n13451), .C(X[41]), .D(Start), .Z(n14478)
         );
    VMW_INV U5426 ( .A(n13151), .Z(n13875) );
    VMW_OAI22 U4779 ( .A(n13641), .B(n14097), .C(n13640), .D(n14102), .Z(
        n14255) );
    VMW_AO21 U5097 ( .A(n13447), .B(n13141), .C(n13736), .Z(n14315) );
    VMW_OR4 U5107 ( .A(n13845), .B(n13882), .C(n13886), .D(n14317), .Z(n14024)
         );
    VMW_FD \temp_reg[12]  ( .D(\arr12639[12] ), .CP(Clk), .Q(\temp[12] ) );
    VMW_FD \OUT_reg[34]  ( .D(\arr12639[11] ), .CP(Clk), .Q(OUT[34]) );
    VMW_OAI21 U4258 ( .A(n13158), .B(n13447), .C(n13738), .Z(n13737) );
    VMW_AND2 U4449 ( .A(n13755), .B(n14011), .Z(n14010) );
    VMW_FD \temp_reg[38]  ( .D(\arr12639[38] ), .CP(Clk), .Q(\temp[38] ) );
    VMW_FD \temp_reg[21]  ( .D(\arr12639[21] ), .CP(Clk), .Q(\temp[21] ) );
    VMW_OAI22 U4662 ( .A(n13621), .B(n14103), .C(n13619), .D(n14112), .Z(
        n14199) );
    VMW_AND3 U5007 ( .A(n13653), .B(n13651), .C(n13655), .Z(n14412) );
    VMW_AND2 U4054 ( .A(\i6749[5] ), .B(n13445), .Z(n14504) );
    VMW_AND2 U4343 ( .A(n13837), .B(n13328), .Z(n13331) );
    VMW_INV U5197 ( .A(n13441), .Z(n13401) );
    VMW_AND2 U4364 ( .A(n13156), .B(n13149), .Z(n13873) );
    VMW_OAI22 U4552 ( .A(n13621), .B(n14090), .C(n13619), .D(n13639), .Z(
        n13080) );
    VMW_OAI2222 U4575 ( .A(n13630), .B(n13640), .C(n13627), .D(n13637), .E(
        n13625), .F(n13635), .G(n13623), .H(n13633), .Z(n13094) );
    VMW_OR4 U4920 ( .A(n14334), .B(n14335), .C(n14332), .D(n14333), .Z(n13391)
         );
    VMW_INV U5337 ( .A(n13123), .Z(n13503) );
    VMW_OAI2222 U4645 ( .A(n13621), .B(n13725), .C(n13619), .D(n13724), .E(
        n13616), .F(n13726), .G(n13644), .H(n13718), .Z(n13130) );
    VMW_OAI211 U4897 ( .A(n14308), .B(n13694), .C(n14309), .D(n14310), .Z(
        n13867) );
    VMW_AND4 U4907 ( .A(n13869), .B(n14325), .C(n14326), .D(n14327), .Z(n14324
        ) );
    VMW_MUX2 U5280 ( .A(n14496), .B(\temp[15] ), .S(n13005), .Z(\arr12639[15] 
        ) );
    VMW_INV U5310 ( .A(\temp[26] ), .Z(n13565) );
    VMW_INV U5491 ( .A(n14475), .Z(n13859) );
    VMW_AND2 U4211 ( .A(n13688), .B(n13685), .Z(n13690) );
    VMW_AND2 U4381 ( .A(n13596), .B(n13603), .Z(n13409) );
    VMW_AND3 U4400 ( .A(n13453), .B(n13660), .C(n13661), .Z(n13932) );
    VMW_AOI211 U4969 ( .A(n13813), .B(n13277), .C(n13411), .D(n13413), .Z(
        n14368) );
    VMW_AND4 U5020 ( .A(n13364), .B(n13424), .C(n13688), .D(n13686), .Z(n13711
        ) );
    VMW_NAND2 U5069 ( .A(n13839), .B(n13584), .Z(n13854) );
    VMW_MUX2 U5265 ( .A(n14488), .B(\temp[21] ), .S(n13005), .Z(\arr12639[21] 
        ) );
    VMW_INV U5359 ( .A(\temp[1] ), .Z(n13541) );
    VMW_INV U5474 ( .A(n14322), .Z(n14439) );
    VMW_OAI22 U4590 ( .A(n13641), .B(n13647), .C(n13640), .D(n13646), .Z(
        n14149) );
    VMW_OAI22 U4872 ( .A(n13631), .B(n14170), .C(n13628), .D(n14166), .Z(
        n14298) );
    VMW_OR4 U5155 ( .A(n13889), .B(n13791), .C(n14376), .D(n14378), .Z(n14068)
         );
    VMW_NOR4 U3976 ( .A(n13129), .B(n13130), .C(n13131), .D(n13132), .Z(n13128
        ) );
    VMW_AO22 U4121 ( .A(n13544), .B(n13595), .C(\temp[3] ), .D(n13380), .Z(
        n13444) );
    VMW_OAI22 U4730 ( .A(n13635), .B(n14160), .C(n13633), .D(n14161), .Z(
        n13231) );
    VMW_INV U5172 ( .A(n13456), .Z(n13651) );
    VMW_AO22 U4096 ( .A(n13462), .B(n13536), .C(\temp[31] ), .D(n13222), .Z(
        n13535) );
    VMW_AO22 U4106 ( .A(\temp[25] ), .B(n13560), .C(n13561), .D(n13251), .Z(
        n13559) );
    VMW_OAI22 U4687 ( .A(n13621), .B(n13623), .C(n13619), .D(n13620), .Z(
        n14212) );
    VMW_AND3 U4203 ( .A(n13351), .B(n13686), .C(n13478), .Z(n13363) );
    VMW_INV U4236 ( .A(KEY[51]), .Z(n13724) );
    VMW_OAI22 U4717 ( .A(n13641), .B(n13716), .C(n13626), .D(n13715), .Z(
        n14227) );
    VMW_AO22 U5242 ( .A(n14023), .B(n13451), .C(X[31]), .D(Start), .Z(n14481)
         );
    VMW_INV U5453 ( .A(n13896), .Z(n14410) );
    VMW_XNOR2 U4427 ( .A(\temp[39] ), .B(n13164), .Z(n13987) );
    VMW_OR4 U4582 ( .A(n14142), .B(n14143), .C(n14140), .D(n14141), .Z(n13073)
         );
    VMW_OAI22 U4855 ( .A(n13619), .B(n14160), .C(n13616), .D(n14161), .Z(
        n13308) );
    VMW_OR4 U4860 ( .A(n14292), .B(n14293), .C(n14290), .D(n14291), .Z(n13290)
         );
    VMW_AO22 U5277 ( .A(n14069), .B(n13451), .C(X[61]), .D(Start), .Z(n14495)
         );
    VMW_INV U5466 ( .A(n13742), .Z(n13747) );
    VMW_NOR2 U4393 ( .A(n13897), .B(n13899), .Z(n13402) );
    VMW_AO22 U4412 ( .A(n13398), .B(n13966), .C(n13967), .D(n13402), .Z(n13965
        ) );
    VMW_NOR4 U3964 ( .A(n13073), .B(n13074), .C(n13075), .D(n13076), .Z(n13072
        ) );
    VMW_INV U4133 ( .A(KEY[38]), .Z(n13615) );
    VMW_OR3 U5147 ( .A(n14456), .B(n13456), .C(n14457), .Z(n13958) );
    VMW_OAI22 U4722 ( .A(n13640), .B(n14160), .C(n13637), .D(n14161), .Z(
        n13216) );
    VMW_AND2 U3981 ( .A(n13151), .B(n13152), .Z(n13150) );
    VMW_AOI211 U4028 ( .A(n13346), .B(n13347), .C(n13348), .D(n13343), .Z(
        n13345) );
    VMW_AO22 U4084 ( .A(n13479), .B(n13508), .C(\temp[19] ), .D(n13169), .Z(
        n13507) );
    VMW_NAND3 U5160 ( .A(n13584), .B(n13604), .C(n13324), .Z(n14388) );
    VMW_AO22 U4114 ( .A(n13579), .B(n13580), .C(\temp[10] ), .D(n13294), .Z(
        n13578) );
    VMW_AO22 U4705 ( .A(X[22]), .B(n13774), .C(n13773), .D(\temp[29] ), .Z(
        n13008) );
    VMW_INV U4224 ( .A(KEY[59]), .Z(n13713) );
    VMW_AND2 U4435 ( .A(n13549), .B(n13356), .Z(n13554) );
    VMW_OAI22 U4695 ( .A(n13623), .B(n13641), .C(n13620), .D(n13640), .Z(
        n14216) );
    VMW_OAI22 U4847 ( .A(n13635), .B(n14173), .C(n13631), .D(n14161), .Z(
        n13303) );
    VMW_AO22 U5250 ( .A(n14033), .B(n13598), .C(n14034), .D(n13443), .Z(n13951
        ) );
    VMW_INV U5441 ( .A(n13815), .Z(n13817) );
    VMW_NOR2 U4288 ( .A(n13437), .B(n13547), .Z(n13549) );
    VMW_OR4 U4509 ( .A(n14098), .B(n14099), .C(n14093), .D(n14095), .Z(n13064)
         );
    VMW_OR3 U4318 ( .A(n13280), .B(n13564), .C(n13808), .Z(n13810) );
    VMW_OAI22 U4499 ( .A(n13625), .B(n13626), .C(n13623), .D(n13624), .Z(
        n14087) );
    VMW_OAI22 U4639 ( .A(n13641), .B(n14160), .C(n13640), .D(n14161), .Z(
        n13117) );
    VMW_FD \temp_reg[35]  ( .D(\arr12639[35] ), .CP(Clk), .Q(\temp[35] ) );
    VMW_FD \OUT_reg[13]  ( .D(\arr12639[54] ), .CP(Clk), .Q(OUT[13]) );
    VMW_AND2 U4061 ( .A(n13443), .B(n13409), .Z(n13449) );
    VMW_OAI22 U4670 ( .A(n13633), .B(n14097), .C(n13609), .D(n14102), .Z(
        n14203) );
    VMW_FD \OUT_reg[39]  ( .D(\arr12639[59] ), .CP(Clk), .Q(OUT[39]) );
    VMW_FD \OUT_reg[20]  ( .D(\arr12639[21] ), .CP(Clk), .Q(OUT[20]) );
    VMW_AO22 U5185 ( .A(n13512), .B(n13505), .C(n13516), .D(n13525), .Z(n13341
        ) );
    VMW_NOR4 U4046 ( .A(n13416), .B(n13417), .C(n13418), .D(n13419), .Z(n13415
        ) );
    VMW_OAI21 U4351 ( .A(n13578), .B(n13841), .C(n13844), .Z(n13843) );
    VMW_OAI22 U4540 ( .A(n13621), .B(n13646), .C(n13619), .D(n14119), .Z(
        n14118) );
    VMW_OAI22 U4932 ( .A(n13626), .B(n14163), .C(n13641), .D(n14164), .Z(
        n14340) );
    VMW_NOR3 U5015 ( .A(n13654), .B(n14413), .C(n14414), .Z(n13675) );
    VMW_FD \OUT_reg[1]  ( .D(\arr12639[39] ), .CP(Clk), .Q(OUT[1]) );
    VMW_OR2 U4376 ( .A(n13443), .B(n13897), .Z(n13896) );
    VMW_AO22 U4885 ( .A(X[24]), .B(n13774), .C(\temp[4] ), .D(n13773), .Z(
        n13033) );
    VMW_INV U5325 ( .A(\temp[18] ), .Z(n13510) );
    VMW_OAI22 U4915 ( .A(n13633), .B(n14160), .C(n13609), .D(n14161), .Z(
        n13369) );
    VMW_OAI2222 U4567 ( .A(n13640), .B(n13645), .C(n13637), .D(n13648), .E(
        n13635), .F(n13647), .G(n13633), .H(n13646), .Z(n13089) );
    VMW_MUX2 U5292 ( .A(n14502), .B(\temp[10] ), .S(n13005), .Z(\arr12639[10] 
        ) );
    VMW_INV U5302 ( .A(\temp[30] ), .Z(n13468) );
    VMW_INV U5483 ( .A(n13706), .Z(n14313) );
    VMW_OR2 U4146 ( .A(n13608), .B(n13617), .Z(n13628) );
    VMW_OR4 U4657 ( .A(n14196), .B(n14197), .C(n14194), .D(n14195), .Z(n13190)
         );
    VMW_OR2 U4757 ( .A(n13537), .B(n13556), .Z(n13800) );
    VMW_AO22 U4829 ( .A(X[42]), .B(n13774), .C(\temp[10] ), .D(n13773), .Z(
        n13027) );
    VMW_AO21 U5032 ( .A(n13139), .B(n13144), .C(n13873), .Z(n14192) );
    VMW_FD \temp_reg[1]  ( .D(\arr12639[1] ), .CP(Clk), .Q(\temp[1] ) );
    VMW_AO21 U5129 ( .A(n13667), .B(n13662), .C(n14444), .Z(n13941) );
    VMW_MUX2 U5219 ( .A(n14470), .B(\temp[6] ), .S(n13005), .Z(\arr12639[6] )
         );
    VMW_INV U5389 ( .A(n13467), .Z(n13470) );
    VMW_INV U5408 ( .A(n13596), .Z(n13904) );
    VMW_AO22 U5132 ( .A(n13662), .B(n13663), .C(n13070), .D(n14360), .Z(n14446
        ) );
    VMW_AO21 U3953 ( .A(\temp[35] ), .B(n13005), .C(n13034), .Z(\arr12639[35] 
        ) );
    VMW_NOR4 U3958 ( .A(n13044), .B(n13045), .C(n13046), .D(n13047), .Z(n13043
        ) );
    VMW_NOR4 U4014 ( .A(n13295), .B(n13296), .C(n13297), .D(n13298), .Z(n13294
        ) );
    VMW_OR2 U4161 ( .A(n13607), .B(n13638), .Z(n13643) );
    VMW_AND2 U4251 ( .A(n13488), .B(n13493), .Z(n13141) );
    VMW_AND2 U4276 ( .A(n13507), .B(n13760), .Z(n13204) );
    VMW_AND2 U4467 ( .A(n13898), .B(n13913), .Z(n14039) );
    VMW_OAI22 U4815 ( .A(n13619), .B(n14090), .C(n13616), .D(n13639), .Z(
        n13244) );
    VMW_AND2 U4985 ( .A(n13447), .B(n14396), .Z(n13930) );
    VMW_OAI22 U4832 ( .A(n13633), .B(n14163), .C(n13644), .D(n14164), .Z(
        n14278) );
    VMW_OR2 U5202 ( .A(n13677), .B(n13660), .Z(n13969) );
    VMW_INV U5392 ( .A(n13493), .Z(n13148) );
    VMW_INV U5413 ( .A(n13667), .Z(n14048) );
    VMW_XOR2 U4440 ( .A(n13998), .B(\temp[37] ), .Z(n13997) );
    VMW_AO22 U5225 ( .A(n13999), .B(n13451), .C(X[25]), .D(Start), .Z(n14472)
         );
    VMW_INV U5434 ( .A(n13781), .Z(n13785) );
    VMW_OR2 U4324 ( .A(n13273), .B(n13803), .Z(n13814) );
    VMW_OAI22 U4770 ( .A(n13615), .B(n13619), .C(n13609), .D(n14096), .Z(
        n14250) );
    VMW_OAI2222 U4929 ( .A(n13616), .B(n13724), .C(n13644), .D(n13726), .E(
        n13642), .F(n13717), .G(n13641), .H(n13723), .Z(n13372) );
    VMW_NAND3 U5029 ( .A(n13425), .B(n13681), .C(n14419), .Z(n13705) );
    VMW_NAND4 U5085 ( .A(n14429), .B(n14428), .C(n14430), .D(n14307), .Z(
        n14016) );
    VMW_NAND4 U5115 ( .A(n13704), .B(n14440), .C(n13429), .D(n14324), .Z(
        n14030) );
    VMW_FD \OUT_reg[8]  ( .D(\arr12639[6] ), .CP(Clk), .Q(OUT[8]) );
    VMW_AO22 U5289 ( .A(n14078), .B(n13451), .C(X[35]), .D(Start), .Z(n14501)
         );
    VMW_INV U5319 ( .A(\temp[21] ), .Z(n13486) );
    VMW_OAI22 U4947 ( .A(n13644), .B(n14173), .C(n13643), .D(n14160), .Z(
        n13379) );
    VMW_INV U5350 ( .A(n13370), .Z(n13594) );
    VMW_FD \temp_reg[8]  ( .D(\arr12639[8] ), .CP(Clk), .Q(\temp[8] ) );
    VMW_OAI22 U4535 ( .A(n13632), .B(n13642), .C(n13618), .D(n13631), .Z(
        n13061) );
    VMW_NAND2 U5060 ( .A(n14275), .B(n13272), .Z(n13827) );
    VMW_AND3 U4033 ( .A(n13362), .B(n13363), .C(n13364), .Z(n13361) );
    VMW_NOR3 U4184 ( .A(n13459), .B(n13456), .C(n13470), .Z(n13664) );
    VMW_OAI22 U4795 ( .A(n13641), .B(n13646), .C(n13640), .D(n14119), .Z(
        n14263) );
    VMW_OAI2222 U4605 ( .A(n13644), .B(n13724), .C(n13641), .D(n13717), .E(
        n13640), .F(n13723), .G(n13637), .H(n13722), .Z(n13135) );
    VMW_OAI22 U4622 ( .A(n13635), .B(n13717), .C(n13633), .D(n13723), .Z(
        n13111) );
    VMW_NAND4 U5047 ( .A(n13769), .B(n13766), .C(n13771), .D(n14219), .Z(
        n13992) );
    VMW_OR2 U4128 ( .A(\i[3] ), .B(\i[2] ), .Z(n13608) );
    VMW_AND2 U4293 ( .A(n13356), .B(n13778), .Z(n13779) );
    VMW_OAI22 U4512 ( .A(n13619), .B(n14091), .C(n14090), .D(n13643), .Z(
        n13067) );
    VMW_OR3 U4960 ( .A(n14316), .B(n13159), .C(n14358), .Z(n13404) );
    VMW_INV U5377 ( .A(KEY[49]), .Z(n14172) );
    VMW_NAND2 U4303 ( .A(n13789), .B(n13790), .Z(n13788) );
    VMW_XOR2 U4482 ( .A(n14060), .B(\temp[52] ), .Z(n14059) );
    VMW_OAI22 U4739 ( .A(n13631), .B(n14163), .C(n13643), .D(n14164), .Z(
        n14237) );
    VMW_FD \temp_reg[16]  ( .D(\arr12639[16] ), .CP(Clk), .Q(\temp[16] ) );
    VMW_FD \OUT_reg[29]  ( .D(\arr12639[52] ), .CP(Clk), .Q(OUT[29]) );
    VMW_FD \OUT_reg[30]  ( .D(\arr12639[28] ), .CP(Clk), .Q(OUT[30]) );
    VMW_NOR4 U3974 ( .A(n13119), .B(n13120), .C(n13121), .D(n13122), .Z(n13118
        ) );
    VMW_AO22 U4094 ( .A(n13532), .B(n13533), .C(\temp[4] ), .D(n13227), .Z(
        n13531) );
    VMW_AO22 U4104 ( .A(n13554), .B(n13540), .C(n13555), .D(n13556), .Z(n13553
        ) );
    VMW_AO22 U4218 ( .A(n13360), .B(n13701), .C(n13702), .D(n13689), .Z(n13700
        ) );
    VMW_OAI211 U4599 ( .A(n14153), .B(n13694), .C(n13704), .D(n13709), .Z(
        n14152) );
    VMW_AND2 U4388 ( .A(n13907), .B(n13440), .Z(n13908) );
    VMW_NAND2 U4409 ( .A(n13958), .B(n13959), .Z(n13957) );
    VMW_FD \temp_reg[25]  ( .D(\arr12639[25] ), .CP(Clk), .Q(\temp[25] ) );
    VMW_OAI22 U4685 ( .A(n13643), .B(n13649), .C(n13631), .D(n14119), .Z(
        n14210) );
    VMW_OAI22 U4715 ( .A(n13643), .B(n14155), .C(n13631), .D(n14166), .Z(
        n14225) );
    VMW_NAND2 U5170 ( .A(n13908), .B(n13901), .Z(n14393) );
    VMW_AO22 U4123 ( .A(n13599), .B(n13600), .C(\temp[5] ), .D(n13375), .Z(
        n13598) );
    VMW_AND2 U4213 ( .A(n13691), .B(n13362), .Z(n13692) );
    VMW_INV U4234 ( .A(KEY[25]), .Z(n13722) );
    VMW_OAI22 U4857 ( .A(n13619), .B(n14166), .C(n13641), .D(n14167), .Z(
        n14291) );
    VMW_AND2 U4383 ( .A(n13440), .B(n13903), .Z(n13400) );
    VMW_NAND5 U4402 ( .A(n13936), .B(n13673), .C(n13937), .D(n13938), .E(
        n13939), .Z(n13935) );
    VMW_NAND2 U4425 ( .A(n13731), .B(n13156), .Z(n13985) );
    VMW_OAI22 U4870 ( .A(n13628), .B(n13726), .C(n13626), .D(n13718), .Z(
        n13297) );
    VMW_AO22 U5240 ( .A(n14021), .B(n13451), .C(X[23]), .D(Start), .Z(n14480)
         );
    VMW_INV U5451 ( .A(n13878), .Z(n13856) );
    VMW_OAI2222 U4592 ( .A(n13609), .B(n13625), .C(n13619), .D(n13649), .E(
        n13643), .F(n13645), .G(n13642), .H(n13648), .Z(n13084) );
    VMW_OAI22 U4732 ( .A(n13644), .B(n14169), .C(n13633), .D(n14167), .Z(
        n14234) );
    VMW_MUX2 U5267 ( .A(n14489), .B(\temp[20] ), .S(n13005), .Z(\arr12639[20] 
        ) );
    VMW_INV U5476 ( .A(n14368), .Z(n13961) );
    VMW_OAI21 U5157 ( .A(n13104), .B(n13690), .C(n13691), .Z(n14382) );
    VMW_NOR4 U3991 ( .A(n13190), .B(n13191), .C(n13192), .D(n13193), .Z(n13189
        ) );
    VMW_NOR4 U4038 ( .A(n13386), .B(n13387), .C(n13388), .D(n13389), .Z(n13385
        ) );
    VMW_AND2 U4298 ( .A(n13437), .B(n13547), .Z(n13238) );
    VMW_NOR2 U4308 ( .A(n13805), .B(n13557), .Z(n13282) );
    VMW_XOR2 U4489 ( .A(n14071), .B(\temp[47] ), .Z(n14070) );
    VMW_FD \temp_reg[34]  ( .D(\arr12639[34] ), .CP(Clk), .Q(\temp[34] ) );
    VMW_FD \OUT_reg[12]  ( .D(\arr12639[22] ), .CP(Clk), .Q(OUT[12]) );
    VMW_OAI22 U4519 ( .A(n13628), .B(n13634), .C(n13626), .D(n13632), .Z(
        n13041) );
    VMW_FD \OUT_reg[38]  ( .D(\arr12639[27] ), .CP(Clk), .Q(OUT[38]) );
    VMW_FD \OUT_reg[21]  ( .D(\arr12639[53] ), .CP(Clk), .Q(OUT[21]) );
    VMW_AND2 U4056 ( .A(\i6749[2] ), .B(n13445), .Z(n14507) );
    VMW_AO22 U4366 ( .A(n13337), .B(n13879), .C(n13833), .D(n13880), .Z(n13878
        ) );
    VMW_OAI22 U4577 ( .A(n13621), .B(n14092), .C(n13619), .D(n14089), .Z(
        n13096) );
    VMW_OAI2222 U4629 ( .A(n13624), .B(n13726), .C(n13621), .D(n13718), .E(
        n13643), .F(n13721), .G(n13642), .H(n13720), .Z(n13125) );
    VMW_NOR3 U4895 ( .A(n13435), .B(n13416), .C(n13960), .Z(n14307) );
    VMW_AOI211 U4905 ( .A(n13540), .B(n14323), .C(n13788), .D(n13588), .Z(
        n14322) );
    VMW_AO22 U5282 ( .A(n14073), .B(n13451), .C(X[11]), .D(Start), .Z(n14498)
         );
    VMW_INV U5312 ( .A(n13251), .Z(n13560) );
    VMW_INV U5493 ( .A(n14497), .Z(n14386) );
    VMW_OAI22 U4647 ( .A(n13609), .B(n14173), .C(n13628), .D(n14160), .Z(
        n13132) );
    VMW_AND3 U5022 ( .A(n13680), .B(n13686), .C(n13424), .Z(n14145) );
    VMW_AND2 U5005 ( .A(n14410), .B(n13409), .Z(n14409) );
    VMW_AO22 U4071 ( .A(n13476), .B(n13477), .C(\temp[20] ), .D(n13087), .Z(
        n13475) );
    VMW_INV U5195 ( .A(n13578), .Z(n13322) );
    VMW_FD \OUT_reg[0]  ( .D(\arr12639[7] ), .CP(Clk), .Q(OUT[0]) );
    VMW_INV U4171 ( .A(\temp[0] ), .Z(n13465) );
    VMW_INV U4241 ( .A(\temp[16] ), .Z(n13500) );
    VMW_AND2 U4341 ( .A(n13329), .B(n13334), .Z(n13324) );
    VMW_OAI22 U4660 ( .A(n13628), .B(n14091), .C(n13632), .D(n13643), .Z(
        n13193) );
    VMW_OAI22 U4922 ( .A(n13642), .B(n13724), .C(n13641), .D(n13726), .Z(
        n13393) );
    VMW_INV U5335 ( .A(\temp[13] ), .Z(n13494) );
    VMW_AND3 U4450 ( .A(n13206), .B(n13754), .C(n13756), .Z(n14012) );
    VMW_OR4 U4550 ( .A(n14126), .B(n14127), .C(n14124), .D(n14125), .Z(n13078)
         );
    VMW_AO22 U4822 ( .A(X[52]), .B(n13774), .C(n13773), .D(\temp[17] ), .Z(
        n13020) );
    VMW_OAI22 U4839 ( .A(n13616), .B(n14173), .C(n13643), .D(n14161), .Z(
        n13313) );
    VMW_AND4 U5139 ( .A(n13842), .B(n13333), .C(n13572), .D(n13328), .Z(n13948
        ) );
    VMW_MUX2 U5209 ( .A(n14465), .B(\temp[9] ), .S(n13005), .Z(\arr12639[9] )
         );
    VMW_INV U5399 ( .A(n13527), .Z(n14011) );
    VMW_INV U5418 ( .A(n14311), .Z(n13868) );
    VMW_FD \temp_reg[0]  ( .D(\arr12639[0] ), .CP(Clk), .Q(\temp[0] ) );
    VMW_AO22 U5235 ( .A(n14015), .B(n13451), .C(X[15]), .D(Start), .Z(n14477)
         );
    VMW_INV U5424 ( .A(n13142), .Z(n13750) );
    VMW_AO22 U4760 ( .A(X[46]), .B(n13774), .C(\temp[26] ), .D(n13773), .Z(
        n13011) );
    VMW_NAND2 U5095 ( .A(n13163), .B(n13141), .Z(n14433) );
    VMW_NAND3 U5105 ( .A(n13833), .B(n13335), .C(n13572), .Z(n14318) );
    VMW_FD \OUT_reg[9]  ( .D(\arr12639[38] ), .CP(Clk), .Q(OUT[9]) );
    VMW_AO21 U3927 ( .A(\temp[61] ), .B(n13005), .C(n13008), .Z(\arr12639[61] 
        ) );
    VMW_AO21 U3928 ( .A(\temp[60] ), .B(n13005), .C(n13009), .Z(\arr12639[60] 
        ) );
    VMW_AO21 U3934 ( .A(\temp[54] ), .B(n13005), .C(n13015), .Z(\arr12639[54] 
        ) );
    VMW_AO21 U3948 ( .A(\temp[40] ), .B(n13005), .C(n13029), .Z(\arr12639[40] 
        ) );
    VMW_NOR4 U4004 ( .A(n13252), .B(n13253), .C(n13254), .D(n13255), .Z(n13251
        ) );
    VMW_AND4 U4023 ( .A(n13333), .B(n13328), .C(n13334), .D(n13335), .Z(n13332
        ) );
    VMW_OR2 U4156 ( .A(n13614), .B(\i[2] ), .Z(n13638) );
    VMW_AO22 U5122 ( .A(n13901), .B(n13443), .C(n13408), .D(n14400), .Z(n14352
        ) );
    VMW_AND2 U4266 ( .A(n13754), .B(n13515), .Z(n13342) );
    VMW_OAI22 U4747 ( .A(n13643), .B(n14163), .C(n13628), .D(n14164), .Z(
        n14241) );
    VMW_OR4 U4805 ( .A(n14267), .B(n14268), .C(n14265), .D(n14266), .Z(n13247)
         );
    VMW_OR4 U4995 ( .A(n13654), .B(n13070), .C(n13453), .D(n14048), .Z(n14122)
         );
    VMW_AO22 U5212 ( .A(n13982), .B(n13451), .C(X[59]), .D(Start), .Z(n14466)
         );
    VMW_INV U5382 ( .A(KEY[17]), .Z(n14167) );
    VMW_INV U5403 ( .A(n13562), .Z(n13280) );
    VMW_XOR2 U4477 ( .A(n14054), .B(\temp[54] ), .Z(n14053) );
    VMW_OAI22 U4939 ( .A(n13642), .B(n14173), .C(n13631), .D(n13726), .Z(
        n13384) );
    VMW_AOI21 U5039 ( .A(n13730), .B(n13732), .C(n14408), .Z(n14193) );
    VMW_FD \temp_reg[9]  ( .D(\arr12639[9] ), .CP(Clk), .Q(\temp[9] ) );
    VMW_INV U5299 ( .A(n13232), .Z(n13534) );
    VMW_INV U5309 ( .A(n13246), .Z(n13568) );
    VMW_INV U5488 ( .A(n14467), .Z(n13752) );
    VMW_INV U4194 ( .A(\temp[23] ), .Z(n13484) );
    VMW_NOR2 U4283 ( .A(n13005), .B(n13451), .Z(n13774) );
    VMW_NAND2 U4313 ( .A(n13557), .B(n13805), .Z(n13284) );
    VMW_XOR2 U4492 ( .A(n14075), .B(\temp[45] ), .Z(n14074) );
    VMW_OAI22 U4632 ( .A(n13643), .B(n13714), .C(n13631), .D(n13713), .Z(
        n14182) );
    VMW_AO22 U4970 ( .A(n13818), .B(n13803), .C(n13816), .D(n13272), .Z(n14369
        ) );
    VMW_AO22 U5057 ( .A(n13344), .B(n13569), .C(n13277), .D(n13412), .Z(n13830
        ) );
    VMW_OAI2222 U4502 ( .A(n13639), .B(n13640), .C(n13636), .D(n13637), .E(
        n13634), .F(n13635), .G(n13632), .H(n13633), .Z(n13055) );
    VMW_OAI211 U4334 ( .A(n13284), .B(n13811), .C(n13827), .D(n13828), .Z(
        n13417) );
    VMW_OR4 U4525 ( .A(n14108), .B(n14109), .C(n14106), .D(n14107), .Z(n13044)
         );
    VMW_OR2 U4957 ( .A(n13396), .B(n13598), .Z(n13926) );
    VMW_INV U5367 ( .A(KEY[47]), .Z(n14097) );
    VMW_INV U5340 ( .A(n13289), .Z(n13585) );
    VMW_OAI22 U4615 ( .A(n13643), .B(n14173), .C(n13631), .D(n13718), .Z(
        n13122) );
    VMW_OAI22 U4785 ( .A(n13642), .B(n14103), .C(n13641), .D(n14112), .Z(
        n14257) );
    VMW_AO21 U5070 ( .A(n13575), .B(n13835), .C(n13842), .Z(n13335) );
    VMW_FD \temp_reg[17]  ( .D(\arr12639[17] ), .CP(Clk), .Q(\temp[17] ) );
    VMW_FD \OUT_reg[31]  ( .D(\arr12639[60] ), .CP(Clk), .Q(OUT[31]) );
    VMW_FD \OUT_reg[28]  ( .D(\arr12639[20] ), .CP(Clk), .Q(OUT[28]) );
    VMW_NOR4 U3998 ( .A(n13223), .B(n13224), .C(n13225), .D(n13226), .Z(n13222
        ) );
    VMW_NOR4 U4016 ( .A(n13305), .B(n13306), .C(n13307), .D(n13308), .Z(n13304
        ) );
    VMW_AND3 U4031 ( .A(n13355), .B(n13356), .C(n13357), .Z(n13354) );
    VMW_INV U4138 ( .A(KEY[6]), .Z(n13620) );
    VMW_OAI22 U4729 ( .A(n13609), .B(n14159), .C(n13619), .D(n13717), .Z(
        n13230) );
    VMW_AND2 U4208 ( .A(n13481), .B(n13364), .Z(n13689) );
    VMW_OAI21 U4398 ( .A(n13925), .B(n13926), .C(n13927), .Z(n13924) );
    VMW_AO21 U4419 ( .A(n13661), .B(n13664), .C(n13665), .Z(n13977) );
    VMW_FD \temp_reg[24]  ( .D(\arr12639[24] ), .CP(Clk), .Q(\temp[24] ) );
    VMW_OAI22 U4589 ( .A(n13637), .B(n14119), .C(n13631), .D(n14096), .Z(
        n14148) );
    VMW_OR4 U4620 ( .A(n14176), .B(n14177), .C(n14174), .D(n14175), .Z(n13109)
         );
    VMW_OAI22 U4879 ( .A(n13637), .B(n14160), .C(n13635), .D(n14161), .Z(
        n13318) );
    VMW_FD \temp_reg[4]  ( .D(\arr12639[4] ), .CP(Clk), .Q(\temp[4] ) );
    VMW_INV U5179 ( .A(n13488), .Z(n13157) );
    VMW_NOR2 U5249 ( .A(n13896), .B(n13911), .Z(n14032) );
    VMW_INV U5458 ( .A(n13676), .Z(n13939) );
    VMW_AND2 U4291 ( .A(n13540), .B(n13550), .Z(n13239) );
    VMW_OAI2222 U4510 ( .A(n13634), .B(n13640), .C(n13632), .D(n13637), .E(
        n13625), .F(n13631), .G(n13623), .H(n13628), .Z(n13065) );
    VMW_NAND3 U5045 ( .A(n13756), .B(n13528), .C(n13341), .Z(n13765) );
    VMW_FD \OUT_reg[4]  ( .D(\arr12639[23] ), .CP(Clk), .Q(OUT[4]) );
    VMW_NOR3 U4301 ( .A(n13546), .B(n13543), .C(n13589), .Z(n13786) );
    VMW_XNOR2 U4480 ( .A(n14057), .B(\temp[53] ), .Z(n14056) );
    VMW_NOR2 U4326 ( .A(n13817), .B(n13814), .Z(n13816) );
    VMW_NOR2 U4962 ( .A(n13459), .B(n13069), .Z(n14360) );
    VMW_INV U5375 ( .A(KEY[3]), .Z(n14161) );
    VMW_OAI22 U4537 ( .A(n13637), .B(n14112), .C(n13631), .D(n14094), .Z(
        n14115) );
    VMW_OAI2222 U4945 ( .A(n13640), .B(n13725), .C(n13637), .D(n13724), .E(
        n13635), .F(n13726), .G(n13633), .H(n13718), .Z(n13377) );
    VMW_INV U5352 ( .A(n13375), .Z(n13600) );
    VMW_AO22 U4078 ( .A(n13494), .B(n13495), .C(\temp[13] ), .D(n13133), .Z(
        n13493) );
    VMW_AO21 U4186 ( .A(n13459), .B(n13651), .C(n13071), .Z(n13667) );
    VMW_OR4 U4797 ( .A(n14263), .B(n14264), .C(n14261), .D(n14262), .Z(n13252)
         );
    VMW_NAND3 U4348 ( .A(n13581), .B(n13572), .C(n13331), .Z(n13841) );
    VMW_OAI2222 U4559 ( .A(n13609), .B(n13636), .C(n13624), .D(n13630), .E(
        n13621), .F(n13627), .G(n13619), .H(n13625), .Z(n13099) );
    VMW_OAI22 U4607 ( .A(n13624), .B(n14160), .C(n13621), .D(n14161), .Z(
        n13137) );
    VMW_AO21 U5062 ( .A(n13807), .B(n13347), .C(n14274), .Z(n13819) );
    VMW_OAI22 U4669 ( .A(n13619), .B(n14094), .C(n14085), .D(n13637), .Z(
        n14202) );
    VMW_FD \temp_reg[30]  ( .D(\arr12639[30] ), .CP(Clk), .Q(\temp[30] ) );
    VMW_FD \temp_reg[29]  ( .D(\arr12639[29] ), .CP(Clk), .Q(\temp[29] ) );
    VMW_FD \OUT_reg[16]  ( .D(\arr12639[5] ), .CP(Clk), .Q(OUT[16]) );
    VMW_INV U4163 ( .A(\temp[28] ), .Z(n13457) );
    VMW_NAND2 U4253 ( .A(n13139), .B(n13152), .Z(n13734) );
    VMW_AO22 U5227 ( .A(n14001), .B(n13572), .C(n14003), .D(n13334), .Z(n14302
        ) );
    VMW_FD \OUT_reg[25]  ( .D(\arr12639[36] ), .CP(Clk), .Q(OUT[25]) );
    VMW_INV U5436 ( .A(n13806), .Z(n13272) );
    VMW_AND2 U4442 ( .A(n13322), .B(n14002), .Z(n14001) );
    VMW_AO22 U4830 ( .A(X[50]), .B(n13774), .C(n13773), .D(\temp[9] ), .Z(
        n13028) );
    VMW_AND2 U5087 ( .A(n13104), .B(n13689), .Z(n13872) );
    VMW_NAND3 U5117 ( .A(n13408), .B(n13899), .C(n13906), .Z(n13923) );
    VMW_OAI22 U4772 ( .A(n13625), .B(n13628), .C(n13623), .D(n13626), .Z(
        n14252) );
    VMW_OR3 U5130 ( .A(n13654), .B(n13467), .C(n14445), .Z(n13936) );
    VMW_AO21 U3941 ( .A(\temp[47] ), .B(n13005), .C(n13022), .Z(\arr12639[47] 
        ) );
    VMW_NOR4 U3966 ( .A(n13083), .B(n13084), .C(n13085), .D(n13086), .Z(n13082
        ) );
    VMW_AND2 U3983 ( .A(n13156), .B(n13157), .Z(n13155) );
    VMW_AND3 U4044 ( .A(n13412), .B(n13288), .C(n13282), .Z(n13411) );
    VMW_OR2 U4144 ( .A(n13608), .B(n13611), .Z(n13626) );
    VMW_AOI21 U4755 ( .A(n13784), .B(n13776), .C(n14245), .Z(n13793) );
    VMW_NAND3 U4178 ( .A(n13659), .B(n13660), .C(n13651), .Z(n13658) );
    VMW_AND2 U4274 ( .A(n13758), .B(n13516), .Z(n13757) );
    VMW_NAND3 U4465 ( .A(n14035), .B(n14036), .C(n14037), .Z(n14034) );
    VMW_INV U5200 ( .A(n13598), .Z(n13443) );
    VMW_INV U5390 ( .A(n13481), .Z(n13686) );
    VMW_INV U5411 ( .A(n14061), .Z(n14490) );
    VMW_AO22 U4817 ( .A(n13818), .B(n13347), .C(n13816), .D(n13277), .Z(n13822
        ) );
    VMW_NAND2 U4987 ( .A(n13334), .B(n14398), .Z(n14319) );
    VMW_AND2 U4248 ( .A(n13496), .B(n13499), .Z(n13154) );
    VMW_OAI22 U4769 ( .A(n13644), .B(n14094), .C(n14085), .D(n13633), .Z(
        n14249) );
    VMW_FD \temp_reg[13]  ( .D(\arr12639[13] ), .CP(Clk), .Q(\temp[13] ) );
    VMW_FD \OUT_reg[35]  ( .D(\arr12639[43] ), .CP(Clk), .Q(OUT[35]) );
    VMW_NOR3 U4374 ( .A(n13358), .B(n13361), .C(n13895), .Z(n13429) );
    VMW_AND3 U4459 ( .A(n13535), .B(n13783), .C(n13355), .Z(n14025) );
    VMW_MUX2 U5290 ( .A(n14501), .B(\temp[11] ), .S(n13005), .Z(\arr12639[11] 
        ) );
    VMW_INV U5300 ( .A(n13048), .Z(n13463) );
    VMW_FD \temp_reg[39]  ( .D(\arr12639[39] ), .CP(Clk), .Q(\temp[39] ) );
    VMW_FD \temp_reg[20]  ( .D(\arr12639[20] ), .CP(Clk), .Q(\temp[20] ) );
    VMW_INV U5481 ( .A(n14151), .Z(n14420) );
    VMW_OAI22 U4565 ( .A(n13609), .B(n14119), .C(n13624), .D(n14096), .Z(
        n14135) );
    VMW_AO22 U4887 ( .A(X[40]), .B(n13774), .C(\temp[2] ), .D(n13773), .Z(
        n13035) );
    VMW_OAI22 U4917 ( .A(n13644), .B(n14170), .C(n13635), .D(n14167), .Z(
        n14333) );
    VMW_NAND3 U5030 ( .A(n13475), .B(n13683), .C(n13104), .Z(n13707) );
    VMW_OAI22 U4655 ( .A(n13640), .B(n14097), .C(n13637), .D(n14102), .Z(
        n14196) );
    VMW_INV U5187 ( .A(n13537), .Z(n13546) );
    VMW_AO22 U4063 ( .A(n13454), .B(n13455), .C(\temp[29] ), .D(n13038), .Z(
        n13453) );
    VMW_OAI22 U4672 ( .A(n13615), .B(n13624), .C(n13616), .D(n13645), .Z(
        n14205) );
    VMW_NAND3 U5017 ( .A(n14048), .B(n13661), .C(n13668), .Z(n14121) );
    VMW_AO22 U4086 ( .A(n13476), .B(n13513), .C(\temp[20] ), .D(n13174), .Z(
        n13512) );
    VMW_NOR2 U4353 ( .A(n13850), .B(n13851), .Z(n13849) );
    VMW_OAI2222 U4542 ( .A(n13635), .B(n13649), .C(n13628), .D(n13645), .E(
        n13626), .F(n13648), .G(n13624), .H(n13647), .Z(n13050) );
    VMW_INV U5327 ( .A(\temp[17] ), .Z(n13518) );
    VMW_OAI22 U4930 ( .A(n13621), .B(n14159), .C(n13619), .D(n13725), .Z(
        n13373) );
    VMW_AO22 U4979 ( .A(n13346), .B(n13814), .C(n14386), .D(n13809), .Z(n13433
        ) );
    VMW_AND4 U5079 ( .A(n13507), .B(n13205), .C(n13512), .D(n13515), .Z(n14009
        ) );
    VMW_INV U5349 ( .A(\temp[6] ), .Z(n13593) );
    VMW_AO22 U4116 ( .A(n13489), .B(n13585), .C(\temp[11] ), .D(n13289), .Z(
        n13584) );
    VMW_OAI22 U4707 ( .A(n13640), .B(n14163), .C(n13621), .D(n14164), .Z(
        n14221) );
    VMW_OR4 U4697 ( .A(n14216), .B(n14217), .C(n14214), .D(n14215), .Z(n13175)
         );
    VMW_NAND2 U4131 ( .A(\i[1] ), .B(n13612), .Z(n13611) );
    VMW_AND2 U4201 ( .A(n13351), .B(n13682), .Z(n13685) );
    VMW_INV U4226 ( .A(KEY[44]), .Z(n13715) );
    VMW_OAI22 U4437 ( .A(n13994), .B(n13546), .C(n13778), .D(n13537), .Z(
        n13993) );
    VMW_NAND4 U5162 ( .A(n13849), .B(n14459), .C(n13947), .D(n14387), .Z(
        n14075) );
    VMW_OAI22 U4580 ( .A(n13624), .B(n13646), .C(n13621), .D(n14119), .Z(
        n14142) );
    VMW_OAI2222 U4845 ( .A(n13624), .B(n13724), .C(n13621), .D(n13726), .E(
        n13619), .F(n13718), .G(n13643), .H(n13722), .Z(n13301) );
    VMW_AO22 U5252 ( .A(n14043), .B(n13451), .C(X[55]), .D(Start), .Z(n14484)
         );
    VMW_INV U5443 ( .A(n13836), .Z(n13879) );
    VMW_AND2 U4391 ( .A(n13911), .B(n13912), .Z(n13410) );
    VMW_OR4 U4410 ( .A(n13829), .B(n13823), .C(n13960), .D(n13961), .Z(n13418)
         );
    VMW_OAI22 U4862 ( .A(n13631), .B(n13727), .C(n13609), .D(n13716), .Z(
        n13292) );
    VMW_AO22 U5275 ( .A(n14067), .B(n13451), .C(X[53]), .D(Start), .Z(n14494)
         );
    VMW_INV U5464 ( .A(n14412), .Z(n14403) );
    VMW_OAI2222 U4720 ( .A(n13609), .B(n13724), .C(n13624), .D(n13717), .E(
        n13621), .F(n13723), .G(n13619), .H(n13722), .Z(n13214) );
    VMW_AO21 U3946 ( .A(\temp[42] ), .B(n13005), .C(n13027), .Z(\arr12639[42] 
        ) );
    VMW_OAI22 U4959 ( .A(n13728), .B(n13749), .C(n13728), .D(n13734), .Z(
        n14358) );
    VMW_NAND3 U5059 ( .A(n13282), .B(n13814), .C(n13274), .Z(n13828) );
    VMW_NAND5 U5145 ( .A(n14453), .B(n14357), .C(n13914), .D(n14454), .E(
        n14455), .Z(n14060) );
    VMW_INV U5369 ( .A(KEY[14]), .Z(n14103) );
    VMW_NOR4 U3961 ( .A(n13059), .B(n13060), .C(n13061), .D(n13062), .Z(n13058
        ) );
    VMW_INV U4136 ( .A(KEY[22]), .Z(n13618) );
    VMW_OR4 U4727 ( .A(n14231), .B(n14232), .C(n14229), .D(n14230), .Z(n13228)
         );
    VMW_AND3 U5142 ( .A(n13603), .B(n13904), .C(n13905), .Z(n14452) );
    VMW_AND2 U4206 ( .A(n13686), .B(n13362), .Z(n13425) );
    VMW_NAND3 U4396 ( .A(n13916), .B(n13914), .C(n13919), .Z(n13918) );
    VMW_OAI22 U4865 ( .A(n13633), .B(n14166), .C(n13621), .D(n14167), .Z(
        n14295) );
    VMW_MUX2 U5272 ( .A(n14492), .B(\temp[19] ), .S(n13005), .Z(\arr12639[19] 
        ) );
    VMW_INV U5463 ( .A(n13954), .Z(n14454) );
    VMW_OR2 U4417 ( .A(n13459), .B(n13070), .Z(n13975) );
    VMW_AOI211 U4221 ( .A(n13681), .B(n13693), .C(n13710), .D(n13711), .Z(
        n13709) );
    VMW_OAI22 U4587 ( .A(n13624), .B(n14103), .C(n13621), .D(n14112), .Z(
        n14146) );
    VMW_OAI22 U4842 ( .A(n13640), .B(n13719), .C(n13637), .D(n13727), .Z(
        n14284) );
    VMW_AO22 U5255 ( .A(n14045), .B(n13451), .C(X[63]), .D(Start), .Z(n14485)
         );
    VMW_INV U5444 ( .A(n13834), .Z(n13880) );
    VMW_AND2 U4430 ( .A(n13516), .B(n13507), .Z(n13523) );
    VMW_AO22 U4081 ( .A(n13502), .B(n13503), .C(\temp[12] ), .D(n13123), .Z(
        n13139) );
    VMW_AO22 U4111 ( .A(n13502), .B(n13571), .C(\temp[12] ), .D(n13309), .Z(
        n13329) );
    VMW_OAI2222 U4690 ( .A(n13635), .B(n13636), .C(n13633), .D(n13634), .E(
        n13609), .F(n13632), .G(n13628), .H(n13630), .Z(n13181) );
    VMW_OR4 U5165 ( .A(n14246), .B(n13891), .C(n13962), .D(n14463), .Z(n14079)
         );
    VMW_OAI22 U4700 ( .A(n13633), .B(n14091), .C(n13631), .D(n14092), .Z(
        n13178) );
    VMW_FD \temp_reg[11]  ( .D(\arr12639[11] ), .CP(Clk), .Q(\temp[11] ) );
    VMW_FD \OUT_reg[37]  ( .D(\arr12639[51] ), .CP(Clk), .Q(OUT[37]) );
    VMW_AO21 U3929 ( .A(\temp[59] ), .B(n13005), .C(n13010), .Z(\arr12639[59] 
        ) );
    VMW_AO21 U3932 ( .A(\temp[56] ), .B(n13005), .C(n13013), .Z(\arr12639[56] 
        ) );
    VMW_AO21 U3933 ( .A(\temp[55] ), .B(n13005), .C(n13014), .Z(\arr12639[55] 
        ) );
    VMW_AOI211 U3984 ( .A(n13143), .B(n13140), .C(n13145), .D(n13159), .Z(
        n13158) );
    VMW_AO22 U4064 ( .A(n13457), .B(n13458), .C(\temp[28] ), .D(n13053), .Z(
        n13456) );
    VMW_OR2 U4158 ( .A(n13622), .B(n13638), .Z(n13640) );
    VMW_NOR2 U4268 ( .A(n13200), .B(n13507), .Z(n13755) );
    VMW_OAI22 U4749 ( .A(n13626), .B(n14169), .C(n13624), .D(n14170), .Z(
        n14243) );
    VMW_FD \temp_reg[22]  ( .D(\arr12639[22] ), .CP(Clk), .Q(\temp[22] ) );
    VMW_OAI211 U4354 ( .A(n13322), .B(n13838), .C(n13853), .D(n13854), .Z(
        n13852) );
    VMW_AO22 U4479 ( .A(n13832), .B(n13880), .C(n13833), .D(n13879), .Z(n14055
        ) );
    VMW_OAI2222 U4937 ( .A(n13609), .B(n13715), .C(n13644), .D(n13714), .E(
        n13633), .F(n13713), .G(n13621), .H(n13712), .Z(n13382) );
    VMW_NAND3 U4545 ( .A(n14121), .B(n14122), .C(n14123), .Z(n14120) );
    VMW_INV U5320 ( .A(n13082), .Z(n13487) );
    VMW_OAI22 U4675 ( .A(n13636), .B(n13642), .C(n13634), .D(n13641), .Z(
        n13172) );
    VMW_AND2 U5010 ( .A(n13402), .B(n13906), .Z(n13952) );
    VMW_INV U5180 ( .A(n13447), .Z(n13161) );
    VMW_AND3 U4043 ( .A(n13408), .B(n13409), .C(n13410), .Z(n13407) );
    VMW_OAI211 U4652 ( .A(n13728), .B(n14193), .C(n13746), .D(n13160), .Z(
        n13168) );
    VMW_AND2 U4058 ( .A(\i6749[0] ), .B(n13445), .Z(n14509) );
    VMW_OAI21 U4368 ( .A(n13883), .B(n13884), .C(n13885), .Z(n13882) );
    VMW_AND2 U4373 ( .A(n13690), .B(n13683), .Z(n13894) );
    VMW_OAI22 U4562 ( .A(n13641), .B(n14094), .C(n14085), .D(n13626), .Z(
        n14132) );
    VMW_AOI211 U4880 ( .A(n13839), .B(n13328), .C(n13843), .D(n14302), .Z(
        n13848) );
    VMW_OAI22 U4910 ( .A(n13640), .B(n14155), .C(n13628), .D(n14169), .Z(
        n14330) );
    VMW_AO22 U5037 ( .A(n13488), .B(n13731), .C(n13152), .D(n13161), .Z(n14190
        ) );
    VMW_OAI22 U4579 ( .A(n13643), .B(n14097), .C(n13642), .D(n14102), .Z(
        n14141) );
    VMW_INV U5297 ( .A(\i[0] ), .Z(n13612) );
    VMW_INV U5307 ( .A(n13261), .Z(n13563) );
    VMW_INV U5486 ( .A(n14464), .Z(n13670) );
    VMW_FD \temp_reg[32]  ( .D(\arr12639[32] ), .CP(Clk), .Q(\temp[32] ) );
    VMW_FD \OUT_reg[14]  ( .D(\arr12639[30] ), .CP(Clk), .Q(OUT[14]) );
    VMW_AOI211 U4649 ( .A(n14190), .B(n13151), .C(n14191), .D(n13737), .Z(
        n13748) );
    VMW_FD \temp_reg[18]  ( .D(\arr12639[18] ), .CP(Clk), .Q(\temp[18] ) );
    VMW_FD \OUT_reg[27]  ( .D(\arr12639[44] ), .CP(Clk), .Q(OUT[27]) );
    VMW_INV U4143 ( .A(KEY[39]), .Z(n13625) );
    VMW_AND3 U4273 ( .A(n13505), .B(n13515), .C(n13517), .Z(n13530) );
    VMW_OAI22 U4810 ( .A(n13643), .B(n13646), .C(n13642), .D(n14119), .Z(
        n14270) );
    VMW_AND3 U4980 ( .A(n13847), .B(n14319), .C(n14388), .Z(n14387) );
    VMW_XOR2 U4462 ( .A(n14030), .B(\temp[58] ), .Z(n14029) );
    VMW_OAI22 U5207 ( .A(n13663), .B(n13471), .C(n13652), .D(n13464), .Z(
        n14414) );
    VMW_INV U5397 ( .A(n13514), .Z(n13206) );
    VMW_INV U5416 ( .A(n13363), .Z(n13106) );
    VMW_OAI2222 U4752 ( .A(n13616), .B(n13715), .C(n13635), .D(n13714), .E(
        n13619), .F(n13713), .G(n13641), .H(n13712), .Z(n13209) );
    VMW_NAND3 U5137 ( .A(n13507), .B(n14447), .C(n13206), .Z(n14448) );
    VMW_AO21 U3954 ( .A(\temp[34] ), .B(n13005), .C(n13035), .Z(\arr12639[34] 
        ) );
    VMW_NOR4 U3968 ( .A(n13093), .B(n13094), .C(n13095), .D(n13096), .Z(n13092
        ) );
    VMW_NOR4 U4003 ( .A(n13247), .B(n13248), .C(n13249), .D(n13250), .Z(n13246
        ) );
    VMW_NOR2 U4011 ( .A(n13284), .B(n13285), .Z(n13283) );
    VMW_INV U4164 ( .A(KEY[21]), .Z(n13645) );
    VMW_OAI22 U4775 ( .A(n14090), .B(n13642), .C(n13639), .D(n13641), .Z(
        n13264) );
    VMW_AND2 U4181 ( .A(n13069), .B(n13471), .Z(n13662) );
    VMW_NAND2 U4254 ( .A(n13156), .B(n13144), .Z(n13735) );
    VMW_AND2 U4445 ( .A(n13835), .B(n13572), .Z(n13587) );
    VMW_OAI2222 U4837 ( .A(n13640), .B(n13724), .C(n13637), .D(n13726), .E(
        n13635), .F(n13718), .G(n13631), .H(n13723), .Z(n13311) );
    VMW_NAND4 U5080 ( .A(n14427), .B(n13771), .C(n13858), .D(n14305), .Z(
        n14014) );
    VMW_AO21 U5110 ( .A(n13535), .B(n13357), .C(n13780), .Z(n14323) );
    VMW_OAI22 U4600 ( .A(n13643), .B(n13713), .C(n13631), .D(n14155), .Z(
        n14154) );
    VMW_OAI22 U4859 ( .A(n13637), .B(n14172), .C(n13635), .D(n14155), .Z(
        n14293) );
    VMW_AO22 U5220 ( .A(n13995), .B(n13535), .C(n13420), .D(n13356), .Z(n14246
        ) );
    VMW_INV U5431 ( .A(n13777), .Z(n13994) );
    VMW_FD \temp_reg[6]  ( .D(\arr12639[6] ), .CP(Clk), .Q(\temp[6] ) );
    VMW_AO21 U5065 ( .A(n13277), .B(n13815), .C(n13818), .Z(n14277) );
    VMW_OR4 U5159 ( .A(n13674), .B(n13935), .C(n13957), .D(n14383), .Z(n14071)
         );
    VMW_AO22 U5269 ( .A(n14062), .B(n13451), .C(X[49]), .D(Start), .Z(n14491)
         );
    VMW_INV U5478 ( .A(n14389), .Z(n14463) );
    VMW_FD \OUT_reg[6]  ( .D(\arr12639[31] ), .CP(Clk), .Q(OUT[6]) );
    VMW_OAI2222 U4790 ( .A(n13621), .B(n13630), .C(n13619), .D(n13627), .E(
        n13616), .F(n13625), .G(n13623), .H(n13644), .Z(n13258) );
    VMW_NOR4 U4036 ( .A(n13376), .B(n13377), .C(n13378), .D(n13379), .Z(n13375
        ) );
    VMW_NOR2 U4296 ( .A(n13546), .B(n13540), .Z(n13355) );
    VMW_OAI211 U4306 ( .A(n13799), .B(n13800), .C(n13801), .D(n13802), .Z(
        n13798) );
    VMW_AND3 U4321 ( .A(n13569), .B(n13564), .C(n13567), .Z(n13812) );
    VMW_OAI22 U4530 ( .A(n13633), .B(n14103), .C(n13609), .D(n14112), .Z(
        n14111) );
    VMW_OAI22 U4942 ( .A(n13626), .B(n13722), .C(n13624), .D(n13721), .Z(
        n14346) );
    VMW_INV U5355 ( .A(n13207), .Z(n13545) );
    VMW_AND2 U4965 ( .A(n14363), .B(n13202), .Z(n13946) );
    VMW_INV U5372 ( .A(KEY[15]), .Z(n14085) );
    VMW_XOR2 U4487 ( .A(n14068), .B(\temp[49] ), .Z(n14067) );
    VMW_OR4 U4517 ( .A(n14104), .B(n14105), .C(n14100), .D(n14101), .Z(n13039)
         );
    VMW_AND3 U5042 ( .A(n13201), .B(n13760), .C(n13202), .Z(n13770) );
    VMW_OAI22 U4627 ( .A(n13641), .B(n13719), .C(n13640), .D(n13727), .Z(
        n14181) );
    VMW_OAI2222 U4782 ( .A(n13626), .B(n13645), .C(n13624), .D(n13648), .E(
        n13621), .F(n13647), .G(n13619), .H(n13646), .Z(n13268) );
    VMW_OAI211 U5077 ( .A(n13326), .B(n13330), .C(n13334), .D(n13320), .Z(
        n13846) );
    VMW_AND3 U4024 ( .A(n13337), .B(n13321), .C(n13322), .Z(n13336) );
    VMW_INV U4193 ( .A(\temp[19] ), .Z(n13479) );
    VMW_OR4 U4612 ( .A(n14168), .B(n14171), .C(n14162), .D(n14165), .Z(n13119)
         );
    VMW_INV U4284 ( .A(\temp[4] ), .Z(n13532) );
    VMW_OR4 U4333 ( .A(n13821), .B(n13432), .C(n13823), .D(n13826), .Z(n13825)
         );
    VMW_INV U5347 ( .A(n13314), .Z(n13583) );
    VMW_OAI22 U4522 ( .A(n13620), .B(n13637), .C(n13618), .D(n13635), .Z(
        n14107) );
    VMW_OAI22 U4950 ( .A(n13635), .B(n14169), .C(n13633), .D(n14170), .Z(
        n14350) );
    VMW_INV U5360 ( .A(n13217), .Z(n13542) );
    VMW_AND2 U4314 ( .A(n13557), .B(n13559), .Z(n13414) );
    VMW_OAI22 U4505 ( .A(n13616), .B(n14094), .C(n14085), .D(n13635), .Z(
        n14093) );
    VMW_XOR2 U4495 ( .A(n14081), .B(\temp[42] ), .Z(n14080) );
    VMW_OAI22 U4635 ( .A(n13621), .B(n13722), .C(n13619), .D(n13721), .Z(
        n14185) );
    VMW_AND3 U4977 ( .A(n14380), .B(n14381), .C(n14382), .Z(n13430) );
    VMW_AO22 U5050 ( .A(n13553), .B(n13537), .C(n13556), .D(n13775), .Z(n14402
        ) );
    VMW_AO22 U4088 ( .A(n13518), .B(n13519), .C(\temp[17] ), .D(n13184), .Z(
        n13517) );
    VMW_OAI22 U4709 ( .A(n13619), .B(n14169), .C(n13616), .D(n14170), .Z(
        n14223) );
    VMW_AOI211 U4118 ( .A(n13589), .B(n13590), .C(n13591), .D(n13537), .Z(
        n13588) );
    VMW_OAI22 U4699 ( .A(n13628), .B(n14089), .C(n13626), .D(n14090), .Z(
        n13177) );
    VMW_NOR4 U3996 ( .A(n13213), .B(n13214), .C(n13215), .D(n13216), .Z(n13212
        ) );
    VMW_AO22 U4076 ( .A(n13489), .B(n13490), .C(\temp[11] ), .D(n13118), .Z(
        n13488) );
    VMW_OR2 U4151 ( .A(n13611), .B(n13629), .Z(n13633) );
    VMW_INV U4228 ( .A(KEY[60]), .Z(n13717) );
    VMW_AND2 U4439 ( .A(n13355), .B(n13779), .Z(n13996) );
    VMW_FD \temp_reg[15]  ( .D(\arr12639[15] ), .CP(Clk), .Q(\temp[15] ) );
    VMW_FD \OUT_reg[33]  ( .D(\arr12639[35] ), .CP(Clk), .Q(OUT[33]) );
    VMW_AND3 U4261 ( .A(n13739), .B(n13747), .C(n13748), .Z(n13746) );
    VMW_XOR2 U4470 ( .A(n14044), .B(\temp[57] ), .Z(n14043) );
    VMW_FD \temp_reg[26]  ( .D(\arr12639[26] ), .CP(Clk), .Q(\temp[26] ) );
    VMW_FD \OUT_reg[19]  ( .D(\arr12639[45] ), .CP(Clk), .Q(OUT[19]) );
    VMW_OAI22 U4740 ( .A(n13640), .B(n14166), .C(n13628), .D(n14167), .Z(
        n14238) );
    VMW_OAI22 U4802 ( .A(n13619), .B(n14103), .C(n13616), .D(n14112), .Z(
        n14266) );
    VMW_AND3 U4992 ( .A(n13548), .B(n13556), .C(n14401), .Z(n14245) );
    VMW_AO22 U5215 ( .A(n13987), .B(n13451), .C(X[1]), .D(Start), .Z(n14468)
         );
    VMW_INV U5385 ( .A(\temp[25] ), .Z(n13561) );
    VMW_INV U5404 ( .A(n13567), .Z(n13808) );
    VMW_AND2 U4176 ( .A(n13069), .B(n13464), .Z(n13656) );
    VMW_OR4 U5125 ( .A(n13918), .B(n13920), .C(n13924), .D(n14353), .Z(n14044)
         );
    VMW_NOR2 U4246 ( .A(n13161), .B(n13493), .Z(n13731) );
    VMW_AO22 U4767 ( .A(X[36]), .B(n13774), .C(n13773), .D(\temp[19] ), .Z(
        n13018) );
    VMW_NAND3 U5092 ( .A(n13732), .B(n13730), .C(n13140), .Z(n13877) );
    VMW_AO21 U5102 ( .A(n13335), .B(n13325), .C(n14438), .Z(n14437) );
    VMW_NOR2 U4346 ( .A(n13836), .B(n13840), .Z(n13839) );
    VMW_XOR2 U4457 ( .A(n14022), .B(\temp[61] ), .Z(n14021) );
    VMW_OAI22 U4557 ( .A(n13616), .B(n13623), .C(n13620), .D(n13644), .Z(
        n14131) );
    VMW_AO22 U4825 ( .A(X[10]), .B(n13774), .C(n13773), .D(\temp[14] ), .Z(
        n13023) );
    VMW_AO22 U4889 ( .A(X[56]), .B(n13774), .C(n13773), .D(\temp[0] ), .Z(
        n13037) );
    VMW_AO22 U5232 ( .A(n14012), .B(n13505), .C(n14010), .D(n13525), .Z(n14475
        ) );
    VMW_INV U5423 ( .A(n13734), .Z(n13143) );
    VMW_OAI22 U4919 ( .A(n13624), .B(n13727), .C(n13633), .D(n13712), .Z(
        n14335) );
    VMW_OR4 U5019 ( .A(n13674), .B(n13669), .C(n13676), .D(n14120), .Z(n13979)
         );
    VMW_INV U5189 ( .A(n13535), .Z(n13356) );
    VMW_INV U5329 ( .A(n13128), .Z(n13501) );
    VMW_OAI22 U4667 ( .A(n13609), .B(n13627), .C(n13616), .D(n13649), .Z(
        n13197) );
    VMW_OAI22 U4925 ( .A(n13609), .B(n13727), .C(n13628), .D(n13716), .Z(
        n14337) );
    VMW_INV U5332 ( .A(n13194), .Z(n13504) );
    VMW_AND4 U4051 ( .A(n13437), .B(n13239), .C(n13438), .D(n13356), .Z(n13436
        ) );
    VMW_NAND3 U5002 ( .A(n13900), .B(n13897), .C(n13902), .Z(n14036) );
    VMW_INV U5192 ( .A(n13329), .Z(n13835) );
    VMW_NOR2 U4361 ( .A(n13867), .B(n13868), .Z(n13427) );
    VMW_OAI22 U4640 ( .A(n13633), .B(n13727), .C(n13631), .D(n13716), .Z(
        n14186) );
    VMW_AO22 U5025 ( .A(n13472), .B(n13363), .C(n13424), .D(n13683), .Z(n13701
        ) );
    VMW_FD \OUT_reg[2]  ( .D(\arr12639[15] ), .CP(Clk), .Q(OUT[2]) );
    VMW_OAI22 U4570 ( .A(n13628), .B(n14103), .C(n13626), .D(n14112), .Z(
        n14136) );
    VMW_AOI211 U4819 ( .A(n14274), .B(n13414), .C(n13279), .D(n13283), .Z(
        n14273) );
    VMW_AND2 U4892 ( .A(n13277), .B(n13814), .Z(n13862) );
    VMW_NAND3 U4902 ( .A(n14318), .B(n14319), .C(n14320), .Z(n14317) );
    VMW_AO22 U5089 ( .A(n13359), .B(n13681), .C(n13685), .D(n14431), .Z(n13865
        ) );
    VMW_AO21 U5119 ( .A(n13897), .B(n13899), .C(n13402), .Z(n14441) );
    VMW_AO22 U5229 ( .A(n14005), .B(n13451), .C(X[33]), .D(Start), .Z(n14473)
         );
    VMW_MUX2 U5285 ( .A(n14499), .B(\temp[13] ), .S(n13005), .Z(\arr12639[13] 
        ) );
    VMW_INV U5315 ( .A(n13072), .Z(n13485) );
    VMW_INV U5494 ( .A(n13341), .Z(n14461) );
    VMW_INV U5438 ( .A(n13275), .Z(n13434) );
    VMW_FD \temp_reg[2]  ( .D(\arr12639[2] ), .CP(Clk), .Q(\temp[2] ) );
    VMW_AND3 U4989 ( .A(n13758), .B(n14363), .C(n14011), .Z(n14220) );
    VMW_NAND3 U5150 ( .A(n13730), .B(n13161), .C(n13873), .Z(n14374) );
    VMW_NOR4 U3973 ( .A(n13114), .B(n13115), .C(n13116), .D(n13117), .Z(n13113
        ) );
    VMW_AO22 U4124 ( .A(n13532), .B(n13601), .C(\temp[4] ), .D(n13390), .Z(
        n13440) );
    VMW_AND2 U4214 ( .A(n13692), .B(n13478), .Z(n13693) );
    VMW_OR4 U4735 ( .A(n14235), .B(n14236), .C(n14233), .D(n14234), .Z(n13223)
         );
    VMW_MUX2 U5260 ( .A(n14486), .B(\temp[23] ), .S(n13005), .Z(\arr12639[23] 
        ) );
    VMW_INV U5471 ( .A(n14273), .Z(n13826) );
    VMW_INV U4233 ( .A(KEY[41]), .Z(n13721) );
    VMW_AND2 U4384 ( .A(n13396), .B(n13441), .Z(n13905) );
    VMW_NAND2 U4595 ( .A(n13103), .B(n13353), .Z(n13699) );
    VMW_AO22 U4405 ( .A(n13524), .B(n13945), .C(n13946), .D(n13757), .Z(n13944
        ) );
    VMW_AO22 U4422 ( .A(n13690), .B(n13475), .C(n13104), .D(n13353), .Z(n13981
        ) );
    VMW_OAI2222 U4877 ( .A(n13621), .B(n13717), .C(n13619), .D(n13723), .E(
        n13616), .F(n13722), .G(n13644), .H(n13721), .Z(n13316) );
    VMW_AO22 U5247 ( .A(n14029), .B(n13451), .C(X[47]), .D(Start), .Z(n14483)
         );
    VMW_INV U5456 ( .A(n13410), .Z(n14400) );
    VMW_OAI22 U4850 ( .A(n13641), .B(n13713), .C(n13631), .D(n13712), .Z(
        n14288) );
    VMW_INV U5177 ( .A(n13362), .Z(n13688) );
    VMW_AND3 U4010 ( .A(n13280), .B(n13281), .C(n13282), .Z(n13279) );
    VMW_NOR4 U4018 ( .A(n13315), .B(n13316), .C(n13317), .D(n13318), .Z(n13314
        ) );
    VMW_AO22 U4093 ( .A(n13529), .B(n13512), .C(n13530), .D(n13516), .Z(n13339
        ) );
    VMW_OAI2222 U4712 ( .A(n13631), .B(n13720), .C(n13628), .D(n13719), .E(
        n13626), .F(n13727), .G(n13635), .H(n13712), .Z(n13219) );
    VMW_AO22 U4103 ( .A(n13552), .B(n13356), .C(n13355), .D(n13535), .Z(n13551
        ) );
    VMW_OAI2222 U4682 ( .A(n13624), .B(n13634), .C(n13621), .D(n13632), .E(
        n13623), .F(n13643), .G(n13620), .H(n13642), .Z(n13186) );
    VMW_AND2 U4328 ( .A(n13562), .B(n13344), .Z(n13818) );
    VMW_OAI22 U4539 ( .A(n13643), .B(n14096), .C(n13642), .D(n14097), .Z(
        n14117) );
    VMW_OAI22 U4799 ( .A(n14090), .B(n13644), .C(n13630), .D(n13637), .Z(
        n13254) );
    VMW_FD \temp_reg[36]  ( .D(\arr12639[36] ), .CP(Clk), .Q(\temp[36] ) );
    VMW_FD \OUT_reg[10]  ( .D(\arr12639[14] ), .CP(Clk), .Q(OUT[10]) );
    VMW_NAND4 U4188 ( .A(n13670), .B(n13671), .C(n13672), .D(n13673), .Z(
        n13669) );
    VMW_OAI22 U4609 ( .A(n13637), .B(n14166), .C(n13626), .D(n14167), .Z(
        n14165) );
    VMW_OAI22 U4858 ( .A(n13624), .B(n14169), .C(n13621), .D(n14170), .Z(
        n14292) );
    VMW_FD \OUT_reg[23]  ( .D(\arr12639[61] ), .CP(Clk), .Q(OUT[23]) );
    VMW_OAI21 U5158 ( .A(n13657), .B(n14411), .C(n13661), .Z(n14385) );
    VMW_OAI22 U5268 ( .A(n14490), .B(n13659), .C(n13655), .D(n13453), .Z(
        n14457) );
    VMW_INV U5479 ( .A(n14364), .Z(n13953) );
    VMW_NOR4 U4037 ( .A(n13381), .B(n13382), .C(n13383), .D(n13384), .Z(n13380
        ) );
    VMW_NOR2 U4180 ( .A(n13651), .B(n13459), .Z(n13071) );
    VMW_OAI22 U4791 ( .A(n13633), .B(n14090), .C(n13609), .D(n13639), .Z(
        n13259) );
    VMW_AND3 U4297 ( .A(n13535), .B(n13783), .C(n13421), .Z(n13782) );
    VMW_OR2 U4320 ( .A(n13804), .B(n13810), .Z(n13811) );
    VMW_OAI22 U4601 ( .A(n13642), .B(n13715), .C(n13628), .D(n13714), .Z(
        n14156) );
    VMW_OAI22 U4943 ( .A(n13631), .B(n13717), .C(n13628), .D(n13723), .Z(
        n14347) );
    VMW_AO21 U5064 ( .A(n13808), .B(n13273), .C(n13812), .Z(n13281) );
    VMW_OAI22 U4516 ( .A(n13633), .B(n13647), .C(n13609), .D(n13646), .Z(
        n14105) );
    VMW_OAI22 U4531 ( .A(n13637), .B(n14097), .C(n13635), .D(n14102), .Z(
        n14113) );
    VMW_OAI211 U4964 ( .A(n13659), .B(n14362), .C(n13670), .D(n14122), .Z(
        n14361) );
    VMW_INV U5354 ( .A(n13390), .Z(n13601) );
    VMW_NOR2 U4307 ( .A(n13804), .B(n13564), .Z(n13803) );
    VMW_XOR2 U4486 ( .A(n14066), .B(\temp[50] ), .Z(n14065) );
    VMW_OAI22 U4626 ( .A(n13644), .B(n13712), .C(n13633), .D(n14169), .Z(
        n14180) );
    VMW_INV U5373 ( .A(KEY[42]), .Z(n14173) );
    VMW_FD \i_reg[0]  ( .D(n14509), .CP(Clk), .Q(\i[0] ) );
    VMW_AND2 U4059 ( .A(n13447), .B(n13156), .Z(n13446) );
    VMW_OAI22 U4369 ( .A(n13881), .B(n13584), .C(n13578), .D(n13887), .Z(
        n13886) );
    VMW_NAND3 U5043 ( .A(n13205), .B(n13515), .C(n13757), .Z(n13990) );
    VMW_OAI22 U4578 ( .A(n13641), .B(n14103), .C(n13640), .D(n14112), .Z(
        n14140) );
    VMW_FD \temp_reg[53]  ( .D(\arr12639[53] ), .CP(Clk), .Q(\temp[53] ) );
    VMW_AND2 U4272 ( .A(n13509), .B(n13754), .Z(n13202) );
    VMW_OAI22 U4463 ( .A(n13901), .B(n13603), .C(n14032), .D(n13440), .Z(
        n14031) );
    VMW_OR2 U4648 ( .A(n13728), .B(n13148), .Z(n13744) );
    VMW_OAI22 U4811 ( .A(n13609), .B(n13618), .C(n13626), .D(n13649), .Z(
        n14271) );
    VMW_AO22 U5206 ( .A(n13977), .B(n13453), .C(n13976), .D(n13659), .Z(n14464
        ) );
    VMW_INV U5396 ( .A(n13509), .Z(n13515) );
    VMW_FD \temp_reg[60]  ( .D(\arr12639[60] ), .CP(Clk), .Q(\temp[60] ) );
    VMW_FD \OUT_reg[46]  ( .D(\arr12639[26] ), .CP(Clk), .Q(OUT[46]) );
    VMW_INV U5417 ( .A(n13689), .Z(n14308) );
    VMW_AOI211 U4981 ( .A(n13782), .B(n13550), .C(n14248), .D(n13436), .Z(
        n14389) );
    VMW_OR2 U4142 ( .A(n13622), .B(n13608), .Z(n13624) );
    VMW_OAI22 U4753 ( .A(n13644), .B(n13717), .C(n13633), .D(n13716), .Z(
        n13210) );
    VMW_AO22 U5136 ( .A(n13200), .B(n13205), .C(n13754), .D(n13943), .Z(n14447
        ) );
    VMW_OR2 U4159 ( .A(n13611), .B(n13638), .Z(n13641) );
    VMW_INV U4165 ( .A(\temp[27] ), .Z(n13460) );
    VMW_AO22 U5081 ( .A(n13272), .B(n13815), .C(n13414), .D(n14306), .Z(n13863
        ) );
    VMW_OR4 U5111 ( .A(n14379), .B(n13795), .C(n13891), .D(n14439), .Z(n14028)
         );
    VMW_AND2 U4255 ( .A(n13139), .B(n13488), .Z(n13147) );
    VMW_OAI2222 U4774 ( .A(n13636), .B(n13640), .C(n13634), .D(n13637), .E(
        n13632), .F(n13635), .G(n13627), .H(n13631), .Z(n13263) );
    VMW_OR4 U4836 ( .A(n14280), .B(n14281), .C(n14278), .D(n14279), .Z(n13310)
         );
    VMW_AO22 U5221 ( .A(n13782), .B(n13543), .C(n13996), .D(n13550), .Z(n13796
        ) );
    VMW_INV U5430 ( .A(n13239), .Z(n13591) );
    VMW_AND2 U4444 ( .A(n13833), .B(n13879), .Z(n14004) );
    VMW_OAI22 U4748 ( .A(n13621), .B(n14166), .C(n13642), .D(n14167), .Z(
        n14242) );
    VMW_FD \OUT_reg[56]  ( .D(\arr12639[0] ), .CP(Clk), .Q(OUT[56]) );
    VMW_AO21 U3947 ( .A(\temp[41] ), .B(n13005), .C(n13028), .Z(\arr12639[41] 
        ) );
    VMW_NAND3 U3985 ( .A(n13161), .B(n13162), .C(n13163), .Z(n13160) );
    VMW_AND2 U4269 ( .A(n13517), .B(n13525), .Z(n13205) );
    VMW_AND2 U4478 ( .A(n13320), .B(n13578), .Z(n13605) );
    VMW_OAI21 U4355 ( .A(n13856), .B(n13322), .C(n13857), .Z(n13855) );
    VMW_OAI22 U4544 ( .A(n13633), .B(n14092), .C(n13609), .D(n14089), .Z(
        n13052) );
    VMW_OR4 U4936 ( .A(n14342), .B(n14343), .C(n14340), .D(n14341), .Z(n13381)
         );
    VMW_INV U5321 ( .A(n13087), .Z(n13477) );
    VMW_FD \temp_reg[43]  ( .D(\arr12639[43] ), .CP(Clk), .Q(\temp[43] ) );
    VMW_NOR4 U4042 ( .A(n13404), .B(n13405), .C(n13167), .D(n13406), .Z(n13403
        ) );
    VMW_AO22 U4065 ( .A(n13460), .B(n13461), .C(\temp[27] ), .D(n13063), .Z(
        n13459) );
    VMW_OAI2222 U4674 ( .A(n13632), .B(n13640), .C(n13623), .D(n13631), .E(
        n13620), .F(n13628), .G(n13618), .H(n13626), .Z(n13171) );
    VMW_AND2 U5011 ( .A(RDY), .B(n13451), .Z(n13452) );
    VMW_INV U5181 ( .A(n13499), .Z(n13729) );
    VMW_NAND3 U5036 ( .A(n13139), .B(n13154), .C(n13733), .Z(n13738) );
    VMW_OR2 U4137 ( .A(n13613), .B(n13617), .Z(n13619) );
    VMW_OR4 U4372 ( .A(n13798), .B(n13892), .C(n13889), .D(n13893), .Z(n13891)
         );
    VMW_OAI22 U4653 ( .A(n13626), .B(n14094), .C(n14085), .D(n13642), .Z(
        n14194) );
    VMW_OR3 U4881 ( .A(n13852), .B(n14304), .C(n13855), .Z(n14303) );
    VMW_INV U5296 ( .A(\i[3] ), .Z(n13614) );
    VMW_INV U5306 ( .A(n13053), .Z(n13458) );
    VMW_INV U5487 ( .A(n13650), .Z(n14413) );
    VMW_OAI22 U4911 ( .A(n13642), .B(n13712), .C(n13641), .D(n14172), .Z(
        n14331) );
    VMW_OAI22 U4563 ( .A(n13616), .B(n14103), .C(n13644), .D(n14112), .Z(
        n14133) );
    VMW_NAND4 U4958 ( .A(n14354), .B(n14355), .C(n14356), .D(n14357), .Z(
        n14353) );
    VMW_AO22 U5058 ( .A(n13272), .B(n13273), .C(n13282), .D(n13803), .Z(n13831
        ) );
    VMW_INV U5368 ( .A(KEY[63]), .Z(n14102) );
    VMW_OAI22 U4726 ( .A(n13640), .B(n13714), .C(n13624), .D(n13713), .Z(
        n14232) );
    VMW_AO21 U5143 ( .A(n13899), .B(n13906), .C(n14452), .Z(n13955) );
    VMW_AO21 U3949 ( .A(\temp[39] ), .B(n13005), .C(n13030), .Z(\arr12639[39] 
        ) );
    VMW_AO21 U3955 ( .A(\temp[33] ), .B(n13005), .C(n13036), .Z(\arr12639[33] 
        ) );
    VMW_NOR4 U3960 ( .A(n13054), .B(n13055), .C(n13056), .D(n13057), .Z(n13053
        ) );
    VMW_AO22 U4080 ( .A(n13500), .B(n13501), .C(\temp[16] ), .D(n13128), .Z(
        n13499) );
    VMW_NOR2 U4207 ( .A(n13475), .B(n13472), .Z(n13364) );
    VMW_AO21 U4586 ( .A(n13684), .B(n13685), .C(n14145), .Z(n14144) );
    VMW_OAI22 U4864 ( .A(n13624), .B(n14163), .C(n13640), .D(n14164), .Z(
        n14294) );
    VMW_AND5 U4220 ( .A(n13705), .B(n13706), .C(n13707), .D(n13708), .E(n13428
        ), .Z(n13704) );
    VMW_OAI211 U4397 ( .A(n13912), .B(n13921), .C(n13922), .D(n13923), .Z(
        n13920) );
    VMW_NAND2 U4416 ( .A(n13070), .B(n13459), .Z(n13974) );
    VMW_NAND2 U4431 ( .A(n13526), .B(n13202), .Z(n13988) );
    VMW_OAI22 U4843 ( .A(n13642), .B(n13721), .C(n13641), .D(n13720), .Z(
        n14285) );
    VMW_AO22 U5273 ( .A(n14065), .B(n13451), .C(X[45]), .D(Start), .Z(n14493)
         );
    VMW_INV U5462 ( .A(n13950), .Z(n14455) );
    VMW_OAI22 U5254 ( .A(n13149), .B(n13157), .C(n13154), .D(n13488), .Z(
        n14443) );
    VMW_INV U5445 ( .A(n13333), .Z(n13840) );
    VMW_AO22 U4110 ( .A(n13484), .B(n13570), .C(\temp[23] ), .D(n13241), .Z(
        n13569) );
    VMW_AOI211 U4701 ( .A(n13755), .B(n13520), .C(n14218), .D(n13199), .Z(
        n13768) );
    VMW_OAI22 U4691 ( .A(n13640), .B(n14090), .C(n13637), .D(n13639), .Z(
        n13182) );
    VMW_NAND5 U5164 ( .A(n13767), .B(n14460), .C(n13769), .D(n14449), .E(
        n13858), .Z(n14077) );
    VMW_AO22 U4125 ( .A(n13603), .B(n13441), .C(n13440), .D(n13401), .Z(n13602
        ) );
    VMW_OAI22 U4734 ( .A(n13626), .B(n13720), .C(n13624), .D(n13719), .Z(
        n14236) );
    VMW_NOR4 U3969 ( .A(n13098), .B(n13099), .C(n13100), .D(n13101), .Z(n13097
        ) );
    VMW_NOR4 U3972 ( .A(n13109), .B(n13110), .C(n13111), .D(n13112), .Z(n13108
        ) );
    VMW_OAI22 U4092 ( .A(n13342), .B(n13512), .C(n13528), .D(n13516), .Z(
        n13527) );
    VMW_AO22 U4102 ( .A(n13356), .B(n13546), .C(n13535), .D(n13537), .Z(n13240
        ) );
    VMW_NOR2 U4215 ( .A(n13362), .B(n13353), .Z(n13360) );
    VMW_NOR2 U4385 ( .A(n13443), .B(n13444), .Z(n13408) );
    VMW_AND2 U4404 ( .A(n13760), .B(n13505), .Z(n13943) );
    VMW_NAND3 U5151 ( .A(n13154), .B(n13731), .C(n13147), .Z(n14373) );
    VMW_OAI22 U4594 ( .A(n13616), .B(n14092), .C(n14089), .D(n13644), .Z(
        n13086) );
    VMW_INV U4232 ( .A(KEY[57]), .Z(n13720) );
    VMW_OR4 U4876 ( .A(n14300), .B(n14301), .C(n14298), .D(n14299), .Z(n13315)
         );
    VMW_AO22 U5261 ( .A(n14053), .B(n13451), .C(X[13]), .D(Start), .Z(n14487)
         );
    VMW_INV U5470 ( .A(n14247), .Z(n14423) );
    VMW_XOR2 U4423 ( .A(n13983), .B(\temp[40] ), .Z(n13982) );
    VMW_OAI22 U4851 ( .A(n13640), .B(n13715), .C(n13624), .D(n13714), .Z(
        n14289) );
    VMW_MUX2 U5246 ( .A(n14482), .B(\temp[27] ), .S(n13005), .Z(\arr12639[27] 
        ) );
    VMW_INV U5457 ( .A(n13928), .Z(n13406) );
    VMW_OAI22 U4683 ( .A(n13628), .B(n13639), .C(n13626), .D(n13636), .Z(
        n13187) );
    VMW_OAI22 U4713 ( .A(n13642), .B(n13726), .C(n13641), .D(n13718), .Z(
        n13220) );
    VMW_NOR4 U3997 ( .A(n13218), .B(n13219), .C(n13220), .D(n13221), .Z(n13217
        ) );
    VMW_AND3 U4019 ( .A(n13320), .B(n13321), .C(n13322), .Z(n13319) );
    VMW_AO21 U4189 ( .A(n13665), .B(n13659), .C(n13675), .Z(n13674) );
    VMW_AND2 U4329 ( .A(n13808), .B(n13569), .Z(n13287) );
    VMW_OAI22 U4538 ( .A(n13641), .B(n14102), .C(n13640), .D(n14103), .Z(
        n14116) );
    VMW_INV U5176 ( .A(n13478), .Z(n13682) );
    VMW_FD \temp_reg[57]  ( .D(\arr12639[57] ), .CP(Clk), .Q(\temp[57] ) );
    VMW_FD \OUT_reg[42]  ( .D(\arr12639[10] ), .CP(Clk), .Q(OUT[42]) );
    VMW_OAI22 U4608 ( .A(n13628), .B(n14163), .C(n13642), .D(n14164), .Z(
        n14162) );
    VMW_NOR2 U4347 ( .A(n13322), .B(n13320), .Z(n13325) );
    VMW_OAI2222 U4798 ( .A(n13627), .B(n13635), .C(n13625), .D(n13633), .E(
        n13609), .F(n13623), .G(n13621), .H(n13649), .Z(n13253) );
    VMW_INV U5333 ( .A(\temp[14] ), .Z(n13491) );
    VMW_FD \i_reg[4]  ( .D(n14505), .CP(Clk), .Q(\i[4] ) );
    VMW_OAI22 U4556 ( .A(n13641), .B(n13649), .C(n13631), .D(n13647), .Z(
        n14130) );
    VMW_OAI22 U4924 ( .A(n13643), .B(n13715), .C(n13631), .D(n13714), .Z(
        n14336) );
    VMW_AND3 U5003 ( .A(n13447), .B(n13156), .C(n13141), .Z(n14408) );
    VMW_INV U5193 ( .A(n13575), .Z(n13606) );
    VMW_NOR4 U4002 ( .A(n13242), .B(n13243), .C(n13244), .D(n13245), .Z(n13241
        ) );
    VMW_NOR5 U4050 ( .A(n13432), .B(n13433), .C(n13418), .D(n13434), .E(n13435
        ), .Z(n13431) );
    VMW_AO22 U4077 ( .A(n13491), .B(n13492), .C(\temp[14] ), .D(n13108), .Z(
        n13447) );
    VMW_OAI22 U4641 ( .A(n13637), .B(n13720), .C(n13635), .D(n13719), .Z(
        n14187) );
    VMW_OAI2222 U4666 ( .A(n13642), .B(n13645), .C(n13641), .D(n13648), .E(
        n13640), .F(n13647), .G(n13637), .H(n13646), .Z(n13196) );
    VMW_AO21 U5024 ( .A(n13478), .B(n13351), .C(n13424), .Z(n14150) );
    VMW_INV U4150 ( .A(KEY[28]), .Z(n13632) );
    VMW_OAI21 U4260 ( .A(n13743), .B(n13744), .C(n13745), .Z(n13742) );
    VMW_AO22 U4360 ( .A(n13687), .B(n13865), .C(n13866), .D(n13104), .Z(n13864
        ) );
    VMW_OAI22 U4571 ( .A(n13641), .B(n14119), .C(n13631), .D(n14102), .Z(
        n14137) );
    VMW_AO22 U5284 ( .A(n14074), .B(n13451), .C(X[19]), .D(Start), .Z(n14499)
         );
    VMW_INV U5314 ( .A(n13256), .Z(n13558) );
    VMW_AND2 U4818 ( .A(n13830), .B(n13562), .Z(n13824) );
    VMW_AND2 U4893 ( .A(n13562), .B(n13567), .Z(n14306) );
    VMW_AO22 U4903 ( .A(n13540), .B(n13786), .C(n13775), .D(n13781), .Z(n13890
        ) );
    VMW_NAND2 U4988 ( .A(n13584), .B(n14399), .Z(n13847) );
    VMW_AO21 U5088 ( .A(n13686), .B(n14418), .C(n13683), .Z(n14431) );
    VMW_AO22 U5228 ( .A(n14407), .B(n13578), .C(n14004), .D(n13322), .Z(n13850
        ) );
    VMW_INV U5439 ( .A(n13285), .Z(n14275) );
    VMW_NAND3 U5118 ( .A(n13444), .B(n14400), .C(n13908), .Z(n13922) );
    VMW_AO22 U5214 ( .A(n13985), .B(n13499), .C(n13986), .D(n13729), .Z(n14467
        ) );
    VMW_INV U5384 ( .A(KEY[58]), .Z(n14164) );
    VMW_INV U5405 ( .A(n13581), .Z(n13320) );
    VMW_XNOR2 U4471 ( .A(\temp[56] ), .B(n13403), .Z(n14045) );
    VMW_OAI22 U4803 ( .A(n13624), .B(n14097), .C(n13621), .D(n14102), .Z(
        n14267) );
    VMW_AND2 U4993 ( .A(n13543), .B(n14402), .Z(n14248) );
    VMW_NAND3 U5124 ( .A(n13441), .B(n14441), .C(n13913), .Z(n14354) );
    VMW_AND2 U4177 ( .A(n13456), .B(n13655), .Z(n13657) );
    VMW_OAI22 U4741 ( .A(n13642), .B(n14169), .C(n13641), .D(n14170), .Z(
        n14239) );
    VMW_AO22 U4766 ( .A(X[28]), .B(n13774), .C(n13773), .D(\temp[20] ), .Z(
        n13017) );
    VMW_OAI21 U5093 ( .A(n13736), .B(n14408), .C(n13154), .Z(n13876) );
    VMW_AO22 U5103 ( .A(n13328), .B(n14437), .C(n13605), .D(n13331), .Z(n14398
        ) );
    VMW_OR2 U4192 ( .A(Reset), .B(n13452), .Z(n13005) );
    VMW_AND2 U4247 ( .A(n13139), .B(n13161), .Z(n13732) );
    VMW_NAND2 U4456 ( .A(n13162), .B(n13499), .Z(n14020) );
    VMW_AO22 U5233 ( .A(n14013), .B(n13451), .C(X[7]), .D(Start), .Z(n14476)
         );
    VMW_INV U5422 ( .A(n13733), .Z(n13749) );
    VMW_AO22 U4824 ( .A(X[2]), .B(n13774), .C(n13773), .D(\temp[15] ), .Z(
        n13022) );
    VMW_AO22 U4888 ( .A(X[48]), .B(n13774), .C(\temp[1] ), .D(n13773), .Z(
        n13036) );
    VMW_OAI22 U4918 ( .A(n13609), .B(n14172), .C(n13616), .D(n14169), .Z(
        n14334) );
    VMW_OAI211 U5018 ( .A(n13664), .B(n13657), .C(n13453), .D(n13653), .Z(
        n14123) );
    VMW_INV U5188 ( .A(n13531), .Z(n13547) );
    VMW_INV U5328 ( .A(n13184), .Z(n13519) );
    VMW_OAI2222 U4613 ( .A(n13633), .B(n13715), .C(n13616), .D(n13714), .E(
        n13635), .F(n13713), .G(n13624), .H(n13712), .Z(n13120) );
    VMW_AND2 U4025 ( .A(n13204), .B(n13339), .Z(n13338) );
    VMW_AND3 U4285 ( .A(n13535), .B(n13776), .C(n13437), .Z(n13775) );
    VMW_AND2 U4315 ( .A(n13808), .B(n13414), .Z(n13344) );
    VMW_AO22 U4332 ( .A(n13816), .B(n13282), .C(n13824), .D(n13564), .Z(n13823
        ) );
    VMW_OAI22 U4523 ( .A(n13625), .B(n13641), .C(n13623), .D(n13640), .Z(
        n14108) );
    VMW_OAI22 U4783 ( .A(n13630), .B(n13644), .C(n13633), .D(n13649), .Z(
        n13269) );
    VMW_AO22 U5076 ( .A(n13335), .B(n13832), .C(n13833), .D(n13842), .Z(n14002
        ) );
    VMW_XOR2 U4494 ( .A(n14079), .B(\temp[43] ), .Z(n14078) );
    VMW_OAI22 U4951 ( .A(n13616), .B(n13712), .C(n13644), .D(n14172), .Z(
        n14351) );
    VMW_INV U5346 ( .A(n13365), .Z(n13592) );
    VMW_OAI22 U4504 ( .A(n14091), .B(n13644), .C(n14092), .D(n13643), .Z(
        n13057) );
    VMW_OR3 U4976 ( .A(n14379), .B(n13420), .C(n13962), .Z(n14378) );
    VMW_INV U5361 ( .A(KEY[54]), .Z(n14091) );
    VMW_OAI22 U4634 ( .A(n13616), .B(n13720), .C(n13644), .D(n13719), .Z(
        n14184) );
    VMW_OR2 U5051 ( .A(n13778), .B(n13994), .Z(n13783) );
    VMW_NOR4 U4005 ( .A(n13257), .B(n13258), .C(n13259), .D(n13260), .Z(n13256
        ) );
    VMW_AND2 U4022 ( .A(n13322), .B(n13331), .Z(n13330) );
    VMW_AO22 U4089 ( .A(n13521), .B(n13512), .C(n13522), .D(n13516), .Z(n13520
        ) );
    VMW_AO22 U4119 ( .A(n13573), .B(n13592), .C(\temp[8] ), .D(n13365), .Z(
        n13441) );
    VMW_FD \OUT_reg[52]  ( .D(\arr12639[17] ), .CP(Clk), .Q(OUT[52]) );
    VMW_OAI2222 U4698 ( .A(n13624), .B(n13639), .C(n13621), .D(n13636), .E(
        n13619), .F(n13634), .G(n13616), .H(n13632), .Z(n13176) );
    VMW_INV U4229 ( .A(KEY[52]), .Z(n13718) );
    VMW_OAI22 U4708 ( .A(n13644), .B(n14166), .C(n13637), .D(n14167), .Z(
        n14222) );
    VMW_FD \temp_reg[47]  ( .D(\arr12639[47] ), .CP(Clk), .Q(\temp[47] ) );
    VMW_FD \OUT_reg[61]  ( .D(\arr12639[48] ), .CP(Clk), .Q(OUT[61]) );
    VMW_NOR2 U4438 ( .A(n13993), .B(n13591), .Z(n13995) );
    VMW_OAI22 U4633 ( .A(n13642), .B(n13716), .C(n13628), .D(n13715), .Z(
        n14183) );
    VMW_OR4 U5056 ( .A(n13795), .B(n13791), .C(n13798), .D(n14423), .Z(n13998)
         );
    VMW_NOR2 U4282 ( .A(n13005), .B(Start), .Z(n13773) );
    VMW_AOI211 U4971 ( .A(n14275), .B(n13414), .C(n14369), .D(n13821), .Z(
        n14370) );
    VMW_INV U5366 ( .A(KEY[31]), .Z(n14096) );
    VMW_AND2 U4312 ( .A(n13567), .B(n13804), .Z(n13412) );
    VMW_OAI22 U4503 ( .A(n14089), .B(n13642), .C(n14090), .D(n13641), .Z(
        n13056) );
    VMW_AO22 U4335 ( .A(n13809), .B(n13830), .C(n13807), .D(n13831), .Z(n13829
        ) );
    VMW_XOR2 U4493 ( .A(n14077), .B(\temp[44] ), .Z(n14076) );
    VMW_AOI211 U4956 ( .A(n13409), .B(n14352), .C(n13951), .D(n13399), .Z(
        n13919) );
    VMW_INV U5341 ( .A(\temp[10] ), .Z(n13579) );
    VMW_OAI22 U4524 ( .A(n13630), .B(n13643), .C(n13627), .D(n13642), .Z(
        n14109) );
    VMW_OAI22 U4784 ( .A(n13631), .B(n14091), .C(n13609), .D(n14092), .Z(
        n13270) );
    VMW_AND4 U5071 ( .A(n13572), .B(n13325), .C(n13328), .D(n13335), .Z(n13851
        ) );
    VMW_OR2 U4139 ( .A(n13607), .B(n13613), .Z(n13621) );
    VMW_INV U4195 ( .A(\temp[24] ), .Z(n13473) );
    VMW_OAI22 U4614 ( .A(n13609), .B(n13717), .C(n13644), .D(n13716), .Z(
        n13121) );
    VMW_OAI2222 U4728 ( .A(n13616), .B(n13723), .C(n13644), .D(n13722), .E(
        n13637), .F(n13716), .G(n13621), .H(n13715), .Z(n13229) );
    VMW_FD \OUT_reg[50]  ( .D(\arr12639[9] ), .CP(Clk), .Q(OUT[50]) );
    VMW_FD \OUT_reg[49]  ( .D(\arr12639[33] ), .CP(Clk), .Q(OUT[49]) );
    VMW_INV U4157 ( .A(KEY[45]), .Z(n13639) );
    VMW_INV U4170 ( .A(\temp[31] ), .Z(n13462) );
    VMW_AND2 U4209 ( .A(n13472), .B(n13686), .Z(n13103) );
    VMW_INV U4240 ( .A(KEY[26]), .Z(n13727) );
    VMW_NOR5 U4399 ( .A(n13929), .B(n13930), .C(n13931), .D(n13166), .E(n13737
        ), .Z(n13928) );
    VMW_OAI22 U4588 ( .A(n13628), .B(n14097), .C(n13626), .D(n14102), .Z(
        n14147) );
    VMW_AND2 U4418 ( .A(n13656), .B(n13657), .Z(n13976) );
    VMW_AO22 U4823 ( .A(X[60]), .B(n13774), .C(n13773), .D(\temp[16] ), .Z(
        n13021) );
    VMW_FD \temp_reg[45]  ( .D(\arr12639[45] ), .CP(Clk), .Q(\temp[45] ) );
    VMW_FD \OUT_reg[63]  ( .D(\arr12639[56] ), .CP(Clk), .Q(OUT[63]) );
    VMW_XOR2 U4451 ( .A(n14014), .B(\temp[63] ), .Z(n14013) );
    VMW_MUX2 U5234 ( .A(n14476), .B(\temp[31] ), .S(n13005), .Z(\arr12639[31] 
        ) );
    VMW_INV U5425 ( .A(n13735), .Z(n13163) );
    VMW_OAI22 U4746 ( .A(n13644), .B(n14160), .C(n13633), .D(n13717), .Z(
        n13236) );
    VMW_AO22 U4761 ( .A(X[54]), .B(n13774), .C(\temp[25] ), .D(n13773), .Z(
        n13012) );
    VMW_NAND3 U5094 ( .A(n13139), .B(n13162), .C(n13149), .Z(n14432) );
    VMW_NAND3 U5104 ( .A(n13586), .B(n13606), .C(n13832), .Z(n13885) );
    VMW_NAND2 U5123 ( .A(n13906), .B(n13408), .Z(n14355) );
    VMW_AO21 U3935 ( .A(\temp[53] ), .B(n13005), .C(n13016), .Z(\arr12639[53] 
        ) );
    VMW_AO21 U3940 ( .A(\temp[48] ), .B(n13005), .C(n13021), .Z(\arr12639[48] 
        ) );
    VMW_AO21 U3952 ( .A(\temp[36] ), .B(n13005), .C(n13033), .Z(\arr12639[36] 
        ) );
    VMW_NOR4 U3975 ( .A(n13124), .B(n13125), .C(n13126), .D(n13127), .Z(n13123
        ) );
    VMW_NOR4 U3990 ( .A(n13185), .B(n13186), .C(n13187), .D(n13188), .Z(n13184
        ) );
    VMW_AND2 U4057 ( .A(\i6749[1] ), .B(n13445), .Z(n14508) );
    VMW_AND2 U4267 ( .A(n13509), .B(n13517), .Z(n13528) );
    VMW_XOR2 U4476 ( .A(n14052), .B(\temp[55] ), .Z(n14051) );
    VMW_OAI22 U4804 ( .A(n13633), .B(n14119), .C(n13626), .D(n14096), .Z(
        n14268) );
    VMW_AO21 U4994 ( .A(n14403), .B(n13968), .C(n13453), .Z(n13673) );
    VMW_NAND2 U4367 ( .A(n13879), .B(n13325), .Z(n13881) );
    VMW_AO22 U4894 ( .A(n14274), .B(n13282), .C(n13276), .D(n13272), .Z(n13348
        ) );
    VMW_OAI22 U4938 ( .A(n13628), .B(n13718), .C(n13643), .D(n13727), .Z(
        n13383) );
    VMW_MUX2 U5213 ( .A(n14466), .B(\temp[8] ), .S(n13005), .Z(\arr12639[8] )
         );
    VMW_INV U5383 ( .A(KEY[1]), .Z(n14163) );
    VMW_INV U5402 ( .A(n13559), .Z(n13805) );
    VMW_AND4 U5038 ( .A(n13447), .B(n13154), .C(n13139), .D(n13162), .Z(n14191
        ) );
    VMW_INV U5298 ( .A(n13043), .Z(n13466) );
    VMW_INV U5308 ( .A(n13063), .Z(n13461) );
    VMW_INV U5489 ( .A(n14469), .Z(n14218) );
    VMW_AOI211 U4904 ( .A(n13784), .B(n13438), .C(n14245), .D(n13354), .Z(
        n14321) );
    VMW_OAI22 U4576 ( .A(n13616), .B(n14090), .C(n13639), .D(n13644), .Z(
        n13095) );
    VMW_MUX2 U5283 ( .A(n14498), .B(\temp[14] ), .S(n13005), .Z(\arr12639[14] 
        ) );
    VMW_INV U5313 ( .A(n13097), .Z(n13474) );
    VMW_INV U5492 ( .A(n13656), .Z(n14456) );
    VMW_AO22 U4070 ( .A(n13473), .B(n13474), .C(\temp[24] ), .D(n13097), .Z(
        n13472) );
    VMW_OAI22 U4646 ( .A(n13626), .B(n14161), .C(n13624), .D(n14159), .Z(
        n13131) );
    VMW_OAI22 U4661 ( .A(n13643), .B(n14094), .C(n14085), .D(n13631), .Z(
        n14198) );
    VMW_AND2 U5023 ( .A(n13359), .B(n13687), .Z(n14405) );
    VMW_INV U5194 ( .A(n13572), .Z(n13334) );
    VMW_NAND3 U4340 ( .A(n13575), .B(n13329), .C(n13572), .Z(n13836) );
    VMW_OAI2222 U4551 ( .A(n13616), .B(n13636), .C(n13634), .D(n13644), .E(
        n13630), .F(n13642), .G(n13627), .H(n13641), .Z(n13079) );
    VMW_OAI22 U4923 ( .A(n13621), .B(n14173), .C(n13643), .D(n13725), .Z(
        n13394) );
    VMW_AND2 U5004 ( .A(n13897), .B(n13400), .Z(n14041) );
    VMW_OAI22 U4838 ( .A(n13642), .B(n14159), .C(n13641), .D(n13725), .Z(
        n13312) );
    VMW_NAND5 U5138 ( .A(n13766), .B(n14448), .C(n13859), .D(n14427), .E(
        n14449), .Z(n14054) );
    VMW_AO22 U5208 ( .A(n13978), .B(n13451), .C(X[51]), .D(Start), .Z(n14465)
         );
    VMW_INV U5334 ( .A(n13108), .Z(n13492) );
    VMW_INV U5398 ( .A(n13517), .Z(n13754) );
    VMW_INV U5419 ( .A(n13696), .Z(n13428) );
    VMW_AO22 U4095 ( .A(n13465), .B(n13534), .C(\temp[0] ), .D(n13232), .Z(
        n13437) );
    VMW_OAI22 U4714 ( .A(n13624), .B(n14173), .C(n13643), .D(n13724), .Z(
        n13221) );
    VMW_OR4 U5171 ( .A(n13918), .B(n13954), .C(n13965), .D(n14392), .Z(n14083)
         );
    VMW_AO22 U4105 ( .A(n13473), .B(n13558), .C(\temp[24] ), .D(n13256), .Z(
        n13557) );
    VMW_OAI22 U4684 ( .A(n13637), .B(n14091), .C(n13631), .D(n14090), .Z(
        n13188) );
    VMW_AND2 U4212 ( .A(n13680), .B(n13481), .Z(n13691) );
    VMW_INV U4235 ( .A(KEY[9]), .Z(n13723) );
    VMW_AO22 U4424 ( .A(n13732), .B(n13488), .C(n13446), .D(n13157), .Z(n13984
        ) );
    VMW_OAI22 U4856 ( .A(n13642), .B(n14163), .C(n13626), .D(n14164), .Z(
        n14290) );
    VMW_MUX2 U5241 ( .A(n14480), .B(\temp[29] ), .S(n13005), .Z(\arr12639[29] 
        ) );
    VMW_INV U5450 ( .A(n13874), .Z(n14435) );
    VMW_OAI22 U4871 ( .A(n13641), .B(n14173), .C(n13631), .D(n13724), .Z(
        n13298) );
    VMW_AO22 U5266 ( .A(n14059), .B(n13451), .C(X[29]), .D(Start), .Z(n14489)
         );
    VMW_INV U5477 ( .A(n14370), .Z(n13419) );
    VMW_AND2 U4382 ( .A(n13904), .B(n13443), .Z(n13903) );
    VMW_OAI22 U4593 ( .A(n13630), .B(n13635), .C(n13627), .D(n13633), .Z(
        n13085) );
    VMW_AO22 U4403 ( .A(n13668), .B(n13941), .C(n13942), .D(n13656), .Z(n13940
        ) );
    VMW_NOR4 U3967 ( .A(n13088), .B(n13089), .C(n13090), .D(n13091), .Z(n13087
        ) );
    VMW_NOR4 U4039 ( .A(n13391), .B(n13392), .C(n13393), .D(n13394), .Z(n13390
        ) );
    VMW_AO22 U4122 ( .A(n13582), .B(n13597), .C(\temp[7] ), .D(n13385), .Z(
        n13596) );
    VMW_OAI211 U5156 ( .A(n13423), .B(n13703), .C(n13353), .D(n13472), .Z(
        n14380) );
    VMW_AND2 U4299 ( .A(n13549), .B(n13550), .Z(n13357) );
    VMW_OAI22 U4733 ( .A(n13621), .B(n13727), .C(n13609), .D(n13712), .Z(
        n14235) );
    VMW_AND2 U4309 ( .A(n13564), .B(n13804), .Z(n13273) );
    VMW_OAI2222 U4518 ( .A(n13618), .B(n13643), .C(n13615), .D(n13642), .E(
        n13637), .F(n13645), .G(n13635), .H(n13648), .Z(n13040) );
    VMW_XNOR2 U4488 ( .A(\temp[48] ), .B(n13426), .Z(n14069) );
    VMW_OR4 U4628 ( .A(n14180), .B(n14181), .C(n14178), .D(n14179), .Z(n13124)
         );
    VMW_FD \temp_reg[55]  ( .D(\arr12639[55] ), .CP(Clk), .Q(\temp[55] ) );
    VMW_OAI211 U4978 ( .A(n14384), .B(n13658), .C(n14385), .D(n13672), .Z(
        n14383) );
    VMW_OR4 U5078 ( .A(n13332), .B(n13336), .C(n13845), .D(n14303), .Z(n14006)
         );
    VMW_FD \OUT_reg[59]  ( .D(\arr12639[40] ), .CP(Clk), .Q(OUT[59]) );
    VMW_FD \OUT_reg[40]  ( .D(\arr12639[2] ), .CP(Clk), .Q(OUT[40]) );
    VMW_INV U5348 ( .A(n13385), .Z(n13597) );
    VMW_OR3 U5163 ( .A(n14461), .B(n13758), .C(n14462), .Z(n14460) );
    VMW_AO22 U4087 ( .A(n13515), .B(n13512), .C(n13509), .D(n13516), .Z(n13514
        ) );
    VMW_AO22 U4117 ( .A(n13587), .B(n13578), .C(n13324), .D(n13322), .Z(n13586
        ) );
    VMW_OAI22 U4696 ( .A(n13627), .B(n13643), .C(n13625), .D(n13642), .Z(
        n14217) );
    VMW_AO22 U4706 ( .A(X[30]), .B(n13774), .C(n13773), .D(\temp[28] ), .Z(
        n13009) );
    VMW_AND2 U4200 ( .A(n13353), .B(n13683), .Z(n13684) );
    VMW_INV U4227 ( .A(KEY[34]), .Z(n13716) );
    VMW_MUX2 U5253 ( .A(n14484), .B(\temp[25] ), .S(n13005), .Z(\arr12639[25] 
        ) );
    VMW_INV U5442 ( .A(n13825), .Z(n14430) );
    VMW_AND2 U4390 ( .A(n13897), .B(n13909), .Z(n13910) );
    VMW_AND2 U4436 ( .A(n13546), .B(n13540), .Z(n13552) );
    VMW_OR4 U4844 ( .A(n14284), .B(n14285), .C(n14282), .D(n14283), .Z(n13300)
         );
    VMW_MUX2 U5274 ( .A(n14493), .B(\temp[18] ), .S(n13005), .Z(\arr12639[18] 
        ) );
    VMW_INV U5465 ( .A(n13981), .Z(n13697) );
    VMW_OAI21 U4411 ( .A(n13785), .B(n13963), .C(n13964), .Z(n13962) );
    VMW_OAI22 U4581 ( .A(n13628), .B(n13648), .C(n13626), .D(n13647), .Z(
        n14143) );
    VMW_OAI22 U4863 ( .A(n13628), .B(n14173), .C(n13643), .D(n13718), .Z(
        n13293) );
    VMW_NAND3 U5144 ( .A(n13397), .B(n14441), .C(n13903), .Z(n14453) );
    VMW_AOI211 U3982 ( .A(n13143), .B(n13154), .C(n13146), .D(n13150), .Z(
        n13153) );
    VMW_AND2 U4045 ( .A(n13414), .B(n13276), .Z(n13413) );
    VMW_NOR3 U4130 ( .A(n13609), .B(\i[5] ), .C(n13610), .Z(RDY) );
    VMW_OAI22 U4721 ( .A(n13635), .B(n14159), .C(n13633), .D(n13725), .Z(
        n13215) );
    VMW_AND2 U4179 ( .A(n13471), .B(n13654), .Z(n13661) );
    VMW_AO22 U4768 ( .A(X[44]), .B(n13774), .C(n13773), .D(\temp[18] ), .Z(
        n13019) );
    VMW_FD \OUT_reg[54]  ( .D(\arr12639[25] ), .CP(Clk), .Q(OUT[54]) );
    VMW_AND3 U4249 ( .A(n13148), .B(n13161), .C(n13488), .Z(n13733) );
    VMW_XOR2 U4458 ( .A(n14024), .B(\temp[60] ), .Z(n14023) );
    VMW_FD \temp_reg[58]  ( .D(\arr12639[58] ), .CP(Clk), .Q(\temp[58] ) );
    VMW_FD \temp_reg[41]  ( .D(\arr12639[41] ), .CP(Clk), .Q(\temp[41] ) );
    VMW_NOR2 U4375 ( .A(n13444), .B(n13598), .Z(n13398) );
    VMW_OAI22 U4564 ( .A(n13621), .B(n14097), .C(n13619), .D(n14102), .Z(
        n14134) );
    VMW_OAI22 U4654 ( .A(n13635), .B(n14103), .C(n13633), .D(n14112), .Z(
        n14195) );
    VMW_AO22 U4886 ( .A(X[32]), .B(n13774), .C(\temp[3] ), .D(n13773), .Z(
        n13034) );
    VMW_OAI22 U4916 ( .A(n13637), .B(n14163), .C(n13619), .D(n14164), .Z(
        n14332) );
    VMW_AO22 U5291 ( .A(n14080), .B(n13451), .C(X[43]), .D(Start), .Z(n14502)
         );
    VMW_INV U5301 ( .A(n13222), .Z(n13536) );
    VMW_INV U5480 ( .A(n14395), .Z(n14365) );
    VMW_AOI211 U4062 ( .A(n13451), .B(\i6749[4] ), .C(n13452), .D(Reset), .Z(
        n13450) );
    VMW_NAND4 U5031 ( .A(n14310), .B(n14381), .C(n14420), .D(n14421), .Z(
        n13983) );
    VMW_OR4 U4673 ( .A(n14204), .B(n14205), .C(n14202), .D(n14203), .Z(n13170)
         );
    VMW_OR3 U5016 ( .A(n13654), .B(n13456), .C(n14415), .Z(n13671) );
    VMW_NOR4 U3999 ( .A(n13228), .B(n13229), .C(n13230), .D(n13231), .Z(n13227
        ) );
    VMW_NOR2 U4349 ( .A(n13322), .B(n13606), .Z(n13327) );
    VMW_NAND4 U4352 ( .A(n13846), .B(n13847), .C(n13841), .D(n13848), .Z(
        n13845) );
    VMW_INV U5186 ( .A(n13540), .Z(n13556) );
    VMW_OAI22 U4543 ( .A(n13616), .B(n13630), .C(n13627), .D(n13644), .Z(
        n13051) );
    VMW_OAI22 U4931 ( .A(n13626), .B(n14160), .C(n13624), .D(n14161), .Z(
        n13374) );
    VMW_INV U5326 ( .A(n13179), .Z(n13511) );
    VMW_FD \temp_reg[51]  ( .D(\arr12639[51] ), .CP(Clk), .Q(\temp[51] ) );
    VMW_FD \temp_reg[48]  ( .D(\arr12639[48] ), .CP(Clk), .Q(\temp[48] ) );
    VMW_OR4 U4558 ( .A(n14130), .B(n14131), .C(n14128), .D(n14129), .Z(n13098)
         );
    VMW_AO22 U4079 ( .A(n13497), .B(n13498), .C(\temp[15] ), .D(n13113), .Z(
        n13496) );
    VMW_FD \temp_reg[62]  ( .D(\arr12639[62] ), .CP(Clk), .Q(\temp[62] ) );
    VMW_FD \OUT_reg[44]  ( .D(\arr12639[18] ), .CP(Clk), .Q(OUT[44]) );
    VMW_INV U4145 ( .A(KEY[23]), .Z(n13627) );
    VMW_OR2 U4162 ( .A(n13613), .B(n13622), .Z(n13644) );
    VMW_AND2 U4252 ( .A(n13493), .B(n13157), .Z(n13152) );
    VMW_AND3 U4443 ( .A(n13578), .B(n13337), .C(n13837), .Z(n14003) );
    VMW_OAI22 U4668 ( .A(n14092), .B(n13644), .C(n13630), .D(n13633), .Z(
        n13198) );
    VMW_OR4 U4773 ( .A(n14251), .B(n14252), .C(n14249), .D(n14250), .Z(n13262)
         );
    VMW_AO22 U4831 ( .A(X[58]), .B(n13774), .C(n13773), .D(\temp[8] ), .Z(
        n13029) );
    VMW_MUX2 U5226 ( .A(n14472), .B(\temp[4] ), .S(n13005), .Z(\arr12639[4] )
         );
    VMW_INV U5437 ( .A(n13284), .Z(n13277) );
    VMW_AND3 U5086 ( .A(n13472), .B(n13363), .C(n13687), .Z(n13871) );
    VMW_OAI21 U5116 ( .A(n14409), .B(n14041), .C(n13905), .Z(n13927) );
    VMW_OAI22 U4754 ( .A(n13631), .B(n14173), .C(n13609), .D(n14160), .Z(
        n13211) );
    VMW_NOR4 U4017 ( .A(n13310), .B(n13311), .C(n13312), .D(n13313), .Z(n13309
        ) );
    VMW_AND3 U4030 ( .A(n13351), .B(n13352), .C(n13353), .Z(n13350) );
    VMW_NOR3 U4275 ( .A(n13760), .B(n13507), .C(n13525), .Z(n13759) );
    VMW_NAND3 U5131 ( .A(n13653), .B(n13659), .C(n13657), .Z(n13937) );
    VMW_AND2 U4464 ( .A(n13901), .B(n13902), .Z(n14033) );
    VMW_OAI22 U4816 ( .A(n13624), .B(n14092), .C(n13621), .D(n14089), .Z(
        n13245) );
    VMW_AND3 U4986 ( .A(n13496), .B(n13139), .C(n14397), .Z(n14316) );
    VMW_OAI22 U4878 ( .A(n13633), .B(n14159), .C(n13609), .D(n13725), .Z(
        n13317) );
    VMW_NAND2 U5201 ( .A(n13656), .B(n13652), .Z(n13970) );
    VMW_INV U5391 ( .A(n13351), .Z(n13681) );
    VMW_INV U5410 ( .A(n13653), .Z(n14384) );
    VMW_NAND3 U5044 ( .A(n13512), .B(n13507), .C(n13530), .Z(n13989) );
    VMW_AO22 U5178 ( .A(n13362), .B(n13478), .C(n13688), .D(n13682), .Z(n13695
        ) );
    VMW_MUX2 U5248 ( .A(n14483), .B(\temp[26] ), .S(n13005), .Z(\arr12639[26] 
        ) );
    VMW_INV U5459 ( .A(n13933), .Z(n13938) );
    VMW_NOR2 U4187 ( .A(n13453), .B(n13470), .Z(n13668) );
    VMW_AND2 U4290 ( .A(n13556), .B(n13546), .Z(n13421) );
    VMW_NOR3 U4300 ( .A(n13356), .B(n13437), .C(n13785), .Z(n13784) );
    VMW_OAI2222 U4621 ( .A(n13609), .B(n13722), .C(n13619), .D(n13716), .E(
        n13637), .F(n13715), .G(n13621), .H(n13714), .Z(n13110) );
    VMW_INV U5374 ( .A(KEY[50]), .Z(n14160) );
    VMW_AO22 U4481 ( .A(n13449), .B(n13444), .C(n13908), .D(n13897), .Z(n14058
        ) );
    VMW_NOR2 U4327 ( .A(n13564), .B(n13569), .Z(n13347) );
    VMW_OAI22 U4511 ( .A(n13639), .B(n13642), .C(n13636), .D(n13641), .Z(
        n13066) );
    VMW_OAI22 U4536 ( .A(n13626), .B(n14091), .C(n13634), .D(n13643), .Z(
        n13062) );
    VMW_AND2 U4963 ( .A(n13650), .B(n13652), .Z(n13942) );
    VMW_INV U5353 ( .A(n13227), .Z(n13533) );
    VMW_FD \i_reg[2]  ( .D(n14507), .CP(Clk), .Q(\i[2] ) );
    VMW_OAI22 U4606 ( .A(n13619), .B(n14159), .C(n13616), .D(n13725), .Z(
        n13136) );
    VMW_OR4 U4944 ( .A(n14346), .B(n14347), .C(n14344), .D(n14345), .Z(n13376)
         );
    VMW_AO22 U5063 ( .A(n13414), .B(n13412), .C(n13287), .D(n13277), .Z(n13820
        ) );
    VMW_OAI22 U4796 ( .A(n13643), .B(n13648), .C(n13642), .D(n13647), .Z(
        n14264) );
endmodule


module DES_Node_WIDTH64_MEMSPACE2_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, key, start, rdy );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [63:0] key;
input  Clk, Reset, RD, WR, ScanEnable, start;
output rdy;
    wire \x[57] , \x[39] , \out[3] , n287, n317, \out[55] , n330, \out[45] , 
        n279, n379, n362, n345, \x[36] , \x[34] , n421, n406, n387, n433, 
        \out[62] , n414, n395, n339, \out[51] , \out[48] , \out[7] , n370, 
        n357, n295, n305, n322, \out[58] , \out[41] , n292, n428, n325, n302, 
        \out[43] , n277, n408, n389, n441, n350, \out[5] , n377, n434, n413, 
        n392, \x[32] , \out[60] , n289, n319, \out[53] , n401, n380, \out[8] , 
        n426, \out[47] , n342, \out[57] , n365, n359, \out[1] , n280, n310, 
        n337, n435, n412, n393, n288, n318, \out[18] , \out[32] , n351, 
        \x[60] , \x[53] , \x[47] , n276, n376, n440, n324, \out[22] , n293, 
        n303, \out[11] , n409, n388, n281, n336, n311, \out[36] , n358, 
        \x[58] , \x[43] , \out[26] , \out[15] , n343, n427, n400, n364, n381, 
        n420, n407, n386, \out[24] , n278, \out[17] , n344, n363, \x[41] , 
        \out[34] , \x[63] , \x[62] , \x[51] , n378, \x[48] , \x[59] , \x[55] , 
        \x[45] , n286, n316, n331, \out[39] , n294, n304, n323, \out[20] , 
        \out[13] , n429, n371, n432, n356, \x[54] , \x[44] , n415, n338, n394, 
        \out[30] , \out[29] , n333, n284, n314, n439, \out[38] , \out[21] , 
        \out[12] , n346, n361, \x[40] , n422, n405, n384, \out[31] , \out[28] , 
        n328, n417, n396, \out[25] , n430, \out[16] , n354, \x[50] , \x[49] , 
        n368, n373, \out[35] , n445, \x[61] , \x[52] , n321, n291, n296, n301, 
        n306, n326, n348, \out[37] , n442, \x[56] , \x[42] , \out[27] , 
        \out[14] , n353, n374, n437, n425, n410, n391, \x[46] , \out[19] , 
        n402, n383, \out[33] , n298, n308, n341, n366, n283, n313, n334, 
        \x[37] , \x[33] , \out[23] , n419, n398, \out[10] , n436, \out[9] , 
        \out[46] , n411, n390, n352, n375, \out[56] , n349, n443, \out[0] , 
        n275, n290, n300, n327, n282, n312, \out[42] , n418, n335, n399, 
        startflag, \out[4] , n424, n340, n367, \x[35] , \out[61] , n403, n382, 
        \out[52] , n299, n309, n404, n385, \out[63] , n423, \out[50] , 
        \out[49] , \out[6] , n329, n347, n360, n332, \x[38] , \out[59] , 
        \out[40] , n285, n438, n315, n320, \out[2] , \out[54] , n297, n307, 
        n369, \out[44] , n444, n355, n372, n416, n397, n431;
    DES_ECB_dummy1 des_module ( .Clk(Clk), .Reset(Reset), .Start(start), .X({
        \x[63] , \x[62] , \x[61] , \x[60] , \x[59] , \x[58] , \x[57] , \x[56] , 
        \x[55] , \x[54] , \x[53] , \x[52] , \x[51] , \x[50] , \x[49] , \x[48] , 
        \x[47] , \x[46] , \x[45] , \x[44] , \x[43] , \x[42] , \x[41] , \x[40] , 
        \x[39] , \x[38] , \x[37] , \x[36] , \x[35] , \x[34] , \x[33] , \x[32] , 
        ScanOut[31], ScanOut[30], ScanOut[29], ScanOut[28], ScanOut[27], 
        ScanOut[26], ScanOut[25], ScanOut[24], ScanOut[23], ScanOut[22], 
        ScanOut[21], ScanOut[20], ScanOut[19], ScanOut[18], ScanOut[17], 
        ScanOut[16], ScanOut[15], ScanOut[14], ScanOut[13], ScanOut[12], 
        ScanOut[11], ScanOut[10], ScanOut[9], ScanOut[8], ScanOut[7], 
        ScanOut[6], ScanOut[5], ScanOut[4], ScanOut[3], ScanOut[2], ScanOut[1], 
        ScanOut[0]}), .KEY(key), .OUT({\out[63] , \out[62] , \out[61] , 
        \out[60] , \out[59] , \out[58] , \out[57] , \out[56] , \out[55] , 
        \out[54] , \out[53] , \out[52] , \out[51] , \out[50] , \out[49] , 
        \out[48] , \out[47] , \out[46] , \out[45] , \out[44] , \out[43] , 
        \out[42] , \out[41] , \out[40] , \out[39] , \out[38] , \out[37] , 
        \out[36] , \out[35] , \out[34] , \out[33] , \out[32] , \out[31] , 
        \out[30] , \out[29] , \out[28] , \out[27] , \out[26] , \out[25] , 
        \out[24] , \out[23] , \out[22] , \out[21] , \out[20] , \out[19] , 
        \out[18] , \out[17] , \out[16] , \out[15] , \out[14] , \out[13] , 
        \out[12] , \out[11] , \out[10] , \out[9] , \out[8] , \out[7] , 
        \out[6] , \out[5] , \out[4] , \out[3] , \out[2] , \out[1] , \out[0] }), 
        .RDY(rdy) );
    VMW_AND2 U48 ( .A(n275), .B(n276), .Z(n445) );
    VMW_OR2 U54 ( .A(n287), .B(n288), .Z(n439) );
    VMW_OR2 U73 ( .A(n325), .B(n326), .Z(n420) );
    VMW_AND2 U113 ( .A(ScanEnable), .B(n375), .Z(n374) );
    VMW_AO22 U134 ( .A(ScanIn[25]), .B(ScanEnable), .C(\out[57] ), .D(n379), 
        .Z(n367) );
    VMW_OR2 U61 ( .A(n301), .B(n302), .Z(n432) );
    VMW_OR2 U68 ( .A(n315), .B(n316), .Z(n425) );
    VMW_AO21 U96 ( .A(\x[47] ), .B(n341), .C(n357), .Z(n397) );
    VMW_AO22 U198 ( .A(n377), .B(\out[48] ), .C(n374), .D(\x[48] ), .Z(n309)
         );
    VMW_AO22 U204 ( .A(n377), .B(\out[45] ), .C(n374), .D(\x[45] ), .Z(n303)
         );
    VMW_FD \x_reg[11]  ( .D(n433), .CP(Clk), .Q(ScanOut[11]) );
    VMW_FD \x_reg[9]  ( .D(n435), .CP(Clk), .Q(ScanOut[9]) );
    VMW_AO21 U108 ( .A(\x[59] ), .B(n341), .C(n369), .Z(n385) );
    VMW_AO22 U141 ( .A(ScanIn[18]), .B(ScanEnable), .C(\out[50] ), .D(n379), 
        .Z(n360) );
    VMW_AO22 U166 ( .A(n377), .B(\out[62] ), .C(n374), .D(\x[62] ), .Z(n337)
         );
    VMW_FD \x_reg[32]  ( .D(n412), .CP(Clk), .Q(\x[32] ) );
    VMW_FD \x_reg[22]  ( .D(n422), .CP(Clk), .Q(ScanOut[22]) );
    VMW_FD \x_reg[18]  ( .D(n426), .CP(Clk), .Q(ScanOut[18]) );
    VMW_AO22 U183 ( .A(ScanOut[23]), .B(n341), .C(\out[23] ), .D(n379), .Z(
        n324) );
    VMW_FD \x_reg[0]  ( .D(n444), .CP(Clk), .Q(ScanOut[0]) );
    VMW_AO21 U84 ( .A(\x[35] ), .B(n341), .C(n345), .Z(n409) );
    VMW_AO22 U148 ( .A(ScanIn[13]), .B(ScanEnable), .C(\out[45] ), .D(n379), 
        .Z(n355) );
    VMW_AO22 U153 ( .A(ScanIn[8]), .B(ScanEnable), .C(\out[40] ), .D(n379), 
        .Z(n350) );
    VMW_AO22 U174 ( .A(n377), .B(\out[59] ), .C(n374), .D(\x[59] ), .Z(n331)
         );
    VMW_AO22 U191 ( .A(ScanOut[1]), .B(n341), .C(\out[1] ), .D(n379), .Z(n280)
         );
    VMW_FD \x_reg[26]  ( .D(n418), .CP(Clk), .Q(ScanOut[26]) );
    VMW_FD \x_reg[15]  ( .D(n429), .CP(Clk), .Q(ScanOut[15]) );
    VMW_FD \x_reg[4]  ( .D(n440), .CP(Clk), .Q(ScanOut[4]) );
    VMW_OR2 U66 ( .A(n311), .B(n312), .Z(n427) );
    VMW_AO21 U101 ( .A(\x[52] ), .B(n341), .C(n362), .Z(n392) );
    VMW_AO21 U106 ( .A(\x[57] ), .B(n341), .C(n367), .Z(n387) );
    VMW_AO22 U121 ( .A(ScanOut[8]), .B(n341), .C(\out[8] ), .D(n379), .Z(n294)
         );
    VMW_AO22 U126 ( .A(ScanIn[31]), .B(ScanEnable), .C(\out[63] ), .D(n379), 
        .Z(n373) );
    VMW_FD \x_reg[36]  ( .D(n408), .CP(Clk), .Q(\x[36] ) );
    VMW_AO22 U211 ( .A(ScanOut[10]), .B(n341), .C(\out[10] ), .D(n379), .Z(
        n298) );
    VMW_INV U216 ( .A(rdy), .Z(n380) );
    VMW_FD \x_reg[34]  ( .D(n410), .CP(Clk), .Q(\x[34] ) );
    VMW_AO21 U83 ( .A(\x[34] ), .B(n341), .C(n344), .Z(n410) );
    VMW_AO22 U168 ( .A(n377), .B(\out[34] ), .C(n374), .D(\x[34] ), .Z(n281)
         );
    VMW_FD \x_reg[6]  ( .D(n438), .CP(Clk), .Q(ScanOut[6]) );
    VMW_AO21 U98 ( .A(\x[49] ), .B(n341), .C(n359), .Z(n395) );
    VMW_AO22 U128 ( .A(ScanIn[29]), .B(ScanEnable), .C(\out[61] ), .D(n379), 
        .Z(n371) );
    VMW_AO22 U154 ( .A(n377), .B(\out[35] ), .C(n374), .D(\x[35] ), .Z(n283)
         );
    VMW_AO22 U173 ( .A(ScanOut[28]), .B(n341), .C(\out[28] ), .D(n379), .Z(
        n334) );
    VMW_AO22 U184 ( .A(n377), .B(\out[54] ), .C(n374), .D(\x[54] ), .Z(n321)
         );
    VMW_AO22 U196 ( .A(n377), .B(\out[49] ), .C(n374), .D(\x[49] ), .Z(n311)
         );
    VMW_FD \x_reg[17]  ( .D(n427), .CP(Clk), .Q(ScanOut[17]) );
    VMW_FD \x_reg[24]  ( .D(n420), .CP(Clk), .Q(ScanOut[24]) );
    VMW_FD \x_reg[2]  ( .D(n442), .CP(Clk), .Q(ScanOut[2]) );
    VMW_OR2 U53 ( .A(n285), .B(n286), .Z(n440) );
    VMW_AO21 U91 ( .A(\x[42] ), .B(n341), .C(n352), .Z(n402) );
    VMW_AO22 U146 ( .A(ScanIn[15]), .B(ScanEnable), .C(\out[47] ), .D(n379), 
        .Z(n357) );
    VMW_INV U218 ( .A(start), .Z(n376) );
    VMW_FD \x_reg[29]  ( .D(n415), .CP(Clk), .Q(ScanOut[29]) );
    VMW_AO22 U161 ( .A(ScanIn[2]), .B(ScanEnable), .C(\out[34] ), .D(n379), 
        .Z(n344) );
    VMW_FD \x_reg[30]  ( .D(n414), .CP(Clk), .Q(ScanOut[30]) );
    VMW_AO22 U203 ( .A(ScanOut[14]), .B(n341), .C(\out[14] ), .D(n379), .Z(
        n306) );
    VMW_FD \x_reg[39]  ( .D(n405), .CP(Clk), .Q(\x[39] ) );
    VMW_FD \x_reg[20]  ( .D(n424), .CP(Clk), .Q(ScanOut[20]) );
    VMW_FD \x_reg[13]  ( .D(n431), .CP(Clk), .Q(ScanOut[13]) );
    VMW_OR2 U74 ( .A(n327), .B(n328), .Z(n419) );
    VMW_NAND4 U114 ( .A(startflag), .B(rdy), .C(n376), .D(n276), .Z(n375) );
    VMW_AO22 U133 ( .A(ScanIn[26]), .B(ScanEnable), .C(\out[58] ), .D(n379), 
        .Z(n368) );
    VMW_AO21 U82 ( .A(\x[33] ), .B(n341), .C(n343), .Z(n411) );
    VMW_AO21 U99 ( .A(\x[50] ), .B(n341), .C(n360), .Z(n394) );
    VMW_AO22 U197 ( .A(ScanOut[17]), .B(n341), .C(\out[17] ), .D(n379), .Z(
        n312) );
    VMW_FD \x_reg[45]  ( .D(n399), .CP(Clk), .Q(\x[45] ) );
    VMW_AO22 U155 ( .A(ScanOut[3]), .B(n341), .C(\out[3] ), .D(n379), .Z(n284)
         );
    VMW_AO22 U169 ( .A(ScanOut[2]), .B(n341), .C(\out[2] ), .D(n379), .Z(n282)
         );
    VMW_AO22 U172 ( .A(n377), .B(\out[60] ), .C(n374), .D(\x[60] ), .Z(n333)
         );
    VMW_OR2 U49 ( .A(n277), .B(n278), .Z(n444) );
    VMW_OR2 U52 ( .A(n283), .B(n284), .Z(n441) );
    VMW_OR2 U67 ( .A(n313), .B(n314), .Z(n426) );
    VMW_AO21 U107 ( .A(\x[58] ), .B(n341), .C(n368), .Z(n386) );
    VMW_AO22 U120 ( .A(n377), .B(\out[40] ), .C(n374), .D(\x[40] ), .Z(n293)
         );
    VMW_AO22 U210 ( .A(n377), .B(\out[42] ), .C(n374), .D(\x[42] ), .Z(n297)
         );
    VMW_FD \x_reg[55]  ( .D(n389), .CP(Clk), .Q(\x[55] ) );
    VMW_OR2 U75 ( .A(n329), .B(n330), .Z(n418) );
    VMW_AND2 U115 ( .A(n378), .B(ScanEnable), .Z(n377) );
    VMW_AO22 U132 ( .A(ScanIn[27]), .B(ScanEnable), .C(\out[59] ), .D(n379), 
        .Z(n369) );
    VMW_AO22 U202 ( .A(n377), .B(\out[46] ), .C(n374), .D(\x[46] ), .Z(n305)
         );
    VMW_AO21 U90 ( .A(n341), .B(\x[41] ), .C(n351), .Z(n403) );
    VMW_AO22 U129 ( .A(ScanIn[28]), .B(ScanEnable), .C(\out[60] ), .D(n379), 
        .Z(n370) );
    VMW_AO22 U147 ( .A(ScanIn[14]), .B(ScanEnable), .C(\out[46] ), .D(n379), 
        .Z(n356) );
    VMW_FD \x_reg[58]  ( .D(n386), .CP(Clk), .Q(\x[58] ) );
    VMW_FD \x_reg[41]  ( .D(n403), .CP(Clk), .Q(\x[41] ) );
    VMW_AO22 U160 ( .A(ScanIn[3]), .B(ScanEnable), .C(\out[35] ), .D(n379), 
        .Z(n345) );
    VMW_FD \x_reg[62]  ( .D(n382), .CP(Clk), .Q(\x[62] ) );
    VMW_FD \x_reg[51]  ( .D(n393), .CP(Clk), .Q(\x[51] ) );
    VMW_FD \x_reg[48]  ( .D(n396), .CP(Clk), .Q(\x[48] ) );
    VMW_AO22 U185 ( .A(ScanOut[22]), .B(n341), .C(\out[22] ), .D(n379), .Z(
        n322) );
    VMW_OR2 U50 ( .A(n279), .B(n280), .Z(n443) );
    VMW_OR2 U55 ( .A(n289), .B(n290), .Z(n438) );
    VMW_OR2 U69 ( .A(n317), .B(n318), .Z(n424) );
    VMW_AO21 U109 ( .A(\x[60] ), .B(n341), .C(n370), .Z(n384) );
    VMW_AO22 U182 ( .A(n377), .B(\out[55] ), .C(n374), .D(\x[55] ), .Z(n323)
         );
    VMW_OR2 U72 ( .A(n323), .B(n324), .Z(n421) );
    VMW_AO21 U97 ( .A(\x[48] ), .B(n341), .C(n358), .Z(n396) );
    VMW_AO22 U140 ( .A(ScanIn[19]), .B(ScanEnable), .C(\out[51] ), .D(n379), 
        .Z(n361) );
    VMW_AO22 U167 ( .A(ScanOut[30]), .B(n341), .C(\out[30] ), .D(n379), .Z(
        n338) );
    VMW_FD \x_reg[60]  ( .D(n384), .CP(Clk), .Q(\x[60] ) );
    VMW_FD \x_reg[53]  ( .D(n391), .CP(Clk), .Q(\x[53] ) );
    VMW_FD \x_reg[43]  ( .D(n401), .CP(Clk), .Q(\x[43] ) );
    VMW_AO21 U112 ( .A(\x[63] ), .B(n341), .C(n373), .Z(n381) );
    VMW_AO22 U135 ( .A(ScanIn[24]), .B(ScanEnable), .C(\out[56] ), .D(n379), 
        .Z(n366) );
    VMW_AO22 U205 ( .A(ScanOut[13]), .B(n341), .C(\out[13] ), .D(n379), .Z(
        n304) );
    VMW_OR2 U57 ( .A(n293), .B(n294), .Z(n436) );
    VMW_OR2 U60 ( .A(n299), .B(n300), .Z(n433) );
    VMW_AO22 U199 ( .A(ScanOut[16]), .B(n341), .C(\out[16] ), .D(n379), .Z(
        n310) );
    VMW_AO21 U85 ( .A(\x[36] ), .B(n341), .C(n346), .Z(n408) );
    VMW_AO21 U100 ( .A(\x[51] ), .B(n341), .C(n361), .Z(n393) );
    VMW_AO22 U127 ( .A(ScanIn[30]), .B(ScanEnable), .C(\out[62] ), .D(n379), 
        .Z(n372) );
    VMW_FD \x_reg[57]  ( .D(n387), .CP(Clk), .Q(\x[57] ) );
    VMW_AO22 U149 ( .A(ScanIn[12]), .B(ScanEnable), .C(\out[44] ), .D(n379), 
        .Z(n354) );
    VMW_INV U217 ( .A(n375), .Z(n378) );
    VMW_AO22 U137 ( .A(ScanIn[22]), .B(ScanEnable), .C(\out[54] ), .D(n379), 
        .Z(n364) );
    VMW_AO22 U152 ( .A(ScanIn[9]), .B(ScanEnable), .C(n379), .D(\out[41] ), 
        .Z(n351) );
    VMW_AO22 U175 ( .A(ScanOut[27]), .B(n341), .C(\out[27] ), .D(n379), .Z(
        n332) );
    VMW_AO22 U190 ( .A(n377), .B(\out[33] ), .C(n374), .D(\x[33] ), .Z(n279)
         );
    VMW_FD \x_reg[47]  ( .D(n397), .CP(Clk), .Q(\x[47] ) );
    VMW_FD \x_reg[56]  ( .D(n388), .CP(Clk), .Q(\x[56] ) );
    VMW_OR2 U59 ( .A(n297), .B(n298), .Z(n434) );
    VMW_OR2 U62 ( .A(n303), .B(n304), .Z(n431) );
    VMW_OR2 U70 ( .A(n319), .B(n320), .Z(n423) );
    VMW_AO22 U207 ( .A(ScanOut[12]), .B(n341), .C(\out[12] ), .D(n379), .Z(
        n302) );
    VMW_OR2 U79 ( .A(n337), .B(n338), .Z(n414) );
    VMW_AO21 U95 ( .A(\x[46] ), .B(n341), .C(n356), .Z(n398) );
    VMW_AO21 U110 ( .A(\x[61] ), .B(n341), .C(n371), .Z(n383) );
    VMW_AO22 U159 ( .A(ScanIn[4]), .B(ScanEnable), .C(\out[36] ), .D(n379), 
        .Z(n346) );
    VMW_AO22 U119 ( .A(ScanOut[9]), .B(n341), .C(\out[9] ), .D(n379), .Z(n296)
         );
    VMW_AO22 U142 ( .A(n377), .B(\out[36] ), .C(n374), .D(\x[36] ), .Z(n285)
         );
    VMW_AO22 U165 ( .A(ScanOut[31]), .B(n341), .C(\out[31] ), .D(n379), .Z(
        n340) );
    VMW_AO22 U180 ( .A(n377), .B(\out[56] ), .C(n374), .D(\x[56] ), .Z(n325)
         );
    VMW_AO22 U192 ( .A(n377), .B(\out[51] ), .C(n374), .D(\x[51] ), .Z(n315)
         );
    VMW_FD \x_reg[46]  ( .D(n398), .CP(Clk), .Q(\x[46] ) );
    VMW_AO21 U87 ( .A(\x[38] ), .B(n341), .C(n348), .Z(n406) );
    VMW_AO22 U150 ( .A(ScanIn[11]), .B(ScanEnable), .C(\out[43] ), .D(n379), 
        .Z(n353) );
    VMW_AO22 U177 ( .A(ScanOut[26]), .B(n341), .C(\out[26] ), .D(n379), .Z(
        n330) );
    VMW_FD \x_reg[52]  ( .D(n392), .CP(Clk), .Q(\x[52] ) );
    VMW_FD \x_reg[61]  ( .D(n383), .CP(Clk), .Q(\x[61] ) );
    VMW_AO22 U125 ( .A(ScanOut[6]), .B(n341), .C(\out[6] ), .D(n379), .Z(n290)
         );
    VMW_FD \x_reg[42]  ( .D(n402), .CP(Clk), .Q(\x[42] ) );
    VMW_INV U215 ( .A(Reset), .Z(n276) );
    VMW_OR2 U65 ( .A(n309), .B(n310), .Z(n428) );
    VMW_AO21 U102 ( .A(\x[53] ), .B(n341), .C(n363), .Z(n391) );
    VMW_AO21 U105 ( .A(\x[56] ), .B(n341), .C(n366), .Z(n388) );
    VMW_AO22 U189 ( .A(ScanOut[20]), .B(n341), .C(\out[20] ), .D(n379), .Z(
        n318) );
    VMW_OR2 U80 ( .A(n339), .B(n340), .Z(n413) );
    VMW_AO22 U122 ( .A(n377), .B(\out[39] ), .C(n374), .D(\x[39] ), .Z(n291)
         );
    VMW_AO22 U212 ( .A(n377), .B(\out[32] ), .C(n374), .D(\x[32] ), .Z(n277)
         );
    VMW_FD \x_reg[59]  ( .D(n385), .CP(Clk), .Q(\x[59] ) );
    VMW_FD \x_reg[40]  ( .D(n404), .CP(Clk), .Q(\x[40] ) );
    VMW_AO22 U139 ( .A(ScanIn[20]), .B(ScanEnable), .C(\out[52] ), .D(n379), 
        .Z(n362) );
    VMW_AO22 U157 ( .A(ScanIn[6]), .B(ScanEnable), .C(\out[38] ), .D(n379), 
        .Z(n348) );
    VMW_AO22 U170 ( .A(n377), .B(\out[61] ), .C(n374), .D(\x[61] ), .Z(n335)
         );
    VMW_FD \x_reg[50]  ( .D(n394), .CP(Clk), .Q(\x[50] ) );
    VMW_AO22 U195 ( .A(ScanOut[18]), .B(n341), .C(\out[18] ), .D(n379), .Z(
        n314) );
    VMW_FD \x_reg[63]  ( .D(n381), .CP(Clk), .Q(\x[63] ) );
    VMW_FD \x_reg[49]  ( .D(n395), .CP(Clk), .Q(\x[49] ) );
    VMW_OR2 U77 ( .A(n333), .B(n334), .Z(n416) );
    VMW_AO21 U89 ( .A(\x[40] ), .B(n341), .C(n350), .Z(n404) );
    VMW_AO22 U187 ( .A(ScanOut[21]), .B(n341), .C(\out[21] ), .D(n379), .Z(
        n320) );
    VMW_AO22 U209 ( .A(ScanOut[11]), .B(n341), .C(\out[11] ), .D(n379), .Z(
        n300) );
    VMW_FD \x_reg[44]  ( .D(n400), .CP(Clk), .Q(\x[44] ) );
    VMW_AO21 U92 ( .A(\x[43] ), .B(n341), .C(n353), .Z(n401) );
    VMW_AO22 U145 ( .A(ScanIn[16]), .B(ScanEnable), .C(\out[48] ), .D(n379), 
        .Z(n358) );
    VMW_AO22 U162 ( .A(ScanIn[1]), .B(ScanEnable), .C(\out[33] ), .D(n379), 
        .Z(n343) );
    VMW_AO22 U179 ( .A(ScanOut[25]), .B(n341), .C(\out[25] ), .D(n379), .Z(
        n328) );
    VMW_NOR2 U117 ( .A(n378), .B(ScanEnable), .Z(n341) );
    VMW_FD \x_reg[54]  ( .D(n390), .CP(Clk), .Q(\x[54] ) );
    VMW_AO22 U200 ( .A(n377), .B(\out[47] ), .C(n374), .D(\x[47] ), .Z(n307)
         );
    VMW_OR2 U51 ( .A(n281), .B(n282), .Z(n442) );
    VMW_OR2 U58 ( .A(n295), .B(n296), .Z(n435) );
    VMW_AO22 U130 ( .A(n377), .B(\out[37] ), .C(n374), .D(\x[37] ), .Z(n287)
         );
    VMW_AO22 U138 ( .A(ScanIn[21]), .B(ScanEnable), .C(\out[53] ), .D(n379), 
        .Z(n363) );
    VMW_AO22 U194 ( .A(n377), .B(\out[50] ), .C(n374), .D(\x[50] ), .Z(n313)
         );
    VMW_AO22 U208 ( .A(n377), .B(\out[43] ), .C(n374), .D(\x[43] ), .Z(n299)
         );
    VMW_FD \x_reg[3]  ( .D(n441), .CP(Clk), .Q(ScanOut[3]) );
    VMW_OR2 U64 ( .A(n307), .B(n308), .Z(n429) );
    VMW_AO21 U81 ( .A(\x[32] ), .B(n341), .C(n342), .Z(n412) );
    VMW_AO22 U156 ( .A(ScanIn[7]), .B(ScanEnable), .C(\out[39] ), .D(n379), 
        .Z(n349) );
    VMW_AO22 U171 ( .A(ScanOut[29]), .B(n341), .C(\out[29] ), .D(n379), .Z(
        n336) );
    VMW_FD \x_reg[38]  ( .D(n406), .CP(Clk), .Q(\x[38] ) );
    VMW_FD \x_reg[31]  ( .D(n413), .CP(Clk), .Q(ScanOut[31]) );
    VMW_FD \x_reg[28]  ( .D(n416), .CP(Clk), .Q(ScanOut[28]) );
    VMW_FD \x_reg[12]  ( .D(n432), .CP(Clk), .Q(ScanOut[12]) );
    VMW_FD \x_reg[21]  ( .D(n423), .CP(Clk), .Q(ScanOut[21]) );
    VMW_AO21 U104 ( .A(\x[55] ), .B(n341), .C(n365), .Z(n389) );
    VMW_OR2 U76 ( .A(n331), .B(n332), .Z(n417) );
    VMW_NOR2 U116 ( .A(n341), .B(ScanEnable), .Z(n379) );
    VMW_AO22 U123 ( .A(ScanOut[7]), .B(n341), .C(\out[7] ), .D(n379), .Z(n292)
         );
    VMW_AO22 U213 ( .A(ScanOut[0]), .B(n341), .C(\out[0] ), .D(n379), .Z(n278)
         );
    VMW_FD startflag_reg ( .D(n445), .CP(Clk), .Q(startflag) );
    VMW_FD \x_reg[35]  ( .D(n409), .CP(Clk), .Q(\x[35] ) );
    VMW_OR2 U56 ( .A(n291), .B(n292), .Z(n437) );
    VMW_AO21 U88 ( .A(\x[39] ), .B(n341), .C(n349), .Z(n405) );
    VMW_AO21 U93 ( .A(\x[44] ), .B(n341), .C(n354), .Z(n400) );
    VMW_AO22 U131 ( .A(ScanOut[5]), .B(n341), .C(\out[5] ), .D(n379), .Z(n288)
         );
    VMW_AO22 U201 ( .A(ScanOut[15]), .B(n341), .C(\out[15] ), .D(n379), .Z(
        n308) );
    VMW_AO22 U178 ( .A(n377), .B(\out[57] ), .C(n374), .D(\x[57] ), .Z(n327)
         );
    VMW_FD \x_reg[7]  ( .D(n437), .CP(Clk), .Q(ScanOut[7]) );
    VMW_AO21 U94 ( .A(\x[45] ), .B(n341), .C(n355), .Z(n399) );
    VMW_AO22 U143 ( .A(ScanOut[4]), .B(n341), .C(\out[4] ), .D(n379), .Z(n286)
         );
    VMW_AO22 U144 ( .A(ScanIn[17]), .B(ScanEnable), .C(\out[49] ), .D(n379), 
        .Z(n359) );
    VMW_AO22 U163 ( .A(ScanIn[0]), .B(ScanEnable), .C(\out[32] ), .D(n379), 
        .Z(n342) );
    VMW_AO22 U181 ( .A(ScanOut[24]), .B(n341), .C(\out[24] ), .D(n379), .Z(
        n326) );
    VMW_AO22 U186 ( .A(n377), .B(\out[53] ), .C(n374), .D(\x[53] ), .Z(n319)
         );
    VMW_FD \x_reg[25]  ( .D(n419), .CP(Clk), .Q(ScanOut[25]) );
    VMW_FD \x_reg[16]  ( .D(n428), .CP(Clk), .Q(ScanOut[16]) );
    VMW_FD \x_reg[27]  ( .D(n417), .CP(Clk), .Q(ScanOut[27]) );
    VMW_FD \x_reg[14]  ( .D(n430), .CP(Clk), .Q(ScanOut[14]) );
    VMW_AO22 U158 ( .A(ScanIn[5]), .B(ScanEnable), .C(\out[37] ), .D(n379), 
        .Z(n347) );
    VMW_AO22 U164 ( .A(n377), .B(\out[63] ), .C(n374), .D(\x[63] ), .Z(n339)
         );
    VMW_FD \x_reg[5]  ( .D(n439), .CP(Clk), .Q(ScanOut[5]) );
    VMW_AO22 U136 ( .A(ScanIn[23]), .B(ScanEnable), .C(\out[55] ), .D(n379), 
        .Z(n365) );
    VMW_FD \x_reg[37]  ( .D(n407), .CP(Clk), .Q(\x[37] ) );
    VMW_AO22 U206 ( .A(n377), .B(\out[44] ), .C(n374), .D(\x[44] ), .Z(n301)
         );
    VMW_OR2 U63 ( .A(n305), .B(n306), .Z(n430) );
    VMW_OR2 U71 ( .A(n321), .B(n322), .Z(n422) );
    VMW_AO21 U111 ( .A(\x[62] ), .B(n341), .C(n372), .Z(n382) );
    VMW_AO22 U124 ( .A(n377), .B(\out[38] ), .C(n374), .D(\x[38] ), .Z(n289)
         );
    VMW_AO21 U214 ( .A(n380), .B(startflag), .C(start), .Z(n275) );
    VMW_OR2 U78 ( .A(n335), .B(n336), .Z(n415) );
    VMW_AO21 U86 ( .A(\x[37] ), .B(n341), .C(n347), .Z(n407) );
    VMW_AO21 U103 ( .A(\x[54] ), .B(n341), .C(n364), .Z(n390) );
    VMW_AO22 U188 ( .A(n377), .B(\out[52] ), .C(n374), .D(\x[52] ), .Z(n317)
         );
    VMW_FD \x_reg[8]  ( .D(n436), .CP(Clk), .Q(ScanOut[8]) );
    VMW_AO22 U118 ( .A(n377), .B(\out[41] ), .C(n374), .D(\x[41] ), .Z(n295)
         );
    VMW_AO22 U151 ( .A(ScanIn[10]), .B(ScanEnable), .C(\out[42] ), .D(n379), 
        .Z(n352) );
    VMW_FD \x_reg[23]  ( .D(n421), .CP(Clk), .Q(ScanOut[23]) );
    VMW_FD \x_reg[10]  ( .D(n434), .CP(Clk), .Q(ScanOut[10]) );
    VMW_AO22 U176 ( .A(n377), .B(\out[58] ), .C(n374), .D(\x[58] ), .Z(n329)
         );
    VMW_FD \x_reg[33]  ( .D(n411), .CP(Clk), .Q(\x[33] ) );
    VMW_AO22 U193 ( .A(ScanOut[19]), .B(n341), .C(\out[19] ), .D(n379), .Z(
        n316) );
    VMW_FD \x_reg[19]  ( .D(n425), .CP(Clk), .Q(ScanOut[19]) );
    VMW_FD \x_reg[1]  ( .D(n443), .CP(Clk), .Q(ScanOut[1]) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \ScanLink0[13] , \key[38] , \ScanLink0[20] , \key[21] , \key[12] , 
        \ScanLink1[19] , \key[2] , \ScanLink1[23] , \ScanLink1[10] , 
        \ScanLink1[7] , \ScanLink0[30] , \ScanLink0[29] , \key[31] , \key[28] , 
        \key[25] , \key[16] , \ScanEnable[0] , \ScanLink0[17] , 
        \ScanLink0[24] , \key[35] , \ScanLink1[27] , \ScanLink1[14] , 
        \ScanLink1[3] , \key[37] , \key[6] , \key[4] , \ScanLink1[25] , 
        \ScanLink1[16] , \ScanLink1[1] , \key[27] , \key[14] , \ScanLink0[15] , 
        \ScanLink0[26] , \ScanLink1[8] , \ScanLink0[18] , \key[33] , \key[19] , 
        \key[9] , \key[0] , \ScanLink1[31] , \ScanLink1[28] , \ScanLink1[21] , 
        \ScanLink1[12] , \ScanLink1[5] , \ScanLink0[11] , \ScanLink0[22] , 
        \key[23] , \key[10] , \key[46] , \ScanLink0[1] , \key[56] , 
        \ScanLink0[8] , \key[42] , \ScanLink0[5] , \key[61] , \key[52] , 
        \key[63] , \key[50] , \key[49] , \key[59] , \key[54] , \key[40] , 
        \ScanLink0[7] , \key[44] , \ScanLink0[3] , \key[55] , \key[45] , 
        \ScanLink0[2] , \key[62] , \key[51] , \key[48] , \key[58] , \key[41] , 
        \ScanLink0[6] , \key[43] , \ScanLink0[4] , \key[60] , \key[53] , rdy1, 
        \key[47] , \ScanLink0[0] , \key[57] , \ScanLink0[9] , \key[32] , 
        \key[18] , \ScanLink0[19] , \key[8] , \key[1] , \ScanLink1[20] , 
        \ScanLink1[13] , \ScanLink1[4] , \ScanLink1[30] , \ScanLink1[29] , 
        \ScanLink0[10] , \key[22] , \ScanLink0[23] , \key[11] , \key[5] , 
        \ScanLink1[24] , \ScanLink1[17] , \ScanLink1[0] , \key[36] , \key[26] , 
        \key[15] , \ScanLink0[14] , \ScanLink0[27] , \ScanLink1[9] , \key[24] , 
        \key[17] , \ScanLink0[16] , \key[34] , \ScanLink0[25] , \key[7] , 
        \ScanLink1[26] , \ScanLink1[15] , \ScanLink1[2] , \ScanLink0[12] , 
        \ScanLink0[21] , \key[39] , \key[20] , \key[13] , \key[30] , \key[29] , 
        \key[3] , \start[0] , \ScanLink1[18] , \ScanLink1[11] , \ScanLink1[6] , 
        \ScanLink1[22] , \ScanLink0[31] , \ScanLink0[28] ;
    DES_Control_WIDTH64_MEMSPACE2_IDWIDTH1_SCAN1 U_DES_Control_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanOut({\ScanLink1[31] , 
        \ScanLink1[30] , \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , 
        \ScanLink1[26] , \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , 
        \ScanLink1[22] , \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , 
        \ScanLink1[18] , \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , 
        \ScanLink1[14] , \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , 
        \ScanLink1[10] , \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , 
        \ScanLink1[6] , \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , 
        \ScanLink1[2] , \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(
        \ScanEnable[0] ), .ScanId(1'b1), .Id(1'b0), .key({\key[63] , \key[62] , 
        \key[61] , \key[60] , \key[59] , \key[58] , \key[57] , \key[56] , 
        \key[55] , \key[54] , \key[53] , \key[52] , \key[51] , \key[50] , 
        \key[49] , \key[48] , \key[47] , \key[46] , \key[45] , \key[44] , 
        \key[43] , \key[42] , \key[41] , \key[40] , \key[39] , \key[38] , 
        \key[37] , \key[36] , \key[35] , \key[34] , \key[33] , \key[32] , 
        \key[31] , \key[30] , \key[29] , \key[28] , \key[27] , \key[26] , 
        \key[25] , \key[24] , \key[23] , \key[22] , \key[21] , \key[20] , 
        \key[19] , \key[18] , \key[17] , \key[16] , \key[15] , \key[14] , 
        \key[13] , \key[12] , \key[11] , \key[10] , \key[9] , \key[8] , 
        \key[7] , \key[6] , \key[5] , \key[4] , \key[3] , \key[2] , \key[1] , 
        \key[0] }), .start(\start[0] ), .rdy(rdy1) );
    DES_Node_WIDTH64_MEMSPACE2_IDWIDTH1_SCAN1 U_DES_Node_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanOut({\ScanLink0[31] , 
        \ScanLink0[30] , \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , 
        \ScanLink0[26] , \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , 
        \ScanLink0[22] , \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , 
        \ScanLink0[18] , \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , 
        \ScanLink0[14] , \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , 
        \ScanLink0[10] , \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , 
        \ScanLink0[6] , \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , 
        \ScanLink0[2] , \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .key({\key[63] , \key[62] , \key[61] , 
        \key[60] , \key[59] , \key[58] , \key[57] , \key[56] , \key[55] , 
        \key[54] , \key[53] , \key[52] , \key[51] , \key[50] , \key[49] , 
        \key[48] , \key[47] , \key[46] , \key[45] , \key[44] , \key[43] , 
        \key[42] , \key[41] , \key[40] , \key[39] , \key[38] , \key[37] , 
        \key[36] , \key[35] , \key[34] , \key[33] , \key[32] , \key[31] , 
        \key[30] , \key[29] , \key[28] , \key[27] , \key[26] , \key[25] , 
        \key[24] , \key[23] , \key[22] , \key[21] , \key[20] , \key[19] , 
        \key[18] , \key[17] , \key[16] , \key[15] , \key[14] , \key[13] , 
        \key[12] , \key[11] , \key[10] , \key[9] , \key[8] , \key[7] , 
        \key[6] , \key[5] , \key[4] , \key[3] , \key[2] , \key[1] , \key[0] }), 
        .start(\start[0] ), .rdy(rdy1) );
endmodule

